module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    reg [161:0] src32;
    reg [161:0] src33;
    reg [161:0] src34;
    reg [161:0] src35;
    reg [161:0] src36;
    reg [161:0] src37;
    reg [161:0] src38;
    reg [161:0] src39;
    reg [161:0] src40;
    reg [161:0] src41;
    reg [161:0] src42;
    reg [161:0] src43;
    reg [161:0] src44;
    reg [161:0] src45;
    reg [161:0] src46;
    reg [161:0] src47;
    reg [161:0] src48;
    reg [161:0] src49;
    reg [161:0] src50;
    reg [161:0] src51;
    reg [161:0] src52;
    reg [161:0] src53;
    reg [161:0] src54;
    reg [161:0] src55;
    reg [161:0] src56;
    reg [161:0] src57;
    reg [161:0] src58;
    reg [161:0] src59;
    reg [161:0] src60;
    reg [161:0] src61;
    reg [161:0] src62;
    reg [161:0] src63;
    compressor2_1_162_64 compressor2_1_162_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
        src12 <= 162'h0;
        src13 <= 162'h0;
        src14 <= 162'h0;
        src15 <= 162'h0;
        src16 <= 162'h0;
        src17 <= 162'h0;
        src18 <= 162'h0;
        src19 <= 162'h0;
        src20 <= 162'h0;
        src21 <= 162'h0;
        src22 <= 162'h0;
        src23 <= 162'h0;
        src24 <= 162'h0;
        src25 <= 162'h0;
        src26 <= 162'h0;
        src27 <= 162'h0;
        src28 <= 162'h0;
        src29 <= 162'h0;
        src30 <= 162'h0;
        src31 <= 162'h0;
        src32 <= 162'h0;
        src33 <= 162'h0;
        src34 <= 162'h0;
        src35 <= 162'h0;
        src36 <= 162'h0;
        src37 <= 162'h0;
        src38 <= 162'h0;
        src39 <= 162'h0;
        src40 <= 162'h0;
        src41 <= 162'h0;
        src42 <= 162'h0;
        src43 <= 162'h0;
        src44 <= 162'h0;
        src45 <= 162'h0;
        src46 <= 162'h0;
        src47 <= 162'h0;
        src48 <= 162'h0;
        src49 <= 162'h0;
        src50 <= 162'h0;
        src51 <= 162'h0;
        src52 <= 162'h0;
        src53 <= 162'h0;
        src54 <= 162'h0;
        src55 <= 162'h0;
        src56 <= 162'h0;
        src57 <= 162'h0;
        src58 <= 162'h0;
        src59 <= 162'h0;
        src60 <= 162'h0;
        src61 <= 162'h0;
        src62 <= 162'h0;
        src63 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor2_1_162_64(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    input [161:0]src12,
    input [161:0]src13,
    input [161:0]src14,
    input [161:0]src15,
    input [161:0]src16,
    input [161:0]src17,
    input [161:0]src18,
    input [161:0]src19,
    input [161:0]src20,
    input [161:0]src21,
    input [161:0]src22,
    input [161:0]src23,
    input [161:0]src24,
    input [161:0]src25,
    input [161:0]src26,
    input [161:0]src27,
    input [161:0]src28,
    input [161:0]src29,
    input [161:0]src30,
    input [161:0]src31,
    input [161:0]src32,
    input [161:0]src33,
    input [161:0]src34,
    input [161:0]src35,
    input [161:0]src36,
    input [161:0]src37,
    input [161:0]src38,
    input [161:0]src39,
    input [161:0]src40,
    input [161:0]src41,
    input [161:0]src42,
    input [161:0]src43,
    input [161:0]src44,
    input [161:0]src45,
    input [161:0]src46,
    input [161:0]src47,
    input [161:0]src48,
    input [161:0]src49,
    input [161:0]src50,
    input [161:0]src51,
    input [161:0]src52,
    input [161:0]src53,
    input [161:0]src54,
    input [161:0]src55,
    input [161:0]src56,
    input [161:0]src57,
    input [161:0]src58,
    input [161:0]src59,
    input [161:0]src60,
    input [161:0]src61,
    input [161:0]src62,
    input [161:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [0:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [0:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [0:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [0:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [0:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [0:0] comp_out70;
    wire [0:0] comp_out71;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71)
    );
    rowadder2_1_72 rowadder2_1inst(
        .src0({comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], 1'h0, comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], 1'h0, comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], 1'h0, comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], 1'h0, comp_out4[1], 1'h0, 1'h0, 1'h0, comp_out0[1]}),
        .dst0({dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      input wire [161:0] src16,
      input wire [161:0] src17,
      input wire [161:0] src18,
      input wire [161:0] src19,
      input wire [161:0] src20,
      input wire [161:0] src21,
      input wire [161:0] src22,
      input wire [161:0] src23,
      input wire [161:0] src24,
      input wire [161:0] src25,
      input wire [161:0] src26,
      input wire [161:0] src27,
      input wire [161:0] src28,
      input wire [161:0] src29,
      input wire [161:0] src30,
      input wire [161:0] src31,
      input wire [161:0] src32,
      input wire [161:0] src33,
      input wire [161:0] src34,
      input wire [161:0] src35,
      input wire [161:0] src36,
      input wire [161:0] src37,
      input wire [161:0] src38,
      input wire [161:0] src39,
      input wire [161:0] src40,
      input wire [161:0] src41,
      input wire [161:0] src42,
      input wire [161:0] src43,
      input wire [161:0] src44,
      input wire [161:0] src45,
      input wire [161:0] src46,
      input wire [161:0] src47,
      input wire [161:0] src48,
      input wire [161:0] src49,
      input wire [161:0] src50,
      input wire [161:0] src51,
      input wire [161:0] src52,
      input wire [161:0] src53,
      input wire [161:0] src54,
      input wire [161:0] src55,
      input wire [161:0] src56,
      input wire [161:0] src57,
      input wire [161:0] src58,
      input wire [161:0] src59,
      input wire [161:0] src60,
      input wire [161:0] src61,
      input wire [161:0] src62,
      input wire [161:0] src63,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [0:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [0:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [0:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [0:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [0:0] dst70,
      output wire [0:0] dst71);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [161:0] stage0_16;
   wire [161:0] stage0_17;
   wire [161:0] stage0_18;
   wire [161:0] stage0_19;
   wire [161:0] stage0_20;
   wire [161:0] stage0_21;
   wire [161:0] stage0_22;
   wire [161:0] stage0_23;
   wire [161:0] stage0_24;
   wire [161:0] stage0_25;
   wire [161:0] stage0_26;
   wire [161:0] stage0_27;
   wire [161:0] stage0_28;
   wire [161:0] stage0_29;
   wire [161:0] stage0_30;
   wire [161:0] stage0_31;
   wire [161:0] stage0_32;
   wire [161:0] stage0_33;
   wire [161:0] stage0_34;
   wire [161:0] stage0_35;
   wire [161:0] stage0_36;
   wire [161:0] stage0_37;
   wire [161:0] stage0_38;
   wire [161:0] stage0_39;
   wire [161:0] stage0_40;
   wire [161:0] stage0_41;
   wire [161:0] stage0_42;
   wire [161:0] stage0_43;
   wire [161:0] stage0_44;
   wire [161:0] stage0_45;
   wire [161:0] stage0_46;
   wire [161:0] stage0_47;
   wire [161:0] stage0_48;
   wire [161:0] stage0_49;
   wire [161:0] stage0_50;
   wire [161:0] stage0_51;
   wire [161:0] stage0_52;
   wire [161:0] stage0_53;
   wire [161:0] stage0_54;
   wire [161:0] stage0_55;
   wire [161:0] stage0_56;
   wire [161:0] stage0_57;
   wire [161:0] stage0_58;
   wire [161:0] stage0_59;
   wire [161:0] stage0_60;
   wire [161:0] stage0_61;
   wire [161:0] stage0_62;
   wire [161:0] stage0_63;
   wire [33:0] stage1_0;
   wire [46:0] stage1_1;
   wire [54:0] stage1_2;
   wire [83:0] stage1_3;
   wire [82:0] stage1_4;
   wire [114:0] stage1_5;
   wire [57:0] stage1_6;
   wire [70:0] stage1_7;
   wire [80:0] stage1_8;
   wire [57:0] stage1_9;
   wire [94:0] stage1_10;
   wire [80:0] stage1_11;
   wire [66:0] stage1_12;
   wire [86:0] stage1_13;
   wire [61:0] stage1_14;
   wire [97:0] stage1_15;
   wire [67:0] stage1_16;
   wire [113:0] stage1_17;
   wire [62:0] stage1_18;
   wire [70:0] stage1_19;
   wire [67:0] stage1_20;
   wire [70:0] stage1_21;
   wire [66:0] stage1_22;
   wire [142:0] stage1_23;
   wire [82:0] stage1_24;
   wire [84:0] stage1_25;
   wire [71:0] stage1_26;
   wire [73:0] stage1_27;
   wire [76:0] stage1_28;
   wire [80:0] stage1_29;
   wire [106:0] stage1_30;
   wire [96:0] stage1_31;
   wire [86:0] stage1_32;
   wire [89:0] stage1_33;
   wire [55:0] stage1_34;
   wire [59:0] stage1_35;
   wire [82:0] stage1_36;
   wire [127:0] stage1_37;
   wire [65:0] stage1_38;
   wire [67:0] stage1_39;
   wire [81:0] stage1_40;
   wire [73:0] stage1_41;
   wire [95:0] stage1_42;
   wire [137:0] stage1_43;
   wire [45:0] stage1_44;
   wire [92:0] stage1_45;
   wire [63:0] stage1_46;
   wire [57:0] stage1_47;
   wire [71:0] stage1_48;
   wire [86:0] stage1_49;
   wire [57:0] stage1_50;
   wire [93:0] stage1_51;
   wire [76:0] stage1_52;
   wire [65:0] stage1_53;
   wire [57:0] stage1_54;
   wire [97:0] stage1_55;
   wire [79:0] stage1_56;
   wire [71:0] stage1_57;
   wire [73:0] stage1_58;
   wire [79:0] stage1_59;
   wire [66:0] stage1_60;
   wire [90:0] stage1_61;
   wire [86:0] stage1_62;
   wire [62:0] stage1_63;
   wire [44:0] stage1_64;
   wire [23:0] stage1_65;
   wire [9:0] stage2_0;
   wire [18:0] stage2_1;
   wire [37:0] stage2_2;
   wire [22:0] stage2_3;
   wire [47:0] stage2_4;
   wire [35:0] stage2_5;
   wire [28:0] stage2_6;
   wire [40:0] stage2_7;
   wire [60:0] stage2_8;
   wire [25:0] stage2_9;
   wire [40:0] stage2_10;
   wire [38:0] stage2_11;
   wire [30:0] stage2_12;
   wire [44:0] stage2_13;
   wire [73:0] stage2_14;
   wire [36:0] stage2_15;
   wire [46:0] stage2_16;
   wire [39:0] stage2_17;
   wire [42:0] stage2_18;
   wire [50:0] stage2_19;
   wire [57:0] stage2_20;
   wire [39:0] stage2_21;
   wire [30:0] stage2_22;
   wire [46:0] stage2_23;
   wire [45:0] stage2_24;
   wire [36:0] stage2_25;
   wire [52:0] stage2_26;
   wire [49:0] stage2_27;
   wire [34:0] stage2_28;
   wire [49:0] stage2_29;
   wire [49:0] stage2_30;
   wire [38:0] stage2_31;
   wire [55:0] stage2_32;
   wire [27:0] stage2_33;
   wire [34:0] stage2_34;
   wire [44:0] stage2_35;
   wire [36:0] stage2_36;
   wire [41:0] stage2_37;
   wire [32:0] stage2_38;
   wire [33:0] stage2_39;
   wire [40:0] stage2_40;
   wire [55:0] stage2_41;
   wire [61:0] stage2_42;
   wire [51:0] stage2_43;
   wire [65:0] stage2_44;
   wire [25:0] stage2_45;
   wire [32:0] stage2_46;
   wire [45:0] stage2_47;
   wire [23:0] stage2_48;
   wire [36:0] stage2_49;
   wire [40:0] stage2_50;
   wire [24:0] stage2_51;
   wire [33:0] stage2_52;
   wire [50:0] stage2_53;
   wire [27:0] stage2_54;
   wire [37:0] stage2_55;
   wire [52:0] stage2_56;
   wire [29:0] stage2_57;
   wire [32:0] stage2_58;
   wire [80:0] stage2_59;
   wire [21:0] stage2_60;
   wire [66:0] stage2_61;
   wire [34:0] stage2_62;
   wire [37:0] stage2_63;
   wire [45:0] stage2_64;
   wire [12:0] stage2_65;
   wire [9:0] stage2_66;
   wire [1:0] stage2_67;
   wire [7:0] stage3_0;
   wire [13:0] stage3_1;
   wire [10:0] stage3_2;
   wire [13:0] stage3_3;
   wire [13:0] stage3_4;
   wire [17:0] stage3_5;
   wire [19:0] stage3_6;
   wire [16:0] stage3_7;
   wire [16:0] stage3_8;
   wire [20:0] stage3_9;
   wire [14:0] stage3_10;
   wire [17:0] stage3_11;
   wire [23:0] stage3_12;
   wire [19:0] stage3_13;
   wire [35:0] stage3_14;
   wire [36:0] stage3_15;
   wire [21:0] stage3_16;
   wire [16:0] stage3_17;
   wire [22:0] stage3_18;
   wire [26:0] stage3_19;
   wire [22:0] stage3_20;
   wire [24:0] stage3_21;
   wire [26:0] stage3_22;
   wire [11:0] stage3_23;
   wire [25:0] stage3_24;
   wire [21:0] stage3_25;
   wire [15:0] stage3_26;
   wire [18:0] stage3_27;
   wire [19:0] stage3_28;
   wire [23:0] stage3_29;
   wire [25:0] stage3_30;
   wire [20:0] stage3_31;
   wire [34:0] stage3_32;
   wire [14:0] stage3_33;
   wire [22:0] stage3_34;
   wire [25:0] stage3_35;
   wire [16:0] stage3_36;
   wire [11:0] stage3_37;
   wire [13:0] stage3_38;
   wire [23:0] stage3_39;
   wire [23:0] stage3_40;
   wire [24:0] stage3_41;
   wire [25:0] stage3_42;
   wire [20:0] stage3_43;
   wire [30:0] stage3_44;
   wire [17:0] stage3_45;
   wire [16:0] stage3_46;
   wire [23:0] stage3_47;
   wire [15:0] stage3_48;
   wire [13:0] stage3_49;
   wire [31:0] stage3_50;
   wire [13:0] stage3_51;
   wire [23:0] stage3_52;
   wire [15:0] stage3_53;
   wire [15:0] stage3_54;
   wire [17:0] stage3_55;
   wire [30:0] stage3_56;
   wire [12:0] stage3_57;
   wire [32:0] stage3_58;
   wire [27:0] stage3_59;
   wire [14:0] stage3_60;
   wire [24:0] stage3_61;
   wire [20:0] stage3_62;
   wire [17:0] stage3_63;
   wire [28:0] stage3_64;
   wire [13:0] stage3_65;
   wire [8:0] stage3_66;
   wire [4:0] stage3_67;
   wire [1:0] stage3_68;
   wire [3:0] stage4_0;
   wire [3:0] stage4_1;
   wire [6:0] stage4_2;
   wire [4:0] stage4_3;
   wire [8:0] stage4_4;
   wire [8:0] stage4_5;
   wire [13:0] stage4_6;
   wire [7:0] stage4_7;
   wire [9:0] stage4_8;
   wire [6:0] stage4_9;
   wire [8:0] stage4_10;
   wire [6:0] stage4_11;
   wire [8:0] stage4_12;
   wire [9:0] stage4_13;
   wire [10:0] stage4_14;
   wire [16:0] stage4_15;
   wire [12:0] stage4_16;
   wire [16:0] stage4_17;
   wire [5:0] stage4_18;
   wire [15:0] stage4_19;
   wire [10:0] stage4_20;
   wire [7:0] stage4_21;
   wire [13:0] stage4_22;
   wire [9:0] stage4_23;
   wire [17:0] stage4_24;
   wire [5:0] stage4_25;
   wire [7:0] stage4_26;
   wire [6:0] stage4_27;
   wire [11:0] stage4_28;
   wire [9:0] stage4_29;
   wire [15:0] stage4_30;
   wire [8:0] stage4_31;
   wire [19:0] stage4_32;
   wire [11:0] stage4_33;
   wire [10:0] stage4_34;
   wire [10:0] stage4_35;
   wire [9:0] stage4_36;
   wire [5:0] stage4_37;
   wire [5:0] stage4_38;
   wire [9:0] stage4_39;
   wire [13:0] stage4_40;
   wire [16:0] stage4_41;
   wire [16:0] stage4_42;
   wire [6:0] stage4_43;
   wire [12:0] stage4_44;
   wire [8:0] stage4_45;
   wire [17:0] stage4_46;
   wire [15:0] stage4_47;
   wire [11:0] stage4_48;
   wire [12:0] stage4_49;
   wire [6:0] stage4_50;
   wire [8:0] stage4_51;
   wire [8:0] stage4_52;
   wire [14:0] stage4_53;
   wire [9:0] stage4_54;
   wire [16:0] stage4_55;
   wire [12:0] stage4_56;
   wire [5:0] stage4_57;
   wire [20:0] stage4_58;
   wire [16:0] stage4_59;
   wire [15:0] stage4_60;
   wire [16:0] stage4_61;
   wire [7:0] stage4_62;
   wire [12:0] stage4_63;
   wire [21:0] stage4_64;
   wire [5:0] stage4_65;
   wire [12:0] stage4_66;
   wire [6:0] stage4_67;
   wire [1:0] stage4_68;
   wire [1:0] stage5_0;
   wire [0:0] stage5_1;
   wire [4:0] stage5_2;
   wire [4:0] stage5_3;
   wire [4:0] stage5_4;
   wire [4:0] stage5_5;
   wire [9:0] stage5_6;
   wire [3:0] stage5_7;
   wire [7:0] stage5_8;
   wire [2:0] stage5_9;
   wire [4:0] stage5_10;
   wire [2:0] stage5_11;
   wire [10:0] stage5_12;
   wire [5:0] stage5_13;
   wire [7:0] stage5_14;
   wire [7:0] stage5_15;
   wire [8:0] stage5_16;
   wire [4:0] stage5_17;
   wire [5:0] stage5_18;
   wire [6:0] stage5_19;
   wire [3:0] stage5_20;
   wire [5:0] stage5_21;
   wire [10:0] stage5_22;
   wire [6:0] stage5_23;
   wire [9:0] stage5_24;
   wire [2:0] stage5_25;
   wire [2:0] stage5_26;
   wire [3:0] stage5_27;
   wire [4:0] stage5_28;
   wire [3:0] stage5_29;
   wire [4:0] stage5_30;
   wire [5:0] stage5_31;
   wire [11:0] stage5_32;
   wire [4:0] stage5_33;
   wire [7:0] stage5_34;
   wire [3:0] stage5_35;
   wire [4:0] stage5_36;
   wire [3:0] stage5_37;
   wire [1:0] stage5_38;
   wire [5:0] stage5_39;
   wire [5:0] stage5_40;
   wire [12:0] stage5_41;
   wire [4:0] stage5_42;
   wire [3:0] stage5_43;
   wire [5:0] stage5_44;
   wire [4:0] stage5_45;
   wire [5:0] stage5_46;
   wire [12:0] stage5_47;
   wire [3:0] stage5_48;
   wire [6:0] stage5_49;
   wire [4:0] stage5_50;
   wire [3:0] stage5_51;
   wire [5:0] stage5_52;
   wire [6:0] stage5_53;
   wire [8:0] stage5_54;
   wire [6:0] stage5_55;
   wire [4:0] stage5_56;
   wire [5:0] stage5_57;
   wire [5:0] stage5_58;
   wire [5:0] stage5_59;
   wire [8:0] stage5_60;
   wire [10:0] stage5_61;
   wire [5:0] stage5_62;
   wire [11:0] stage5_63;
   wire [10:0] stage5_64;
   wire [3:0] stage5_65;
   wire [4:0] stage5_66;
   wire [3:0] stage5_67;
   wire [4:0] stage5_68;
   wire [0:0] stage5_69;
   wire [1:0] stage6_0;
   wire [0:0] stage6_1;
   wire [4:0] stage6_2;
   wire [0:0] stage6_3;
   wire [4:0] stage6_4;
   wire [0:0] stage6_5;
   wire [2:0] stage6_6;
   wire [4:0] stage6_7;
   wire [1:0] stage6_8;
   wire [2:0] stage6_9;
   wire [6:0] stage6_10;
   wire [2:0] stage6_11;
   wire [5:0] stage6_12;
   wire [1:0] stage6_13;
   wire [3:0] stage6_14;
   wire [3:0] stage6_15;
   wire [5:0] stage6_16;
   wire [6:0] stage6_17;
   wire [0:0] stage6_18;
   wire [3:0] stage6_19;
   wire [2:0] stage6_20;
   wire [5:0] stage6_21;
   wire [3:0] stage6_22;
   wire [2:0] stage6_23;
   wire [2:0] stage6_24;
   wire [2:0] stage6_25;
   wire [2:0] stage6_26;
   wire [1:0] stage6_27;
   wire [2:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [8:0] stage6_32;
   wire [2:0] stage6_33;
   wire [2:0] stage6_34;
   wire [1:0] stage6_35;
   wire [6:0] stage6_36;
   wire [4:0] stage6_37;
   wire [0:0] stage6_38;
   wire [1:0] stage6_39;
   wire [1:0] stage6_40;
   wire [3:0] stage6_41;
   wire [7:0] stage6_42;
   wire [1:0] stage6_43;
   wire [1:0] stage6_44;
   wire [2:0] stage6_45;
   wire [1:0] stage6_46;
   wire [4:0] stage6_47;
   wire [5:0] stage6_48;
   wire [2:0] stage6_49;
   wire [3:0] stage6_50;
   wire [1:0] stage6_51;
   wire [3:0] stage6_52;
   wire [4:0] stage6_53;
   wire [2:0] stage6_54;
   wire [2:0] stage6_55;
   wire [4:0] stage6_56;
   wire [1:0] stage6_57;
   wire [1:0] stage6_58;
   wire [2:0] stage6_59;
   wire [4:0] stage6_60;
   wire [2:0] stage6_61;
   wire [3:0] stage6_62;
   wire [3:0] stage6_63;
   wire [3:0] stage6_64;
   wire [3:0] stage6_65;
   wire [2:0] stage6_66;
   wire [5:0] stage6_67;
   wire [5:0] stage6_68;
   wire [0:0] stage6_69;
   wire [1:0] stage7_0;
   wire [0:0] stage7_1;
   wire [0:0] stage7_2;
   wire [0:0] stage7_3;
   wire [1:0] stage7_4;
   wire [0:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage7_24;
   wire [1:0] stage7_25;
   wire [0:0] stage7_26;
   wire [1:0] stage7_27;
   wire [1:0] stage7_28;
   wire [1:0] stage7_29;
   wire [1:0] stage7_30;
   wire [1:0] stage7_31;
   wire [1:0] stage7_32;
   wire [1:0] stage7_33;
   wire [1:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [1:0] stage7_38;
   wire [1:0] stage7_39;
   wire [0:0] stage7_40;
   wire [1:0] stage7_41;
   wire [1:0] stage7_42;
   wire [1:0] stage7_43;
   wire [1:0] stage7_44;
   wire [1:0] stage7_45;
   wire [1:0] stage7_46;
   wire [1:0] stage7_47;
   wire [1:0] stage7_48;
   wire [1:0] stage7_49;
   wire [1:0] stage7_50;
   wire [1:0] stage7_51;
   wire [1:0] stage7_52;
   wire [1:0] stage7_53;
   wire [1:0] stage7_54;
   wire [1:0] stage7_55;
   wire [1:0] stage7_56;
   wire [1:0] stage7_57;
   wire [1:0] stage7_58;
   wire [1:0] stage7_59;
   wire [1:0] stage7_60;
   wire [0:0] stage7_61;
   wire [1:0] stage7_62;
   wire [1:0] stage7_63;
   wire [1:0] stage7_64;
   wire [1:0] stage7_65;
   wire [1:0] stage7_66;
   wire [1:0] stage7_67;
   wire [1:0] stage7_68;
   wire [1:0] stage7_69;
   wire [0:0] stage7_70;
   wire [0:0] stage7_71;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;
   assign dst25 = stage7_25;
   assign dst26 = stage7_26;
   assign dst27 = stage7_27;
   assign dst28 = stage7_28;
   assign dst29 = stage7_29;
   assign dst30 = stage7_30;
   assign dst31 = stage7_31;
   assign dst32 = stage7_32;
   assign dst33 = stage7_33;
   assign dst34 = stage7_34;
   assign dst35 = stage7_35;
   assign dst36 = stage7_36;
   assign dst37 = stage7_37;
   assign dst38 = stage7_38;
   assign dst39 = stage7_39;
   assign dst40 = stage7_40;
   assign dst41 = stage7_41;
   assign dst42 = stage7_42;
   assign dst43 = stage7_43;
   assign dst44 = stage7_44;
   assign dst45 = stage7_45;
   assign dst46 = stage7_46;
   assign dst47 = stage7_47;
   assign dst48 = stage7_48;
   assign dst49 = stage7_49;
   assign dst50 = stage7_50;
   assign dst51 = stage7_51;
   assign dst52 = stage7_52;
   assign dst53 = stage7_53;
   assign dst54 = stage7_54;
   assign dst55 = stage7_55;
   assign dst56 = stage7_56;
   assign dst57 = stage7_57;
   assign dst58 = stage7_58;
   assign dst59 = stage7_59;
   assign dst60 = stage7_60;
   assign dst61 = stage7_61;
   assign dst62 = stage7_62;
   assign dst63 = stage7_63;
   assign dst64 = stage7_64;
   assign dst65 = stage7_65;
   assign dst66 = stage7_66;
   assign dst67 = stage7_67;
   assign dst68 = stage7_68;
   assign dst69 = stage7_69;
   assign dst70 = stage7_70;
   assign dst71 = stage7_71;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7]},
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[1]},
      {stage0_3[2]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[2]},
      {stage0_3[3]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[3]},
      {stage0_3[4]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[4]},
      {stage0_3[5]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[5]},
      {stage0_3[6]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[20], stage0_0[21], stage0_0[22]},
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_2[6]},
      {stage0_3[7]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_2[7]},
      {stage0_3[8]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_2[8]},
      {stage0_3[9]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[29], stage0_0[30], stage0_0[31]},
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_2[9]},
      {stage0_3[10]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_2[10]},
      {stage0_3[11]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_2[11]},
      {stage0_3[12]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[38], stage0_0[39], stage0_0[40]},
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_2[12]},
      {stage0_3[13]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_2[13]},
      {stage0_3[14]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc207_4 gpc14 (
      {stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[14], stage0_2[15]},
      {stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21]},
      {stage1_4[14],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27]},
      {stage1_4[15],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33]},
      {stage1_4[16],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39]},
      {stage1_4[17],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45]},
      {stage1_4[18],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51]},
      {stage1_4[19],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57]},
      {stage1_4[20],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage1_4[21],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69]},
      {stage1_4[22],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75]},
      {stage1_4[23],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage1_4[24],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122]},
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87]},
      {stage1_4[25],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128]},
      {stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93]},
      {stage1_4[26],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134]},
      {stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99]},
      {stage1_4[27],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140]},
      {stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105]},
      {stage1_4[28],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage1_4[29],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc615_5 gpc31 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151]},
      {stage0_1[81]},
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117]},
      {stage1_4[30],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc615_5 gpc32 (
      {stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[82]},
      {stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123]},
      {stage1_4[31],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc615_5 gpc33 (
      {stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161]},
      {stage0_1[83]},
      {stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129]},
      {stage1_4[32],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[0],stage1_4[33],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[1],stage1_4[34],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[2],stage1_4[35],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[3],stage1_4[36],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[4],stage1_4[37],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[5],stage1_4[38],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[6],stage1_4[39],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[7],stage1_4[40],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[8],stage1_4[41],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[9],stage1_4[42],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[10],stage1_4[43],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[11],stage1_4[44],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[12],stage1_4[45],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc615_5 gpc47 (
      {stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage0_3[93]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[13],stage1_4[46],stage1_3[47],stage1_2[47]}
   );
   gpc615_5 gpc48 (
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139]},
      {stage0_3[94]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[14],stage1_4[47],stage1_3[48],stage1_2[48]}
   );
   gpc615_5 gpc49 (
      {stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage0_3[95]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[15],stage1_4[48],stage1_3[49],stage1_2[49]}
   );
   gpc615_5 gpc50 (
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage0_3[96]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[16],stage1_4[49],stage1_3[50],stage1_2[50]}
   );
   gpc615_5 gpc51 (
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154]},
      {stage0_3[97]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[17],stage1_4[50],stage1_3[51],stage1_2[51]}
   );
   gpc615_5 gpc52 (
      {stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159]},
      {stage0_3[98]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[18],stage1_4[51],stage1_3[52],stage1_2[52]}
   );
   gpc615_5 gpc53 (
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage0_4[36]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[6],stage1_5[19],stage1_4[52],stage1_3[53]}
   );
   gpc615_5 gpc54 (
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108]},
      {stage0_4[37]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[7],stage1_5[20],stage1_4[53],stage1_3[54]}
   );
   gpc615_5 gpc55 (
      {stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113]},
      {stage0_4[38]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[8],stage1_5[21],stage1_4[54],stage1_3[55]}
   );
   gpc615_5 gpc56 (
      {stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118]},
      {stage0_4[39]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[9],stage1_5[22],stage1_4[55],stage1_3[56]}
   );
   gpc615_5 gpc57 (
      {stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage0_4[40]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[10],stage1_5[23],stage1_4[56],stage1_3[57]}
   );
   gpc615_5 gpc58 (
      {stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage0_4[41]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[11],stage1_5[24],stage1_4[57],stage1_3[58]}
   );
   gpc615_5 gpc59 (
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage0_4[42]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[12],stage1_5[25],stage1_4[58],stage1_3[59]}
   );
   gpc615_5 gpc60 (
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138]},
      {stage0_4[43]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[13],stage1_5[26],stage1_4[59],stage1_3[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[8],stage1_6[14],stage1_5[27],stage1_4[60]}
   );
   gpc606_5 gpc62 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[9],stage1_6[15],stage1_5[28],stage1_4[61]}
   );
   gpc606_5 gpc63 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[10],stage1_6[16],stage1_5[29],stage1_4[62]}
   );
   gpc606_5 gpc64 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[11],stage1_6[17],stage1_5[30],stage1_4[63]}
   );
   gpc606_5 gpc65 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[12],stage1_6[18],stage1_5[31],stage1_4[64]}
   );
   gpc606_5 gpc66 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[13],stage1_6[19],stage1_5[32],stage1_4[65]}
   );
   gpc606_5 gpc67 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[14],stage1_6[20],stage1_5[33],stage1_4[66]}
   );
   gpc606_5 gpc68 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[15],stage1_6[21],stage1_5[34],stage1_4[67]}
   );
   gpc606_5 gpc69 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[16],stage1_6[22],stage1_5[35],stage1_4[68]}
   );
   gpc606_5 gpc70 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[17],stage1_6[23],stage1_5[36],stage1_4[69]}
   );
   gpc606_5 gpc71 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[18],stage1_6[24],stage1_5[37],stage1_4[70]}
   );
   gpc606_5 gpc72 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[19],stage1_6[25],stage1_5[38],stage1_4[71]}
   );
   gpc606_5 gpc73 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[20],stage1_6[26],stage1_5[39],stage1_4[72]}
   );
   gpc606_5 gpc74 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[21],stage1_6[27],stage1_5[40],stage1_4[73]}
   );
   gpc606_5 gpc75 (
      {stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[22],stage1_6[28],stage1_5[41],stage1_4[74]}
   );
   gpc606_5 gpc76 (
      {stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[23],stage1_6[29],stage1_5[42],stage1_4[75]}
   );
   gpc606_5 gpc77 (
      {stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[24],stage1_6[30],stage1_5[43],stage1_4[76]}
   );
   gpc606_5 gpc78 (
      {stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[25],stage1_6[31],stage1_5[44],stage1_4[77]}
   );
   gpc606_5 gpc79 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[26],stage1_6[32],stage1_5[45],stage1_4[78]}
   );
   gpc606_5 gpc80 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[19],stage1_7[27],stage1_6[33],stage1_5[46]}
   );
   gpc606_5 gpc81 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[20],stage1_7[28],stage1_6[34],stage1_5[47]}
   );
   gpc606_5 gpc82 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[21],stage1_7[29],stage1_6[35],stage1_5[48]}
   );
   gpc606_5 gpc83 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[22],stage1_7[30],stage1_6[36],stage1_5[49]}
   );
   gpc606_5 gpc84 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[23],stage1_7[31],stage1_6[37],stage1_5[50]}
   );
   gpc606_5 gpc85 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[24],stage1_7[32],stage1_6[38],stage1_5[51]}
   );
   gpc606_5 gpc86 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[25],stage1_7[33],stage1_6[39],stage1_5[52]}
   );
   gpc606_5 gpc87 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[26],stage1_7[34],stage1_6[40],stage1_5[53]}
   );
   gpc606_5 gpc88 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[27],stage1_7[35],stage1_6[41],stage1_5[54]}
   );
   gpc615_5 gpc89 (
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118]},
      {stage0_7[54]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[28],stage1_7[36],stage1_6[42]}
   );
   gpc615_5 gpc90 (
      {stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123]},
      {stage0_7[55]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[29],stage1_7[37],stage1_6[43]}
   );
   gpc615_5 gpc91 (
      {stage0_6[124], stage0_6[125], stage0_6[126], stage0_6[127], stage0_6[128]},
      {stage0_7[56]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[11],stage1_8[30],stage1_7[38],stage1_6[44]}
   );
   gpc615_5 gpc92 (
      {stage0_6[129], stage0_6[130], stage0_6[131], stage0_6[132], stage0_6[133]},
      {stage0_7[57]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[12],stage1_8[31],stage1_7[39],stage1_6[45]}
   );
   gpc615_5 gpc93 (
      {stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137], stage0_6[138]},
      {stage0_7[58]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[13],stage1_8[32],stage1_7[40],stage1_6[46]}
   );
   gpc615_5 gpc94 (
      {stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage0_7[59]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[14],stage1_8[33],stage1_7[41],stage1_6[47]}
   );
   gpc615_5 gpc95 (
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148]},
      {stage0_7[60]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[15],stage1_8[34],stage1_7[42],stage1_6[48]}
   );
   gpc615_5 gpc96 (
      {stage0_6[149], stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153]},
      {stage0_7[61]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[16],stage1_8[35],stage1_7[43],stage1_6[49]}
   );
   gpc606_5 gpc97 (
      {stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65], stage0_7[66], stage0_7[67]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[8],stage1_9[17],stage1_8[36],stage1_7[44]}
   );
   gpc615_5 gpc98 (
      {stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71], stage0_7[72]},
      {stage0_8[48]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[9],stage1_9[18],stage1_8[37],stage1_7[45]}
   );
   gpc615_5 gpc99 (
      {stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage0_8[49]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[10],stage1_9[19],stage1_8[38],stage1_7[46]}
   );
   gpc615_5 gpc100 (
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82]},
      {stage0_8[50]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[11],stage1_9[20],stage1_8[39],stage1_7[47]}
   );
   gpc615_5 gpc101 (
      {stage0_7[83], stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87]},
      {stage0_8[51]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[12],stage1_9[21],stage1_8[40],stage1_7[48]}
   );
   gpc615_5 gpc102 (
      {stage0_7[88], stage0_7[89], stage0_7[90], stage0_7[91], stage0_7[92]},
      {stage0_8[52]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[13],stage1_9[22],stage1_8[41],stage1_7[49]}
   );
   gpc615_5 gpc103 (
      {stage0_7[93], stage0_7[94], stage0_7[95], stage0_7[96], stage0_7[97]},
      {stage0_8[53]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[14],stage1_9[23],stage1_8[42],stage1_7[50]}
   );
   gpc615_5 gpc104 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[54]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[15],stage1_9[24],stage1_8[43],stage1_7[51]}
   );
   gpc615_5 gpc105 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[55]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[16],stage1_9[25],stage1_8[44],stage1_7[52]}
   );
   gpc615_5 gpc106 (
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112]},
      {stage0_8[56]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[17],stage1_9[26],stage1_8[45],stage1_7[53]}
   );
   gpc615_5 gpc107 (
      {stage0_7[113], stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117]},
      {stage0_8[57]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[18],stage1_9[27],stage1_8[46],stage1_7[54]}
   );
   gpc615_5 gpc108 (
      {stage0_7[118], stage0_7[119], stage0_7[120], stage0_7[121], stage0_7[122]},
      {stage0_8[58]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[19],stage1_9[28],stage1_8[47],stage1_7[55]}
   );
   gpc615_5 gpc109 (
      {stage0_7[123], stage0_7[124], stage0_7[125], stage0_7[126], stage0_7[127]},
      {stage0_8[59]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[20],stage1_9[29],stage1_8[48],stage1_7[56]}
   );
   gpc615_5 gpc110 (
      {stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131], stage0_7[132]},
      {stage0_8[60]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[21],stage1_9[30],stage1_8[49],stage1_7[57]}
   );
   gpc615_5 gpc111 (
      {stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage0_8[61]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[22],stage1_9[31],stage1_8[50],stage1_7[58]}
   );
   gpc615_5 gpc112 (
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142]},
      {stage0_8[62]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[23],stage1_9[32],stage1_8[51],stage1_7[59]}
   );
   gpc615_5 gpc113 (
      {stage0_7[143], stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147]},
      {stage0_8[63]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[24],stage1_9[33],stage1_8[52],stage1_7[60]}
   );
   gpc615_5 gpc114 (
      {stage0_7[148], stage0_7[149], stage0_7[150], stage0_7[151], stage0_7[152]},
      {stage0_8[64]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[25],stage1_9[34],stage1_8[53],stage1_7[61]}
   );
   gpc606_5 gpc115 (
      {stage0_8[65], stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[18],stage1_10[26],stage1_9[35],stage1_8[54]}
   );
   gpc606_5 gpc116 (
      {stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[19],stage1_10[27],stage1_9[36],stage1_8[55]}
   );
   gpc606_5 gpc117 (
      {stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[20],stage1_10[28],stage1_9[37],stage1_8[56]}
   );
   gpc606_5 gpc118 (
      {stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[21],stage1_10[29],stage1_9[38],stage1_8[57]}
   );
   gpc606_5 gpc119 (
      {stage0_8[89], stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[22],stage1_10[30],stage1_9[39],stage1_8[58]}
   );
   gpc606_5 gpc120 (
      {stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[23],stage1_10[31],stage1_9[40],stage1_8[59]}
   );
   gpc606_5 gpc121 (
      {stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[24],stage1_10[32],stage1_9[41],stage1_8[60]}
   );
   gpc606_5 gpc122 (
      {stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[25],stage1_10[33],stage1_9[42],stage1_8[61]}
   );
   gpc606_5 gpc123 (
      {stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[26],stage1_10[34],stage1_9[43],stage1_8[62]}
   );
   gpc606_5 gpc124 (
      {stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[27],stage1_10[35],stage1_9[44],stage1_8[63]}
   );
   gpc606_5 gpc125 (
      {stage0_8[125], stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[28],stage1_10[36],stage1_9[45],stage1_8[64]}
   );
   gpc606_5 gpc126 (
      {stage0_8[131], stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[29],stage1_10[37],stage1_9[46],stage1_8[65]}
   );
   gpc606_5 gpc127 (
      {stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[30],stage1_10[38],stage1_9[47],stage1_8[66]}
   );
   gpc606_5 gpc128 (
      {stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[31],stage1_10[39],stage1_9[48],stage1_8[67]}
   );
   gpc606_5 gpc129 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[14],stage1_11[32],stage1_10[40],stage1_9[49]}
   );
   gpc606_5 gpc130 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[15],stage1_11[33],stage1_10[41],stage1_9[50]}
   );
   gpc606_5 gpc131 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[16],stage1_11[34],stage1_10[42],stage1_9[51]}
   );
   gpc606_5 gpc132 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[17],stage1_11[35],stage1_10[43],stage1_9[52]}
   );
   gpc606_5 gpc133 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[18],stage1_11[36],stage1_10[44],stage1_9[53]}
   );
   gpc606_5 gpc134 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[19],stage1_11[37],stage1_10[45],stage1_9[54]}
   );
   gpc606_5 gpc135 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[20],stage1_11[38],stage1_10[46],stage1_9[55]}
   );
   gpc606_5 gpc136 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[21],stage1_11[39],stage1_10[47],stage1_9[56]}
   );
   gpc606_5 gpc137 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[22],stage1_11[40],stage1_10[48],stage1_9[57]}
   );
   gpc615_5 gpc138 (
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88]},
      {stage0_11[54]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[9],stage1_12[23],stage1_11[41],stage1_10[49]}
   );
   gpc615_5 gpc139 (
      {stage0_10[89], stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93]},
      {stage0_11[55]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[10],stage1_12[24],stage1_11[42],stage1_10[50]}
   );
   gpc615_5 gpc140 (
      {stage0_10[94], stage0_10[95], stage0_10[96], stage0_10[97], stage0_10[98]},
      {stage0_11[56]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[11],stage1_12[25],stage1_11[43],stage1_10[51]}
   );
   gpc615_5 gpc141 (
      {stage0_10[99], stage0_10[100], stage0_10[101], stage0_10[102], stage0_10[103]},
      {stage0_11[57]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[12],stage1_12[26],stage1_11[44],stage1_10[52]}
   );
   gpc615_5 gpc142 (
      {stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107], stage0_10[108]},
      {stage0_11[58]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[13],stage1_12[27],stage1_11[45],stage1_10[53]}
   );
   gpc615_5 gpc143 (
      {stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage0_11[59]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[14],stage1_12[28],stage1_11[46],stage1_10[54]}
   );
   gpc615_5 gpc144 (
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118]},
      {stage0_11[60]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[15],stage1_12[29],stage1_11[47],stage1_10[55]}
   );
   gpc615_5 gpc145 (
      {stage0_10[119], stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123]},
      {stage0_11[61]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[16],stage1_12[30],stage1_11[48],stage1_10[56]}
   );
   gpc606_5 gpc146 (
      {stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65], stage0_11[66], stage0_11[67]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[8],stage1_13[17],stage1_12[31],stage1_11[49]}
   );
   gpc606_5 gpc147 (
      {stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71], stage0_11[72], stage0_11[73]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[9],stage1_13[18],stage1_12[32],stage1_11[50]}
   );
   gpc606_5 gpc148 (
      {stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77], stage0_11[78], stage0_11[79]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[10],stage1_13[19],stage1_12[33],stage1_11[51]}
   );
   gpc606_5 gpc149 (
      {stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83], stage0_11[84], stage0_11[85]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[11],stage1_13[20],stage1_12[34],stage1_11[52]}
   );
   gpc606_5 gpc150 (
      {stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89], stage0_11[90], stage0_11[91]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[12],stage1_13[21],stage1_12[35],stage1_11[53]}
   );
   gpc606_5 gpc151 (
      {stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95], stage0_11[96], stage0_11[97]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[13],stage1_13[22],stage1_12[36],stage1_11[54]}
   );
   gpc606_5 gpc152 (
      {stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101], stage0_11[102], stage0_11[103]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[14],stage1_13[23],stage1_12[37],stage1_11[55]}
   );
   gpc606_5 gpc153 (
      {stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107], stage0_11[108], stage0_11[109]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[15],stage1_13[24],stage1_12[38],stage1_11[56]}
   );
   gpc606_5 gpc154 (
      {stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113], stage0_11[114], stage0_11[115]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[16],stage1_13[25],stage1_12[39],stage1_11[57]}
   );
   gpc606_5 gpc155 (
      {stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119], stage0_11[120], stage0_11[121]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[17],stage1_13[26],stage1_12[40],stage1_11[58]}
   );
   gpc606_5 gpc156 (
      {stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125], stage0_11[126], stage0_11[127]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[18],stage1_13[27],stage1_12[41],stage1_11[59]}
   );
   gpc606_5 gpc157 (
      {stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[19],stage1_13[28],stage1_12[42],stage1_11[60]}
   );
   gpc615_5 gpc158 (
      {stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137], stage0_11[138]},
      {stage0_12[48]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[20],stage1_13[29],stage1_12[43],stage1_11[61]}
   );
   gpc615_5 gpc159 (
      {stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage0_12[49]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[21],stage1_13[30],stage1_12[44],stage1_11[62]}
   );
   gpc606_5 gpc160 (
      {stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[14],stage1_14[22],stage1_13[31],stage1_12[45]}
   );
   gpc606_5 gpc161 (
      {stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[15],stage1_14[23],stage1_13[32],stage1_12[46]}
   );
   gpc606_5 gpc162 (
      {stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[16],stage1_14[24],stage1_13[33],stage1_12[47]}
   );
   gpc606_5 gpc163 (
      {stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[17],stage1_14[25],stage1_13[34],stage1_12[48]}
   );
   gpc606_5 gpc164 (
      {stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[18],stage1_14[26],stage1_13[35],stage1_12[49]}
   );
   gpc606_5 gpc165 (
      {stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[19],stage1_14[27],stage1_13[36],stage1_12[50]}
   );
   gpc606_5 gpc166 (
      {stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[20],stage1_14[28],stage1_13[37],stage1_12[51]}
   );
   gpc606_5 gpc167 (
      {stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[21],stage1_14[29],stage1_13[38],stage1_12[52]}
   );
   gpc606_5 gpc168 (
      {stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[22],stage1_14[30],stage1_13[39],stage1_12[53]}
   );
   gpc606_5 gpc169 (
      {stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[23],stage1_14[31],stage1_13[40],stage1_12[54]}
   );
   gpc606_5 gpc170 (
      {stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[24],stage1_14[32],stage1_13[41],stage1_12[55]}
   );
   gpc606_5 gpc171 (
      {stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[25],stage1_14[33],stage1_13[42],stage1_12[56]}
   );
   gpc606_5 gpc172 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[26],stage1_14[34],stage1_13[43],stage1_12[57]}
   );
   gpc606_5 gpc173 (
      {stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[27],stage1_14[35],stage1_13[44],stage1_12[58]}
   );
   gpc606_5 gpc174 (
      {stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[28],stage1_14[36],stage1_13[45],stage1_12[59]}
   );
   gpc606_5 gpc175 (
      {stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[29],stage1_14[37],stage1_13[46],stage1_12[60]}
   );
   gpc606_5 gpc176 (
      {stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[30],stage1_14[38],stage1_13[47],stage1_12[61]}
   );
   gpc606_5 gpc177 (
      {stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[31],stage1_14[39],stage1_13[48],stage1_12[62]}
   );
   gpc606_5 gpc178 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[18],stage1_15[32],stage1_14[40],stage1_13[49]}
   );
   gpc606_5 gpc179 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[19],stage1_15[33],stage1_14[41],stage1_13[50]}
   );
   gpc606_5 gpc180 (
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[20],stage1_15[34],stage1_14[42],stage1_13[51]}
   );
   gpc606_5 gpc181 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[21],stage1_15[35],stage1_14[43],stage1_13[52]}
   );
   gpc606_5 gpc182 (
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[22],stage1_15[36],stage1_14[44],stage1_13[53]}
   );
   gpc606_5 gpc183 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[23],stage1_15[37],stage1_14[45],stage1_13[54]}
   );
   gpc606_5 gpc184 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[24],stage1_15[38],stage1_14[46],stage1_13[55]}
   );
   gpc606_5 gpc185 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[25],stage1_15[39],stage1_14[47],stage1_13[56]}
   );
   gpc615_5 gpc186 (
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112]},
      {stage0_15[48]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[8],stage1_16[26],stage1_15[40],stage1_14[48]}
   );
   gpc615_5 gpc187 (
      {stage0_14[113], stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117]},
      {stage0_15[49]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[9],stage1_16[27],stage1_15[41],stage1_14[49]}
   );
   gpc615_5 gpc188 (
      {stage0_14[118], stage0_14[119], stage0_14[120], stage0_14[121], stage0_14[122]},
      {stage0_15[50]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[10],stage1_16[28],stage1_15[42],stage1_14[50]}
   );
   gpc615_5 gpc189 (
      {stage0_14[123], stage0_14[124], stage0_14[125], stage0_14[126], stage0_14[127]},
      {stage0_15[51]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[11],stage1_16[29],stage1_15[43],stage1_14[51]}
   );
   gpc615_5 gpc190 (
      {stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_15[52]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[12],stage1_16[30],stage1_15[44],stage1_14[52]}
   );
   gpc615_5 gpc191 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage0_15[53]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[13],stage1_16[31],stage1_15[45],stage1_14[53]}
   );
   gpc615_5 gpc192 (
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142]},
      {stage0_15[54]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[14],stage1_16[32],stage1_15[46],stage1_14[54]}
   );
   gpc615_5 gpc193 (
      {stage0_14[143], stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147]},
      {stage0_15[55]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[15],stage1_16[33],stage1_15[47],stage1_14[55]}
   );
   gpc615_5 gpc194 (
      {stage0_14[148], stage0_14[149], stage0_14[150], stage0_14[151], stage0_14[152]},
      {stage0_15[56]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[16],stage1_16[34],stage1_15[48],stage1_14[56]}
   );
   gpc615_5 gpc195 (
      {stage0_14[153], stage0_14[154], stage0_14[155], stage0_14[156], stage0_14[157]},
      {stage0_15[57]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[17],stage1_16[35],stage1_15[49],stage1_14[57]}
   );
   gpc615_5 gpc196 (
      {stage0_15[58], stage0_15[59], stage0_15[60], stage0_15[61], stage0_15[62]},
      {stage0_16[60]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[10],stage1_17[18],stage1_16[36],stage1_15[50]}
   );
   gpc615_5 gpc197 (
      {stage0_15[63], stage0_15[64], stage0_15[65], stage0_15[66], stage0_15[67]},
      {stage0_16[61]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[11],stage1_17[19],stage1_16[37],stage1_15[51]}
   );
   gpc615_5 gpc198 (
      {stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71], stage0_15[72]},
      {stage0_16[62]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[12],stage1_17[20],stage1_16[38],stage1_15[52]}
   );
   gpc615_5 gpc199 (
      {stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage0_16[63]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[13],stage1_17[21],stage1_16[39],stage1_15[53]}
   );
   gpc615_5 gpc200 (
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82]},
      {stage0_16[64]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[14],stage1_17[22],stage1_16[40],stage1_15[54]}
   );
   gpc615_5 gpc201 (
      {stage0_15[83], stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87]},
      {stage0_16[65]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[15],stage1_17[23],stage1_16[41],stage1_15[55]}
   );
   gpc615_5 gpc202 (
      {stage0_15[88], stage0_15[89], stage0_15[90], stage0_15[91], stage0_15[92]},
      {stage0_16[66]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[16],stage1_17[24],stage1_16[42],stage1_15[56]}
   );
   gpc615_5 gpc203 (
      {stage0_15[93], stage0_15[94], stage0_15[95], stage0_15[96], stage0_15[97]},
      {stage0_16[67]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[17],stage1_17[25],stage1_16[43],stage1_15[57]}
   );
   gpc615_5 gpc204 (
      {stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101], stage0_15[102]},
      {stage0_16[68]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[18],stage1_17[26],stage1_16[44],stage1_15[58]}
   );
   gpc615_5 gpc205 (
      {stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage0_16[69]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[19],stage1_17[27],stage1_16[45],stage1_15[59]}
   );
   gpc615_5 gpc206 (
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112]},
      {stage0_16[70]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[20],stage1_17[28],stage1_16[46],stage1_15[60]}
   );
   gpc615_5 gpc207 (
      {stage0_15[113], stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117]},
      {stage0_16[71]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[21],stage1_17[29],stage1_16[47],stage1_15[61]}
   );
   gpc615_5 gpc208 (
      {stage0_15[118], stage0_15[119], stage0_15[120], stage0_15[121], stage0_15[122]},
      {stage0_16[72]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[22],stage1_17[30],stage1_16[48],stage1_15[62]}
   );
   gpc615_5 gpc209 (
      {stage0_15[123], stage0_15[124], stage0_15[125], stage0_15[126], stage0_15[127]},
      {stage0_16[73]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[23],stage1_17[31],stage1_16[49],stage1_15[63]}
   );
   gpc606_5 gpc210 (
      {stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78], stage0_16[79]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[14],stage1_18[24],stage1_17[32],stage1_16[50]}
   );
   gpc606_5 gpc211 (
      {stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84], stage0_16[85]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[15],stage1_18[25],stage1_17[33],stage1_16[51]}
   );
   gpc606_5 gpc212 (
      {stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[16],stage1_18[26],stage1_17[34],stage1_16[52]}
   );
   gpc606_5 gpc213 (
      {stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[17],stage1_18[27],stage1_17[35],stage1_16[53]}
   );
   gpc606_5 gpc214 (
      {stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[18],stage1_18[28],stage1_17[36],stage1_16[54]}
   );
   gpc606_5 gpc215 (
      {stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[19],stage1_18[29],stage1_17[37],stage1_16[55]}
   );
   gpc606_5 gpc216 (
      {stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114], stage0_16[115]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[20],stage1_18[30],stage1_17[38],stage1_16[56]}
   );
   gpc606_5 gpc217 (
      {stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120], stage0_16[121]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[21],stage1_18[31],stage1_17[39],stage1_16[57]}
   );
   gpc606_5 gpc218 (
      {stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[22],stage1_18[32],stage1_17[40],stage1_16[58]}
   );
   gpc606_5 gpc219 (
      {stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[23],stage1_18[33],stage1_17[41],stage1_16[59]}
   );
   gpc606_5 gpc220 (
      {stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[24],stage1_18[34],stage1_17[42],stage1_16[60]}
   );
   gpc606_5 gpc221 (
      {stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[25],stage1_18[35],stage1_17[43],stage1_16[61]}
   );
   gpc606_5 gpc222 (
      {stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[26],stage1_18[36],stage1_17[44],stage1_16[62]}
   );
   gpc606_5 gpc223 (
      {stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[27],stage1_18[37],stage1_17[45],stage1_16[63]}
   );
   gpc606_5 gpc224 (
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[14],stage1_19[28],stage1_18[38],stage1_17[46]}
   );
   gpc606_5 gpc225 (
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[15],stage1_19[29],stage1_18[39],stage1_17[47]}
   );
   gpc606_5 gpc226 (
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[2],stage1_20[16],stage1_19[30],stage1_18[40]}
   );
   gpc606_5 gpc227 (
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[3],stage1_20[17],stage1_19[31],stage1_18[41]}
   );
   gpc606_5 gpc228 (
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[4],stage1_20[18],stage1_19[32],stage1_18[42]}
   );
   gpc606_5 gpc229 (
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[5],stage1_20[19],stage1_19[33],stage1_18[43]}
   );
   gpc606_5 gpc230 (
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[6],stage1_20[20],stage1_19[34],stage1_18[44]}
   );
   gpc606_5 gpc231 (
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[7],stage1_20[21],stage1_19[35],stage1_18[45]}
   );
   gpc606_5 gpc232 (
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[8],stage1_20[22],stage1_19[36],stage1_18[46]}
   );
   gpc615_5 gpc233 (
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130]},
      {stage0_19[12]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[9],stage1_20[23],stage1_19[37],stage1_18[47]}
   );
   gpc615_5 gpc234 (
      {stage0_18[131], stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135]},
      {stage0_19[13]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[10],stage1_20[24],stage1_19[38],stage1_18[48]}
   );
   gpc615_5 gpc235 (
      {stage0_18[136], stage0_18[137], stage0_18[138], stage0_18[139], stage0_18[140]},
      {stage0_19[14]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[11],stage1_20[25],stage1_19[39],stage1_18[49]}
   );
   gpc615_5 gpc236 (
      {stage0_18[141], stage0_18[142], stage0_18[143], stage0_18[144], stage0_18[145]},
      {stage0_19[15]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[12],stage1_20[26],stage1_19[40],stage1_18[50]}
   );
   gpc615_5 gpc237 (
      {stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149], stage0_18[150]},
      {stage0_19[16]},
      {stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71]},
      {stage1_22[11],stage1_21[13],stage1_20[27],stage1_19[41],stage1_18[51]}
   );
   gpc207_4 gpc238 (
      {stage0_19[17], stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage0_21[0], stage0_21[1]},
      {stage1_22[12],stage1_21[14],stage1_20[28],stage1_19[42]}
   );
   gpc207_4 gpc239 (
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29], stage0_19[30]},
      {stage0_21[2], stage0_21[3]},
      {stage1_22[13],stage1_21[15],stage1_20[29],stage1_19[43]}
   );
   gpc207_4 gpc240 (
      {stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35], stage0_19[36], stage0_19[37]},
      {stage0_21[4], stage0_21[5]},
      {stage1_22[14],stage1_21[16],stage1_20[30],stage1_19[44]}
   );
   gpc207_4 gpc241 (
      {stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41], stage0_19[42], stage0_19[43], stage0_19[44]},
      {stage0_21[6], stage0_21[7]},
      {stage1_22[15],stage1_21[17],stage1_20[31],stage1_19[45]}
   );
   gpc606_5 gpc242 (
      {stage0_19[45], stage0_19[46], stage0_19[47], stage0_19[48], stage0_19[49], stage0_19[50]},
      {stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13]},
      {stage1_23[0],stage1_22[16],stage1_21[18],stage1_20[32],stage1_19[46]}
   );
   gpc606_5 gpc243 (
      {stage0_19[51], stage0_19[52], stage0_19[53], stage0_19[54], stage0_19[55], stage0_19[56]},
      {stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19]},
      {stage1_23[1],stage1_22[17],stage1_21[19],stage1_20[33],stage1_19[47]}
   );
   gpc606_5 gpc244 (
      {stage0_19[57], stage0_19[58], stage0_19[59], stage0_19[60], stage0_19[61], stage0_19[62]},
      {stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25]},
      {stage1_23[2],stage1_22[18],stage1_21[20],stage1_20[34],stage1_19[48]}
   );
   gpc606_5 gpc245 (
      {stage0_19[63], stage0_19[64], stage0_19[65], stage0_19[66], stage0_19[67], stage0_19[68]},
      {stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31]},
      {stage1_23[3],stage1_22[19],stage1_21[21],stage1_20[35],stage1_19[49]}
   );
   gpc606_5 gpc246 (
      {stage0_19[69], stage0_19[70], stage0_19[71], stage0_19[72], stage0_19[73], stage0_19[74]},
      {stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36], stage0_21[37]},
      {stage1_23[4],stage1_22[20],stage1_21[22],stage1_20[36],stage1_19[50]}
   );
   gpc606_5 gpc247 (
      {stage0_19[75], stage0_19[76], stage0_19[77], stage0_19[78], stage0_19[79], stage0_19[80]},
      {stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43]},
      {stage1_23[5],stage1_22[21],stage1_21[23],stage1_20[37],stage1_19[51]}
   );
   gpc606_5 gpc248 (
      {stage0_19[81], stage0_19[82], stage0_19[83], stage0_19[84], stage0_19[85], stage0_19[86]},
      {stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48], stage0_21[49]},
      {stage1_23[6],stage1_22[22],stage1_21[24],stage1_20[38],stage1_19[52]}
   );
   gpc606_5 gpc249 (
      {stage0_19[87], stage0_19[88], stage0_19[89], stage0_19[90], stage0_19[91], stage0_19[92]},
      {stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53], stage0_21[54], stage0_21[55]},
      {stage1_23[7],stage1_22[23],stage1_21[25],stage1_20[39],stage1_19[53]}
   );
   gpc606_5 gpc250 (
      {stage0_19[93], stage0_19[94], stage0_19[95], stage0_19[96], stage0_19[97], stage0_19[98]},
      {stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59], stage0_21[60], stage0_21[61]},
      {stage1_23[8],stage1_22[24],stage1_21[26],stage1_20[40],stage1_19[54]}
   );
   gpc606_5 gpc251 (
      {stage0_19[99], stage0_19[100], stage0_19[101], stage0_19[102], stage0_19[103], stage0_19[104]},
      {stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65], stage0_21[66], stage0_21[67]},
      {stage1_23[9],stage1_22[25],stage1_21[27],stage1_20[41],stage1_19[55]}
   );
   gpc606_5 gpc252 (
      {stage0_19[105], stage0_19[106], stage0_19[107], stage0_19[108], stage0_19[109], stage0_19[110]},
      {stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71], stage0_21[72], stage0_21[73]},
      {stage1_23[10],stage1_22[26],stage1_21[28],stage1_20[42],stage1_19[56]}
   );
   gpc606_5 gpc253 (
      {stage0_19[111], stage0_19[112], stage0_19[113], stage0_19[114], stage0_19[115], stage0_19[116]},
      {stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77], stage0_21[78], stage0_21[79]},
      {stage1_23[11],stage1_22[27],stage1_21[29],stage1_20[43],stage1_19[57]}
   );
   gpc606_5 gpc254 (
      {stage0_19[117], stage0_19[118], stage0_19[119], stage0_19[120], stage0_19[121], stage0_19[122]},
      {stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83], stage0_21[84], stage0_21[85]},
      {stage1_23[12],stage1_22[28],stage1_21[30],stage1_20[44],stage1_19[58]}
   );
   gpc606_5 gpc255 (
      {stage0_19[123], stage0_19[124], stage0_19[125], stage0_19[126], stage0_19[127], stage0_19[128]},
      {stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89], stage0_21[90], stage0_21[91]},
      {stage1_23[13],stage1_22[29],stage1_21[31],stage1_20[45],stage1_19[59]}
   );
   gpc606_5 gpc256 (
      {stage0_19[129], stage0_19[130], stage0_19[131], stage0_19[132], stage0_19[133], stage0_19[134]},
      {stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95], stage0_21[96], stage0_21[97]},
      {stage1_23[14],stage1_22[30],stage1_21[32],stage1_20[46],stage1_19[60]}
   );
   gpc606_5 gpc257 (
      {stage0_19[135], stage0_19[136], stage0_19[137], stage0_19[138], stage0_19[139], stage0_19[140]},
      {stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101], stage0_21[102], stage0_21[103]},
      {stage1_23[15],stage1_22[31],stage1_21[33],stage1_20[47],stage1_19[61]}
   );
   gpc615_5 gpc258 (
      {stage0_19[141], stage0_19[142], stage0_19[143], stage0_19[144], stage0_19[145]},
      {stage0_20[72]},
      {stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107], stage0_21[108], stage0_21[109]},
      {stage1_23[16],stage1_22[32],stage1_21[34],stage1_20[48],stage1_19[62]}
   );
   gpc615_5 gpc259 (
      {stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149], stage0_19[150]},
      {stage0_20[73]},
      {stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115]},
      {stage1_23[17],stage1_22[33],stage1_21[35],stage1_20[49],stage1_19[63]}
   );
   gpc615_5 gpc260 (
      {stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage0_20[74]},
      {stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119], stage0_21[120], stage0_21[121]},
      {stage1_23[18],stage1_22[34],stage1_21[36],stage1_20[50],stage1_19[64]}
   );
   gpc606_5 gpc261 (
      {stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[19],stage1_22[35],stage1_21[37],stage1_20[51]}
   );
   gpc606_5 gpc262 (
      {stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[20],stage1_22[36],stage1_21[38],stage1_20[52]}
   );
   gpc606_5 gpc263 (
      {stage0_20[87], stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[21],stage1_22[37],stage1_21[39],stage1_20[53]}
   );
   gpc606_5 gpc264 (
      {stage0_20[93], stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[22],stage1_22[38],stage1_21[40],stage1_20[54]}
   );
   gpc606_5 gpc265 (
      {stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[23],stage1_22[39],stage1_21[41],stage1_20[55]}
   );
   gpc606_5 gpc266 (
      {stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[24],stage1_22[40],stage1_21[42],stage1_20[56]}
   );
   gpc606_5 gpc267 (
      {stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[25],stage1_22[41],stage1_21[43],stage1_20[57]}
   );
   gpc606_5 gpc268 (
      {stage0_20[117], stage0_20[118], stage0_20[119], stage0_20[120], stage0_20[121], stage0_20[122]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[26],stage1_22[42],stage1_21[44],stage1_20[58]}
   );
   gpc606_5 gpc269 (
      {stage0_20[123], stage0_20[124], stage0_20[125], stage0_20[126], stage0_20[127], stage0_20[128]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[27],stage1_22[43],stage1_21[45],stage1_20[59]}
   );
   gpc606_5 gpc270 (
      {stage0_20[129], stage0_20[130], stage0_20[131], stage0_20[132], stage0_20[133], stage0_20[134]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[28],stage1_22[44],stage1_21[46],stage1_20[60]}
   );
   gpc606_5 gpc271 (
      {stage0_20[135], stage0_20[136], stage0_20[137], stage0_20[138], stage0_20[139], stage0_20[140]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[29],stage1_22[45],stage1_21[47],stage1_20[61]}
   );
   gpc606_5 gpc272 (
      {stage0_20[141], stage0_20[142], stage0_20[143], stage0_20[144], stage0_20[145], stage0_20[146]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[30],stage1_22[46],stage1_21[48],stage1_20[62]}
   );
   gpc606_5 gpc273 (
      {stage0_20[147], stage0_20[148], stage0_20[149], stage0_20[150], stage0_20[151], stage0_20[152]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[31],stage1_22[47],stage1_21[49],stage1_20[63]}
   );
   gpc606_5 gpc274 (
      {stage0_20[153], stage0_20[154], stage0_20[155], stage0_20[156], stage0_20[157], stage0_20[158]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[32],stage1_22[48],stage1_21[50],stage1_20[64]}
   );
   gpc615_5 gpc275 (
      {stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125], stage0_21[126]},
      {stage0_22[84]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[14],stage1_23[33],stage1_22[49],stage1_21[51]}
   );
   gpc615_5 gpc276 (
      {stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_22[85]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[15],stage1_23[34],stage1_22[50],stage1_21[52]}
   );
   gpc615_5 gpc277 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136]},
      {stage0_22[86]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[16],stage1_23[35],stage1_22[51],stage1_21[53]}
   );
   gpc615_5 gpc278 (
      {stage0_21[137], stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141]},
      {stage0_22[87]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[17],stage1_23[36],stage1_22[52],stage1_21[54]}
   );
   gpc615_5 gpc279 (
      {stage0_21[142], stage0_21[143], stage0_21[144], stage0_21[145], stage0_21[146]},
      {stage0_22[88]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[18],stage1_23[37],stage1_22[53],stage1_21[55]}
   );
   gpc606_5 gpc280 (
      {stage0_22[89], stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[5],stage1_24[19],stage1_23[38],stage1_22[54]}
   );
   gpc606_5 gpc281 (
      {stage0_22[95], stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[6],stage1_24[20],stage1_23[39],stage1_22[55]}
   );
   gpc606_5 gpc282 (
      {stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[7],stage1_24[21],stage1_23[40],stage1_22[56]}
   );
   gpc606_5 gpc283 (
      {stage0_22[107], stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[8],stage1_24[22],stage1_23[41],stage1_22[57]}
   );
   gpc606_5 gpc284 (
      {stage0_22[113], stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[9],stage1_24[23],stage1_23[42],stage1_22[58]}
   );
   gpc606_5 gpc285 (
      {stage0_22[119], stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[10],stage1_24[24],stage1_23[43],stage1_22[59]}
   );
   gpc606_5 gpc286 (
      {stage0_22[125], stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[11],stage1_24[25],stage1_23[44],stage1_22[60]}
   );
   gpc606_5 gpc287 (
      {stage0_22[131], stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[12],stage1_24[26],stage1_23[45],stage1_22[61]}
   );
   gpc615_5 gpc288 (
      {stage0_22[137], stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141]},
      {stage0_23[30]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[13],stage1_24[27],stage1_23[46],stage1_22[62]}
   );
   gpc615_5 gpc289 (
      {stage0_22[142], stage0_22[143], stage0_22[144], stage0_22[145], stage0_22[146]},
      {stage0_23[31]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[14],stage1_24[28],stage1_23[47],stage1_22[63]}
   );
   gpc615_5 gpc290 (
      {stage0_22[147], stage0_22[148], stage0_22[149], stage0_22[150], stage0_22[151]},
      {stage0_23[32]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[15],stage1_24[29],stage1_23[48],stage1_22[64]}
   );
   gpc615_5 gpc291 (
      {stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155], stage0_22[156]},
      {stage0_23[33]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[16],stage1_24[30],stage1_23[49],stage1_22[65]}
   );
   gpc615_5 gpc292 (
      {stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage0_23[34]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[17],stage1_24[31],stage1_23[50],stage1_22[66]}
   );
   gpc606_5 gpc293 (
      {stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[13],stage1_25[18],stage1_24[32],stage1_23[51]}
   );
   gpc606_5 gpc294 (
      {stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[14],stage1_25[19],stage1_24[33],stage1_23[52]}
   );
   gpc606_5 gpc295 (
      {stage0_23[47], stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[15],stage1_25[20],stage1_24[34],stage1_23[53]}
   );
   gpc606_5 gpc296 (
      {stage0_23[53], stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[16],stage1_25[21],stage1_24[35],stage1_23[54]}
   );
   gpc606_5 gpc297 (
      {stage0_23[59], stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[17],stage1_25[22],stage1_24[36],stage1_23[55]}
   );
   gpc606_5 gpc298 (
      {stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[18],stage1_25[23],stage1_24[37],stage1_23[56]}
   );
   gpc606_5 gpc299 (
      {stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[19],stage1_25[24],stage1_24[38],stage1_23[57]}
   );
   gpc606_5 gpc300 (
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[7],stage1_26[20],stage1_25[25],stage1_24[39]}
   );
   gpc606_5 gpc301 (
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[8],stage1_26[21],stage1_25[26],stage1_24[40]}
   );
   gpc606_5 gpc302 (
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[9],stage1_26[22],stage1_25[27],stage1_24[41]}
   );
   gpc606_5 gpc303 (
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[10],stage1_26[23],stage1_25[28],stage1_24[42]}
   );
   gpc606_5 gpc304 (
      {stage0_24[102], stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[11],stage1_26[24],stage1_25[29],stage1_24[43]}
   );
   gpc606_5 gpc305 (
      {stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[12],stage1_26[25],stage1_25[30],stage1_24[44]}
   );
   gpc606_5 gpc306 (
      {stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[13],stage1_26[26],stage1_25[31],stage1_24[45]}
   );
   gpc606_5 gpc307 (
      {stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[14],stage1_26[27],stage1_25[32],stage1_24[46]}
   );
   gpc615_5 gpc308 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46]},
      {stage0_26[48]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[8],stage1_27[15],stage1_26[28],stage1_25[33]}
   );
   gpc615_5 gpc309 (
      {stage0_25[47], stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51]},
      {stage0_26[49]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[9],stage1_27[16],stage1_26[29],stage1_25[34]}
   );
   gpc615_5 gpc310 (
      {stage0_25[52], stage0_25[53], stage0_25[54], stage0_25[55], stage0_25[56]},
      {stage0_26[50]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[10],stage1_27[17],stage1_26[30],stage1_25[35]}
   );
   gpc615_5 gpc311 (
      {stage0_25[57], stage0_25[58], stage0_25[59], stage0_25[60], stage0_25[61]},
      {stage0_26[51]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[11],stage1_27[18],stage1_26[31],stage1_25[36]}
   );
   gpc615_5 gpc312 (
      {stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65], stage0_25[66]},
      {stage0_26[52]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[12],stage1_27[19],stage1_26[32],stage1_25[37]}
   );
   gpc615_5 gpc313 (
      {stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_26[53]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[13],stage1_27[20],stage1_26[33],stage1_25[38]}
   );
   gpc615_5 gpc314 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76]},
      {stage0_26[54]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[14],stage1_27[21],stage1_26[34],stage1_25[39]}
   );
   gpc615_5 gpc315 (
      {stage0_25[77], stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81]},
      {stage0_26[55]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[15],stage1_27[22],stage1_26[35],stage1_25[40]}
   );
   gpc615_5 gpc316 (
      {stage0_25[82], stage0_25[83], stage0_25[84], stage0_25[85], stage0_25[86]},
      {stage0_26[56]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[16],stage1_27[23],stage1_26[36],stage1_25[41]}
   );
   gpc615_5 gpc317 (
      {stage0_25[87], stage0_25[88], stage0_25[89], stage0_25[90], stage0_25[91]},
      {stage0_26[57]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[17],stage1_27[24],stage1_26[37],stage1_25[42]}
   );
   gpc615_5 gpc318 (
      {stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95], stage0_25[96]},
      {stage0_26[58]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[18],stage1_27[25],stage1_26[38],stage1_25[43]}
   );
   gpc615_5 gpc319 (
      {stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_26[59]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[19],stage1_27[26],stage1_26[39],stage1_25[44]}
   );
   gpc615_5 gpc320 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106]},
      {stage0_26[60]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[20],stage1_27[27],stage1_26[40],stage1_25[45]}
   );
   gpc615_5 gpc321 (
      {stage0_25[107], stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111]},
      {stage0_26[61]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[21],stage1_27[28],stage1_26[41],stage1_25[46]}
   );
   gpc615_5 gpc322 (
      {stage0_25[112], stage0_25[113], stage0_25[114], stage0_25[115], stage0_25[116]},
      {stage0_26[62]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[22],stage1_27[29],stage1_26[42],stage1_25[47]}
   );
   gpc615_5 gpc323 (
      {stage0_25[117], stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121]},
      {stage0_26[63]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[23],stage1_27[30],stage1_26[43],stage1_25[48]}
   );
   gpc615_5 gpc324 (
      {stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125], stage0_25[126]},
      {stage0_26[64]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[24],stage1_27[31],stage1_26[44],stage1_25[49]}
   );
   gpc606_5 gpc325 (
      {stage0_26[65], stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[17],stage1_28[25],stage1_27[32],stage1_26[45]}
   );
   gpc606_5 gpc326 (
      {stage0_26[71], stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[18],stage1_28[26],stage1_27[33],stage1_26[46]}
   );
   gpc606_5 gpc327 (
      {stage0_26[77], stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[19],stage1_28[27],stage1_27[34],stage1_26[47]}
   );
   gpc606_5 gpc328 (
      {stage0_26[83], stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[20],stage1_28[28],stage1_27[35],stage1_26[48]}
   );
   gpc606_5 gpc329 (
      {stage0_26[89], stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[21],stage1_28[29],stage1_27[36],stage1_26[49]}
   );
   gpc606_5 gpc330 (
      {stage0_26[95], stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100]},
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage1_30[5],stage1_29[22],stage1_28[30],stage1_27[37],stage1_26[50]}
   );
   gpc606_5 gpc331 (
      {stage0_26[101], stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106]},
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage1_30[6],stage1_29[23],stage1_28[31],stage1_27[38],stage1_26[51]}
   );
   gpc606_5 gpc332 (
      {stage0_26[107], stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112]},
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage1_30[7],stage1_29[24],stage1_28[32],stage1_27[39],stage1_26[52]}
   );
   gpc606_5 gpc333 (
      {stage0_26[113], stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118]},
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage1_30[8],stage1_29[25],stage1_28[33],stage1_27[40],stage1_26[53]}
   );
   gpc606_5 gpc334 (
      {stage0_26[119], stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124]},
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage1_30[9],stage1_29[26],stage1_28[34],stage1_27[41],stage1_26[54]}
   );
   gpc606_5 gpc335 (
      {stage0_26[125], stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130]},
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage1_30[10],stage1_29[27],stage1_28[35],stage1_27[42],stage1_26[55]}
   );
   gpc606_5 gpc336 (
      {stage0_26[131], stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136]},
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage1_30[11],stage1_29[28],stage1_28[36],stage1_27[43],stage1_26[56]}
   );
   gpc606_5 gpc337 (
      {stage0_26[137], stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142]},
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage1_30[12],stage1_29[29],stage1_28[37],stage1_27[44],stage1_26[57]}
   );
   gpc606_5 gpc338 (
      {stage0_26[143], stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148]},
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage1_30[13],stage1_29[30],stage1_28[38],stage1_27[45],stage1_26[58]}
   );
   gpc615_5 gpc339 (
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106]},
      {stage0_28[84]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[14],stage1_29[31],stage1_28[39],stage1_27[46]}
   );
   gpc615_5 gpc340 (
      {stage0_27[107], stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111]},
      {stage0_28[85]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[15],stage1_29[32],stage1_28[40],stage1_27[47]}
   );
   gpc615_5 gpc341 (
      {stage0_27[112], stage0_27[113], stage0_27[114], stage0_27[115], stage0_27[116]},
      {stage0_28[86]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[16],stage1_29[33],stage1_28[41],stage1_27[48]}
   );
   gpc615_5 gpc342 (
      {stage0_27[117], stage0_27[118], stage0_27[119], stage0_27[120], stage0_27[121]},
      {stage0_28[87]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[17],stage1_29[34],stage1_28[42],stage1_27[49]}
   );
   gpc615_5 gpc343 (
      {stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125], stage0_27[126]},
      {stage0_28[88]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[18],stage1_29[35],stage1_28[43],stage1_27[50]}
   );
   gpc615_5 gpc344 (
      {stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage0_28[89]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[19],stage1_29[36],stage1_28[44],stage1_27[51]}
   );
   gpc615_5 gpc345 (
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136]},
      {stage0_28[90]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[20],stage1_29[37],stage1_28[45],stage1_27[52]}
   );
   gpc615_5 gpc346 (
      {stage0_27[137], stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141]},
      {stage0_28[91]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[21],stage1_29[38],stage1_28[46],stage1_27[53]}
   );
   gpc606_5 gpc347 (
      {stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96], stage0_28[97]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[8],stage1_30[22],stage1_29[39],stage1_28[47]}
   );
   gpc606_5 gpc348 (
      {stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102], stage0_28[103]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[9],stage1_30[23],stage1_29[40],stage1_28[48]}
   );
   gpc606_5 gpc349 (
      {stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108], stage0_28[109]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[10],stage1_30[24],stage1_29[41],stage1_28[49]}
   );
   gpc606_5 gpc350 (
      {stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114], stage0_28[115]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[11],stage1_30[25],stage1_29[42],stage1_28[50]}
   );
   gpc606_5 gpc351 (
      {stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120], stage0_28[121]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[12],stage1_30[26],stage1_29[43],stage1_28[51]}
   );
   gpc606_5 gpc352 (
      {stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126], stage0_28[127]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[13],stage1_30[27],stage1_29[44],stage1_28[52]}
   );
   gpc606_5 gpc353 (
      {stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132], stage0_28[133]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[14],stage1_30[28],stage1_29[45],stage1_28[53]}
   );
   gpc606_5 gpc354 (
      {stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138], stage0_28[139]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[15],stage1_30[29],stage1_29[46],stage1_28[54]}
   );
   gpc606_5 gpc355 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[8],stage1_31[16],stage1_30[30],stage1_29[47]}
   );
   gpc606_5 gpc356 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[9],stage1_31[17],stage1_30[31],stage1_29[48]}
   );
   gpc606_5 gpc357 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[10],stage1_31[18],stage1_30[32],stage1_29[49]}
   );
   gpc606_5 gpc358 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[11],stage1_31[19],stage1_30[33],stage1_29[50]}
   );
   gpc606_5 gpc359 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[12],stage1_31[20],stage1_30[34],stage1_29[51]}
   );
   gpc606_5 gpc360 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[13],stage1_31[21],stage1_30[35],stage1_29[52]}
   );
   gpc606_5 gpc361 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[14],stage1_31[22],stage1_30[36],stage1_29[53]}
   );
   gpc606_5 gpc362 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[15],stage1_31[23],stage1_30[37],stage1_29[54]}
   );
   gpc606_5 gpc363 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[16],stage1_31[24],stage1_30[38],stage1_29[55]}
   );
   gpc606_5 gpc364 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[17],stage1_31[25],stage1_30[39],stage1_29[56]}
   );
   gpc606_5 gpc365 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[18],stage1_31[26],stage1_30[40],stage1_29[57]}
   );
   gpc606_5 gpc366 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[19],stage1_31[27],stage1_30[41],stage1_29[58]}
   );
   gpc606_5 gpc367 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[20],stage1_31[28],stage1_30[42],stage1_29[59]}
   );
   gpc606_5 gpc368 (
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[21],stage1_31[29],stage1_30[43],stage1_29[60]}
   );
   gpc606_5 gpc369 (
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[22],stage1_31[30],stage1_30[44],stage1_29[61]}
   );
   gpc606_5 gpc370 (
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[23],stage1_31[31],stage1_30[45],stage1_29[62]}
   );
   gpc1406_5 gpc371 (
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3]},
      {stage0_33[0]},
      {stage1_34[0],stage1_33[16],stage1_32[24],stage1_31[32],stage1_30[46]}
   );
   gpc207_4 gpc372 (
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60]},
      {stage0_32[4], stage0_32[5]},
      {stage1_33[17],stage1_32[25],stage1_31[33],stage1_30[47]}
   );
   gpc207_4 gpc373 (
      {stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66], stage0_30[67]},
      {stage0_32[6], stage0_32[7]},
      {stage1_33[18],stage1_32[26],stage1_31[34],stage1_30[48]}
   );
   gpc207_4 gpc374 (
      {stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72], stage0_30[73], stage0_30[74]},
      {stage0_32[8], stage0_32[9]},
      {stage1_33[19],stage1_32[27],stage1_31[35],stage1_30[49]}
   );
   gpc207_4 gpc375 (
      {stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81]},
      {stage0_32[10], stage0_32[11]},
      {stage1_33[20],stage1_32[28],stage1_31[36],stage1_30[50]}
   );
   gpc207_4 gpc376 (
      {stage0_30[82], stage0_30[83], stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88]},
      {stage0_32[12], stage0_32[13]},
      {stage1_33[21],stage1_32[29],stage1_31[37],stage1_30[51]}
   );
   gpc207_4 gpc377 (
      {stage0_30[89], stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage0_32[14], stage0_32[15]},
      {stage1_33[22],stage1_32[30],stage1_31[38],stage1_30[52]}
   );
   gpc615_5 gpc378 (
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100]},
      {stage0_31[96]},
      {stage0_32[16], stage0_32[17], stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21]},
      {stage1_34[1],stage1_33[23],stage1_32[31],stage1_31[39],stage1_30[53]}
   );
   gpc615_5 gpc379 (
      {stage0_30[101], stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105]},
      {stage0_31[97]},
      {stage0_32[22], stage0_32[23], stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27]},
      {stage1_34[2],stage1_33[24],stage1_32[32],stage1_31[40],stage1_30[54]}
   );
   gpc615_5 gpc380 (
      {stage0_30[106], stage0_30[107], stage0_30[108], stage0_30[109], stage0_30[110]},
      {stage0_31[98]},
      {stage0_32[28], stage0_32[29], stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33]},
      {stage1_34[3],stage1_33[25],stage1_32[33],stage1_31[41],stage1_30[55]}
   );
   gpc615_5 gpc381 (
      {stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage0_32[34]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[0],stage1_34[4],stage1_33[26],stage1_32[34],stage1_31[42]}
   );
   gpc615_5 gpc382 (
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108]},
      {stage0_32[35]},
      {stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage1_35[1],stage1_34[5],stage1_33[27],stage1_32[35],stage1_31[43]}
   );
   gpc606_5 gpc383 (
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[2],stage1_34[6],stage1_33[28],stage1_32[36]}
   );
   gpc606_5 gpc384 (
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[3],stage1_34[7],stage1_33[29],stage1_32[37]}
   );
   gpc606_5 gpc385 (
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52], stage0_32[53]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[4],stage1_34[8],stage1_33[30],stage1_32[38]}
   );
   gpc615_5 gpc386 (
      {stage0_32[54], stage0_32[55], stage0_32[56], stage0_32[57], stage0_32[58]},
      {stage0_33[13]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[5],stage1_34[9],stage1_33[31],stage1_32[39]}
   );
   gpc615_5 gpc387 (
      {stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62], stage0_32[63]},
      {stage0_33[14]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[6],stage1_34[10],stage1_33[32],stage1_32[40]}
   );
   gpc615_5 gpc388 (
      {stage0_32[64], stage0_32[65], stage0_32[66], stage0_32[67], stage0_32[68]},
      {stage0_33[15]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[7],stage1_34[11],stage1_33[33],stage1_32[41]}
   );
   gpc615_5 gpc389 (
      {stage0_32[69], stage0_32[70], stage0_32[71], stage0_32[72], stage0_32[73]},
      {stage0_33[16]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[8],stage1_34[12],stage1_33[34],stage1_32[42]}
   );
   gpc615_5 gpc390 (
      {stage0_32[74], stage0_32[75], stage0_32[76], stage0_32[77], stage0_32[78]},
      {stage0_33[17]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[9],stage1_34[13],stage1_33[35],stage1_32[43]}
   );
   gpc615_5 gpc391 (
      {stage0_32[79], stage0_32[80], stage0_32[81], stage0_32[82], stage0_32[83]},
      {stage0_33[18]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[10],stage1_34[14],stage1_33[36],stage1_32[44]}
   );
   gpc615_5 gpc392 (
      {stage0_32[84], stage0_32[85], stage0_32[86], stage0_32[87], stage0_32[88]},
      {stage0_33[19]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[11],stage1_34[15],stage1_33[37],stage1_32[45]}
   );
   gpc615_5 gpc393 (
      {stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92], stage0_32[93]},
      {stage0_33[20]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[12],stage1_34[16],stage1_33[38],stage1_32[46]}
   );
   gpc615_5 gpc394 (
      {stage0_32[94], stage0_32[95], stage0_32[96], stage0_32[97], stage0_32[98]},
      {stage0_33[21]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[13],stage1_34[17],stage1_33[39],stage1_32[47]}
   );
   gpc615_5 gpc395 (
      {stage0_32[99], stage0_32[100], stage0_32[101], stage0_32[102], stage0_32[103]},
      {stage0_33[22]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[14],stage1_34[18],stage1_33[40],stage1_32[48]}
   );
   gpc615_5 gpc396 (
      {stage0_32[104], stage0_32[105], stage0_32[106], stage0_32[107], stage0_32[108]},
      {stage0_33[23]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[15],stage1_34[19],stage1_33[41],stage1_32[49]}
   );
   gpc615_5 gpc397 (
      {stage0_32[109], stage0_32[110], stage0_32[111], stage0_32[112], stage0_32[113]},
      {stage0_33[24]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[16],stage1_34[20],stage1_33[42],stage1_32[50]}
   );
   gpc615_5 gpc398 (
      {stage0_32[114], stage0_32[115], stage0_32[116], stage0_32[117], stage0_32[118]},
      {stage0_33[25]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[17],stage1_34[21],stage1_33[43],stage1_32[51]}
   );
   gpc615_5 gpc399 (
      {stage0_32[119], stage0_32[120], stage0_32[121], stage0_32[122], stage0_32[123]},
      {stage0_33[26]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[18],stage1_34[22],stage1_33[44],stage1_32[52]}
   );
   gpc615_5 gpc400 (
      {stage0_32[124], stage0_32[125], stage0_32[126], stage0_32[127], stage0_32[128]},
      {stage0_33[27]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[19],stage1_34[23],stage1_33[45],stage1_32[53]}
   );
   gpc606_5 gpc401 (
      {stage0_33[28], stage0_33[29], stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[18],stage1_35[20],stage1_34[24],stage1_33[46]}
   );
   gpc606_5 gpc402 (
      {stage0_33[34], stage0_33[35], stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[19],stage1_35[21],stage1_34[25],stage1_33[47]}
   );
   gpc606_5 gpc403 (
      {stage0_33[40], stage0_33[41], stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[20],stage1_35[22],stage1_34[26],stage1_33[48]}
   );
   gpc606_5 gpc404 (
      {stage0_33[46], stage0_33[47], stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[21],stage1_35[23],stage1_34[27],stage1_33[49]}
   );
   gpc606_5 gpc405 (
      {stage0_33[52], stage0_33[53], stage0_33[54], stage0_33[55], stage0_33[56], stage0_33[57]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[22],stage1_35[24],stage1_34[28],stage1_33[50]}
   );
   gpc606_5 gpc406 (
      {stage0_33[58], stage0_33[59], stage0_33[60], stage0_33[61], stage0_33[62], stage0_33[63]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[23],stage1_35[25],stage1_34[29],stage1_33[51]}
   );
   gpc606_5 gpc407 (
      {stage0_33[64], stage0_33[65], stage0_33[66], stage0_33[67], stage0_33[68], stage0_33[69]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[24],stage1_35[26],stage1_34[30],stage1_33[52]}
   );
   gpc606_5 gpc408 (
      {stage0_33[70], stage0_33[71], stage0_33[72], stage0_33[73], stage0_33[74], stage0_33[75]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[25],stage1_35[27],stage1_34[31],stage1_33[53]}
   );
   gpc606_5 gpc409 (
      {stage0_33[76], stage0_33[77], stage0_33[78], stage0_33[79], stage0_33[80], stage0_33[81]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[26],stage1_35[28],stage1_34[32],stage1_33[54]}
   );
   gpc606_5 gpc410 (
      {stage0_33[82], stage0_33[83], stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[27],stage1_35[29],stage1_34[33],stage1_33[55]}
   );
   gpc606_5 gpc411 (
      {stage0_33[88], stage0_33[89], stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[28],stage1_35[30],stage1_34[34],stage1_33[56]}
   );
   gpc606_5 gpc412 (
      {stage0_33[94], stage0_33[95], stage0_33[96], stage0_33[97], stage0_33[98], stage0_33[99]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[29],stage1_35[31],stage1_34[35],stage1_33[57]}
   );
   gpc606_5 gpc413 (
      {stage0_33[100], stage0_33[101], stage0_33[102], stage0_33[103], stage0_33[104], stage0_33[105]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage1_37[12],stage1_36[30],stage1_35[32],stage1_34[36],stage1_33[58]}
   );
   gpc606_5 gpc414 (
      {stage0_33[106], stage0_33[107], stage0_33[108], stage0_33[109], stage0_33[110], stage0_33[111]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage1_37[13],stage1_36[31],stage1_35[33],stage1_34[37],stage1_33[59]}
   );
   gpc606_5 gpc415 (
      {stage0_33[112], stage0_33[113], stage0_33[114], stage0_33[115], stage0_33[116], stage0_33[117]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage1_37[14],stage1_36[32],stage1_35[34],stage1_34[38],stage1_33[60]}
   );
   gpc606_5 gpc416 (
      {stage0_33[118], stage0_33[119], stage0_33[120], stage0_33[121], stage0_33[122], stage0_33[123]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage1_37[15],stage1_36[33],stage1_35[35],stage1_34[39],stage1_33[61]}
   );
   gpc606_5 gpc417 (
      {stage0_33[124], stage0_33[125], stage0_33[126], stage0_33[127], stage0_33[128], stage0_33[129]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage1_37[16],stage1_36[34],stage1_35[36],stage1_34[40],stage1_33[62]}
   );
   gpc606_5 gpc418 (
      {stage0_33[130], stage0_33[131], stage0_33[132], stage0_33[133], stage0_33[134], stage0_33[135]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage1_37[17],stage1_36[35],stage1_35[37],stage1_34[41],stage1_33[63]}
   );
   gpc615_5 gpc419 (
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112]},
      {stage0_35[108]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[18],stage1_36[36],stage1_35[38],stage1_34[42]}
   );
   gpc615_5 gpc420 (
      {stage0_34[113], stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117]},
      {stage0_35[109]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[19],stage1_36[37],stage1_35[39],stage1_34[43]}
   );
   gpc615_5 gpc421 (
      {stage0_34[118], stage0_34[119], stage0_34[120], stage0_34[121], stage0_34[122]},
      {stage0_35[110]},
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17]},
      {stage1_38[2],stage1_37[20],stage1_36[38],stage1_35[40],stage1_34[44]}
   );
   gpc615_5 gpc422 (
      {stage0_34[123], stage0_34[124], stage0_34[125], stage0_34[126], stage0_34[127]},
      {stage0_35[111]},
      {stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23]},
      {stage1_38[3],stage1_37[21],stage1_36[39],stage1_35[41],stage1_34[45]}
   );
   gpc615_5 gpc423 (
      {stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131], stage0_34[132]},
      {stage0_35[112]},
      {stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29]},
      {stage1_38[4],stage1_37[22],stage1_36[40],stage1_35[42],stage1_34[46]}
   );
   gpc615_5 gpc424 (
      {stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage0_35[113]},
      {stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35]},
      {stage1_38[5],stage1_37[23],stage1_36[41],stage1_35[43],stage1_34[47]}
   );
   gpc615_5 gpc425 (
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142]},
      {stage0_35[114]},
      {stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41]},
      {stage1_38[6],stage1_37[24],stage1_36[42],stage1_35[44],stage1_34[48]}
   );
   gpc615_5 gpc426 (
      {stage0_34[143], stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147]},
      {stage0_35[115]},
      {stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47]},
      {stage1_38[7],stage1_37[25],stage1_36[43],stage1_35[45],stage1_34[49]}
   );
   gpc615_5 gpc427 (
      {stage0_34[148], stage0_34[149], stage0_34[150], stage0_34[151], stage0_34[152]},
      {stage0_35[116]},
      {stage0_36[48], stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53]},
      {stage1_38[8],stage1_37[26],stage1_36[44],stage1_35[46],stage1_34[50]}
   );
   gpc615_5 gpc428 (
      {stage0_34[153], stage0_34[154], stage0_34[155], stage0_34[156], stage0_34[157]},
      {stage0_35[117]},
      {stage0_36[54], stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59]},
      {stage1_38[9],stage1_37[27],stage1_36[45],stage1_35[47],stage1_34[51]}
   );
   gpc615_5 gpc429 (
      {stage0_35[118], stage0_35[119], stage0_35[120], stage0_35[121], stage0_35[122]},
      {stage0_36[60]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[10],stage1_37[28],stage1_36[46],stage1_35[48]}
   );
   gpc615_5 gpc430 (
      {stage0_35[123], stage0_35[124], stage0_35[125], stage0_35[126], stage0_35[127]},
      {stage0_36[61]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[11],stage1_37[29],stage1_36[47],stage1_35[49]}
   );
   gpc615_5 gpc431 (
      {stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131], stage0_35[132]},
      {stage0_36[62]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[12],stage1_37[30],stage1_36[48],stage1_35[50]}
   );
   gpc615_5 gpc432 (
      {stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage0_36[63]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[13],stage1_37[31],stage1_36[49],stage1_35[51]}
   );
   gpc615_5 gpc433 (
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142]},
      {stage0_36[64]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[14],stage1_37[32],stage1_36[50],stage1_35[52]}
   );
   gpc615_5 gpc434 (
      {stage0_35[143], stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147]},
      {stage0_36[65]},
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage1_39[5],stage1_38[15],stage1_37[33],stage1_36[51],stage1_35[53]}
   );
   gpc615_5 gpc435 (
      {stage0_35[148], stage0_35[149], stage0_35[150], stage0_35[151], stage0_35[152]},
      {stage0_36[66]},
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage1_39[6],stage1_38[16],stage1_37[34],stage1_36[52],stage1_35[54]}
   );
   gpc615_5 gpc436 (
      {stage0_35[153], stage0_35[154], stage0_35[155], stage0_35[156], stage0_35[157]},
      {stage0_36[67]},
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage1_39[7],stage1_38[17],stage1_37[35],stage1_36[53],stage1_35[55]}
   );
   gpc606_5 gpc437 (
      {stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71], stage0_36[72], stage0_36[73]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[8],stage1_38[18],stage1_37[36],stage1_36[54]}
   );
   gpc606_5 gpc438 (
      {stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77], stage0_36[78], stage0_36[79]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[9],stage1_38[19],stage1_37[37],stage1_36[55]}
   );
   gpc606_5 gpc439 (
      {stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83], stage0_36[84], stage0_36[85]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[10],stage1_38[20],stage1_37[38],stage1_36[56]}
   );
   gpc606_5 gpc440 (
      {stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89], stage0_36[90], stage0_36[91]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[11],stage1_38[21],stage1_37[39],stage1_36[57]}
   );
   gpc606_5 gpc441 (
      {stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95], stage0_36[96], stage0_36[97]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[12],stage1_38[22],stage1_37[40],stage1_36[58]}
   );
   gpc606_5 gpc442 (
      {stage0_36[98], stage0_36[99], stage0_36[100], stage0_36[101], stage0_36[102], stage0_36[103]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[13],stage1_38[23],stage1_37[41],stage1_36[59]}
   );
   gpc606_5 gpc443 (
      {stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107], stage0_36[108], stage0_36[109]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[14],stage1_38[24],stage1_37[42],stage1_36[60]}
   );
   gpc606_5 gpc444 (
      {stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113], stage0_36[114], stage0_36[115]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[15],stage1_38[25],stage1_37[43],stage1_36[61]}
   );
   gpc606_5 gpc445 (
      {stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119], stage0_36[120], stage0_36[121]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[16],stage1_38[26],stage1_37[44],stage1_36[62]}
   );
   gpc606_5 gpc446 (
      {stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126], stage0_36[127]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[17],stage1_38[27],stage1_37[45],stage1_36[63]}
   );
   gpc606_5 gpc447 (
      {stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132], stage0_36[133]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[18],stage1_38[28],stage1_37[46],stage1_36[64]}
   );
   gpc606_5 gpc448 (
      {stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138], stage0_36[139]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[19],stage1_38[29],stage1_37[47],stage1_36[65]}
   );
   gpc606_5 gpc449 (
      {stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144], stage0_36[145]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[20],stage1_38[30],stage1_37[48],stage1_36[66]}
   );
   gpc606_5 gpc450 (
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[13],stage1_39[21],stage1_38[31],stage1_37[49]}
   );
   gpc606_5 gpc451 (
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[14],stage1_39[22],stage1_38[32],stage1_37[50]}
   );
   gpc606_5 gpc452 (
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[15],stage1_39[23],stage1_38[33],stage1_37[51]}
   );
   gpc606_5 gpc453 (
      {stage0_37[66], stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[16],stage1_39[24],stage1_38[34],stage1_37[52]}
   );
   gpc606_5 gpc454 (
      {stage0_37[72], stage0_37[73], stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[17],stage1_39[25],stage1_38[35],stage1_37[53]}
   );
   gpc606_5 gpc455 (
      {stage0_37[78], stage0_37[79], stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[18],stage1_39[26],stage1_38[36],stage1_37[54]}
   );
   gpc606_5 gpc456 (
      {stage0_37[84], stage0_37[85], stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[19],stage1_39[27],stage1_38[37],stage1_37[55]}
   );
   gpc615_5 gpc457 (
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82]},
      {stage0_39[42]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[7],stage1_40[20],stage1_39[28],stage1_38[38]}
   );
   gpc615_5 gpc458 (
      {stage0_38[83], stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87]},
      {stage0_39[43]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[8],stage1_40[21],stage1_39[29],stage1_38[39]}
   );
   gpc615_5 gpc459 (
      {stage0_38[88], stage0_38[89], stage0_38[90], stage0_38[91], stage0_38[92]},
      {stage0_39[44]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[9],stage1_40[22],stage1_39[30],stage1_38[40]}
   );
   gpc615_5 gpc460 (
      {stage0_38[93], stage0_38[94], stage0_38[95], stage0_38[96], stage0_38[97]},
      {stage0_39[45]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[10],stage1_40[23],stage1_39[31],stage1_38[41]}
   );
   gpc615_5 gpc461 (
      {stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101], stage0_38[102]},
      {stage0_39[46]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[11],stage1_40[24],stage1_39[32],stage1_38[42]}
   );
   gpc615_5 gpc462 (
      {stage0_38[103], stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107]},
      {stage0_39[47]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[12],stage1_40[25],stage1_39[33],stage1_38[43]}
   );
   gpc615_5 gpc463 (
      {stage0_38[108], stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112]},
      {stage0_39[48]},
      {stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39], stage0_40[40], stage0_40[41]},
      {stage1_42[6],stage1_41[13],stage1_40[26],stage1_39[34],stage1_38[44]}
   );
   gpc615_5 gpc464 (
      {stage0_38[113], stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117]},
      {stage0_39[49]},
      {stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45], stage0_40[46], stage0_40[47]},
      {stage1_42[7],stage1_41[14],stage1_40[27],stage1_39[35],stage1_38[45]}
   );
   gpc615_5 gpc465 (
      {stage0_38[118], stage0_38[119], stage0_38[120], stage0_38[121], stage0_38[122]},
      {stage0_39[50]},
      {stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51], stage0_40[52], stage0_40[53]},
      {stage1_42[8],stage1_41[15],stage1_40[28],stage1_39[36],stage1_38[46]}
   );
   gpc615_5 gpc466 (
      {stage0_38[123], stage0_38[124], stage0_38[125], stage0_38[126], stage0_38[127]},
      {stage0_39[51]},
      {stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57], stage0_40[58], stage0_40[59]},
      {stage1_42[9],stage1_41[16],stage1_40[29],stage1_39[37],stage1_38[47]}
   );
   gpc615_5 gpc467 (
      {stage0_38[128], stage0_38[129], stage0_38[130], stage0_38[131], stage0_38[132]},
      {stage0_39[52]},
      {stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63], stage0_40[64], stage0_40[65]},
      {stage1_42[10],stage1_41[17],stage1_40[30],stage1_39[38],stage1_38[48]}
   );
   gpc615_5 gpc468 (
      {stage0_38[133], stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137]},
      {stage0_39[53]},
      {stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69], stage0_40[70], stage0_40[71]},
      {stage1_42[11],stage1_41[18],stage1_40[31],stage1_39[39],stage1_38[49]}
   );
   gpc615_5 gpc469 (
      {stage0_38[138], stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142]},
      {stage0_39[54]},
      {stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75], stage0_40[76], stage0_40[77]},
      {stage1_42[12],stage1_41[19],stage1_40[32],stage1_39[40],stage1_38[50]}
   );
   gpc615_5 gpc470 (
      {stage0_38[143], stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147]},
      {stage0_39[55]},
      {stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81], stage0_40[82], stage0_40[83]},
      {stage1_42[13],stage1_41[20],stage1_40[33],stage1_39[41],stage1_38[51]}
   );
   gpc615_5 gpc471 (
      {stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59], stage0_39[60]},
      {stage0_40[84]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[14],stage1_41[21],stage1_40[34],stage1_39[42]}
   );
   gpc615_5 gpc472 (
      {stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage0_40[85]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[15],stage1_41[22],stage1_40[35],stage1_39[43]}
   );
   gpc615_5 gpc473 (
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70]},
      {stage0_40[86]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[16],stage1_41[23],stage1_40[36],stage1_39[44]}
   );
   gpc615_5 gpc474 (
      {stage0_39[71], stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75]},
      {stage0_40[87]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[17],stage1_41[24],stage1_40[37],stage1_39[45]}
   );
   gpc615_5 gpc475 (
      {stage0_39[76], stage0_39[77], stage0_39[78], stage0_39[79], stage0_39[80]},
      {stage0_40[88]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[18],stage1_41[25],stage1_40[38],stage1_39[46]}
   );
   gpc615_5 gpc476 (
      {stage0_39[81], stage0_39[82], stage0_39[83], stage0_39[84], stage0_39[85]},
      {stage0_40[89]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[19],stage1_41[26],stage1_40[39],stage1_39[47]}
   );
   gpc615_5 gpc477 (
      {stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89], stage0_39[90]},
      {stage0_40[90]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[20],stage1_41[27],stage1_40[40],stage1_39[48]}
   );
   gpc615_5 gpc478 (
      {stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage0_40[91]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[21],stage1_41[28],stage1_40[41],stage1_39[49]}
   );
   gpc615_5 gpc479 (
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100]},
      {stage0_40[92]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[22],stage1_41[29],stage1_40[42],stage1_39[50]}
   );
   gpc615_5 gpc480 (
      {stage0_39[101], stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105]},
      {stage0_40[93]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[23],stage1_41[30],stage1_40[43],stage1_39[51]}
   );
   gpc615_5 gpc481 (
      {stage0_39[106], stage0_39[107], stage0_39[108], stage0_39[109], stage0_39[110]},
      {stage0_40[94]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[24],stage1_41[31],stage1_40[44],stage1_39[52]}
   );
   gpc615_5 gpc482 (
      {stage0_39[111], stage0_39[112], stage0_39[113], stage0_39[114], stage0_39[115]},
      {stage0_40[95]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[25],stage1_41[32],stage1_40[45],stage1_39[53]}
   );
   gpc615_5 gpc483 (
      {stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119], stage0_39[120]},
      {stage0_40[96]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[26],stage1_41[33],stage1_40[46],stage1_39[54]}
   );
   gpc615_5 gpc484 (
      {stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage0_40[97]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[27],stage1_41[34],stage1_40[47],stage1_39[55]}
   );
   gpc615_5 gpc485 (
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130]},
      {stage0_40[98]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[28],stage1_41[35],stage1_40[48],stage1_39[56]}
   );
   gpc615_5 gpc486 (
      {stage0_39[131], stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135]},
      {stage0_40[99]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage1_43[15],stage1_42[29],stage1_41[36],stage1_40[49],stage1_39[57]}
   );
   gpc615_5 gpc487 (
      {stage0_39[136], stage0_39[137], stage0_39[138], stage0_39[139], stage0_39[140]},
      {stage0_40[100]},
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage1_43[16],stage1_42[30],stage1_41[37],stage1_40[50],stage1_39[58]}
   );
   gpc615_5 gpc488 (
      {stage0_39[141], stage0_39[142], stage0_39[143], stage0_39[144], stage0_39[145]},
      {stage0_40[101]},
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage1_43[17],stage1_42[31],stage1_41[38],stage1_40[51],stage1_39[59]}
   );
   gpc615_5 gpc489 (
      {stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149], stage0_39[150]},
      {stage0_40[102]},
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage1_43[18],stage1_42[32],stage1_41[39],stage1_40[52],stage1_39[60]}
   );
   gpc615_5 gpc490 (
      {stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage0_40[103]},
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage1_43[19],stage1_42[33],stage1_41[40],stage1_40[53],stage1_39[61]}
   );
   gpc606_5 gpc491 (
      {stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107], stage0_40[108], stage0_40[109]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[20],stage1_42[34],stage1_41[41],stage1_40[54]}
   );
   gpc606_5 gpc492 (
      {stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113], stage0_40[114], stage0_40[115]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[21],stage1_42[35],stage1_41[42],stage1_40[55]}
   );
   gpc606_5 gpc493 (
      {stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119], stage0_40[120], stage0_40[121]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[22],stage1_42[36],stage1_41[43],stage1_40[56]}
   );
   gpc606_5 gpc494 (
      {stage0_40[122], stage0_40[123], stage0_40[124], stage0_40[125], stage0_40[126], stage0_40[127]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[23],stage1_42[37],stage1_41[44],stage1_40[57]}
   );
   gpc606_5 gpc495 (
      {stage0_40[128], stage0_40[129], stage0_40[130], stage0_40[131], stage0_40[132], stage0_40[133]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[24],stage1_42[38],stage1_41[45],stage1_40[58]}
   );
   gpc606_5 gpc496 (
      {stage0_40[134], stage0_40[135], stage0_40[136], stage0_40[137], stage0_40[138], stage0_40[139]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[25],stage1_42[39],stage1_41[46],stage1_40[59]}
   );
   gpc606_5 gpc497 (
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[6],stage1_43[26],stage1_42[40],stage1_41[47]}
   );
   gpc606_5 gpc498 (
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[7],stage1_43[27],stage1_42[41],stage1_41[48]}
   );
   gpc606_5 gpc499 (
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[8],stage1_43[28],stage1_42[42],stage1_41[49]}
   );
   gpc606_5 gpc500 (
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[3],stage1_44[9],stage1_43[29],stage1_42[43]}
   );
   gpc606_5 gpc501 (
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[4],stage1_44[10],stage1_43[30],stage1_42[44]}
   );
   gpc606_5 gpc502 (
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[5],stage1_44[11],stage1_43[31],stage1_42[45]}
   );
   gpc606_5 gpc503 (
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[6],stage1_44[12],stage1_43[32],stage1_42[46]}
   );
   gpc606_5 gpc504 (
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[7],stage1_44[13],stage1_43[33],stage1_42[47]}
   );
   gpc615_5 gpc505 (
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70]},
      {stage0_43[18]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[8],stage1_44[14],stage1_43[34],stage1_42[48]}
   );
   gpc615_5 gpc506 (
      {stage0_42[71], stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75]},
      {stage0_43[19]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[9],stage1_44[15],stage1_43[35],stage1_42[49]}
   );
   gpc615_5 gpc507 (
      {stage0_42[76], stage0_42[77], stage0_42[78], stage0_42[79], stage0_42[80]},
      {stage0_43[20]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[10],stage1_44[16],stage1_43[36],stage1_42[50]}
   );
   gpc615_5 gpc508 (
      {stage0_42[81], stage0_42[82], stage0_42[83], stage0_42[84], stage0_42[85]},
      {stage0_43[21]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[11],stage1_44[17],stage1_43[37],stage1_42[51]}
   );
   gpc615_5 gpc509 (
      {stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89], stage0_42[90]},
      {stage0_43[22]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[12],stage1_44[18],stage1_43[38],stage1_42[52]}
   );
   gpc615_5 gpc510 (
      {stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage0_43[23]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[13],stage1_44[19],stage1_43[39],stage1_42[53]}
   );
   gpc615_5 gpc511 (
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100]},
      {stage0_43[24]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[14],stage1_44[20],stage1_43[40],stage1_42[54]}
   );
   gpc615_5 gpc512 (
      {stage0_42[101], stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105]},
      {stage0_43[25]},
      {stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76], stage0_44[77]},
      {stage1_46[12],stage1_45[15],stage1_44[21],stage1_43[41],stage1_42[55]}
   );
   gpc615_5 gpc513 (
      {stage0_42[106], stage0_42[107], stage0_42[108], stage0_42[109], stage0_42[110]},
      {stage0_43[26]},
      {stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82], stage0_44[83]},
      {stage1_46[13],stage1_45[16],stage1_44[22],stage1_43[42],stage1_42[56]}
   );
   gpc615_5 gpc514 (
      {stage0_42[111], stage0_42[112], stage0_42[113], stage0_42[114], stage0_42[115]},
      {stage0_43[27]},
      {stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88], stage0_44[89]},
      {stage1_46[14],stage1_45[17],stage1_44[23],stage1_43[43],stage1_42[57]}
   );
   gpc615_5 gpc515 (
      {stage0_42[116], stage0_42[117], stage0_42[118], stage0_42[119], stage0_42[120]},
      {stage0_43[28]},
      {stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94], stage0_44[95]},
      {stage1_46[15],stage1_45[18],stage1_44[24],stage1_43[44],stage1_42[58]}
   );
   gpc615_5 gpc516 (
      {stage0_42[121], stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125]},
      {stage0_43[29]},
      {stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100], stage0_44[101]},
      {stage1_46[16],stage1_45[19],stage1_44[25],stage1_43[45],stage1_42[59]}
   );
   gpc606_5 gpc517 (
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[17],stage1_45[20],stage1_44[26],stage1_43[46]}
   );
   gpc606_5 gpc518 (
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[18],stage1_45[21],stage1_44[27],stage1_43[47]}
   );
   gpc606_5 gpc519 (
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[19],stage1_45[22],stage1_44[28],stage1_43[48]}
   );
   gpc606_5 gpc520 (
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[20],stage1_45[23],stage1_44[29],stage1_43[49]}
   );
   gpc606_5 gpc521 (
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[21],stage1_45[24],stage1_44[30],stage1_43[50]}
   );
   gpc606_5 gpc522 (
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[22],stage1_45[25],stage1_44[31],stage1_43[51]}
   );
   gpc606_5 gpc523 (
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[23],stage1_45[26],stage1_44[32],stage1_43[52]}
   );
   gpc606_5 gpc524 (
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[24],stage1_45[27],stage1_44[33],stage1_43[53]}
   );
   gpc606_5 gpc525 (
      {stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106], stage0_44[107]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[8],stage1_46[25],stage1_45[28],stage1_44[34]}
   );
   gpc606_5 gpc526 (
      {stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112], stage0_44[113]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[9],stage1_46[26],stage1_45[29],stage1_44[35]}
   );
   gpc606_5 gpc527 (
      {stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118], stage0_44[119]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[10],stage1_46[27],stage1_45[30],stage1_44[36]}
   );
   gpc606_5 gpc528 (
      {stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124], stage0_44[125]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[11],stage1_46[28],stage1_45[31],stage1_44[37]}
   );
   gpc606_5 gpc529 (
      {stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130], stage0_44[131]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[12],stage1_46[29],stage1_45[32],stage1_44[38]}
   );
   gpc606_5 gpc530 (
      {stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136], stage0_44[137]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[13],stage1_46[30],stage1_45[33],stage1_44[39]}
   );
   gpc606_5 gpc531 (
      {stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142], stage0_44[143]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[14],stage1_46[31],stage1_45[34],stage1_44[40]}
   );
   gpc606_5 gpc532 (
      {stage0_44[144], stage0_44[145], stage0_44[146], stage0_44[147], stage0_44[148], stage0_44[149]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[15],stage1_46[32],stage1_45[35],stage1_44[41]}
   );
   gpc615_5 gpc533 (
      {stage0_44[150], stage0_44[151], stage0_44[152], stage0_44[153], stage0_44[154]},
      {stage0_45[48]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[16],stage1_46[33],stage1_45[36],stage1_44[42]}
   );
   gpc615_5 gpc534 (
      {stage0_44[155], stage0_44[156], stage0_44[157], stage0_44[158], stage0_44[159]},
      {stage0_45[49]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[17],stage1_46[34],stage1_45[37],stage1_44[43]}
   );
   gpc606_5 gpc535 (
      {stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53], stage0_45[54], stage0_45[55]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[10],stage1_47[18],stage1_46[35],stage1_45[38]}
   );
   gpc615_5 gpc536 (
      {stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59], stage0_45[60]},
      {stage0_46[60]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[11],stage1_47[19],stage1_46[36],stage1_45[39]}
   );
   gpc615_5 gpc537 (
      {stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage0_46[61]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[12],stage1_47[20],stage1_46[37],stage1_45[40]}
   );
   gpc615_5 gpc538 (
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70]},
      {stage0_46[62]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[13],stage1_47[21],stage1_46[38],stage1_45[41]}
   );
   gpc615_5 gpc539 (
      {stage0_45[71], stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75]},
      {stage0_46[63]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[14],stage1_47[22],stage1_46[39],stage1_45[42]}
   );
   gpc615_5 gpc540 (
      {stage0_45[76], stage0_45[77], stage0_45[78], stage0_45[79], stage0_45[80]},
      {stage0_46[64]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[15],stage1_47[23],stage1_46[40],stage1_45[43]}
   );
   gpc615_5 gpc541 (
      {stage0_45[81], stage0_45[82], stage0_45[83], stage0_45[84], stage0_45[85]},
      {stage0_46[65]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[16],stage1_47[24],stage1_46[41],stage1_45[44]}
   );
   gpc615_5 gpc542 (
      {stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89], stage0_45[90]},
      {stage0_46[66]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[17],stage1_47[25],stage1_46[42],stage1_45[45]}
   );
   gpc615_5 gpc543 (
      {stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage0_46[67]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[18],stage1_47[26],stage1_46[43],stage1_45[46]}
   );
   gpc615_5 gpc544 (
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100]},
      {stage0_46[68]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[19],stage1_47[27],stage1_46[44],stage1_45[47]}
   );
   gpc615_5 gpc545 (
      {stage0_45[101], stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105]},
      {stage0_46[69]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[20],stage1_47[28],stage1_46[45],stage1_45[48]}
   );
   gpc615_5 gpc546 (
      {stage0_45[106], stage0_45[107], stage0_45[108], stage0_45[109], stage0_45[110]},
      {stage0_46[70]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[21],stage1_47[29],stage1_46[46],stage1_45[49]}
   );
   gpc615_5 gpc547 (
      {stage0_45[111], stage0_45[112], stage0_45[113], stage0_45[114], stage0_45[115]},
      {stage0_46[71]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[22],stage1_47[30],stage1_46[47],stage1_45[50]}
   );
   gpc615_5 gpc548 (
      {stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119], stage0_45[120]},
      {stage0_46[72]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[23],stage1_47[31],stage1_46[48],stage1_45[51]}
   );
   gpc117_4 gpc549 (
      {stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77], stage0_46[78], stage0_46[79]},
      {stage0_47[84]},
      {stage0_48[0]},
      {stage1_49[14],stage1_48[24],stage1_47[32],stage1_46[49]}
   );
   gpc117_4 gpc550 (
      {stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83], stage0_46[84], stage0_46[85], stage0_46[86]},
      {stage0_47[85]},
      {stage0_48[1]},
      {stage1_49[15],stage1_48[25],stage1_47[33],stage1_46[50]}
   );
   gpc117_4 gpc551 (
      {stage0_46[87], stage0_46[88], stage0_46[89], stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93]},
      {stage0_47[86]},
      {stage0_48[2]},
      {stage1_49[16],stage1_48[26],stage1_47[34],stage1_46[51]}
   );
   gpc117_4 gpc552 (
      {stage0_46[94], stage0_46[95], stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100]},
      {stage0_47[87]},
      {stage0_48[3]},
      {stage1_49[17],stage1_48[27],stage1_47[35],stage1_46[52]}
   );
   gpc117_4 gpc553 (
      {stage0_46[101], stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage0_47[88]},
      {stage0_48[4]},
      {stage1_49[18],stage1_48[28],stage1_47[36],stage1_46[53]}
   );
   gpc117_4 gpc554 (
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113], stage0_46[114]},
      {stage0_47[89]},
      {stage0_48[5]},
      {stage1_49[19],stage1_48[29],stage1_47[37],stage1_46[54]}
   );
   gpc117_4 gpc555 (
      {stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119], stage0_46[120], stage0_46[121]},
      {stage0_47[90]},
      {stage0_48[6]},
      {stage1_49[20],stage1_48[30],stage1_47[38],stage1_46[55]}
   );
   gpc606_5 gpc556 (
      {stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125], stage0_46[126], stage0_46[127]},
      {stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11], stage0_48[12]},
      {stage1_50[0],stage1_49[21],stage1_48[31],stage1_47[39],stage1_46[56]}
   );
   gpc606_5 gpc557 (
      {stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131], stage0_46[132], stage0_46[133]},
      {stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17], stage0_48[18]},
      {stage1_50[1],stage1_49[22],stage1_48[32],stage1_47[40],stage1_46[57]}
   );
   gpc606_5 gpc558 (
      {stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137], stage0_46[138], stage0_46[139]},
      {stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23], stage0_48[24]},
      {stage1_50[2],stage1_49[23],stage1_48[33],stage1_47[41],stage1_46[58]}
   );
   gpc606_5 gpc559 (
      {stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143], stage0_46[144], stage0_46[145]},
      {stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29], stage0_48[30]},
      {stage1_50[3],stage1_49[24],stage1_48[34],stage1_47[42],stage1_46[59]}
   );
   gpc615_5 gpc560 (
      {stage0_46[146], stage0_46[147], stage0_46[148], stage0_46[149], stage0_46[150]},
      {stage0_47[91]},
      {stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35], stage0_48[36]},
      {stage1_50[4],stage1_49[25],stage1_48[35],stage1_47[43],stage1_46[60]}
   );
   gpc615_5 gpc561 (
      {stage0_46[151], stage0_46[152], stage0_46[153], stage0_46[154], stage0_46[155]},
      {stage0_47[92]},
      {stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41], stage0_48[42]},
      {stage1_50[5],stage1_49[26],stage1_48[36],stage1_47[44],stage1_46[61]}
   );
   gpc615_5 gpc562 (
      {stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159], stage0_46[160]},
      {stage0_47[93]},
      {stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47], stage0_48[48]},
      {stage1_50[6],stage1_49[27],stage1_48[37],stage1_47[45],stage1_46[62]}
   );
   gpc606_5 gpc563 (
      {stage0_47[94], stage0_47[95], stage0_47[96], stage0_47[97], stage0_47[98], stage0_47[99]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[7],stage1_49[28],stage1_48[38],stage1_47[46]}
   );
   gpc606_5 gpc564 (
      {stage0_47[100], stage0_47[101], stage0_47[102], stage0_47[103], stage0_47[104], stage0_47[105]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[8],stage1_49[29],stage1_48[39],stage1_47[47]}
   );
   gpc606_5 gpc565 (
      {stage0_47[106], stage0_47[107], stage0_47[108], stage0_47[109], stage0_47[110], stage0_47[111]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[9],stage1_49[30],stage1_48[40],stage1_47[48]}
   );
   gpc606_5 gpc566 (
      {stage0_47[112], stage0_47[113], stage0_47[114], stage0_47[115], stage0_47[116], stage0_47[117]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[10],stage1_49[31],stage1_48[41],stage1_47[49]}
   );
   gpc606_5 gpc567 (
      {stage0_47[118], stage0_47[119], stage0_47[120], stage0_47[121], stage0_47[122], stage0_47[123]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[11],stage1_49[32],stage1_48[42],stage1_47[50]}
   );
   gpc606_5 gpc568 (
      {stage0_47[124], stage0_47[125], stage0_47[126], stage0_47[127], stage0_47[128], stage0_47[129]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[12],stage1_49[33],stage1_48[43],stage1_47[51]}
   );
   gpc606_5 gpc569 (
      {stage0_47[130], stage0_47[131], stage0_47[132], stage0_47[133], stage0_47[134], stage0_47[135]},
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage1_51[6],stage1_50[13],stage1_49[34],stage1_48[44],stage1_47[52]}
   );
   gpc606_5 gpc570 (
      {stage0_47[136], stage0_47[137], stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141]},
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage1_51[7],stage1_50[14],stage1_49[35],stage1_48[45],stage1_47[53]}
   );
   gpc615_5 gpc571 (
      {stage0_47[142], stage0_47[143], stage0_47[144], stage0_47[145], stage0_47[146]},
      {stage0_48[49]},
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage1_51[8],stage1_50[15],stage1_49[36],stage1_48[46],stage1_47[54]}
   );
   gpc615_5 gpc572 (
      {stage0_47[147], stage0_47[148], stage0_47[149], stage0_47[150], stage0_47[151]},
      {stage0_48[50]},
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage1_51[9],stage1_50[16],stage1_49[37],stage1_48[47],stage1_47[55]}
   );
   gpc615_5 gpc573 (
      {stage0_47[152], stage0_47[153], stage0_47[154], stage0_47[155], stage0_47[156]},
      {stage0_48[51]},
      {stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64], stage0_49[65]},
      {stage1_51[10],stage1_50[17],stage1_49[38],stage1_48[48],stage1_47[56]}
   );
   gpc615_5 gpc574 (
      {stage0_47[157], stage0_47[158], stage0_47[159], stage0_47[160], stage0_47[161]},
      {stage0_48[52]},
      {stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70], stage0_49[71]},
      {stage1_51[11],stage1_50[18],stage1_49[39],stage1_48[49],stage1_47[57]}
   );
   gpc606_5 gpc575 (
      {stage0_48[53], stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57], stage0_48[58]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[12],stage1_50[19],stage1_49[40],stage1_48[50]}
   );
   gpc606_5 gpc576 (
      {stage0_48[59], stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63], stage0_48[64]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[13],stage1_50[20],stage1_49[41],stage1_48[51]}
   );
   gpc606_5 gpc577 (
      {stage0_48[65], stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69], stage0_48[70]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[14],stage1_50[21],stage1_49[42],stage1_48[52]}
   );
   gpc615_5 gpc578 (
      {stage0_48[71], stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75]},
      {stage0_49[72]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[15],stage1_50[22],stage1_49[43],stage1_48[53]}
   );
   gpc615_5 gpc579 (
      {stage0_48[76], stage0_48[77], stage0_48[78], stage0_48[79], stage0_48[80]},
      {stage0_49[73]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[16],stage1_50[23],stage1_49[44],stage1_48[54]}
   );
   gpc615_5 gpc580 (
      {stage0_48[81], stage0_48[82], stage0_48[83], stage0_48[84], stage0_48[85]},
      {stage0_49[74]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[17],stage1_50[24],stage1_49[45],stage1_48[55]}
   );
   gpc615_5 gpc581 (
      {stage0_48[86], stage0_48[87], stage0_48[88], stage0_48[89], stage0_48[90]},
      {stage0_49[75]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[18],stage1_50[25],stage1_49[46],stage1_48[56]}
   );
   gpc615_5 gpc582 (
      {stage0_48[91], stage0_48[92], stage0_48[93], stage0_48[94], stage0_48[95]},
      {stage0_49[76]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[19],stage1_50[26],stage1_49[47],stage1_48[57]}
   );
   gpc615_5 gpc583 (
      {stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99], stage0_48[100]},
      {stage0_49[77]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[20],stage1_50[27],stage1_49[48],stage1_48[58]}
   );
   gpc615_5 gpc584 (
      {stage0_48[101], stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105]},
      {stage0_49[78]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[21],stage1_50[28],stage1_49[49],stage1_48[59]}
   );
   gpc615_5 gpc585 (
      {stage0_48[106], stage0_48[107], stage0_48[108], stage0_48[109], stage0_48[110]},
      {stage0_49[79]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[22],stage1_50[29],stage1_49[50],stage1_48[60]}
   );
   gpc615_5 gpc586 (
      {stage0_48[111], stage0_48[112], stage0_48[113], stage0_48[114], stage0_48[115]},
      {stage0_49[80]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[23],stage1_50[30],stage1_49[51],stage1_48[61]}
   );
   gpc615_5 gpc587 (
      {stage0_48[116], stage0_48[117], stage0_48[118], stage0_48[119], stage0_48[120]},
      {stage0_49[81]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[24],stage1_50[31],stage1_49[52],stage1_48[62]}
   );
   gpc615_5 gpc588 (
      {stage0_48[121], stage0_48[122], stage0_48[123], stage0_48[124], stage0_48[125]},
      {stage0_49[82]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[25],stage1_50[32],stage1_49[53],stage1_48[63]}
   );
   gpc615_5 gpc589 (
      {stage0_48[126], stage0_48[127], stage0_48[128], stage0_48[129], stage0_48[130]},
      {stage0_49[83]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[26],stage1_50[33],stage1_49[54],stage1_48[64]}
   );
   gpc615_5 gpc590 (
      {stage0_48[131], stage0_48[132], stage0_48[133], stage0_48[134], stage0_48[135]},
      {stage0_49[84]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[27],stage1_50[34],stage1_49[55],stage1_48[65]}
   );
   gpc615_5 gpc591 (
      {stage0_48[136], stage0_48[137], stage0_48[138], stage0_48[139], stage0_48[140]},
      {stage0_49[85]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[28],stage1_50[35],stage1_49[56],stage1_48[66]}
   );
   gpc615_5 gpc592 (
      {stage0_48[141], stage0_48[142], stage0_48[143], stage0_48[144], stage0_48[145]},
      {stage0_49[86]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[29],stage1_50[36],stage1_49[57],stage1_48[67]}
   );
   gpc615_5 gpc593 (
      {stage0_48[146], stage0_48[147], stage0_48[148], stage0_48[149], stage0_48[150]},
      {stage0_49[87]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[30],stage1_50[37],stage1_49[58],stage1_48[68]}
   );
   gpc615_5 gpc594 (
      {stage0_48[151], stage0_48[152], stage0_48[153], stage0_48[154], stage0_48[155]},
      {stage0_49[88]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[31],stage1_50[38],stage1_49[59],stage1_48[69]}
   );
   gpc615_5 gpc595 (
      {stage0_48[156], stage0_48[157], stage0_48[158], stage0_48[159], stage0_48[160]},
      {stage0_49[89]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[32],stage1_50[39],stage1_49[60],stage1_48[70]}
   );
   gpc606_5 gpc596 (
      {stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94], stage0_49[95]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[21],stage1_51[33],stage1_50[40],stage1_49[61]}
   );
   gpc606_5 gpc597 (
      {stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100], stage0_49[101]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[22],stage1_51[34],stage1_50[41],stage1_49[62]}
   );
   gpc615_5 gpc598 (
      {stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106]},
      {stage0_50[126]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[23],stage1_51[35],stage1_50[42],stage1_49[63]}
   );
   gpc615_5 gpc599 (
      {stage0_49[107], stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111]},
      {stage0_50[127]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[24],stage1_51[36],stage1_50[43],stage1_49[64]}
   );
   gpc615_5 gpc600 (
      {stage0_49[112], stage0_49[113], stage0_49[114], stage0_49[115], stage0_49[116]},
      {stage0_50[128]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[25],stage1_51[37],stage1_50[44],stage1_49[65]}
   );
   gpc615_5 gpc601 (
      {stage0_49[117], stage0_49[118], stage0_49[119], stage0_49[120], stage0_49[121]},
      {stage0_50[129]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[26],stage1_51[38],stage1_50[45],stage1_49[66]}
   );
   gpc615_5 gpc602 (
      {stage0_49[122], stage0_49[123], stage0_49[124], stage0_49[125], stage0_49[126]},
      {stage0_50[130]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[27],stage1_51[39],stage1_50[46],stage1_49[67]}
   );
   gpc615_5 gpc603 (
      {stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130], stage0_49[131]},
      {stage0_50[131]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[28],stage1_51[40],stage1_50[47],stage1_49[68]}
   );
   gpc615_5 gpc604 (
      {stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136]},
      {stage0_50[132]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[29],stage1_51[41],stage1_50[48],stage1_49[69]}
   );
   gpc615_5 gpc605 (
      {stage0_49[137], stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141]},
      {stage0_50[133]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[30],stage1_51[42],stage1_50[49],stage1_49[70]}
   );
   gpc615_5 gpc606 (
      {stage0_49[142], stage0_49[143], stage0_49[144], stage0_49[145], stage0_49[146]},
      {stage0_50[134]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[31],stage1_51[43],stage1_50[50],stage1_49[71]}
   );
   gpc606_5 gpc607 (
      {stage0_50[135], stage0_50[136], stage0_50[137], stage0_50[138], stage0_50[139], stage0_50[140]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[11],stage1_52[32],stage1_51[44],stage1_50[51]}
   );
   gpc606_5 gpc608 (
      {stage0_50[141], stage0_50[142], stage0_50[143], stage0_50[144], stage0_50[145], stage0_50[146]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[12],stage1_52[33],stage1_51[45],stage1_50[52]}
   );
   gpc606_5 gpc609 (
      {stage0_50[147], stage0_50[148], stage0_50[149], stage0_50[150], stage0_50[151], stage0_50[152]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[13],stage1_52[34],stage1_51[46],stage1_50[53]}
   );
   gpc606_5 gpc610 (
      {stage0_50[153], stage0_50[154], stage0_50[155], stage0_50[156], stage0_50[157], stage0_50[158]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[14],stage1_52[35],stage1_51[47],stage1_50[54]}
   );
   gpc606_5 gpc611 (
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[4],stage1_53[15],stage1_52[36],stage1_51[48]}
   );
   gpc606_5 gpc612 (
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[5],stage1_53[16],stage1_52[37],stage1_51[49]}
   );
   gpc606_5 gpc613 (
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[6],stage1_53[17],stage1_52[38],stage1_51[50]}
   );
   gpc606_5 gpc614 (
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[7],stage1_53[18],stage1_52[39],stage1_51[51]}
   );
   gpc606_5 gpc615 (
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[8],stage1_53[19],stage1_52[40],stage1_51[52]}
   );
   gpc606_5 gpc616 (
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[9],stage1_53[20],stage1_52[41],stage1_51[53]}
   );
   gpc606_5 gpc617 (
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[10],stage1_53[21],stage1_52[42],stage1_51[54]}
   );
   gpc606_5 gpc618 (
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[11],stage1_53[22],stage1_52[43],stage1_51[55]}
   );
   gpc606_5 gpc619 (
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[12],stage1_53[23],stage1_52[44],stage1_51[56]}
   );
   gpc606_5 gpc620 (
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[13],stage1_53[24],stage1_52[45],stage1_51[57]}
   );
   gpc606_5 gpc621 (
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[10],stage1_54[14],stage1_53[25],stage1_52[46]}
   );
   gpc606_5 gpc622 (
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[11],stage1_54[15],stage1_53[26],stage1_52[47]}
   );
   gpc606_5 gpc623 (
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[12],stage1_54[16],stage1_53[27],stage1_52[48]}
   );
   gpc606_5 gpc624 (
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[13],stage1_54[17],stage1_53[28],stage1_52[49]}
   );
   gpc606_5 gpc625 (
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[14],stage1_54[18],stage1_53[29],stage1_52[50]}
   );
   gpc606_5 gpc626 (
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[15],stage1_54[19],stage1_53[30],stage1_52[51]}
   );
   gpc606_5 gpc627 (
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[16],stage1_54[20],stage1_53[31],stage1_52[52]}
   );
   gpc606_5 gpc628 (
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[17],stage1_54[21],stage1_53[32],stage1_52[53]}
   );
   gpc606_5 gpc629 (
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[18],stage1_54[22],stage1_53[33],stage1_52[54]}
   );
   gpc606_5 gpc630 (
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[19],stage1_54[23],stage1_53[34],stage1_52[55]}
   );
   gpc606_5 gpc631 (
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[20],stage1_54[24],stage1_53[35],stage1_52[56]}
   );
   gpc606_5 gpc632 (
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[21],stage1_54[25],stage1_53[36],stage1_52[57]}
   );
   gpc606_5 gpc633 (
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[22],stage1_54[26],stage1_53[37],stage1_52[58]}
   );
   gpc606_5 gpc634 (
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[23],stage1_54[27],stage1_53[38],stage1_52[59]}
   );
   gpc606_5 gpc635 (
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[24],stage1_54[28],stage1_53[39],stage1_52[60]}
   );
   gpc606_5 gpc636 (
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[25],stage1_54[29],stage1_53[40],stage1_52[61]}
   );
   gpc606_5 gpc637 (
      {stage0_52[120], stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[26],stage1_54[30],stage1_53[41],stage1_52[62]}
   );
   gpc606_5 gpc638 (
      {stage0_52[126], stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[27],stage1_54[31],stage1_53[42],stage1_52[63]}
   );
   gpc606_5 gpc639 (
      {stage0_52[132], stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[28],stage1_54[32],stage1_53[43],stage1_52[64]}
   );
   gpc615_5 gpc640 (
      {stage0_52[138], stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142]},
      {stage0_53[60]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[29],stage1_54[33],stage1_53[44],stage1_52[65]}
   );
   gpc615_5 gpc641 (
      {stage0_52[143], stage0_52[144], stage0_52[145], stage0_52[146], stage0_52[147]},
      {stage0_53[61]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[30],stage1_54[34],stage1_53[45],stage1_52[66]}
   );
   gpc615_5 gpc642 (
      {stage0_52[148], stage0_52[149], stage0_52[150], stage0_52[151], stage0_52[152]},
      {stage0_53[62]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[31],stage1_54[35],stage1_53[46],stage1_52[67]}
   );
   gpc606_5 gpc643 (
      {stage0_53[63], stage0_53[64], stage0_53[65], stage0_53[66], stage0_53[67], stage0_53[68]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[22],stage1_55[32],stage1_54[36],stage1_53[47]}
   );
   gpc606_5 gpc644 (
      {stage0_53[69], stage0_53[70], stage0_53[71], stage0_53[72], stage0_53[73], stage0_53[74]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[23],stage1_55[33],stage1_54[37],stage1_53[48]}
   );
   gpc606_5 gpc645 (
      {stage0_53[75], stage0_53[76], stage0_53[77], stage0_53[78], stage0_53[79], stage0_53[80]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[24],stage1_55[34],stage1_54[38],stage1_53[49]}
   );
   gpc606_5 gpc646 (
      {stage0_53[81], stage0_53[82], stage0_53[83], stage0_53[84], stage0_53[85], stage0_53[86]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[25],stage1_55[35],stage1_54[39],stage1_53[50]}
   );
   gpc606_5 gpc647 (
      {stage0_53[87], stage0_53[88], stage0_53[89], stage0_53[90], stage0_53[91], stage0_53[92]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[26],stage1_55[36],stage1_54[40],stage1_53[51]}
   );
   gpc606_5 gpc648 (
      {stage0_53[93], stage0_53[94], stage0_53[95], stage0_53[96], stage0_53[97], stage0_53[98]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[27],stage1_55[37],stage1_54[41],stage1_53[52]}
   );
   gpc606_5 gpc649 (
      {stage0_53[99], stage0_53[100], stage0_53[101], stage0_53[102], stage0_53[103], stage0_53[104]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[28],stage1_55[38],stage1_54[42],stage1_53[53]}
   );
   gpc606_5 gpc650 (
      {stage0_53[105], stage0_53[106], stage0_53[107], stage0_53[108], stage0_53[109], stage0_53[110]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[29],stage1_55[39],stage1_54[43],stage1_53[54]}
   );
   gpc606_5 gpc651 (
      {stage0_53[111], stage0_53[112], stage0_53[113], stage0_53[114], stage0_53[115], stage0_53[116]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[30],stage1_55[40],stage1_54[44],stage1_53[55]}
   );
   gpc606_5 gpc652 (
      {stage0_53[117], stage0_53[118], stage0_53[119], stage0_53[120], stage0_53[121], stage0_53[122]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[31],stage1_55[41],stage1_54[45],stage1_53[56]}
   );
   gpc606_5 gpc653 (
      {stage0_53[123], stage0_53[124], stage0_53[125], stage0_53[126], stage0_53[127], stage0_53[128]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[32],stage1_55[42],stage1_54[46],stage1_53[57]}
   );
   gpc606_5 gpc654 (
      {stage0_53[129], stage0_53[130], stage0_53[131], stage0_53[132], stage0_53[133], stage0_53[134]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[33],stage1_55[43],stage1_54[47],stage1_53[58]}
   );
   gpc606_5 gpc655 (
      {stage0_53[135], stage0_53[136], stage0_53[137], stage0_53[138], stage0_53[139], stage0_53[140]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[34],stage1_55[44],stage1_54[48],stage1_53[59]}
   );
   gpc606_5 gpc656 (
      {stage0_53[141], stage0_53[142], stage0_53[143], stage0_53[144], stage0_53[145], stage0_53[146]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[35],stage1_55[45],stage1_54[49],stage1_53[60]}
   );
   gpc606_5 gpc657 (
      {stage0_53[147], stage0_53[148], stage0_53[149], stage0_53[150], stage0_53[151], stage0_53[152]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[36],stage1_55[46],stage1_54[50],stage1_53[61]}
   );
   gpc606_5 gpc658 (
      {stage0_53[153], stage0_53[154], stage0_53[155], stage0_53[156], stage0_53[157], stage0_53[158]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[37],stage1_55[47],stage1_54[51],stage1_53[62]}
   );
   gpc615_5 gpc659 (
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136]},
      {stage0_55[96]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[16],stage1_56[38],stage1_55[48],stage1_54[52]}
   );
   gpc615_5 gpc660 (
      {stage0_54[137], stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141]},
      {stage0_55[97]},
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage1_58[1],stage1_57[17],stage1_56[39],stage1_55[49],stage1_54[53]}
   );
   gpc615_5 gpc661 (
      {stage0_54[142], stage0_54[143], stage0_54[144], stage0_54[145], stage0_54[146]},
      {stage0_55[98]},
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage1_58[2],stage1_57[18],stage1_56[40],stage1_55[50],stage1_54[54]}
   );
   gpc615_5 gpc662 (
      {stage0_54[147], stage0_54[148], stage0_54[149], stage0_54[150], stage0_54[151]},
      {stage0_55[99]},
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage1_58[3],stage1_57[19],stage1_56[41],stage1_55[51],stage1_54[55]}
   );
   gpc615_5 gpc663 (
      {stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155], stage0_54[156]},
      {stage0_55[100]},
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage1_58[4],stage1_57[20],stage1_56[42],stage1_55[52],stage1_54[56]}
   );
   gpc615_5 gpc664 (
      {stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage0_55[101]},
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage1_58[5],stage1_57[21],stage1_56[43],stage1_55[53],stage1_54[57]}
   );
   gpc615_5 gpc665 (
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106]},
      {stage0_56[36]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[6],stage1_57[22],stage1_56[44],stage1_55[54]}
   );
   gpc615_5 gpc666 (
      {stage0_55[107], stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111]},
      {stage0_56[37]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[7],stage1_57[23],stage1_56[45],stage1_55[55]}
   );
   gpc615_5 gpc667 (
      {stage0_55[112], stage0_55[113], stage0_55[114], stage0_55[115], stage0_55[116]},
      {stage0_56[38]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[8],stage1_57[24],stage1_56[46],stage1_55[56]}
   );
   gpc615_5 gpc668 (
      {stage0_55[117], stage0_55[118], stage0_55[119], stage0_55[120], stage0_55[121]},
      {stage0_56[39]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[9],stage1_57[25],stage1_56[47],stage1_55[57]}
   );
   gpc606_5 gpc669 (
      {stage0_56[40], stage0_56[41], stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[4],stage1_58[10],stage1_57[26],stage1_56[48]}
   );
   gpc606_5 gpc670 (
      {stage0_56[46], stage0_56[47], stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[5],stage1_58[11],stage1_57[27],stage1_56[49]}
   );
   gpc606_5 gpc671 (
      {stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55], stage0_56[56], stage0_56[57]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[6],stage1_58[12],stage1_57[28],stage1_56[50]}
   );
   gpc606_5 gpc672 (
      {stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61], stage0_56[62], stage0_56[63]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[7],stage1_58[13],stage1_57[29],stage1_56[51]}
   );
   gpc606_5 gpc673 (
      {stage0_56[64], stage0_56[65], stage0_56[66], stage0_56[67], stage0_56[68], stage0_56[69]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[8],stage1_58[14],stage1_57[30],stage1_56[52]}
   );
   gpc606_5 gpc674 (
      {stage0_56[70], stage0_56[71], stage0_56[72], stage0_56[73], stage0_56[74], stage0_56[75]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[9],stage1_58[15],stage1_57[31],stage1_56[53]}
   );
   gpc606_5 gpc675 (
      {stage0_56[76], stage0_56[77], stage0_56[78], stage0_56[79], stage0_56[80], stage0_56[81]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[10],stage1_58[16],stage1_57[32],stage1_56[54]}
   );
   gpc606_5 gpc676 (
      {stage0_56[82], stage0_56[83], stage0_56[84], stage0_56[85], stage0_56[86], stage0_56[87]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[11],stage1_58[17],stage1_57[33],stage1_56[55]}
   );
   gpc606_5 gpc677 (
      {stage0_56[88], stage0_56[89], stage0_56[90], stage0_56[91], stage0_56[92], stage0_56[93]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[12],stage1_58[18],stage1_57[34],stage1_56[56]}
   );
   gpc606_5 gpc678 (
      {stage0_56[94], stage0_56[95], stage0_56[96], stage0_56[97], stage0_56[98], stage0_56[99]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[13],stage1_58[19],stage1_57[35],stage1_56[57]}
   );
   gpc606_5 gpc679 (
      {stage0_56[100], stage0_56[101], stage0_56[102], stage0_56[103], stage0_56[104], stage0_56[105]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[14],stage1_58[20],stage1_57[36],stage1_56[58]}
   );
   gpc606_5 gpc680 (
      {stage0_56[106], stage0_56[107], stage0_56[108], stage0_56[109], stage0_56[110], stage0_56[111]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[15],stage1_58[21],stage1_57[37],stage1_56[59]}
   );
   gpc606_5 gpc681 (
      {stage0_56[112], stage0_56[113], stage0_56[114], stage0_56[115], stage0_56[116], stage0_56[117]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[16],stage1_58[22],stage1_57[38],stage1_56[60]}
   );
   gpc606_5 gpc682 (
      {stage0_56[118], stage0_56[119], stage0_56[120], stage0_56[121], stage0_56[122], stage0_56[123]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[17],stage1_58[23],stage1_57[39],stage1_56[61]}
   );
   gpc606_5 gpc683 (
      {stage0_56[124], stage0_56[125], stage0_56[126], stage0_56[127], stage0_56[128], stage0_56[129]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[18],stage1_58[24],stage1_57[40],stage1_56[62]}
   );
   gpc606_5 gpc684 (
      {stage0_56[130], stage0_56[131], stage0_56[132], stage0_56[133], stage0_56[134], stage0_56[135]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[19],stage1_58[25],stage1_57[41],stage1_56[63]}
   );
   gpc606_5 gpc685 (
      {stage0_56[136], stage0_56[137], stage0_56[138], stage0_56[139], stage0_56[140], stage0_56[141]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[20],stage1_58[26],stage1_57[42],stage1_56[64]}
   );
   gpc606_5 gpc686 (
      {stage0_56[142], stage0_56[143], stage0_56[144], stage0_56[145], stage0_56[146], stage0_56[147]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[21],stage1_58[27],stage1_57[43],stage1_56[65]}
   );
   gpc606_5 gpc687 (
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[18],stage1_59[22],stage1_58[28],stage1_57[44]}
   );
   gpc606_5 gpc688 (
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[19],stage1_59[23],stage1_58[29],stage1_57[45]}
   );
   gpc606_5 gpc689 (
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[20],stage1_59[24],stage1_58[30],stage1_57[46]}
   );
   gpc606_5 gpc690 (
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[21],stage1_59[25],stage1_58[31],stage1_57[47]}
   );
   gpc606_5 gpc691 (
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[22],stage1_59[26],stage1_58[32],stage1_57[48]}
   );
   gpc606_5 gpc692 (
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[23],stage1_59[27],stage1_58[33],stage1_57[49]}
   );
   gpc606_5 gpc693 (
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[24],stage1_59[28],stage1_58[34],stage1_57[50]}
   );
   gpc606_5 gpc694 (
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[25],stage1_59[29],stage1_58[35],stage1_57[51]}
   );
   gpc606_5 gpc695 (
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[26],stage1_59[30],stage1_58[36],stage1_57[52]}
   );
   gpc606_5 gpc696 (
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[27],stage1_59[31],stage1_58[37],stage1_57[53]}
   );
   gpc606_5 gpc697 (
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[28],stage1_59[32],stage1_58[38],stage1_57[54]}
   );
   gpc606_5 gpc698 (
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[29],stage1_59[33],stage1_58[39],stage1_57[55]}
   );
   gpc606_5 gpc699 (
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[30],stage1_59[34],stage1_58[40],stage1_57[56]}
   );
   gpc606_5 gpc700 (
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[31],stage1_59[35],stage1_58[41],stage1_57[57]}
   );
   gpc606_5 gpc701 (
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[32],stage1_59[36],stage1_58[42],stage1_57[58]}
   );
   gpc606_5 gpc702 (
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[33],stage1_59[37],stage1_58[43],stage1_57[59]}
   );
   gpc606_5 gpc703 (
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[34],stage1_59[38],stage1_58[44],stage1_57[60]}
   );
   gpc606_5 gpc704 (
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[35],stage1_59[39],stage1_58[45],stage1_57[61]}
   );
   gpc606_5 gpc705 (
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[36],stage1_59[40],stage1_58[46],stage1_57[62]}
   );
   gpc606_5 gpc706 (
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[37],stage1_59[41],stage1_58[47],stage1_57[63]}
   );
   gpc606_5 gpc707 (
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[38],stage1_59[42],stage1_58[48],stage1_57[64]}
   );
   gpc606_5 gpc708 (
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[39],stage1_59[43],stage1_58[49],stage1_57[65]}
   );
   gpc606_5 gpc709 (
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[22],stage1_60[40],stage1_59[44],stage1_58[50]}
   );
   gpc606_5 gpc710 (
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[23],stage1_60[41],stage1_59[45],stage1_58[51]}
   );
   gpc606_5 gpc711 (
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[24],stage1_60[42],stage1_59[46],stage1_58[52]}
   );
   gpc606_5 gpc712 (
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[25],stage1_60[43],stage1_59[47],stage1_58[53]}
   );
   gpc606_5 gpc713 (
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[26],stage1_60[44],stage1_59[48],stage1_58[54]}
   );
   gpc606_5 gpc714 (
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[27],stage1_60[45],stage1_59[49],stage1_58[55]}
   );
   gpc606_5 gpc715 (
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[0],stage1_62[6],stage1_61[28],stage1_60[46]}
   );
   gpc606_5 gpc716 (
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[1],stage1_62[7],stage1_61[29],stage1_60[47]}
   );
   gpc606_5 gpc717 (
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[2],stage1_62[8],stage1_61[30],stage1_60[48]}
   );
   gpc606_5 gpc718 (
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[3],stage1_62[9],stage1_61[31],stage1_60[49]}
   );
   gpc606_5 gpc719 (
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[4],stage1_62[10],stage1_61[32],stage1_60[50]}
   );
   gpc606_5 gpc720 (
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[5],stage1_62[11],stage1_61[33],stage1_60[51]}
   );
   gpc606_5 gpc721 (
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[6],stage1_62[12],stage1_61[34],stage1_60[52]}
   );
   gpc606_5 gpc722 (
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[7],stage1_62[13],stage1_61[35],stage1_60[53]}
   );
   gpc606_5 gpc723 (
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[8],stage1_62[14],stage1_61[36],stage1_60[54]}
   );
   gpc606_5 gpc724 (
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[9],stage1_62[15],stage1_61[37],stage1_60[55]}
   );
   gpc606_5 gpc725 (
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[10],stage1_62[16],stage1_61[38],stage1_60[56]}
   );
   gpc606_5 gpc726 (
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[11],stage1_62[17],stage1_61[39],stage1_60[57]}
   );
   gpc606_5 gpc727 (
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage0_62[72], stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77]},
      {stage1_64[12],stage1_63[12],stage1_62[18],stage1_61[40],stage1_60[58]}
   );
   gpc606_5 gpc728 (
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage0_62[78], stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83]},
      {stage1_64[13],stage1_63[13],stage1_62[19],stage1_61[41],stage1_60[59]}
   );
   gpc606_5 gpc729 (
      {stage0_60[120], stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125]},
      {stage0_62[84], stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89]},
      {stage1_64[14],stage1_63[14],stage1_62[20],stage1_61[42],stage1_60[60]}
   );
   gpc606_5 gpc730 (
      {stage0_60[126], stage0_60[127], stage0_60[128], stage0_60[129], stage0_60[130], stage0_60[131]},
      {stage0_62[90], stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95]},
      {stage1_64[15],stage1_63[15],stage1_62[21],stage1_61[43],stage1_60[61]}
   );
   gpc606_5 gpc731 (
      {stage0_60[132], stage0_60[133], stage0_60[134], stage0_60[135], stage0_60[136], stage0_60[137]},
      {stage0_62[96], stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101]},
      {stage1_64[16],stage1_63[16],stage1_62[22],stage1_61[44],stage1_60[62]}
   );
   gpc606_5 gpc732 (
      {stage0_60[138], stage0_60[139], stage0_60[140], stage0_60[141], stage0_60[142], stage0_60[143]},
      {stage0_62[102], stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107]},
      {stage1_64[17],stage1_63[17],stage1_62[23],stage1_61[45],stage1_60[63]}
   );
   gpc606_5 gpc733 (
      {stage0_60[144], stage0_60[145], stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149]},
      {stage0_62[108], stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113]},
      {stage1_64[18],stage1_63[18],stage1_62[24],stage1_61[46],stage1_60[64]}
   );
   gpc606_5 gpc734 (
      {stage0_60[150], stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155]},
      {stage0_62[114], stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119]},
      {stage1_64[19],stage1_63[19],stage1_62[25],stage1_61[47],stage1_60[65]}
   );
   gpc606_5 gpc735 (
      {stage0_60[156], stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160], stage0_60[161]},
      {stage0_62[120], stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125]},
      {stage1_64[20],stage1_63[20],stage1_62[26],stage1_61[48],stage1_60[66]}
   );
   gpc606_5 gpc736 (
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[21],stage1_63[21],stage1_62[27],stage1_61[49]}
   );
   gpc606_5 gpc737 (
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[22],stage1_63[22],stage1_62[28],stage1_61[50]}
   );
   gpc606_5 gpc738 (
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[23],stage1_63[23],stage1_62[29],stage1_61[51]}
   );
   gpc606_5 gpc739 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22], stage0_61[23]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[24],stage1_63[24],stage1_62[30],stage1_61[52]}
   );
   gpc606_5 gpc740 (
      {stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27], stage0_61[28], stage0_61[29]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[25],stage1_63[25],stage1_62[31],stage1_61[53]}
   );
   gpc606_5 gpc741 (
      {stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33], stage0_61[34], stage0_61[35]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[26],stage1_63[26],stage1_62[32],stage1_61[54]}
   );
   gpc606_5 gpc742 (
      {stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[27],stage1_63[27],stage1_62[33],stage1_61[55]}
   );
   gpc606_5 gpc743 (
      {stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[28],stage1_63[28],stage1_62[34],stage1_61[56]}
   );
   gpc606_5 gpc744 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52], stage0_61[53]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[29],stage1_63[29],stage1_62[35],stage1_61[57]}
   );
   gpc606_5 gpc745 (
      {stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57], stage0_61[58], stage0_61[59]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[30],stage1_63[30],stage1_62[36],stage1_61[58]}
   );
   gpc606_5 gpc746 (
      {stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63], stage0_61[64], stage0_61[65]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[31],stage1_63[31],stage1_62[37],stage1_61[59]}
   );
   gpc606_5 gpc747 (
      {stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69], stage0_61[70], stage0_61[71]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[32],stage1_63[32],stage1_62[38],stage1_61[60]}
   );
   gpc606_5 gpc748 (
      {stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75], stage0_61[76], stage0_61[77]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[33],stage1_63[33],stage1_62[39],stage1_61[61]}
   );
   gpc606_5 gpc749 (
      {stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81], stage0_61[82], stage0_61[83]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[34],stage1_63[34],stage1_62[40],stage1_61[62]}
   );
   gpc606_5 gpc750 (
      {stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87], stage0_61[88], stage0_61[89]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[35],stage1_63[35],stage1_62[41],stage1_61[63]}
   );
   gpc606_5 gpc751 (
      {stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93], stage0_61[94], stage0_61[95]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[36],stage1_63[36],stage1_62[42],stage1_61[64]}
   );
   gpc606_5 gpc752 (
      {stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99], stage0_61[100], stage0_61[101]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[37],stage1_63[37],stage1_62[43],stage1_61[65]}
   );
   gpc606_5 gpc753 (
      {stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105], stage0_61[106], stage0_61[107]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[38],stage1_63[38],stage1_62[44],stage1_61[66]}
   );
   gpc606_5 gpc754 (
      {stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111], stage0_61[112], stage0_61[113]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[39],stage1_63[39],stage1_62[45],stage1_61[67]}
   );
   gpc606_5 gpc755 (
      {stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117], stage0_61[118], stage0_61[119]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[40],stage1_63[40],stage1_62[46],stage1_61[68]}
   );
   gpc606_5 gpc756 (
      {stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123], stage0_61[124], stage0_61[125]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[41],stage1_63[41],stage1_62[47],stage1_61[69]}
   );
   gpc606_5 gpc757 (
      {stage0_61[126], stage0_61[127], stage0_61[128], stage0_61[129], stage0_61[130], stage0_61[131]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[42],stage1_63[42],stage1_62[48],stage1_61[70]}
   );
   gpc606_5 gpc758 (
      {stage0_61[132], stage0_61[133], stage0_61[134], stage0_61[135], stage0_61[136], stage0_61[137]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[43],stage1_63[43],stage1_62[49],stage1_61[71]}
   );
   gpc606_5 gpc759 (
      {stage0_61[138], stage0_61[139], stage0_61[140], stage0_61[141], stage0_61[142], stage0_61[143]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[44],stage1_63[44],stage1_62[50],stage1_61[72]}
   );
   gpc1_1 gpc760 (
      {stage0_2[160]},
      {stage1_2[53]}
   );
   gpc1_1 gpc761 (
      {stage0_2[161]},
      {stage1_2[54]}
   );
   gpc1_1 gpc762 (
      {stage0_3[139]},
      {stage1_3[61]}
   );
   gpc1_1 gpc763 (
      {stage0_3[140]},
      {stage1_3[62]}
   );
   gpc1_1 gpc764 (
      {stage0_3[141]},
      {stage1_3[63]}
   );
   gpc1_1 gpc765 (
      {stage0_3[142]},
      {stage1_3[64]}
   );
   gpc1_1 gpc766 (
      {stage0_3[143]},
      {stage1_3[65]}
   );
   gpc1_1 gpc767 (
      {stage0_3[144]},
      {stage1_3[66]}
   );
   gpc1_1 gpc768 (
      {stage0_3[145]},
      {stage1_3[67]}
   );
   gpc1_1 gpc769 (
      {stage0_3[146]},
      {stage1_3[68]}
   );
   gpc1_1 gpc770 (
      {stage0_3[147]},
      {stage1_3[69]}
   );
   gpc1_1 gpc771 (
      {stage0_3[148]},
      {stage1_3[70]}
   );
   gpc1_1 gpc772 (
      {stage0_3[149]},
      {stage1_3[71]}
   );
   gpc1_1 gpc773 (
      {stage0_3[150]},
      {stage1_3[72]}
   );
   gpc1_1 gpc774 (
      {stage0_3[151]},
      {stage1_3[73]}
   );
   gpc1_1 gpc775 (
      {stage0_3[152]},
      {stage1_3[74]}
   );
   gpc1_1 gpc776 (
      {stage0_3[153]},
      {stage1_3[75]}
   );
   gpc1_1 gpc777 (
      {stage0_3[154]},
      {stage1_3[76]}
   );
   gpc1_1 gpc778 (
      {stage0_3[155]},
      {stage1_3[77]}
   );
   gpc1_1 gpc779 (
      {stage0_3[156]},
      {stage1_3[78]}
   );
   gpc1_1 gpc780 (
      {stage0_3[157]},
      {stage1_3[79]}
   );
   gpc1_1 gpc781 (
      {stage0_3[158]},
      {stage1_3[80]}
   );
   gpc1_1 gpc782 (
      {stage0_3[159]},
      {stage1_3[81]}
   );
   gpc1_1 gpc783 (
      {stage0_3[160]},
      {stage1_3[82]}
   );
   gpc1_1 gpc784 (
      {stage0_3[161]},
      {stage1_3[83]}
   );
   gpc1_1 gpc785 (
      {stage0_4[158]},
      {stage1_4[79]}
   );
   gpc1_1 gpc786 (
      {stage0_4[159]},
      {stage1_4[80]}
   );
   gpc1_1 gpc787 (
      {stage0_4[160]},
      {stage1_4[81]}
   );
   gpc1_1 gpc788 (
      {stage0_4[161]},
      {stage1_4[82]}
   );
   gpc1_1 gpc789 (
      {stage0_5[102]},
      {stage1_5[55]}
   );
   gpc1_1 gpc790 (
      {stage0_5[103]},
      {stage1_5[56]}
   );
   gpc1_1 gpc791 (
      {stage0_5[104]},
      {stage1_5[57]}
   );
   gpc1_1 gpc792 (
      {stage0_5[105]},
      {stage1_5[58]}
   );
   gpc1_1 gpc793 (
      {stage0_5[106]},
      {stage1_5[59]}
   );
   gpc1_1 gpc794 (
      {stage0_5[107]},
      {stage1_5[60]}
   );
   gpc1_1 gpc795 (
      {stage0_5[108]},
      {stage1_5[61]}
   );
   gpc1_1 gpc796 (
      {stage0_5[109]},
      {stage1_5[62]}
   );
   gpc1_1 gpc797 (
      {stage0_5[110]},
      {stage1_5[63]}
   );
   gpc1_1 gpc798 (
      {stage0_5[111]},
      {stage1_5[64]}
   );
   gpc1_1 gpc799 (
      {stage0_5[112]},
      {stage1_5[65]}
   );
   gpc1_1 gpc800 (
      {stage0_5[113]},
      {stage1_5[66]}
   );
   gpc1_1 gpc801 (
      {stage0_5[114]},
      {stage1_5[67]}
   );
   gpc1_1 gpc802 (
      {stage0_5[115]},
      {stage1_5[68]}
   );
   gpc1_1 gpc803 (
      {stage0_5[116]},
      {stage1_5[69]}
   );
   gpc1_1 gpc804 (
      {stage0_5[117]},
      {stage1_5[70]}
   );
   gpc1_1 gpc805 (
      {stage0_5[118]},
      {stage1_5[71]}
   );
   gpc1_1 gpc806 (
      {stage0_5[119]},
      {stage1_5[72]}
   );
   gpc1_1 gpc807 (
      {stage0_5[120]},
      {stage1_5[73]}
   );
   gpc1_1 gpc808 (
      {stage0_5[121]},
      {stage1_5[74]}
   );
   gpc1_1 gpc809 (
      {stage0_5[122]},
      {stage1_5[75]}
   );
   gpc1_1 gpc810 (
      {stage0_5[123]},
      {stage1_5[76]}
   );
   gpc1_1 gpc811 (
      {stage0_5[124]},
      {stage1_5[77]}
   );
   gpc1_1 gpc812 (
      {stage0_5[125]},
      {stage1_5[78]}
   );
   gpc1_1 gpc813 (
      {stage0_5[126]},
      {stage1_5[79]}
   );
   gpc1_1 gpc814 (
      {stage0_5[127]},
      {stage1_5[80]}
   );
   gpc1_1 gpc815 (
      {stage0_5[128]},
      {stage1_5[81]}
   );
   gpc1_1 gpc816 (
      {stage0_5[129]},
      {stage1_5[82]}
   );
   gpc1_1 gpc817 (
      {stage0_5[130]},
      {stage1_5[83]}
   );
   gpc1_1 gpc818 (
      {stage0_5[131]},
      {stage1_5[84]}
   );
   gpc1_1 gpc819 (
      {stage0_5[132]},
      {stage1_5[85]}
   );
   gpc1_1 gpc820 (
      {stage0_5[133]},
      {stage1_5[86]}
   );
   gpc1_1 gpc821 (
      {stage0_5[134]},
      {stage1_5[87]}
   );
   gpc1_1 gpc822 (
      {stage0_5[135]},
      {stage1_5[88]}
   );
   gpc1_1 gpc823 (
      {stage0_5[136]},
      {stage1_5[89]}
   );
   gpc1_1 gpc824 (
      {stage0_5[137]},
      {stage1_5[90]}
   );
   gpc1_1 gpc825 (
      {stage0_5[138]},
      {stage1_5[91]}
   );
   gpc1_1 gpc826 (
      {stage0_5[139]},
      {stage1_5[92]}
   );
   gpc1_1 gpc827 (
      {stage0_5[140]},
      {stage1_5[93]}
   );
   gpc1_1 gpc828 (
      {stage0_5[141]},
      {stage1_5[94]}
   );
   gpc1_1 gpc829 (
      {stage0_5[142]},
      {stage1_5[95]}
   );
   gpc1_1 gpc830 (
      {stage0_5[143]},
      {stage1_5[96]}
   );
   gpc1_1 gpc831 (
      {stage0_5[144]},
      {stage1_5[97]}
   );
   gpc1_1 gpc832 (
      {stage0_5[145]},
      {stage1_5[98]}
   );
   gpc1_1 gpc833 (
      {stage0_5[146]},
      {stage1_5[99]}
   );
   gpc1_1 gpc834 (
      {stage0_5[147]},
      {stage1_5[100]}
   );
   gpc1_1 gpc835 (
      {stage0_5[148]},
      {stage1_5[101]}
   );
   gpc1_1 gpc836 (
      {stage0_5[149]},
      {stage1_5[102]}
   );
   gpc1_1 gpc837 (
      {stage0_5[150]},
      {stage1_5[103]}
   );
   gpc1_1 gpc838 (
      {stage0_5[151]},
      {stage1_5[104]}
   );
   gpc1_1 gpc839 (
      {stage0_5[152]},
      {stage1_5[105]}
   );
   gpc1_1 gpc840 (
      {stage0_5[153]},
      {stage1_5[106]}
   );
   gpc1_1 gpc841 (
      {stage0_5[154]},
      {stage1_5[107]}
   );
   gpc1_1 gpc842 (
      {stage0_5[155]},
      {stage1_5[108]}
   );
   gpc1_1 gpc843 (
      {stage0_5[156]},
      {stage1_5[109]}
   );
   gpc1_1 gpc844 (
      {stage0_5[157]},
      {stage1_5[110]}
   );
   gpc1_1 gpc845 (
      {stage0_5[158]},
      {stage1_5[111]}
   );
   gpc1_1 gpc846 (
      {stage0_5[159]},
      {stage1_5[112]}
   );
   gpc1_1 gpc847 (
      {stage0_5[160]},
      {stage1_5[113]}
   );
   gpc1_1 gpc848 (
      {stage0_5[161]},
      {stage1_5[114]}
   );
   gpc1_1 gpc849 (
      {stage0_6[154]},
      {stage1_6[50]}
   );
   gpc1_1 gpc850 (
      {stage0_6[155]},
      {stage1_6[51]}
   );
   gpc1_1 gpc851 (
      {stage0_6[156]},
      {stage1_6[52]}
   );
   gpc1_1 gpc852 (
      {stage0_6[157]},
      {stage1_6[53]}
   );
   gpc1_1 gpc853 (
      {stage0_6[158]},
      {stage1_6[54]}
   );
   gpc1_1 gpc854 (
      {stage0_6[159]},
      {stage1_6[55]}
   );
   gpc1_1 gpc855 (
      {stage0_6[160]},
      {stage1_6[56]}
   );
   gpc1_1 gpc856 (
      {stage0_6[161]},
      {stage1_6[57]}
   );
   gpc1_1 gpc857 (
      {stage0_7[153]},
      {stage1_7[62]}
   );
   gpc1_1 gpc858 (
      {stage0_7[154]},
      {stage1_7[63]}
   );
   gpc1_1 gpc859 (
      {stage0_7[155]},
      {stage1_7[64]}
   );
   gpc1_1 gpc860 (
      {stage0_7[156]},
      {stage1_7[65]}
   );
   gpc1_1 gpc861 (
      {stage0_7[157]},
      {stage1_7[66]}
   );
   gpc1_1 gpc862 (
      {stage0_7[158]},
      {stage1_7[67]}
   );
   gpc1_1 gpc863 (
      {stage0_7[159]},
      {stage1_7[68]}
   );
   gpc1_1 gpc864 (
      {stage0_7[160]},
      {stage1_7[69]}
   );
   gpc1_1 gpc865 (
      {stage0_7[161]},
      {stage1_7[70]}
   );
   gpc1_1 gpc866 (
      {stage0_8[149]},
      {stage1_8[68]}
   );
   gpc1_1 gpc867 (
      {stage0_8[150]},
      {stage1_8[69]}
   );
   gpc1_1 gpc868 (
      {stage0_8[151]},
      {stage1_8[70]}
   );
   gpc1_1 gpc869 (
      {stage0_8[152]},
      {stage1_8[71]}
   );
   gpc1_1 gpc870 (
      {stage0_8[153]},
      {stage1_8[72]}
   );
   gpc1_1 gpc871 (
      {stage0_8[154]},
      {stage1_8[73]}
   );
   gpc1_1 gpc872 (
      {stage0_8[155]},
      {stage1_8[74]}
   );
   gpc1_1 gpc873 (
      {stage0_8[156]},
      {stage1_8[75]}
   );
   gpc1_1 gpc874 (
      {stage0_8[157]},
      {stage1_8[76]}
   );
   gpc1_1 gpc875 (
      {stage0_8[158]},
      {stage1_8[77]}
   );
   gpc1_1 gpc876 (
      {stage0_8[159]},
      {stage1_8[78]}
   );
   gpc1_1 gpc877 (
      {stage0_8[160]},
      {stage1_8[79]}
   );
   gpc1_1 gpc878 (
      {stage0_8[161]},
      {stage1_8[80]}
   );
   gpc1_1 gpc879 (
      {stage0_10[124]},
      {stage1_10[57]}
   );
   gpc1_1 gpc880 (
      {stage0_10[125]},
      {stage1_10[58]}
   );
   gpc1_1 gpc881 (
      {stage0_10[126]},
      {stage1_10[59]}
   );
   gpc1_1 gpc882 (
      {stage0_10[127]},
      {stage1_10[60]}
   );
   gpc1_1 gpc883 (
      {stage0_10[128]},
      {stage1_10[61]}
   );
   gpc1_1 gpc884 (
      {stage0_10[129]},
      {stage1_10[62]}
   );
   gpc1_1 gpc885 (
      {stage0_10[130]},
      {stage1_10[63]}
   );
   gpc1_1 gpc886 (
      {stage0_10[131]},
      {stage1_10[64]}
   );
   gpc1_1 gpc887 (
      {stage0_10[132]},
      {stage1_10[65]}
   );
   gpc1_1 gpc888 (
      {stage0_10[133]},
      {stage1_10[66]}
   );
   gpc1_1 gpc889 (
      {stage0_10[134]},
      {stage1_10[67]}
   );
   gpc1_1 gpc890 (
      {stage0_10[135]},
      {stage1_10[68]}
   );
   gpc1_1 gpc891 (
      {stage0_10[136]},
      {stage1_10[69]}
   );
   gpc1_1 gpc892 (
      {stage0_10[137]},
      {stage1_10[70]}
   );
   gpc1_1 gpc893 (
      {stage0_10[138]},
      {stage1_10[71]}
   );
   gpc1_1 gpc894 (
      {stage0_10[139]},
      {stage1_10[72]}
   );
   gpc1_1 gpc895 (
      {stage0_10[140]},
      {stage1_10[73]}
   );
   gpc1_1 gpc896 (
      {stage0_10[141]},
      {stage1_10[74]}
   );
   gpc1_1 gpc897 (
      {stage0_10[142]},
      {stage1_10[75]}
   );
   gpc1_1 gpc898 (
      {stage0_10[143]},
      {stage1_10[76]}
   );
   gpc1_1 gpc899 (
      {stage0_10[144]},
      {stage1_10[77]}
   );
   gpc1_1 gpc900 (
      {stage0_10[145]},
      {stage1_10[78]}
   );
   gpc1_1 gpc901 (
      {stage0_10[146]},
      {stage1_10[79]}
   );
   gpc1_1 gpc902 (
      {stage0_10[147]},
      {stage1_10[80]}
   );
   gpc1_1 gpc903 (
      {stage0_10[148]},
      {stage1_10[81]}
   );
   gpc1_1 gpc904 (
      {stage0_10[149]},
      {stage1_10[82]}
   );
   gpc1_1 gpc905 (
      {stage0_10[150]},
      {stage1_10[83]}
   );
   gpc1_1 gpc906 (
      {stage0_10[151]},
      {stage1_10[84]}
   );
   gpc1_1 gpc907 (
      {stage0_10[152]},
      {stage1_10[85]}
   );
   gpc1_1 gpc908 (
      {stage0_10[153]},
      {stage1_10[86]}
   );
   gpc1_1 gpc909 (
      {stage0_10[154]},
      {stage1_10[87]}
   );
   gpc1_1 gpc910 (
      {stage0_10[155]},
      {stage1_10[88]}
   );
   gpc1_1 gpc911 (
      {stage0_10[156]},
      {stage1_10[89]}
   );
   gpc1_1 gpc912 (
      {stage0_10[157]},
      {stage1_10[90]}
   );
   gpc1_1 gpc913 (
      {stage0_10[158]},
      {stage1_10[91]}
   );
   gpc1_1 gpc914 (
      {stage0_10[159]},
      {stage1_10[92]}
   );
   gpc1_1 gpc915 (
      {stage0_10[160]},
      {stage1_10[93]}
   );
   gpc1_1 gpc916 (
      {stage0_10[161]},
      {stage1_10[94]}
   );
   gpc1_1 gpc917 (
      {stage0_11[144]},
      {stage1_11[63]}
   );
   gpc1_1 gpc918 (
      {stage0_11[145]},
      {stage1_11[64]}
   );
   gpc1_1 gpc919 (
      {stage0_11[146]},
      {stage1_11[65]}
   );
   gpc1_1 gpc920 (
      {stage0_11[147]},
      {stage1_11[66]}
   );
   gpc1_1 gpc921 (
      {stage0_11[148]},
      {stage1_11[67]}
   );
   gpc1_1 gpc922 (
      {stage0_11[149]},
      {stage1_11[68]}
   );
   gpc1_1 gpc923 (
      {stage0_11[150]},
      {stage1_11[69]}
   );
   gpc1_1 gpc924 (
      {stage0_11[151]},
      {stage1_11[70]}
   );
   gpc1_1 gpc925 (
      {stage0_11[152]},
      {stage1_11[71]}
   );
   gpc1_1 gpc926 (
      {stage0_11[153]},
      {stage1_11[72]}
   );
   gpc1_1 gpc927 (
      {stage0_11[154]},
      {stage1_11[73]}
   );
   gpc1_1 gpc928 (
      {stage0_11[155]},
      {stage1_11[74]}
   );
   gpc1_1 gpc929 (
      {stage0_11[156]},
      {stage1_11[75]}
   );
   gpc1_1 gpc930 (
      {stage0_11[157]},
      {stage1_11[76]}
   );
   gpc1_1 gpc931 (
      {stage0_11[158]},
      {stage1_11[77]}
   );
   gpc1_1 gpc932 (
      {stage0_11[159]},
      {stage1_11[78]}
   );
   gpc1_1 gpc933 (
      {stage0_11[160]},
      {stage1_11[79]}
   );
   gpc1_1 gpc934 (
      {stage0_11[161]},
      {stage1_11[80]}
   );
   gpc1_1 gpc935 (
      {stage0_12[158]},
      {stage1_12[63]}
   );
   gpc1_1 gpc936 (
      {stage0_12[159]},
      {stage1_12[64]}
   );
   gpc1_1 gpc937 (
      {stage0_12[160]},
      {stage1_12[65]}
   );
   gpc1_1 gpc938 (
      {stage0_12[161]},
      {stage1_12[66]}
   );
   gpc1_1 gpc939 (
      {stage0_13[132]},
      {stage1_13[57]}
   );
   gpc1_1 gpc940 (
      {stage0_13[133]},
      {stage1_13[58]}
   );
   gpc1_1 gpc941 (
      {stage0_13[134]},
      {stage1_13[59]}
   );
   gpc1_1 gpc942 (
      {stage0_13[135]},
      {stage1_13[60]}
   );
   gpc1_1 gpc943 (
      {stage0_13[136]},
      {stage1_13[61]}
   );
   gpc1_1 gpc944 (
      {stage0_13[137]},
      {stage1_13[62]}
   );
   gpc1_1 gpc945 (
      {stage0_13[138]},
      {stage1_13[63]}
   );
   gpc1_1 gpc946 (
      {stage0_13[139]},
      {stage1_13[64]}
   );
   gpc1_1 gpc947 (
      {stage0_13[140]},
      {stage1_13[65]}
   );
   gpc1_1 gpc948 (
      {stage0_13[141]},
      {stage1_13[66]}
   );
   gpc1_1 gpc949 (
      {stage0_13[142]},
      {stage1_13[67]}
   );
   gpc1_1 gpc950 (
      {stage0_13[143]},
      {stage1_13[68]}
   );
   gpc1_1 gpc951 (
      {stage0_13[144]},
      {stage1_13[69]}
   );
   gpc1_1 gpc952 (
      {stage0_13[145]},
      {stage1_13[70]}
   );
   gpc1_1 gpc953 (
      {stage0_13[146]},
      {stage1_13[71]}
   );
   gpc1_1 gpc954 (
      {stage0_13[147]},
      {stage1_13[72]}
   );
   gpc1_1 gpc955 (
      {stage0_13[148]},
      {stage1_13[73]}
   );
   gpc1_1 gpc956 (
      {stage0_13[149]},
      {stage1_13[74]}
   );
   gpc1_1 gpc957 (
      {stage0_13[150]},
      {stage1_13[75]}
   );
   gpc1_1 gpc958 (
      {stage0_13[151]},
      {stage1_13[76]}
   );
   gpc1_1 gpc959 (
      {stage0_13[152]},
      {stage1_13[77]}
   );
   gpc1_1 gpc960 (
      {stage0_13[153]},
      {stage1_13[78]}
   );
   gpc1_1 gpc961 (
      {stage0_13[154]},
      {stage1_13[79]}
   );
   gpc1_1 gpc962 (
      {stage0_13[155]},
      {stage1_13[80]}
   );
   gpc1_1 gpc963 (
      {stage0_13[156]},
      {stage1_13[81]}
   );
   gpc1_1 gpc964 (
      {stage0_13[157]},
      {stage1_13[82]}
   );
   gpc1_1 gpc965 (
      {stage0_13[158]},
      {stage1_13[83]}
   );
   gpc1_1 gpc966 (
      {stage0_13[159]},
      {stage1_13[84]}
   );
   gpc1_1 gpc967 (
      {stage0_13[160]},
      {stage1_13[85]}
   );
   gpc1_1 gpc968 (
      {stage0_13[161]},
      {stage1_13[86]}
   );
   gpc1_1 gpc969 (
      {stage0_14[158]},
      {stage1_14[58]}
   );
   gpc1_1 gpc970 (
      {stage0_14[159]},
      {stage1_14[59]}
   );
   gpc1_1 gpc971 (
      {stage0_14[160]},
      {stage1_14[60]}
   );
   gpc1_1 gpc972 (
      {stage0_14[161]},
      {stage1_14[61]}
   );
   gpc1_1 gpc973 (
      {stage0_15[128]},
      {stage1_15[64]}
   );
   gpc1_1 gpc974 (
      {stage0_15[129]},
      {stage1_15[65]}
   );
   gpc1_1 gpc975 (
      {stage0_15[130]},
      {stage1_15[66]}
   );
   gpc1_1 gpc976 (
      {stage0_15[131]},
      {stage1_15[67]}
   );
   gpc1_1 gpc977 (
      {stage0_15[132]},
      {stage1_15[68]}
   );
   gpc1_1 gpc978 (
      {stage0_15[133]},
      {stage1_15[69]}
   );
   gpc1_1 gpc979 (
      {stage0_15[134]},
      {stage1_15[70]}
   );
   gpc1_1 gpc980 (
      {stage0_15[135]},
      {stage1_15[71]}
   );
   gpc1_1 gpc981 (
      {stage0_15[136]},
      {stage1_15[72]}
   );
   gpc1_1 gpc982 (
      {stage0_15[137]},
      {stage1_15[73]}
   );
   gpc1_1 gpc983 (
      {stage0_15[138]},
      {stage1_15[74]}
   );
   gpc1_1 gpc984 (
      {stage0_15[139]},
      {stage1_15[75]}
   );
   gpc1_1 gpc985 (
      {stage0_15[140]},
      {stage1_15[76]}
   );
   gpc1_1 gpc986 (
      {stage0_15[141]},
      {stage1_15[77]}
   );
   gpc1_1 gpc987 (
      {stage0_15[142]},
      {stage1_15[78]}
   );
   gpc1_1 gpc988 (
      {stage0_15[143]},
      {stage1_15[79]}
   );
   gpc1_1 gpc989 (
      {stage0_15[144]},
      {stage1_15[80]}
   );
   gpc1_1 gpc990 (
      {stage0_15[145]},
      {stage1_15[81]}
   );
   gpc1_1 gpc991 (
      {stage0_15[146]},
      {stage1_15[82]}
   );
   gpc1_1 gpc992 (
      {stage0_15[147]},
      {stage1_15[83]}
   );
   gpc1_1 gpc993 (
      {stage0_15[148]},
      {stage1_15[84]}
   );
   gpc1_1 gpc994 (
      {stage0_15[149]},
      {stage1_15[85]}
   );
   gpc1_1 gpc995 (
      {stage0_15[150]},
      {stage1_15[86]}
   );
   gpc1_1 gpc996 (
      {stage0_15[151]},
      {stage1_15[87]}
   );
   gpc1_1 gpc997 (
      {stage0_15[152]},
      {stage1_15[88]}
   );
   gpc1_1 gpc998 (
      {stage0_15[153]},
      {stage1_15[89]}
   );
   gpc1_1 gpc999 (
      {stage0_15[154]},
      {stage1_15[90]}
   );
   gpc1_1 gpc1000 (
      {stage0_15[155]},
      {stage1_15[91]}
   );
   gpc1_1 gpc1001 (
      {stage0_15[156]},
      {stage1_15[92]}
   );
   gpc1_1 gpc1002 (
      {stage0_15[157]},
      {stage1_15[93]}
   );
   gpc1_1 gpc1003 (
      {stage0_15[158]},
      {stage1_15[94]}
   );
   gpc1_1 gpc1004 (
      {stage0_15[159]},
      {stage1_15[95]}
   );
   gpc1_1 gpc1005 (
      {stage0_15[160]},
      {stage1_15[96]}
   );
   gpc1_1 gpc1006 (
      {stage0_15[161]},
      {stage1_15[97]}
   );
   gpc1_1 gpc1007 (
      {stage0_16[158]},
      {stage1_16[64]}
   );
   gpc1_1 gpc1008 (
      {stage0_16[159]},
      {stage1_16[65]}
   );
   gpc1_1 gpc1009 (
      {stage0_16[160]},
      {stage1_16[66]}
   );
   gpc1_1 gpc1010 (
      {stage0_16[161]},
      {stage1_16[67]}
   );
   gpc1_1 gpc1011 (
      {stage0_17[96]},
      {stage1_17[48]}
   );
   gpc1_1 gpc1012 (
      {stage0_17[97]},
      {stage1_17[49]}
   );
   gpc1_1 gpc1013 (
      {stage0_17[98]},
      {stage1_17[50]}
   );
   gpc1_1 gpc1014 (
      {stage0_17[99]},
      {stage1_17[51]}
   );
   gpc1_1 gpc1015 (
      {stage0_17[100]},
      {stage1_17[52]}
   );
   gpc1_1 gpc1016 (
      {stage0_17[101]},
      {stage1_17[53]}
   );
   gpc1_1 gpc1017 (
      {stage0_17[102]},
      {stage1_17[54]}
   );
   gpc1_1 gpc1018 (
      {stage0_17[103]},
      {stage1_17[55]}
   );
   gpc1_1 gpc1019 (
      {stage0_17[104]},
      {stage1_17[56]}
   );
   gpc1_1 gpc1020 (
      {stage0_17[105]},
      {stage1_17[57]}
   );
   gpc1_1 gpc1021 (
      {stage0_17[106]},
      {stage1_17[58]}
   );
   gpc1_1 gpc1022 (
      {stage0_17[107]},
      {stage1_17[59]}
   );
   gpc1_1 gpc1023 (
      {stage0_17[108]},
      {stage1_17[60]}
   );
   gpc1_1 gpc1024 (
      {stage0_17[109]},
      {stage1_17[61]}
   );
   gpc1_1 gpc1025 (
      {stage0_17[110]},
      {stage1_17[62]}
   );
   gpc1_1 gpc1026 (
      {stage0_17[111]},
      {stage1_17[63]}
   );
   gpc1_1 gpc1027 (
      {stage0_17[112]},
      {stage1_17[64]}
   );
   gpc1_1 gpc1028 (
      {stage0_17[113]},
      {stage1_17[65]}
   );
   gpc1_1 gpc1029 (
      {stage0_17[114]},
      {stage1_17[66]}
   );
   gpc1_1 gpc1030 (
      {stage0_17[115]},
      {stage1_17[67]}
   );
   gpc1_1 gpc1031 (
      {stage0_17[116]},
      {stage1_17[68]}
   );
   gpc1_1 gpc1032 (
      {stage0_17[117]},
      {stage1_17[69]}
   );
   gpc1_1 gpc1033 (
      {stage0_17[118]},
      {stage1_17[70]}
   );
   gpc1_1 gpc1034 (
      {stage0_17[119]},
      {stage1_17[71]}
   );
   gpc1_1 gpc1035 (
      {stage0_17[120]},
      {stage1_17[72]}
   );
   gpc1_1 gpc1036 (
      {stage0_17[121]},
      {stage1_17[73]}
   );
   gpc1_1 gpc1037 (
      {stage0_17[122]},
      {stage1_17[74]}
   );
   gpc1_1 gpc1038 (
      {stage0_17[123]},
      {stage1_17[75]}
   );
   gpc1_1 gpc1039 (
      {stage0_17[124]},
      {stage1_17[76]}
   );
   gpc1_1 gpc1040 (
      {stage0_17[125]},
      {stage1_17[77]}
   );
   gpc1_1 gpc1041 (
      {stage0_17[126]},
      {stage1_17[78]}
   );
   gpc1_1 gpc1042 (
      {stage0_17[127]},
      {stage1_17[79]}
   );
   gpc1_1 gpc1043 (
      {stage0_17[128]},
      {stage1_17[80]}
   );
   gpc1_1 gpc1044 (
      {stage0_17[129]},
      {stage1_17[81]}
   );
   gpc1_1 gpc1045 (
      {stage0_17[130]},
      {stage1_17[82]}
   );
   gpc1_1 gpc1046 (
      {stage0_17[131]},
      {stage1_17[83]}
   );
   gpc1_1 gpc1047 (
      {stage0_17[132]},
      {stage1_17[84]}
   );
   gpc1_1 gpc1048 (
      {stage0_17[133]},
      {stage1_17[85]}
   );
   gpc1_1 gpc1049 (
      {stage0_17[134]},
      {stage1_17[86]}
   );
   gpc1_1 gpc1050 (
      {stage0_17[135]},
      {stage1_17[87]}
   );
   gpc1_1 gpc1051 (
      {stage0_17[136]},
      {stage1_17[88]}
   );
   gpc1_1 gpc1052 (
      {stage0_17[137]},
      {stage1_17[89]}
   );
   gpc1_1 gpc1053 (
      {stage0_17[138]},
      {stage1_17[90]}
   );
   gpc1_1 gpc1054 (
      {stage0_17[139]},
      {stage1_17[91]}
   );
   gpc1_1 gpc1055 (
      {stage0_17[140]},
      {stage1_17[92]}
   );
   gpc1_1 gpc1056 (
      {stage0_17[141]},
      {stage1_17[93]}
   );
   gpc1_1 gpc1057 (
      {stage0_17[142]},
      {stage1_17[94]}
   );
   gpc1_1 gpc1058 (
      {stage0_17[143]},
      {stage1_17[95]}
   );
   gpc1_1 gpc1059 (
      {stage0_17[144]},
      {stage1_17[96]}
   );
   gpc1_1 gpc1060 (
      {stage0_17[145]},
      {stage1_17[97]}
   );
   gpc1_1 gpc1061 (
      {stage0_17[146]},
      {stage1_17[98]}
   );
   gpc1_1 gpc1062 (
      {stage0_17[147]},
      {stage1_17[99]}
   );
   gpc1_1 gpc1063 (
      {stage0_17[148]},
      {stage1_17[100]}
   );
   gpc1_1 gpc1064 (
      {stage0_17[149]},
      {stage1_17[101]}
   );
   gpc1_1 gpc1065 (
      {stage0_17[150]},
      {stage1_17[102]}
   );
   gpc1_1 gpc1066 (
      {stage0_17[151]},
      {stage1_17[103]}
   );
   gpc1_1 gpc1067 (
      {stage0_17[152]},
      {stage1_17[104]}
   );
   gpc1_1 gpc1068 (
      {stage0_17[153]},
      {stage1_17[105]}
   );
   gpc1_1 gpc1069 (
      {stage0_17[154]},
      {stage1_17[106]}
   );
   gpc1_1 gpc1070 (
      {stage0_17[155]},
      {stage1_17[107]}
   );
   gpc1_1 gpc1071 (
      {stage0_17[156]},
      {stage1_17[108]}
   );
   gpc1_1 gpc1072 (
      {stage0_17[157]},
      {stage1_17[109]}
   );
   gpc1_1 gpc1073 (
      {stage0_17[158]},
      {stage1_17[110]}
   );
   gpc1_1 gpc1074 (
      {stage0_17[159]},
      {stage1_17[111]}
   );
   gpc1_1 gpc1075 (
      {stage0_17[160]},
      {stage1_17[112]}
   );
   gpc1_1 gpc1076 (
      {stage0_17[161]},
      {stage1_17[113]}
   );
   gpc1_1 gpc1077 (
      {stage0_18[151]},
      {stage1_18[52]}
   );
   gpc1_1 gpc1078 (
      {stage0_18[152]},
      {stage1_18[53]}
   );
   gpc1_1 gpc1079 (
      {stage0_18[153]},
      {stage1_18[54]}
   );
   gpc1_1 gpc1080 (
      {stage0_18[154]},
      {stage1_18[55]}
   );
   gpc1_1 gpc1081 (
      {stage0_18[155]},
      {stage1_18[56]}
   );
   gpc1_1 gpc1082 (
      {stage0_18[156]},
      {stage1_18[57]}
   );
   gpc1_1 gpc1083 (
      {stage0_18[157]},
      {stage1_18[58]}
   );
   gpc1_1 gpc1084 (
      {stage0_18[158]},
      {stage1_18[59]}
   );
   gpc1_1 gpc1085 (
      {stage0_18[159]},
      {stage1_18[60]}
   );
   gpc1_1 gpc1086 (
      {stage0_18[160]},
      {stage1_18[61]}
   );
   gpc1_1 gpc1087 (
      {stage0_18[161]},
      {stage1_18[62]}
   );
   gpc1_1 gpc1088 (
      {stage0_19[156]},
      {stage1_19[65]}
   );
   gpc1_1 gpc1089 (
      {stage0_19[157]},
      {stage1_19[66]}
   );
   gpc1_1 gpc1090 (
      {stage0_19[158]},
      {stage1_19[67]}
   );
   gpc1_1 gpc1091 (
      {stage0_19[159]},
      {stage1_19[68]}
   );
   gpc1_1 gpc1092 (
      {stage0_19[160]},
      {stage1_19[69]}
   );
   gpc1_1 gpc1093 (
      {stage0_19[161]},
      {stage1_19[70]}
   );
   gpc1_1 gpc1094 (
      {stage0_20[159]},
      {stage1_20[65]}
   );
   gpc1_1 gpc1095 (
      {stage0_20[160]},
      {stage1_20[66]}
   );
   gpc1_1 gpc1096 (
      {stage0_20[161]},
      {stage1_20[67]}
   );
   gpc1_1 gpc1097 (
      {stage0_21[147]},
      {stage1_21[56]}
   );
   gpc1_1 gpc1098 (
      {stage0_21[148]},
      {stage1_21[57]}
   );
   gpc1_1 gpc1099 (
      {stage0_21[149]},
      {stage1_21[58]}
   );
   gpc1_1 gpc1100 (
      {stage0_21[150]},
      {stage1_21[59]}
   );
   gpc1_1 gpc1101 (
      {stage0_21[151]},
      {stage1_21[60]}
   );
   gpc1_1 gpc1102 (
      {stage0_21[152]},
      {stage1_21[61]}
   );
   gpc1_1 gpc1103 (
      {stage0_21[153]},
      {stage1_21[62]}
   );
   gpc1_1 gpc1104 (
      {stage0_21[154]},
      {stage1_21[63]}
   );
   gpc1_1 gpc1105 (
      {stage0_21[155]},
      {stage1_21[64]}
   );
   gpc1_1 gpc1106 (
      {stage0_21[156]},
      {stage1_21[65]}
   );
   gpc1_1 gpc1107 (
      {stage0_21[157]},
      {stage1_21[66]}
   );
   gpc1_1 gpc1108 (
      {stage0_21[158]},
      {stage1_21[67]}
   );
   gpc1_1 gpc1109 (
      {stage0_21[159]},
      {stage1_21[68]}
   );
   gpc1_1 gpc1110 (
      {stage0_21[160]},
      {stage1_21[69]}
   );
   gpc1_1 gpc1111 (
      {stage0_21[161]},
      {stage1_21[70]}
   );
   gpc1_1 gpc1112 (
      {stage0_23[77]},
      {stage1_23[58]}
   );
   gpc1_1 gpc1113 (
      {stage0_23[78]},
      {stage1_23[59]}
   );
   gpc1_1 gpc1114 (
      {stage0_23[79]},
      {stage1_23[60]}
   );
   gpc1_1 gpc1115 (
      {stage0_23[80]},
      {stage1_23[61]}
   );
   gpc1_1 gpc1116 (
      {stage0_23[81]},
      {stage1_23[62]}
   );
   gpc1_1 gpc1117 (
      {stage0_23[82]},
      {stage1_23[63]}
   );
   gpc1_1 gpc1118 (
      {stage0_23[83]},
      {stage1_23[64]}
   );
   gpc1_1 gpc1119 (
      {stage0_23[84]},
      {stage1_23[65]}
   );
   gpc1_1 gpc1120 (
      {stage0_23[85]},
      {stage1_23[66]}
   );
   gpc1_1 gpc1121 (
      {stage0_23[86]},
      {stage1_23[67]}
   );
   gpc1_1 gpc1122 (
      {stage0_23[87]},
      {stage1_23[68]}
   );
   gpc1_1 gpc1123 (
      {stage0_23[88]},
      {stage1_23[69]}
   );
   gpc1_1 gpc1124 (
      {stage0_23[89]},
      {stage1_23[70]}
   );
   gpc1_1 gpc1125 (
      {stage0_23[90]},
      {stage1_23[71]}
   );
   gpc1_1 gpc1126 (
      {stage0_23[91]},
      {stage1_23[72]}
   );
   gpc1_1 gpc1127 (
      {stage0_23[92]},
      {stage1_23[73]}
   );
   gpc1_1 gpc1128 (
      {stage0_23[93]},
      {stage1_23[74]}
   );
   gpc1_1 gpc1129 (
      {stage0_23[94]},
      {stage1_23[75]}
   );
   gpc1_1 gpc1130 (
      {stage0_23[95]},
      {stage1_23[76]}
   );
   gpc1_1 gpc1131 (
      {stage0_23[96]},
      {stage1_23[77]}
   );
   gpc1_1 gpc1132 (
      {stage0_23[97]},
      {stage1_23[78]}
   );
   gpc1_1 gpc1133 (
      {stage0_23[98]},
      {stage1_23[79]}
   );
   gpc1_1 gpc1134 (
      {stage0_23[99]},
      {stage1_23[80]}
   );
   gpc1_1 gpc1135 (
      {stage0_23[100]},
      {stage1_23[81]}
   );
   gpc1_1 gpc1136 (
      {stage0_23[101]},
      {stage1_23[82]}
   );
   gpc1_1 gpc1137 (
      {stage0_23[102]},
      {stage1_23[83]}
   );
   gpc1_1 gpc1138 (
      {stage0_23[103]},
      {stage1_23[84]}
   );
   gpc1_1 gpc1139 (
      {stage0_23[104]},
      {stage1_23[85]}
   );
   gpc1_1 gpc1140 (
      {stage0_23[105]},
      {stage1_23[86]}
   );
   gpc1_1 gpc1141 (
      {stage0_23[106]},
      {stage1_23[87]}
   );
   gpc1_1 gpc1142 (
      {stage0_23[107]},
      {stage1_23[88]}
   );
   gpc1_1 gpc1143 (
      {stage0_23[108]},
      {stage1_23[89]}
   );
   gpc1_1 gpc1144 (
      {stage0_23[109]},
      {stage1_23[90]}
   );
   gpc1_1 gpc1145 (
      {stage0_23[110]},
      {stage1_23[91]}
   );
   gpc1_1 gpc1146 (
      {stage0_23[111]},
      {stage1_23[92]}
   );
   gpc1_1 gpc1147 (
      {stage0_23[112]},
      {stage1_23[93]}
   );
   gpc1_1 gpc1148 (
      {stage0_23[113]},
      {stage1_23[94]}
   );
   gpc1_1 gpc1149 (
      {stage0_23[114]},
      {stage1_23[95]}
   );
   gpc1_1 gpc1150 (
      {stage0_23[115]},
      {stage1_23[96]}
   );
   gpc1_1 gpc1151 (
      {stage0_23[116]},
      {stage1_23[97]}
   );
   gpc1_1 gpc1152 (
      {stage0_23[117]},
      {stage1_23[98]}
   );
   gpc1_1 gpc1153 (
      {stage0_23[118]},
      {stage1_23[99]}
   );
   gpc1_1 gpc1154 (
      {stage0_23[119]},
      {stage1_23[100]}
   );
   gpc1_1 gpc1155 (
      {stage0_23[120]},
      {stage1_23[101]}
   );
   gpc1_1 gpc1156 (
      {stage0_23[121]},
      {stage1_23[102]}
   );
   gpc1_1 gpc1157 (
      {stage0_23[122]},
      {stage1_23[103]}
   );
   gpc1_1 gpc1158 (
      {stage0_23[123]},
      {stage1_23[104]}
   );
   gpc1_1 gpc1159 (
      {stage0_23[124]},
      {stage1_23[105]}
   );
   gpc1_1 gpc1160 (
      {stage0_23[125]},
      {stage1_23[106]}
   );
   gpc1_1 gpc1161 (
      {stage0_23[126]},
      {stage1_23[107]}
   );
   gpc1_1 gpc1162 (
      {stage0_23[127]},
      {stage1_23[108]}
   );
   gpc1_1 gpc1163 (
      {stage0_23[128]},
      {stage1_23[109]}
   );
   gpc1_1 gpc1164 (
      {stage0_23[129]},
      {stage1_23[110]}
   );
   gpc1_1 gpc1165 (
      {stage0_23[130]},
      {stage1_23[111]}
   );
   gpc1_1 gpc1166 (
      {stage0_23[131]},
      {stage1_23[112]}
   );
   gpc1_1 gpc1167 (
      {stage0_23[132]},
      {stage1_23[113]}
   );
   gpc1_1 gpc1168 (
      {stage0_23[133]},
      {stage1_23[114]}
   );
   gpc1_1 gpc1169 (
      {stage0_23[134]},
      {stage1_23[115]}
   );
   gpc1_1 gpc1170 (
      {stage0_23[135]},
      {stage1_23[116]}
   );
   gpc1_1 gpc1171 (
      {stage0_23[136]},
      {stage1_23[117]}
   );
   gpc1_1 gpc1172 (
      {stage0_23[137]},
      {stage1_23[118]}
   );
   gpc1_1 gpc1173 (
      {stage0_23[138]},
      {stage1_23[119]}
   );
   gpc1_1 gpc1174 (
      {stage0_23[139]},
      {stage1_23[120]}
   );
   gpc1_1 gpc1175 (
      {stage0_23[140]},
      {stage1_23[121]}
   );
   gpc1_1 gpc1176 (
      {stage0_23[141]},
      {stage1_23[122]}
   );
   gpc1_1 gpc1177 (
      {stage0_23[142]},
      {stage1_23[123]}
   );
   gpc1_1 gpc1178 (
      {stage0_23[143]},
      {stage1_23[124]}
   );
   gpc1_1 gpc1179 (
      {stage0_23[144]},
      {stage1_23[125]}
   );
   gpc1_1 gpc1180 (
      {stage0_23[145]},
      {stage1_23[126]}
   );
   gpc1_1 gpc1181 (
      {stage0_23[146]},
      {stage1_23[127]}
   );
   gpc1_1 gpc1182 (
      {stage0_23[147]},
      {stage1_23[128]}
   );
   gpc1_1 gpc1183 (
      {stage0_23[148]},
      {stage1_23[129]}
   );
   gpc1_1 gpc1184 (
      {stage0_23[149]},
      {stage1_23[130]}
   );
   gpc1_1 gpc1185 (
      {stage0_23[150]},
      {stage1_23[131]}
   );
   gpc1_1 gpc1186 (
      {stage0_23[151]},
      {stage1_23[132]}
   );
   gpc1_1 gpc1187 (
      {stage0_23[152]},
      {stage1_23[133]}
   );
   gpc1_1 gpc1188 (
      {stage0_23[153]},
      {stage1_23[134]}
   );
   gpc1_1 gpc1189 (
      {stage0_23[154]},
      {stage1_23[135]}
   );
   gpc1_1 gpc1190 (
      {stage0_23[155]},
      {stage1_23[136]}
   );
   gpc1_1 gpc1191 (
      {stage0_23[156]},
      {stage1_23[137]}
   );
   gpc1_1 gpc1192 (
      {stage0_23[157]},
      {stage1_23[138]}
   );
   gpc1_1 gpc1193 (
      {stage0_23[158]},
      {stage1_23[139]}
   );
   gpc1_1 gpc1194 (
      {stage0_23[159]},
      {stage1_23[140]}
   );
   gpc1_1 gpc1195 (
      {stage0_23[160]},
      {stage1_23[141]}
   );
   gpc1_1 gpc1196 (
      {stage0_23[161]},
      {stage1_23[142]}
   );
   gpc1_1 gpc1197 (
      {stage0_24[126]},
      {stage1_24[47]}
   );
   gpc1_1 gpc1198 (
      {stage0_24[127]},
      {stage1_24[48]}
   );
   gpc1_1 gpc1199 (
      {stage0_24[128]},
      {stage1_24[49]}
   );
   gpc1_1 gpc1200 (
      {stage0_24[129]},
      {stage1_24[50]}
   );
   gpc1_1 gpc1201 (
      {stage0_24[130]},
      {stage1_24[51]}
   );
   gpc1_1 gpc1202 (
      {stage0_24[131]},
      {stage1_24[52]}
   );
   gpc1_1 gpc1203 (
      {stage0_24[132]},
      {stage1_24[53]}
   );
   gpc1_1 gpc1204 (
      {stage0_24[133]},
      {stage1_24[54]}
   );
   gpc1_1 gpc1205 (
      {stage0_24[134]},
      {stage1_24[55]}
   );
   gpc1_1 gpc1206 (
      {stage0_24[135]},
      {stage1_24[56]}
   );
   gpc1_1 gpc1207 (
      {stage0_24[136]},
      {stage1_24[57]}
   );
   gpc1_1 gpc1208 (
      {stage0_24[137]},
      {stage1_24[58]}
   );
   gpc1_1 gpc1209 (
      {stage0_24[138]},
      {stage1_24[59]}
   );
   gpc1_1 gpc1210 (
      {stage0_24[139]},
      {stage1_24[60]}
   );
   gpc1_1 gpc1211 (
      {stage0_24[140]},
      {stage1_24[61]}
   );
   gpc1_1 gpc1212 (
      {stage0_24[141]},
      {stage1_24[62]}
   );
   gpc1_1 gpc1213 (
      {stage0_24[142]},
      {stage1_24[63]}
   );
   gpc1_1 gpc1214 (
      {stage0_24[143]},
      {stage1_24[64]}
   );
   gpc1_1 gpc1215 (
      {stage0_24[144]},
      {stage1_24[65]}
   );
   gpc1_1 gpc1216 (
      {stage0_24[145]},
      {stage1_24[66]}
   );
   gpc1_1 gpc1217 (
      {stage0_24[146]},
      {stage1_24[67]}
   );
   gpc1_1 gpc1218 (
      {stage0_24[147]},
      {stage1_24[68]}
   );
   gpc1_1 gpc1219 (
      {stage0_24[148]},
      {stage1_24[69]}
   );
   gpc1_1 gpc1220 (
      {stage0_24[149]},
      {stage1_24[70]}
   );
   gpc1_1 gpc1221 (
      {stage0_24[150]},
      {stage1_24[71]}
   );
   gpc1_1 gpc1222 (
      {stage0_24[151]},
      {stage1_24[72]}
   );
   gpc1_1 gpc1223 (
      {stage0_24[152]},
      {stage1_24[73]}
   );
   gpc1_1 gpc1224 (
      {stage0_24[153]},
      {stage1_24[74]}
   );
   gpc1_1 gpc1225 (
      {stage0_24[154]},
      {stage1_24[75]}
   );
   gpc1_1 gpc1226 (
      {stage0_24[155]},
      {stage1_24[76]}
   );
   gpc1_1 gpc1227 (
      {stage0_24[156]},
      {stage1_24[77]}
   );
   gpc1_1 gpc1228 (
      {stage0_24[157]},
      {stage1_24[78]}
   );
   gpc1_1 gpc1229 (
      {stage0_24[158]},
      {stage1_24[79]}
   );
   gpc1_1 gpc1230 (
      {stage0_24[159]},
      {stage1_24[80]}
   );
   gpc1_1 gpc1231 (
      {stage0_24[160]},
      {stage1_24[81]}
   );
   gpc1_1 gpc1232 (
      {stage0_24[161]},
      {stage1_24[82]}
   );
   gpc1_1 gpc1233 (
      {stage0_25[127]},
      {stage1_25[50]}
   );
   gpc1_1 gpc1234 (
      {stage0_25[128]},
      {stage1_25[51]}
   );
   gpc1_1 gpc1235 (
      {stage0_25[129]},
      {stage1_25[52]}
   );
   gpc1_1 gpc1236 (
      {stage0_25[130]},
      {stage1_25[53]}
   );
   gpc1_1 gpc1237 (
      {stage0_25[131]},
      {stage1_25[54]}
   );
   gpc1_1 gpc1238 (
      {stage0_25[132]},
      {stage1_25[55]}
   );
   gpc1_1 gpc1239 (
      {stage0_25[133]},
      {stage1_25[56]}
   );
   gpc1_1 gpc1240 (
      {stage0_25[134]},
      {stage1_25[57]}
   );
   gpc1_1 gpc1241 (
      {stage0_25[135]},
      {stage1_25[58]}
   );
   gpc1_1 gpc1242 (
      {stage0_25[136]},
      {stage1_25[59]}
   );
   gpc1_1 gpc1243 (
      {stage0_25[137]},
      {stage1_25[60]}
   );
   gpc1_1 gpc1244 (
      {stage0_25[138]},
      {stage1_25[61]}
   );
   gpc1_1 gpc1245 (
      {stage0_25[139]},
      {stage1_25[62]}
   );
   gpc1_1 gpc1246 (
      {stage0_25[140]},
      {stage1_25[63]}
   );
   gpc1_1 gpc1247 (
      {stage0_25[141]},
      {stage1_25[64]}
   );
   gpc1_1 gpc1248 (
      {stage0_25[142]},
      {stage1_25[65]}
   );
   gpc1_1 gpc1249 (
      {stage0_25[143]},
      {stage1_25[66]}
   );
   gpc1_1 gpc1250 (
      {stage0_25[144]},
      {stage1_25[67]}
   );
   gpc1_1 gpc1251 (
      {stage0_25[145]},
      {stage1_25[68]}
   );
   gpc1_1 gpc1252 (
      {stage0_25[146]},
      {stage1_25[69]}
   );
   gpc1_1 gpc1253 (
      {stage0_25[147]},
      {stage1_25[70]}
   );
   gpc1_1 gpc1254 (
      {stage0_25[148]},
      {stage1_25[71]}
   );
   gpc1_1 gpc1255 (
      {stage0_25[149]},
      {stage1_25[72]}
   );
   gpc1_1 gpc1256 (
      {stage0_25[150]},
      {stage1_25[73]}
   );
   gpc1_1 gpc1257 (
      {stage0_25[151]},
      {stage1_25[74]}
   );
   gpc1_1 gpc1258 (
      {stage0_25[152]},
      {stage1_25[75]}
   );
   gpc1_1 gpc1259 (
      {stage0_25[153]},
      {stage1_25[76]}
   );
   gpc1_1 gpc1260 (
      {stage0_25[154]},
      {stage1_25[77]}
   );
   gpc1_1 gpc1261 (
      {stage0_25[155]},
      {stage1_25[78]}
   );
   gpc1_1 gpc1262 (
      {stage0_25[156]},
      {stage1_25[79]}
   );
   gpc1_1 gpc1263 (
      {stage0_25[157]},
      {stage1_25[80]}
   );
   gpc1_1 gpc1264 (
      {stage0_25[158]},
      {stage1_25[81]}
   );
   gpc1_1 gpc1265 (
      {stage0_25[159]},
      {stage1_25[82]}
   );
   gpc1_1 gpc1266 (
      {stage0_25[160]},
      {stage1_25[83]}
   );
   gpc1_1 gpc1267 (
      {stage0_25[161]},
      {stage1_25[84]}
   );
   gpc1_1 gpc1268 (
      {stage0_26[149]},
      {stage1_26[59]}
   );
   gpc1_1 gpc1269 (
      {stage0_26[150]},
      {stage1_26[60]}
   );
   gpc1_1 gpc1270 (
      {stage0_26[151]},
      {stage1_26[61]}
   );
   gpc1_1 gpc1271 (
      {stage0_26[152]},
      {stage1_26[62]}
   );
   gpc1_1 gpc1272 (
      {stage0_26[153]},
      {stage1_26[63]}
   );
   gpc1_1 gpc1273 (
      {stage0_26[154]},
      {stage1_26[64]}
   );
   gpc1_1 gpc1274 (
      {stage0_26[155]},
      {stage1_26[65]}
   );
   gpc1_1 gpc1275 (
      {stage0_26[156]},
      {stage1_26[66]}
   );
   gpc1_1 gpc1276 (
      {stage0_26[157]},
      {stage1_26[67]}
   );
   gpc1_1 gpc1277 (
      {stage0_26[158]},
      {stage1_26[68]}
   );
   gpc1_1 gpc1278 (
      {stage0_26[159]},
      {stage1_26[69]}
   );
   gpc1_1 gpc1279 (
      {stage0_26[160]},
      {stage1_26[70]}
   );
   gpc1_1 gpc1280 (
      {stage0_26[161]},
      {stage1_26[71]}
   );
   gpc1_1 gpc1281 (
      {stage0_27[142]},
      {stage1_27[54]}
   );
   gpc1_1 gpc1282 (
      {stage0_27[143]},
      {stage1_27[55]}
   );
   gpc1_1 gpc1283 (
      {stage0_27[144]},
      {stage1_27[56]}
   );
   gpc1_1 gpc1284 (
      {stage0_27[145]},
      {stage1_27[57]}
   );
   gpc1_1 gpc1285 (
      {stage0_27[146]},
      {stage1_27[58]}
   );
   gpc1_1 gpc1286 (
      {stage0_27[147]},
      {stage1_27[59]}
   );
   gpc1_1 gpc1287 (
      {stage0_27[148]},
      {stage1_27[60]}
   );
   gpc1_1 gpc1288 (
      {stage0_27[149]},
      {stage1_27[61]}
   );
   gpc1_1 gpc1289 (
      {stage0_27[150]},
      {stage1_27[62]}
   );
   gpc1_1 gpc1290 (
      {stage0_27[151]},
      {stage1_27[63]}
   );
   gpc1_1 gpc1291 (
      {stage0_27[152]},
      {stage1_27[64]}
   );
   gpc1_1 gpc1292 (
      {stage0_27[153]},
      {stage1_27[65]}
   );
   gpc1_1 gpc1293 (
      {stage0_27[154]},
      {stage1_27[66]}
   );
   gpc1_1 gpc1294 (
      {stage0_27[155]},
      {stage1_27[67]}
   );
   gpc1_1 gpc1295 (
      {stage0_27[156]},
      {stage1_27[68]}
   );
   gpc1_1 gpc1296 (
      {stage0_27[157]},
      {stage1_27[69]}
   );
   gpc1_1 gpc1297 (
      {stage0_27[158]},
      {stage1_27[70]}
   );
   gpc1_1 gpc1298 (
      {stage0_27[159]},
      {stage1_27[71]}
   );
   gpc1_1 gpc1299 (
      {stage0_27[160]},
      {stage1_27[72]}
   );
   gpc1_1 gpc1300 (
      {stage0_27[161]},
      {stage1_27[73]}
   );
   gpc1_1 gpc1301 (
      {stage0_28[140]},
      {stage1_28[55]}
   );
   gpc1_1 gpc1302 (
      {stage0_28[141]},
      {stage1_28[56]}
   );
   gpc1_1 gpc1303 (
      {stage0_28[142]},
      {stage1_28[57]}
   );
   gpc1_1 gpc1304 (
      {stage0_28[143]},
      {stage1_28[58]}
   );
   gpc1_1 gpc1305 (
      {stage0_28[144]},
      {stage1_28[59]}
   );
   gpc1_1 gpc1306 (
      {stage0_28[145]},
      {stage1_28[60]}
   );
   gpc1_1 gpc1307 (
      {stage0_28[146]},
      {stage1_28[61]}
   );
   gpc1_1 gpc1308 (
      {stage0_28[147]},
      {stage1_28[62]}
   );
   gpc1_1 gpc1309 (
      {stage0_28[148]},
      {stage1_28[63]}
   );
   gpc1_1 gpc1310 (
      {stage0_28[149]},
      {stage1_28[64]}
   );
   gpc1_1 gpc1311 (
      {stage0_28[150]},
      {stage1_28[65]}
   );
   gpc1_1 gpc1312 (
      {stage0_28[151]},
      {stage1_28[66]}
   );
   gpc1_1 gpc1313 (
      {stage0_28[152]},
      {stage1_28[67]}
   );
   gpc1_1 gpc1314 (
      {stage0_28[153]},
      {stage1_28[68]}
   );
   gpc1_1 gpc1315 (
      {stage0_28[154]},
      {stage1_28[69]}
   );
   gpc1_1 gpc1316 (
      {stage0_28[155]},
      {stage1_28[70]}
   );
   gpc1_1 gpc1317 (
      {stage0_28[156]},
      {stage1_28[71]}
   );
   gpc1_1 gpc1318 (
      {stage0_28[157]},
      {stage1_28[72]}
   );
   gpc1_1 gpc1319 (
      {stage0_28[158]},
      {stage1_28[73]}
   );
   gpc1_1 gpc1320 (
      {stage0_28[159]},
      {stage1_28[74]}
   );
   gpc1_1 gpc1321 (
      {stage0_28[160]},
      {stage1_28[75]}
   );
   gpc1_1 gpc1322 (
      {stage0_28[161]},
      {stage1_28[76]}
   );
   gpc1_1 gpc1323 (
      {stage0_29[144]},
      {stage1_29[63]}
   );
   gpc1_1 gpc1324 (
      {stage0_29[145]},
      {stage1_29[64]}
   );
   gpc1_1 gpc1325 (
      {stage0_29[146]},
      {stage1_29[65]}
   );
   gpc1_1 gpc1326 (
      {stage0_29[147]},
      {stage1_29[66]}
   );
   gpc1_1 gpc1327 (
      {stage0_29[148]},
      {stage1_29[67]}
   );
   gpc1_1 gpc1328 (
      {stage0_29[149]},
      {stage1_29[68]}
   );
   gpc1_1 gpc1329 (
      {stage0_29[150]},
      {stage1_29[69]}
   );
   gpc1_1 gpc1330 (
      {stage0_29[151]},
      {stage1_29[70]}
   );
   gpc1_1 gpc1331 (
      {stage0_29[152]},
      {stage1_29[71]}
   );
   gpc1_1 gpc1332 (
      {stage0_29[153]},
      {stage1_29[72]}
   );
   gpc1_1 gpc1333 (
      {stage0_29[154]},
      {stage1_29[73]}
   );
   gpc1_1 gpc1334 (
      {stage0_29[155]},
      {stage1_29[74]}
   );
   gpc1_1 gpc1335 (
      {stage0_29[156]},
      {stage1_29[75]}
   );
   gpc1_1 gpc1336 (
      {stage0_29[157]},
      {stage1_29[76]}
   );
   gpc1_1 gpc1337 (
      {stage0_29[158]},
      {stage1_29[77]}
   );
   gpc1_1 gpc1338 (
      {stage0_29[159]},
      {stage1_29[78]}
   );
   gpc1_1 gpc1339 (
      {stage0_29[160]},
      {stage1_29[79]}
   );
   gpc1_1 gpc1340 (
      {stage0_29[161]},
      {stage1_29[80]}
   );
   gpc1_1 gpc1341 (
      {stage0_30[111]},
      {stage1_30[56]}
   );
   gpc1_1 gpc1342 (
      {stage0_30[112]},
      {stage1_30[57]}
   );
   gpc1_1 gpc1343 (
      {stage0_30[113]},
      {stage1_30[58]}
   );
   gpc1_1 gpc1344 (
      {stage0_30[114]},
      {stage1_30[59]}
   );
   gpc1_1 gpc1345 (
      {stage0_30[115]},
      {stage1_30[60]}
   );
   gpc1_1 gpc1346 (
      {stage0_30[116]},
      {stage1_30[61]}
   );
   gpc1_1 gpc1347 (
      {stage0_30[117]},
      {stage1_30[62]}
   );
   gpc1_1 gpc1348 (
      {stage0_30[118]},
      {stage1_30[63]}
   );
   gpc1_1 gpc1349 (
      {stage0_30[119]},
      {stage1_30[64]}
   );
   gpc1_1 gpc1350 (
      {stage0_30[120]},
      {stage1_30[65]}
   );
   gpc1_1 gpc1351 (
      {stage0_30[121]},
      {stage1_30[66]}
   );
   gpc1_1 gpc1352 (
      {stage0_30[122]},
      {stage1_30[67]}
   );
   gpc1_1 gpc1353 (
      {stage0_30[123]},
      {stage1_30[68]}
   );
   gpc1_1 gpc1354 (
      {stage0_30[124]},
      {stage1_30[69]}
   );
   gpc1_1 gpc1355 (
      {stage0_30[125]},
      {stage1_30[70]}
   );
   gpc1_1 gpc1356 (
      {stage0_30[126]},
      {stage1_30[71]}
   );
   gpc1_1 gpc1357 (
      {stage0_30[127]},
      {stage1_30[72]}
   );
   gpc1_1 gpc1358 (
      {stage0_30[128]},
      {stage1_30[73]}
   );
   gpc1_1 gpc1359 (
      {stage0_30[129]},
      {stage1_30[74]}
   );
   gpc1_1 gpc1360 (
      {stage0_30[130]},
      {stage1_30[75]}
   );
   gpc1_1 gpc1361 (
      {stage0_30[131]},
      {stage1_30[76]}
   );
   gpc1_1 gpc1362 (
      {stage0_30[132]},
      {stage1_30[77]}
   );
   gpc1_1 gpc1363 (
      {stage0_30[133]},
      {stage1_30[78]}
   );
   gpc1_1 gpc1364 (
      {stage0_30[134]},
      {stage1_30[79]}
   );
   gpc1_1 gpc1365 (
      {stage0_30[135]},
      {stage1_30[80]}
   );
   gpc1_1 gpc1366 (
      {stage0_30[136]},
      {stage1_30[81]}
   );
   gpc1_1 gpc1367 (
      {stage0_30[137]},
      {stage1_30[82]}
   );
   gpc1_1 gpc1368 (
      {stage0_30[138]},
      {stage1_30[83]}
   );
   gpc1_1 gpc1369 (
      {stage0_30[139]},
      {stage1_30[84]}
   );
   gpc1_1 gpc1370 (
      {stage0_30[140]},
      {stage1_30[85]}
   );
   gpc1_1 gpc1371 (
      {stage0_30[141]},
      {stage1_30[86]}
   );
   gpc1_1 gpc1372 (
      {stage0_30[142]},
      {stage1_30[87]}
   );
   gpc1_1 gpc1373 (
      {stage0_30[143]},
      {stage1_30[88]}
   );
   gpc1_1 gpc1374 (
      {stage0_30[144]},
      {stage1_30[89]}
   );
   gpc1_1 gpc1375 (
      {stage0_30[145]},
      {stage1_30[90]}
   );
   gpc1_1 gpc1376 (
      {stage0_30[146]},
      {stage1_30[91]}
   );
   gpc1_1 gpc1377 (
      {stage0_30[147]},
      {stage1_30[92]}
   );
   gpc1_1 gpc1378 (
      {stage0_30[148]},
      {stage1_30[93]}
   );
   gpc1_1 gpc1379 (
      {stage0_30[149]},
      {stage1_30[94]}
   );
   gpc1_1 gpc1380 (
      {stage0_30[150]},
      {stage1_30[95]}
   );
   gpc1_1 gpc1381 (
      {stage0_30[151]},
      {stage1_30[96]}
   );
   gpc1_1 gpc1382 (
      {stage0_30[152]},
      {stage1_30[97]}
   );
   gpc1_1 gpc1383 (
      {stage0_30[153]},
      {stage1_30[98]}
   );
   gpc1_1 gpc1384 (
      {stage0_30[154]},
      {stage1_30[99]}
   );
   gpc1_1 gpc1385 (
      {stage0_30[155]},
      {stage1_30[100]}
   );
   gpc1_1 gpc1386 (
      {stage0_30[156]},
      {stage1_30[101]}
   );
   gpc1_1 gpc1387 (
      {stage0_30[157]},
      {stage1_30[102]}
   );
   gpc1_1 gpc1388 (
      {stage0_30[158]},
      {stage1_30[103]}
   );
   gpc1_1 gpc1389 (
      {stage0_30[159]},
      {stage1_30[104]}
   );
   gpc1_1 gpc1390 (
      {stage0_30[160]},
      {stage1_30[105]}
   );
   gpc1_1 gpc1391 (
      {stage0_30[161]},
      {stage1_30[106]}
   );
   gpc1_1 gpc1392 (
      {stage0_31[109]},
      {stage1_31[44]}
   );
   gpc1_1 gpc1393 (
      {stage0_31[110]},
      {stage1_31[45]}
   );
   gpc1_1 gpc1394 (
      {stage0_31[111]},
      {stage1_31[46]}
   );
   gpc1_1 gpc1395 (
      {stage0_31[112]},
      {stage1_31[47]}
   );
   gpc1_1 gpc1396 (
      {stage0_31[113]},
      {stage1_31[48]}
   );
   gpc1_1 gpc1397 (
      {stage0_31[114]},
      {stage1_31[49]}
   );
   gpc1_1 gpc1398 (
      {stage0_31[115]},
      {stage1_31[50]}
   );
   gpc1_1 gpc1399 (
      {stage0_31[116]},
      {stage1_31[51]}
   );
   gpc1_1 gpc1400 (
      {stage0_31[117]},
      {stage1_31[52]}
   );
   gpc1_1 gpc1401 (
      {stage0_31[118]},
      {stage1_31[53]}
   );
   gpc1_1 gpc1402 (
      {stage0_31[119]},
      {stage1_31[54]}
   );
   gpc1_1 gpc1403 (
      {stage0_31[120]},
      {stage1_31[55]}
   );
   gpc1_1 gpc1404 (
      {stage0_31[121]},
      {stage1_31[56]}
   );
   gpc1_1 gpc1405 (
      {stage0_31[122]},
      {stage1_31[57]}
   );
   gpc1_1 gpc1406 (
      {stage0_31[123]},
      {stage1_31[58]}
   );
   gpc1_1 gpc1407 (
      {stage0_31[124]},
      {stage1_31[59]}
   );
   gpc1_1 gpc1408 (
      {stage0_31[125]},
      {stage1_31[60]}
   );
   gpc1_1 gpc1409 (
      {stage0_31[126]},
      {stage1_31[61]}
   );
   gpc1_1 gpc1410 (
      {stage0_31[127]},
      {stage1_31[62]}
   );
   gpc1_1 gpc1411 (
      {stage0_31[128]},
      {stage1_31[63]}
   );
   gpc1_1 gpc1412 (
      {stage0_31[129]},
      {stage1_31[64]}
   );
   gpc1_1 gpc1413 (
      {stage0_31[130]},
      {stage1_31[65]}
   );
   gpc1_1 gpc1414 (
      {stage0_31[131]},
      {stage1_31[66]}
   );
   gpc1_1 gpc1415 (
      {stage0_31[132]},
      {stage1_31[67]}
   );
   gpc1_1 gpc1416 (
      {stage0_31[133]},
      {stage1_31[68]}
   );
   gpc1_1 gpc1417 (
      {stage0_31[134]},
      {stage1_31[69]}
   );
   gpc1_1 gpc1418 (
      {stage0_31[135]},
      {stage1_31[70]}
   );
   gpc1_1 gpc1419 (
      {stage0_31[136]},
      {stage1_31[71]}
   );
   gpc1_1 gpc1420 (
      {stage0_31[137]},
      {stage1_31[72]}
   );
   gpc1_1 gpc1421 (
      {stage0_31[138]},
      {stage1_31[73]}
   );
   gpc1_1 gpc1422 (
      {stage0_31[139]},
      {stage1_31[74]}
   );
   gpc1_1 gpc1423 (
      {stage0_31[140]},
      {stage1_31[75]}
   );
   gpc1_1 gpc1424 (
      {stage0_31[141]},
      {stage1_31[76]}
   );
   gpc1_1 gpc1425 (
      {stage0_31[142]},
      {stage1_31[77]}
   );
   gpc1_1 gpc1426 (
      {stage0_31[143]},
      {stage1_31[78]}
   );
   gpc1_1 gpc1427 (
      {stage0_31[144]},
      {stage1_31[79]}
   );
   gpc1_1 gpc1428 (
      {stage0_31[145]},
      {stage1_31[80]}
   );
   gpc1_1 gpc1429 (
      {stage0_31[146]},
      {stage1_31[81]}
   );
   gpc1_1 gpc1430 (
      {stage0_31[147]},
      {stage1_31[82]}
   );
   gpc1_1 gpc1431 (
      {stage0_31[148]},
      {stage1_31[83]}
   );
   gpc1_1 gpc1432 (
      {stage0_31[149]},
      {stage1_31[84]}
   );
   gpc1_1 gpc1433 (
      {stage0_31[150]},
      {stage1_31[85]}
   );
   gpc1_1 gpc1434 (
      {stage0_31[151]},
      {stage1_31[86]}
   );
   gpc1_1 gpc1435 (
      {stage0_31[152]},
      {stage1_31[87]}
   );
   gpc1_1 gpc1436 (
      {stage0_31[153]},
      {stage1_31[88]}
   );
   gpc1_1 gpc1437 (
      {stage0_31[154]},
      {stage1_31[89]}
   );
   gpc1_1 gpc1438 (
      {stage0_31[155]},
      {stage1_31[90]}
   );
   gpc1_1 gpc1439 (
      {stage0_31[156]},
      {stage1_31[91]}
   );
   gpc1_1 gpc1440 (
      {stage0_31[157]},
      {stage1_31[92]}
   );
   gpc1_1 gpc1441 (
      {stage0_31[158]},
      {stage1_31[93]}
   );
   gpc1_1 gpc1442 (
      {stage0_31[159]},
      {stage1_31[94]}
   );
   gpc1_1 gpc1443 (
      {stage0_31[160]},
      {stage1_31[95]}
   );
   gpc1_1 gpc1444 (
      {stage0_31[161]},
      {stage1_31[96]}
   );
   gpc1_1 gpc1445 (
      {stage0_32[129]},
      {stage1_32[54]}
   );
   gpc1_1 gpc1446 (
      {stage0_32[130]},
      {stage1_32[55]}
   );
   gpc1_1 gpc1447 (
      {stage0_32[131]},
      {stage1_32[56]}
   );
   gpc1_1 gpc1448 (
      {stage0_32[132]},
      {stage1_32[57]}
   );
   gpc1_1 gpc1449 (
      {stage0_32[133]},
      {stage1_32[58]}
   );
   gpc1_1 gpc1450 (
      {stage0_32[134]},
      {stage1_32[59]}
   );
   gpc1_1 gpc1451 (
      {stage0_32[135]},
      {stage1_32[60]}
   );
   gpc1_1 gpc1452 (
      {stage0_32[136]},
      {stage1_32[61]}
   );
   gpc1_1 gpc1453 (
      {stage0_32[137]},
      {stage1_32[62]}
   );
   gpc1_1 gpc1454 (
      {stage0_32[138]},
      {stage1_32[63]}
   );
   gpc1_1 gpc1455 (
      {stage0_32[139]},
      {stage1_32[64]}
   );
   gpc1_1 gpc1456 (
      {stage0_32[140]},
      {stage1_32[65]}
   );
   gpc1_1 gpc1457 (
      {stage0_32[141]},
      {stage1_32[66]}
   );
   gpc1_1 gpc1458 (
      {stage0_32[142]},
      {stage1_32[67]}
   );
   gpc1_1 gpc1459 (
      {stage0_32[143]},
      {stage1_32[68]}
   );
   gpc1_1 gpc1460 (
      {stage0_32[144]},
      {stage1_32[69]}
   );
   gpc1_1 gpc1461 (
      {stage0_32[145]},
      {stage1_32[70]}
   );
   gpc1_1 gpc1462 (
      {stage0_32[146]},
      {stage1_32[71]}
   );
   gpc1_1 gpc1463 (
      {stage0_32[147]},
      {stage1_32[72]}
   );
   gpc1_1 gpc1464 (
      {stage0_32[148]},
      {stage1_32[73]}
   );
   gpc1_1 gpc1465 (
      {stage0_32[149]},
      {stage1_32[74]}
   );
   gpc1_1 gpc1466 (
      {stage0_32[150]},
      {stage1_32[75]}
   );
   gpc1_1 gpc1467 (
      {stage0_32[151]},
      {stage1_32[76]}
   );
   gpc1_1 gpc1468 (
      {stage0_32[152]},
      {stage1_32[77]}
   );
   gpc1_1 gpc1469 (
      {stage0_32[153]},
      {stage1_32[78]}
   );
   gpc1_1 gpc1470 (
      {stage0_32[154]},
      {stage1_32[79]}
   );
   gpc1_1 gpc1471 (
      {stage0_32[155]},
      {stage1_32[80]}
   );
   gpc1_1 gpc1472 (
      {stage0_32[156]},
      {stage1_32[81]}
   );
   gpc1_1 gpc1473 (
      {stage0_32[157]},
      {stage1_32[82]}
   );
   gpc1_1 gpc1474 (
      {stage0_32[158]},
      {stage1_32[83]}
   );
   gpc1_1 gpc1475 (
      {stage0_32[159]},
      {stage1_32[84]}
   );
   gpc1_1 gpc1476 (
      {stage0_32[160]},
      {stage1_32[85]}
   );
   gpc1_1 gpc1477 (
      {stage0_32[161]},
      {stage1_32[86]}
   );
   gpc1_1 gpc1478 (
      {stage0_33[136]},
      {stage1_33[64]}
   );
   gpc1_1 gpc1479 (
      {stage0_33[137]},
      {stage1_33[65]}
   );
   gpc1_1 gpc1480 (
      {stage0_33[138]},
      {stage1_33[66]}
   );
   gpc1_1 gpc1481 (
      {stage0_33[139]},
      {stage1_33[67]}
   );
   gpc1_1 gpc1482 (
      {stage0_33[140]},
      {stage1_33[68]}
   );
   gpc1_1 gpc1483 (
      {stage0_33[141]},
      {stage1_33[69]}
   );
   gpc1_1 gpc1484 (
      {stage0_33[142]},
      {stage1_33[70]}
   );
   gpc1_1 gpc1485 (
      {stage0_33[143]},
      {stage1_33[71]}
   );
   gpc1_1 gpc1486 (
      {stage0_33[144]},
      {stage1_33[72]}
   );
   gpc1_1 gpc1487 (
      {stage0_33[145]},
      {stage1_33[73]}
   );
   gpc1_1 gpc1488 (
      {stage0_33[146]},
      {stage1_33[74]}
   );
   gpc1_1 gpc1489 (
      {stage0_33[147]},
      {stage1_33[75]}
   );
   gpc1_1 gpc1490 (
      {stage0_33[148]},
      {stage1_33[76]}
   );
   gpc1_1 gpc1491 (
      {stage0_33[149]},
      {stage1_33[77]}
   );
   gpc1_1 gpc1492 (
      {stage0_33[150]},
      {stage1_33[78]}
   );
   gpc1_1 gpc1493 (
      {stage0_33[151]},
      {stage1_33[79]}
   );
   gpc1_1 gpc1494 (
      {stage0_33[152]},
      {stage1_33[80]}
   );
   gpc1_1 gpc1495 (
      {stage0_33[153]},
      {stage1_33[81]}
   );
   gpc1_1 gpc1496 (
      {stage0_33[154]},
      {stage1_33[82]}
   );
   gpc1_1 gpc1497 (
      {stage0_33[155]},
      {stage1_33[83]}
   );
   gpc1_1 gpc1498 (
      {stage0_33[156]},
      {stage1_33[84]}
   );
   gpc1_1 gpc1499 (
      {stage0_33[157]},
      {stage1_33[85]}
   );
   gpc1_1 gpc1500 (
      {stage0_33[158]},
      {stage1_33[86]}
   );
   gpc1_1 gpc1501 (
      {stage0_33[159]},
      {stage1_33[87]}
   );
   gpc1_1 gpc1502 (
      {stage0_33[160]},
      {stage1_33[88]}
   );
   gpc1_1 gpc1503 (
      {stage0_33[161]},
      {stage1_33[89]}
   );
   gpc1_1 gpc1504 (
      {stage0_34[158]},
      {stage1_34[52]}
   );
   gpc1_1 gpc1505 (
      {stage0_34[159]},
      {stage1_34[53]}
   );
   gpc1_1 gpc1506 (
      {stage0_34[160]},
      {stage1_34[54]}
   );
   gpc1_1 gpc1507 (
      {stage0_34[161]},
      {stage1_34[55]}
   );
   gpc1_1 gpc1508 (
      {stage0_35[158]},
      {stage1_35[56]}
   );
   gpc1_1 gpc1509 (
      {stage0_35[159]},
      {stage1_35[57]}
   );
   gpc1_1 gpc1510 (
      {stage0_35[160]},
      {stage1_35[58]}
   );
   gpc1_1 gpc1511 (
      {stage0_35[161]},
      {stage1_35[59]}
   );
   gpc1_1 gpc1512 (
      {stage0_36[146]},
      {stage1_36[67]}
   );
   gpc1_1 gpc1513 (
      {stage0_36[147]},
      {stage1_36[68]}
   );
   gpc1_1 gpc1514 (
      {stage0_36[148]},
      {stage1_36[69]}
   );
   gpc1_1 gpc1515 (
      {stage0_36[149]},
      {stage1_36[70]}
   );
   gpc1_1 gpc1516 (
      {stage0_36[150]},
      {stage1_36[71]}
   );
   gpc1_1 gpc1517 (
      {stage0_36[151]},
      {stage1_36[72]}
   );
   gpc1_1 gpc1518 (
      {stage0_36[152]},
      {stage1_36[73]}
   );
   gpc1_1 gpc1519 (
      {stage0_36[153]},
      {stage1_36[74]}
   );
   gpc1_1 gpc1520 (
      {stage0_36[154]},
      {stage1_36[75]}
   );
   gpc1_1 gpc1521 (
      {stage0_36[155]},
      {stage1_36[76]}
   );
   gpc1_1 gpc1522 (
      {stage0_36[156]},
      {stage1_36[77]}
   );
   gpc1_1 gpc1523 (
      {stage0_36[157]},
      {stage1_36[78]}
   );
   gpc1_1 gpc1524 (
      {stage0_36[158]},
      {stage1_36[79]}
   );
   gpc1_1 gpc1525 (
      {stage0_36[159]},
      {stage1_36[80]}
   );
   gpc1_1 gpc1526 (
      {stage0_36[160]},
      {stage1_36[81]}
   );
   gpc1_1 gpc1527 (
      {stage0_36[161]},
      {stage1_36[82]}
   );
   gpc1_1 gpc1528 (
      {stage0_37[90]},
      {stage1_37[56]}
   );
   gpc1_1 gpc1529 (
      {stage0_37[91]},
      {stage1_37[57]}
   );
   gpc1_1 gpc1530 (
      {stage0_37[92]},
      {stage1_37[58]}
   );
   gpc1_1 gpc1531 (
      {stage0_37[93]},
      {stage1_37[59]}
   );
   gpc1_1 gpc1532 (
      {stage0_37[94]},
      {stage1_37[60]}
   );
   gpc1_1 gpc1533 (
      {stage0_37[95]},
      {stage1_37[61]}
   );
   gpc1_1 gpc1534 (
      {stage0_37[96]},
      {stage1_37[62]}
   );
   gpc1_1 gpc1535 (
      {stage0_37[97]},
      {stage1_37[63]}
   );
   gpc1_1 gpc1536 (
      {stage0_37[98]},
      {stage1_37[64]}
   );
   gpc1_1 gpc1537 (
      {stage0_37[99]},
      {stage1_37[65]}
   );
   gpc1_1 gpc1538 (
      {stage0_37[100]},
      {stage1_37[66]}
   );
   gpc1_1 gpc1539 (
      {stage0_37[101]},
      {stage1_37[67]}
   );
   gpc1_1 gpc1540 (
      {stage0_37[102]},
      {stage1_37[68]}
   );
   gpc1_1 gpc1541 (
      {stage0_37[103]},
      {stage1_37[69]}
   );
   gpc1_1 gpc1542 (
      {stage0_37[104]},
      {stage1_37[70]}
   );
   gpc1_1 gpc1543 (
      {stage0_37[105]},
      {stage1_37[71]}
   );
   gpc1_1 gpc1544 (
      {stage0_37[106]},
      {stage1_37[72]}
   );
   gpc1_1 gpc1545 (
      {stage0_37[107]},
      {stage1_37[73]}
   );
   gpc1_1 gpc1546 (
      {stage0_37[108]},
      {stage1_37[74]}
   );
   gpc1_1 gpc1547 (
      {stage0_37[109]},
      {stage1_37[75]}
   );
   gpc1_1 gpc1548 (
      {stage0_37[110]},
      {stage1_37[76]}
   );
   gpc1_1 gpc1549 (
      {stage0_37[111]},
      {stage1_37[77]}
   );
   gpc1_1 gpc1550 (
      {stage0_37[112]},
      {stage1_37[78]}
   );
   gpc1_1 gpc1551 (
      {stage0_37[113]},
      {stage1_37[79]}
   );
   gpc1_1 gpc1552 (
      {stage0_37[114]},
      {stage1_37[80]}
   );
   gpc1_1 gpc1553 (
      {stage0_37[115]},
      {stage1_37[81]}
   );
   gpc1_1 gpc1554 (
      {stage0_37[116]},
      {stage1_37[82]}
   );
   gpc1_1 gpc1555 (
      {stage0_37[117]},
      {stage1_37[83]}
   );
   gpc1_1 gpc1556 (
      {stage0_37[118]},
      {stage1_37[84]}
   );
   gpc1_1 gpc1557 (
      {stage0_37[119]},
      {stage1_37[85]}
   );
   gpc1_1 gpc1558 (
      {stage0_37[120]},
      {stage1_37[86]}
   );
   gpc1_1 gpc1559 (
      {stage0_37[121]},
      {stage1_37[87]}
   );
   gpc1_1 gpc1560 (
      {stage0_37[122]},
      {stage1_37[88]}
   );
   gpc1_1 gpc1561 (
      {stage0_37[123]},
      {stage1_37[89]}
   );
   gpc1_1 gpc1562 (
      {stage0_37[124]},
      {stage1_37[90]}
   );
   gpc1_1 gpc1563 (
      {stage0_37[125]},
      {stage1_37[91]}
   );
   gpc1_1 gpc1564 (
      {stage0_37[126]},
      {stage1_37[92]}
   );
   gpc1_1 gpc1565 (
      {stage0_37[127]},
      {stage1_37[93]}
   );
   gpc1_1 gpc1566 (
      {stage0_37[128]},
      {stage1_37[94]}
   );
   gpc1_1 gpc1567 (
      {stage0_37[129]},
      {stage1_37[95]}
   );
   gpc1_1 gpc1568 (
      {stage0_37[130]},
      {stage1_37[96]}
   );
   gpc1_1 gpc1569 (
      {stage0_37[131]},
      {stage1_37[97]}
   );
   gpc1_1 gpc1570 (
      {stage0_37[132]},
      {stage1_37[98]}
   );
   gpc1_1 gpc1571 (
      {stage0_37[133]},
      {stage1_37[99]}
   );
   gpc1_1 gpc1572 (
      {stage0_37[134]},
      {stage1_37[100]}
   );
   gpc1_1 gpc1573 (
      {stage0_37[135]},
      {stage1_37[101]}
   );
   gpc1_1 gpc1574 (
      {stage0_37[136]},
      {stage1_37[102]}
   );
   gpc1_1 gpc1575 (
      {stage0_37[137]},
      {stage1_37[103]}
   );
   gpc1_1 gpc1576 (
      {stage0_37[138]},
      {stage1_37[104]}
   );
   gpc1_1 gpc1577 (
      {stage0_37[139]},
      {stage1_37[105]}
   );
   gpc1_1 gpc1578 (
      {stage0_37[140]},
      {stage1_37[106]}
   );
   gpc1_1 gpc1579 (
      {stage0_37[141]},
      {stage1_37[107]}
   );
   gpc1_1 gpc1580 (
      {stage0_37[142]},
      {stage1_37[108]}
   );
   gpc1_1 gpc1581 (
      {stage0_37[143]},
      {stage1_37[109]}
   );
   gpc1_1 gpc1582 (
      {stage0_37[144]},
      {stage1_37[110]}
   );
   gpc1_1 gpc1583 (
      {stage0_37[145]},
      {stage1_37[111]}
   );
   gpc1_1 gpc1584 (
      {stage0_37[146]},
      {stage1_37[112]}
   );
   gpc1_1 gpc1585 (
      {stage0_37[147]},
      {stage1_37[113]}
   );
   gpc1_1 gpc1586 (
      {stage0_37[148]},
      {stage1_37[114]}
   );
   gpc1_1 gpc1587 (
      {stage0_37[149]},
      {stage1_37[115]}
   );
   gpc1_1 gpc1588 (
      {stage0_37[150]},
      {stage1_37[116]}
   );
   gpc1_1 gpc1589 (
      {stage0_37[151]},
      {stage1_37[117]}
   );
   gpc1_1 gpc1590 (
      {stage0_37[152]},
      {stage1_37[118]}
   );
   gpc1_1 gpc1591 (
      {stage0_37[153]},
      {stage1_37[119]}
   );
   gpc1_1 gpc1592 (
      {stage0_37[154]},
      {stage1_37[120]}
   );
   gpc1_1 gpc1593 (
      {stage0_37[155]},
      {stage1_37[121]}
   );
   gpc1_1 gpc1594 (
      {stage0_37[156]},
      {stage1_37[122]}
   );
   gpc1_1 gpc1595 (
      {stage0_37[157]},
      {stage1_37[123]}
   );
   gpc1_1 gpc1596 (
      {stage0_37[158]},
      {stage1_37[124]}
   );
   gpc1_1 gpc1597 (
      {stage0_37[159]},
      {stage1_37[125]}
   );
   gpc1_1 gpc1598 (
      {stage0_37[160]},
      {stage1_37[126]}
   );
   gpc1_1 gpc1599 (
      {stage0_37[161]},
      {stage1_37[127]}
   );
   gpc1_1 gpc1600 (
      {stage0_38[148]},
      {stage1_38[52]}
   );
   gpc1_1 gpc1601 (
      {stage0_38[149]},
      {stage1_38[53]}
   );
   gpc1_1 gpc1602 (
      {stage0_38[150]},
      {stage1_38[54]}
   );
   gpc1_1 gpc1603 (
      {stage0_38[151]},
      {stage1_38[55]}
   );
   gpc1_1 gpc1604 (
      {stage0_38[152]},
      {stage1_38[56]}
   );
   gpc1_1 gpc1605 (
      {stage0_38[153]},
      {stage1_38[57]}
   );
   gpc1_1 gpc1606 (
      {stage0_38[154]},
      {stage1_38[58]}
   );
   gpc1_1 gpc1607 (
      {stage0_38[155]},
      {stage1_38[59]}
   );
   gpc1_1 gpc1608 (
      {stage0_38[156]},
      {stage1_38[60]}
   );
   gpc1_1 gpc1609 (
      {stage0_38[157]},
      {stage1_38[61]}
   );
   gpc1_1 gpc1610 (
      {stage0_38[158]},
      {stage1_38[62]}
   );
   gpc1_1 gpc1611 (
      {stage0_38[159]},
      {stage1_38[63]}
   );
   gpc1_1 gpc1612 (
      {stage0_38[160]},
      {stage1_38[64]}
   );
   gpc1_1 gpc1613 (
      {stage0_38[161]},
      {stage1_38[65]}
   );
   gpc1_1 gpc1614 (
      {stage0_39[156]},
      {stage1_39[62]}
   );
   gpc1_1 gpc1615 (
      {stage0_39[157]},
      {stage1_39[63]}
   );
   gpc1_1 gpc1616 (
      {stage0_39[158]},
      {stage1_39[64]}
   );
   gpc1_1 gpc1617 (
      {stage0_39[159]},
      {stage1_39[65]}
   );
   gpc1_1 gpc1618 (
      {stage0_39[160]},
      {stage1_39[66]}
   );
   gpc1_1 gpc1619 (
      {stage0_39[161]},
      {stage1_39[67]}
   );
   gpc1_1 gpc1620 (
      {stage0_40[140]},
      {stage1_40[60]}
   );
   gpc1_1 gpc1621 (
      {stage0_40[141]},
      {stage1_40[61]}
   );
   gpc1_1 gpc1622 (
      {stage0_40[142]},
      {stage1_40[62]}
   );
   gpc1_1 gpc1623 (
      {stage0_40[143]},
      {stage1_40[63]}
   );
   gpc1_1 gpc1624 (
      {stage0_40[144]},
      {stage1_40[64]}
   );
   gpc1_1 gpc1625 (
      {stage0_40[145]},
      {stage1_40[65]}
   );
   gpc1_1 gpc1626 (
      {stage0_40[146]},
      {stage1_40[66]}
   );
   gpc1_1 gpc1627 (
      {stage0_40[147]},
      {stage1_40[67]}
   );
   gpc1_1 gpc1628 (
      {stage0_40[148]},
      {stage1_40[68]}
   );
   gpc1_1 gpc1629 (
      {stage0_40[149]},
      {stage1_40[69]}
   );
   gpc1_1 gpc1630 (
      {stage0_40[150]},
      {stage1_40[70]}
   );
   gpc1_1 gpc1631 (
      {stage0_40[151]},
      {stage1_40[71]}
   );
   gpc1_1 gpc1632 (
      {stage0_40[152]},
      {stage1_40[72]}
   );
   gpc1_1 gpc1633 (
      {stage0_40[153]},
      {stage1_40[73]}
   );
   gpc1_1 gpc1634 (
      {stage0_40[154]},
      {stage1_40[74]}
   );
   gpc1_1 gpc1635 (
      {stage0_40[155]},
      {stage1_40[75]}
   );
   gpc1_1 gpc1636 (
      {stage0_40[156]},
      {stage1_40[76]}
   );
   gpc1_1 gpc1637 (
      {stage0_40[157]},
      {stage1_40[77]}
   );
   gpc1_1 gpc1638 (
      {stage0_40[158]},
      {stage1_40[78]}
   );
   gpc1_1 gpc1639 (
      {stage0_40[159]},
      {stage1_40[79]}
   );
   gpc1_1 gpc1640 (
      {stage0_40[160]},
      {stage1_40[80]}
   );
   gpc1_1 gpc1641 (
      {stage0_40[161]},
      {stage1_40[81]}
   );
   gpc1_1 gpc1642 (
      {stage0_41[138]},
      {stage1_41[50]}
   );
   gpc1_1 gpc1643 (
      {stage0_41[139]},
      {stage1_41[51]}
   );
   gpc1_1 gpc1644 (
      {stage0_41[140]},
      {stage1_41[52]}
   );
   gpc1_1 gpc1645 (
      {stage0_41[141]},
      {stage1_41[53]}
   );
   gpc1_1 gpc1646 (
      {stage0_41[142]},
      {stage1_41[54]}
   );
   gpc1_1 gpc1647 (
      {stage0_41[143]},
      {stage1_41[55]}
   );
   gpc1_1 gpc1648 (
      {stage0_41[144]},
      {stage1_41[56]}
   );
   gpc1_1 gpc1649 (
      {stage0_41[145]},
      {stage1_41[57]}
   );
   gpc1_1 gpc1650 (
      {stage0_41[146]},
      {stage1_41[58]}
   );
   gpc1_1 gpc1651 (
      {stage0_41[147]},
      {stage1_41[59]}
   );
   gpc1_1 gpc1652 (
      {stage0_41[148]},
      {stage1_41[60]}
   );
   gpc1_1 gpc1653 (
      {stage0_41[149]},
      {stage1_41[61]}
   );
   gpc1_1 gpc1654 (
      {stage0_41[150]},
      {stage1_41[62]}
   );
   gpc1_1 gpc1655 (
      {stage0_41[151]},
      {stage1_41[63]}
   );
   gpc1_1 gpc1656 (
      {stage0_41[152]},
      {stage1_41[64]}
   );
   gpc1_1 gpc1657 (
      {stage0_41[153]},
      {stage1_41[65]}
   );
   gpc1_1 gpc1658 (
      {stage0_41[154]},
      {stage1_41[66]}
   );
   gpc1_1 gpc1659 (
      {stage0_41[155]},
      {stage1_41[67]}
   );
   gpc1_1 gpc1660 (
      {stage0_41[156]},
      {stage1_41[68]}
   );
   gpc1_1 gpc1661 (
      {stage0_41[157]},
      {stage1_41[69]}
   );
   gpc1_1 gpc1662 (
      {stage0_41[158]},
      {stage1_41[70]}
   );
   gpc1_1 gpc1663 (
      {stage0_41[159]},
      {stage1_41[71]}
   );
   gpc1_1 gpc1664 (
      {stage0_41[160]},
      {stage1_41[72]}
   );
   gpc1_1 gpc1665 (
      {stage0_41[161]},
      {stage1_41[73]}
   );
   gpc1_1 gpc1666 (
      {stage0_42[126]},
      {stage1_42[60]}
   );
   gpc1_1 gpc1667 (
      {stage0_42[127]},
      {stage1_42[61]}
   );
   gpc1_1 gpc1668 (
      {stage0_42[128]},
      {stage1_42[62]}
   );
   gpc1_1 gpc1669 (
      {stage0_42[129]},
      {stage1_42[63]}
   );
   gpc1_1 gpc1670 (
      {stage0_42[130]},
      {stage1_42[64]}
   );
   gpc1_1 gpc1671 (
      {stage0_42[131]},
      {stage1_42[65]}
   );
   gpc1_1 gpc1672 (
      {stage0_42[132]},
      {stage1_42[66]}
   );
   gpc1_1 gpc1673 (
      {stage0_42[133]},
      {stage1_42[67]}
   );
   gpc1_1 gpc1674 (
      {stage0_42[134]},
      {stage1_42[68]}
   );
   gpc1_1 gpc1675 (
      {stage0_42[135]},
      {stage1_42[69]}
   );
   gpc1_1 gpc1676 (
      {stage0_42[136]},
      {stage1_42[70]}
   );
   gpc1_1 gpc1677 (
      {stage0_42[137]},
      {stage1_42[71]}
   );
   gpc1_1 gpc1678 (
      {stage0_42[138]},
      {stage1_42[72]}
   );
   gpc1_1 gpc1679 (
      {stage0_42[139]},
      {stage1_42[73]}
   );
   gpc1_1 gpc1680 (
      {stage0_42[140]},
      {stage1_42[74]}
   );
   gpc1_1 gpc1681 (
      {stage0_42[141]},
      {stage1_42[75]}
   );
   gpc1_1 gpc1682 (
      {stage0_42[142]},
      {stage1_42[76]}
   );
   gpc1_1 gpc1683 (
      {stage0_42[143]},
      {stage1_42[77]}
   );
   gpc1_1 gpc1684 (
      {stage0_42[144]},
      {stage1_42[78]}
   );
   gpc1_1 gpc1685 (
      {stage0_42[145]},
      {stage1_42[79]}
   );
   gpc1_1 gpc1686 (
      {stage0_42[146]},
      {stage1_42[80]}
   );
   gpc1_1 gpc1687 (
      {stage0_42[147]},
      {stage1_42[81]}
   );
   gpc1_1 gpc1688 (
      {stage0_42[148]},
      {stage1_42[82]}
   );
   gpc1_1 gpc1689 (
      {stage0_42[149]},
      {stage1_42[83]}
   );
   gpc1_1 gpc1690 (
      {stage0_42[150]},
      {stage1_42[84]}
   );
   gpc1_1 gpc1691 (
      {stage0_42[151]},
      {stage1_42[85]}
   );
   gpc1_1 gpc1692 (
      {stage0_42[152]},
      {stage1_42[86]}
   );
   gpc1_1 gpc1693 (
      {stage0_42[153]},
      {stage1_42[87]}
   );
   gpc1_1 gpc1694 (
      {stage0_42[154]},
      {stage1_42[88]}
   );
   gpc1_1 gpc1695 (
      {stage0_42[155]},
      {stage1_42[89]}
   );
   gpc1_1 gpc1696 (
      {stage0_42[156]},
      {stage1_42[90]}
   );
   gpc1_1 gpc1697 (
      {stage0_42[157]},
      {stage1_42[91]}
   );
   gpc1_1 gpc1698 (
      {stage0_42[158]},
      {stage1_42[92]}
   );
   gpc1_1 gpc1699 (
      {stage0_42[159]},
      {stage1_42[93]}
   );
   gpc1_1 gpc1700 (
      {stage0_42[160]},
      {stage1_42[94]}
   );
   gpc1_1 gpc1701 (
      {stage0_42[161]},
      {stage1_42[95]}
   );
   gpc1_1 gpc1702 (
      {stage0_43[78]},
      {stage1_43[54]}
   );
   gpc1_1 gpc1703 (
      {stage0_43[79]},
      {stage1_43[55]}
   );
   gpc1_1 gpc1704 (
      {stage0_43[80]},
      {stage1_43[56]}
   );
   gpc1_1 gpc1705 (
      {stage0_43[81]},
      {stage1_43[57]}
   );
   gpc1_1 gpc1706 (
      {stage0_43[82]},
      {stage1_43[58]}
   );
   gpc1_1 gpc1707 (
      {stage0_43[83]},
      {stage1_43[59]}
   );
   gpc1_1 gpc1708 (
      {stage0_43[84]},
      {stage1_43[60]}
   );
   gpc1_1 gpc1709 (
      {stage0_43[85]},
      {stage1_43[61]}
   );
   gpc1_1 gpc1710 (
      {stage0_43[86]},
      {stage1_43[62]}
   );
   gpc1_1 gpc1711 (
      {stage0_43[87]},
      {stage1_43[63]}
   );
   gpc1_1 gpc1712 (
      {stage0_43[88]},
      {stage1_43[64]}
   );
   gpc1_1 gpc1713 (
      {stage0_43[89]},
      {stage1_43[65]}
   );
   gpc1_1 gpc1714 (
      {stage0_43[90]},
      {stage1_43[66]}
   );
   gpc1_1 gpc1715 (
      {stage0_43[91]},
      {stage1_43[67]}
   );
   gpc1_1 gpc1716 (
      {stage0_43[92]},
      {stage1_43[68]}
   );
   gpc1_1 gpc1717 (
      {stage0_43[93]},
      {stage1_43[69]}
   );
   gpc1_1 gpc1718 (
      {stage0_43[94]},
      {stage1_43[70]}
   );
   gpc1_1 gpc1719 (
      {stage0_43[95]},
      {stage1_43[71]}
   );
   gpc1_1 gpc1720 (
      {stage0_43[96]},
      {stage1_43[72]}
   );
   gpc1_1 gpc1721 (
      {stage0_43[97]},
      {stage1_43[73]}
   );
   gpc1_1 gpc1722 (
      {stage0_43[98]},
      {stage1_43[74]}
   );
   gpc1_1 gpc1723 (
      {stage0_43[99]},
      {stage1_43[75]}
   );
   gpc1_1 gpc1724 (
      {stage0_43[100]},
      {stage1_43[76]}
   );
   gpc1_1 gpc1725 (
      {stage0_43[101]},
      {stage1_43[77]}
   );
   gpc1_1 gpc1726 (
      {stage0_43[102]},
      {stage1_43[78]}
   );
   gpc1_1 gpc1727 (
      {stage0_43[103]},
      {stage1_43[79]}
   );
   gpc1_1 gpc1728 (
      {stage0_43[104]},
      {stage1_43[80]}
   );
   gpc1_1 gpc1729 (
      {stage0_43[105]},
      {stage1_43[81]}
   );
   gpc1_1 gpc1730 (
      {stage0_43[106]},
      {stage1_43[82]}
   );
   gpc1_1 gpc1731 (
      {stage0_43[107]},
      {stage1_43[83]}
   );
   gpc1_1 gpc1732 (
      {stage0_43[108]},
      {stage1_43[84]}
   );
   gpc1_1 gpc1733 (
      {stage0_43[109]},
      {stage1_43[85]}
   );
   gpc1_1 gpc1734 (
      {stage0_43[110]},
      {stage1_43[86]}
   );
   gpc1_1 gpc1735 (
      {stage0_43[111]},
      {stage1_43[87]}
   );
   gpc1_1 gpc1736 (
      {stage0_43[112]},
      {stage1_43[88]}
   );
   gpc1_1 gpc1737 (
      {stage0_43[113]},
      {stage1_43[89]}
   );
   gpc1_1 gpc1738 (
      {stage0_43[114]},
      {stage1_43[90]}
   );
   gpc1_1 gpc1739 (
      {stage0_43[115]},
      {stage1_43[91]}
   );
   gpc1_1 gpc1740 (
      {stage0_43[116]},
      {stage1_43[92]}
   );
   gpc1_1 gpc1741 (
      {stage0_43[117]},
      {stage1_43[93]}
   );
   gpc1_1 gpc1742 (
      {stage0_43[118]},
      {stage1_43[94]}
   );
   gpc1_1 gpc1743 (
      {stage0_43[119]},
      {stage1_43[95]}
   );
   gpc1_1 gpc1744 (
      {stage0_43[120]},
      {stage1_43[96]}
   );
   gpc1_1 gpc1745 (
      {stage0_43[121]},
      {stage1_43[97]}
   );
   gpc1_1 gpc1746 (
      {stage0_43[122]},
      {stage1_43[98]}
   );
   gpc1_1 gpc1747 (
      {stage0_43[123]},
      {stage1_43[99]}
   );
   gpc1_1 gpc1748 (
      {stage0_43[124]},
      {stage1_43[100]}
   );
   gpc1_1 gpc1749 (
      {stage0_43[125]},
      {stage1_43[101]}
   );
   gpc1_1 gpc1750 (
      {stage0_43[126]},
      {stage1_43[102]}
   );
   gpc1_1 gpc1751 (
      {stage0_43[127]},
      {stage1_43[103]}
   );
   gpc1_1 gpc1752 (
      {stage0_43[128]},
      {stage1_43[104]}
   );
   gpc1_1 gpc1753 (
      {stage0_43[129]},
      {stage1_43[105]}
   );
   gpc1_1 gpc1754 (
      {stage0_43[130]},
      {stage1_43[106]}
   );
   gpc1_1 gpc1755 (
      {stage0_43[131]},
      {stage1_43[107]}
   );
   gpc1_1 gpc1756 (
      {stage0_43[132]},
      {stage1_43[108]}
   );
   gpc1_1 gpc1757 (
      {stage0_43[133]},
      {stage1_43[109]}
   );
   gpc1_1 gpc1758 (
      {stage0_43[134]},
      {stage1_43[110]}
   );
   gpc1_1 gpc1759 (
      {stage0_43[135]},
      {stage1_43[111]}
   );
   gpc1_1 gpc1760 (
      {stage0_43[136]},
      {stage1_43[112]}
   );
   gpc1_1 gpc1761 (
      {stage0_43[137]},
      {stage1_43[113]}
   );
   gpc1_1 gpc1762 (
      {stage0_43[138]},
      {stage1_43[114]}
   );
   gpc1_1 gpc1763 (
      {stage0_43[139]},
      {stage1_43[115]}
   );
   gpc1_1 gpc1764 (
      {stage0_43[140]},
      {stage1_43[116]}
   );
   gpc1_1 gpc1765 (
      {stage0_43[141]},
      {stage1_43[117]}
   );
   gpc1_1 gpc1766 (
      {stage0_43[142]},
      {stage1_43[118]}
   );
   gpc1_1 gpc1767 (
      {stage0_43[143]},
      {stage1_43[119]}
   );
   gpc1_1 gpc1768 (
      {stage0_43[144]},
      {stage1_43[120]}
   );
   gpc1_1 gpc1769 (
      {stage0_43[145]},
      {stage1_43[121]}
   );
   gpc1_1 gpc1770 (
      {stage0_43[146]},
      {stage1_43[122]}
   );
   gpc1_1 gpc1771 (
      {stage0_43[147]},
      {stage1_43[123]}
   );
   gpc1_1 gpc1772 (
      {stage0_43[148]},
      {stage1_43[124]}
   );
   gpc1_1 gpc1773 (
      {stage0_43[149]},
      {stage1_43[125]}
   );
   gpc1_1 gpc1774 (
      {stage0_43[150]},
      {stage1_43[126]}
   );
   gpc1_1 gpc1775 (
      {stage0_43[151]},
      {stage1_43[127]}
   );
   gpc1_1 gpc1776 (
      {stage0_43[152]},
      {stage1_43[128]}
   );
   gpc1_1 gpc1777 (
      {stage0_43[153]},
      {stage1_43[129]}
   );
   gpc1_1 gpc1778 (
      {stage0_43[154]},
      {stage1_43[130]}
   );
   gpc1_1 gpc1779 (
      {stage0_43[155]},
      {stage1_43[131]}
   );
   gpc1_1 gpc1780 (
      {stage0_43[156]},
      {stage1_43[132]}
   );
   gpc1_1 gpc1781 (
      {stage0_43[157]},
      {stage1_43[133]}
   );
   gpc1_1 gpc1782 (
      {stage0_43[158]},
      {stage1_43[134]}
   );
   gpc1_1 gpc1783 (
      {stage0_43[159]},
      {stage1_43[135]}
   );
   gpc1_1 gpc1784 (
      {stage0_43[160]},
      {stage1_43[136]}
   );
   gpc1_1 gpc1785 (
      {stage0_43[161]},
      {stage1_43[137]}
   );
   gpc1_1 gpc1786 (
      {stage0_44[160]},
      {stage1_44[44]}
   );
   gpc1_1 gpc1787 (
      {stage0_44[161]},
      {stage1_44[45]}
   );
   gpc1_1 gpc1788 (
      {stage0_45[121]},
      {stage1_45[52]}
   );
   gpc1_1 gpc1789 (
      {stage0_45[122]},
      {stage1_45[53]}
   );
   gpc1_1 gpc1790 (
      {stage0_45[123]},
      {stage1_45[54]}
   );
   gpc1_1 gpc1791 (
      {stage0_45[124]},
      {stage1_45[55]}
   );
   gpc1_1 gpc1792 (
      {stage0_45[125]},
      {stage1_45[56]}
   );
   gpc1_1 gpc1793 (
      {stage0_45[126]},
      {stage1_45[57]}
   );
   gpc1_1 gpc1794 (
      {stage0_45[127]},
      {stage1_45[58]}
   );
   gpc1_1 gpc1795 (
      {stage0_45[128]},
      {stage1_45[59]}
   );
   gpc1_1 gpc1796 (
      {stage0_45[129]},
      {stage1_45[60]}
   );
   gpc1_1 gpc1797 (
      {stage0_45[130]},
      {stage1_45[61]}
   );
   gpc1_1 gpc1798 (
      {stage0_45[131]},
      {stage1_45[62]}
   );
   gpc1_1 gpc1799 (
      {stage0_45[132]},
      {stage1_45[63]}
   );
   gpc1_1 gpc1800 (
      {stage0_45[133]},
      {stage1_45[64]}
   );
   gpc1_1 gpc1801 (
      {stage0_45[134]},
      {stage1_45[65]}
   );
   gpc1_1 gpc1802 (
      {stage0_45[135]},
      {stage1_45[66]}
   );
   gpc1_1 gpc1803 (
      {stage0_45[136]},
      {stage1_45[67]}
   );
   gpc1_1 gpc1804 (
      {stage0_45[137]},
      {stage1_45[68]}
   );
   gpc1_1 gpc1805 (
      {stage0_45[138]},
      {stage1_45[69]}
   );
   gpc1_1 gpc1806 (
      {stage0_45[139]},
      {stage1_45[70]}
   );
   gpc1_1 gpc1807 (
      {stage0_45[140]},
      {stage1_45[71]}
   );
   gpc1_1 gpc1808 (
      {stage0_45[141]},
      {stage1_45[72]}
   );
   gpc1_1 gpc1809 (
      {stage0_45[142]},
      {stage1_45[73]}
   );
   gpc1_1 gpc1810 (
      {stage0_45[143]},
      {stage1_45[74]}
   );
   gpc1_1 gpc1811 (
      {stage0_45[144]},
      {stage1_45[75]}
   );
   gpc1_1 gpc1812 (
      {stage0_45[145]},
      {stage1_45[76]}
   );
   gpc1_1 gpc1813 (
      {stage0_45[146]},
      {stage1_45[77]}
   );
   gpc1_1 gpc1814 (
      {stage0_45[147]},
      {stage1_45[78]}
   );
   gpc1_1 gpc1815 (
      {stage0_45[148]},
      {stage1_45[79]}
   );
   gpc1_1 gpc1816 (
      {stage0_45[149]},
      {stage1_45[80]}
   );
   gpc1_1 gpc1817 (
      {stage0_45[150]},
      {stage1_45[81]}
   );
   gpc1_1 gpc1818 (
      {stage0_45[151]},
      {stage1_45[82]}
   );
   gpc1_1 gpc1819 (
      {stage0_45[152]},
      {stage1_45[83]}
   );
   gpc1_1 gpc1820 (
      {stage0_45[153]},
      {stage1_45[84]}
   );
   gpc1_1 gpc1821 (
      {stage0_45[154]},
      {stage1_45[85]}
   );
   gpc1_1 gpc1822 (
      {stage0_45[155]},
      {stage1_45[86]}
   );
   gpc1_1 gpc1823 (
      {stage0_45[156]},
      {stage1_45[87]}
   );
   gpc1_1 gpc1824 (
      {stage0_45[157]},
      {stage1_45[88]}
   );
   gpc1_1 gpc1825 (
      {stage0_45[158]},
      {stage1_45[89]}
   );
   gpc1_1 gpc1826 (
      {stage0_45[159]},
      {stage1_45[90]}
   );
   gpc1_1 gpc1827 (
      {stage0_45[160]},
      {stage1_45[91]}
   );
   gpc1_1 gpc1828 (
      {stage0_45[161]},
      {stage1_45[92]}
   );
   gpc1_1 gpc1829 (
      {stage0_46[161]},
      {stage1_46[63]}
   );
   gpc1_1 gpc1830 (
      {stage0_48[161]},
      {stage1_48[71]}
   );
   gpc1_1 gpc1831 (
      {stage0_49[147]},
      {stage1_49[72]}
   );
   gpc1_1 gpc1832 (
      {stage0_49[148]},
      {stage1_49[73]}
   );
   gpc1_1 gpc1833 (
      {stage0_49[149]},
      {stage1_49[74]}
   );
   gpc1_1 gpc1834 (
      {stage0_49[150]},
      {stage1_49[75]}
   );
   gpc1_1 gpc1835 (
      {stage0_49[151]},
      {stage1_49[76]}
   );
   gpc1_1 gpc1836 (
      {stage0_49[152]},
      {stage1_49[77]}
   );
   gpc1_1 gpc1837 (
      {stage0_49[153]},
      {stage1_49[78]}
   );
   gpc1_1 gpc1838 (
      {stage0_49[154]},
      {stage1_49[79]}
   );
   gpc1_1 gpc1839 (
      {stage0_49[155]},
      {stage1_49[80]}
   );
   gpc1_1 gpc1840 (
      {stage0_49[156]},
      {stage1_49[81]}
   );
   gpc1_1 gpc1841 (
      {stage0_49[157]},
      {stage1_49[82]}
   );
   gpc1_1 gpc1842 (
      {stage0_49[158]},
      {stage1_49[83]}
   );
   gpc1_1 gpc1843 (
      {stage0_49[159]},
      {stage1_49[84]}
   );
   gpc1_1 gpc1844 (
      {stage0_49[160]},
      {stage1_49[85]}
   );
   gpc1_1 gpc1845 (
      {stage0_49[161]},
      {stage1_49[86]}
   );
   gpc1_1 gpc1846 (
      {stage0_50[159]},
      {stage1_50[55]}
   );
   gpc1_1 gpc1847 (
      {stage0_50[160]},
      {stage1_50[56]}
   );
   gpc1_1 gpc1848 (
      {stage0_50[161]},
      {stage1_50[57]}
   );
   gpc1_1 gpc1849 (
      {stage0_51[126]},
      {stage1_51[58]}
   );
   gpc1_1 gpc1850 (
      {stage0_51[127]},
      {stage1_51[59]}
   );
   gpc1_1 gpc1851 (
      {stage0_51[128]},
      {stage1_51[60]}
   );
   gpc1_1 gpc1852 (
      {stage0_51[129]},
      {stage1_51[61]}
   );
   gpc1_1 gpc1853 (
      {stage0_51[130]},
      {stage1_51[62]}
   );
   gpc1_1 gpc1854 (
      {stage0_51[131]},
      {stage1_51[63]}
   );
   gpc1_1 gpc1855 (
      {stage0_51[132]},
      {stage1_51[64]}
   );
   gpc1_1 gpc1856 (
      {stage0_51[133]},
      {stage1_51[65]}
   );
   gpc1_1 gpc1857 (
      {stage0_51[134]},
      {stage1_51[66]}
   );
   gpc1_1 gpc1858 (
      {stage0_51[135]},
      {stage1_51[67]}
   );
   gpc1_1 gpc1859 (
      {stage0_51[136]},
      {stage1_51[68]}
   );
   gpc1_1 gpc1860 (
      {stage0_51[137]},
      {stage1_51[69]}
   );
   gpc1_1 gpc1861 (
      {stage0_51[138]},
      {stage1_51[70]}
   );
   gpc1_1 gpc1862 (
      {stage0_51[139]},
      {stage1_51[71]}
   );
   gpc1_1 gpc1863 (
      {stage0_51[140]},
      {stage1_51[72]}
   );
   gpc1_1 gpc1864 (
      {stage0_51[141]},
      {stage1_51[73]}
   );
   gpc1_1 gpc1865 (
      {stage0_51[142]},
      {stage1_51[74]}
   );
   gpc1_1 gpc1866 (
      {stage0_51[143]},
      {stage1_51[75]}
   );
   gpc1_1 gpc1867 (
      {stage0_51[144]},
      {stage1_51[76]}
   );
   gpc1_1 gpc1868 (
      {stage0_51[145]},
      {stage1_51[77]}
   );
   gpc1_1 gpc1869 (
      {stage0_51[146]},
      {stage1_51[78]}
   );
   gpc1_1 gpc1870 (
      {stage0_51[147]},
      {stage1_51[79]}
   );
   gpc1_1 gpc1871 (
      {stage0_51[148]},
      {stage1_51[80]}
   );
   gpc1_1 gpc1872 (
      {stage0_51[149]},
      {stage1_51[81]}
   );
   gpc1_1 gpc1873 (
      {stage0_51[150]},
      {stage1_51[82]}
   );
   gpc1_1 gpc1874 (
      {stage0_51[151]},
      {stage1_51[83]}
   );
   gpc1_1 gpc1875 (
      {stage0_51[152]},
      {stage1_51[84]}
   );
   gpc1_1 gpc1876 (
      {stage0_51[153]},
      {stage1_51[85]}
   );
   gpc1_1 gpc1877 (
      {stage0_51[154]},
      {stage1_51[86]}
   );
   gpc1_1 gpc1878 (
      {stage0_51[155]},
      {stage1_51[87]}
   );
   gpc1_1 gpc1879 (
      {stage0_51[156]},
      {stage1_51[88]}
   );
   gpc1_1 gpc1880 (
      {stage0_51[157]},
      {stage1_51[89]}
   );
   gpc1_1 gpc1881 (
      {stage0_51[158]},
      {stage1_51[90]}
   );
   gpc1_1 gpc1882 (
      {stage0_51[159]},
      {stage1_51[91]}
   );
   gpc1_1 gpc1883 (
      {stage0_51[160]},
      {stage1_51[92]}
   );
   gpc1_1 gpc1884 (
      {stage0_51[161]},
      {stage1_51[93]}
   );
   gpc1_1 gpc1885 (
      {stage0_52[153]},
      {stage1_52[68]}
   );
   gpc1_1 gpc1886 (
      {stage0_52[154]},
      {stage1_52[69]}
   );
   gpc1_1 gpc1887 (
      {stage0_52[155]},
      {stage1_52[70]}
   );
   gpc1_1 gpc1888 (
      {stage0_52[156]},
      {stage1_52[71]}
   );
   gpc1_1 gpc1889 (
      {stage0_52[157]},
      {stage1_52[72]}
   );
   gpc1_1 gpc1890 (
      {stage0_52[158]},
      {stage1_52[73]}
   );
   gpc1_1 gpc1891 (
      {stage0_52[159]},
      {stage1_52[74]}
   );
   gpc1_1 gpc1892 (
      {stage0_52[160]},
      {stage1_52[75]}
   );
   gpc1_1 gpc1893 (
      {stage0_52[161]},
      {stage1_52[76]}
   );
   gpc1_1 gpc1894 (
      {stage0_53[159]},
      {stage1_53[63]}
   );
   gpc1_1 gpc1895 (
      {stage0_53[160]},
      {stage1_53[64]}
   );
   gpc1_1 gpc1896 (
      {stage0_53[161]},
      {stage1_53[65]}
   );
   gpc1_1 gpc1897 (
      {stage0_55[122]},
      {stage1_55[58]}
   );
   gpc1_1 gpc1898 (
      {stage0_55[123]},
      {stage1_55[59]}
   );
   gpc1_1 gpc1899 (
      {stage0_55[124]},
      {stage1_55[60]}
   );
   gpc1_1 gpc1900 (
      {stage0_55[125]},
      {stage1_55[61]}
   );
   gpc1_1 gpc1901 (
      {stage0_55[126]},
      {stage1_55[62]}
   );
   gpc1_1 gpc1902 (
      {stage0_55[127]},
      {stage1_55[63]}
   );
   gpc1_1 gpc1903 (
      {stage0_55[128]},
      {stage1_55[64]}
   );
   gpc1_1 gpc1904 (
      {stage0_55[129]},
      {stage1_55[65]}
   );
   gpc1_1 gpc1905 (
      {stage0_55[130]},
      {stage1_55[66]}
   );
   gpc1_1 gpc1906 (
      {stage0_55[131]},
      {stage1_55[67]}
   );
   gpc1_1 gpc1907 (
      {stage0_55[132]},
      {stage1_55[68]}
   );
   gpc1_1 gpc1908 (
      {stage0_55[133]},
      {stage1_55[69]}
   );
   gpc1_1 gpc1909 (
      {stage0_55[134]},
      {stage1_55[70]}
   );
   gpc1_1 gpc1910 (
      {stage0_55[135]},
      {stage1_55[71]}
   );
   gpc1_1 gpc1911 (
      {stage0_55[136]},
      {stage1_55[72]}
   );
   gpc1_1 gpc1912 (
      {stage0_55[137]},
      {stage1_55[73]}
   );
   gpc1_1 gpc1913 (
      {stage0_55[138]},
      {stage1_55[74]}
   );
   gpc1_1 gpc1914 (
      {stage0_55[139]},
      {stage1_55[75]}
   );
   gpc1_1 gpc1915 (
      {stage0_55[140]},
      {stage1_55[76]}
   );
   gpc1_1 gpc1916 (
      {stage0_55[141]},
      {stage1_55[77]}
   );
   gpc1_1 gpc1917 (
      {stage0_55[142]},
      {stage1_55[78]}
   );
   gpc1_1 gpc1918 (
      {stage0_55[143]},
      {stage1_55[79]}
   );
   gpc1_1 gpc1919 (
      {stage0_55[144]},
      {stage1_55[80]}
   );
   gpc1_1 gpc1920 (
      {stage0_55[145]},
      {stage1_55[81]}
   );
   gpc1_1 gpc1921 (
      {stage0_55[146]},
      {stage1_55[82]}
   );
   gpc1_1 gpc1922 (
      {stage0_55[147]},
      {stage1_55[83]}
   );
   gpc1_1 gpc1923 (
      {stage0_55[148]},
      {stage1_55[84]}
   );
   gpc1_1 gpc1924 (
      {stage0_55[149]},
      {stage1_55[85]}
   );
   gpc1_1 gpc1925 (
      {stage0_55[150]},
      {stage1_55[86]}
   );
   gpc1_1 gpc1926 (
      {stage0_55[151]},
      {stage1_55[87]}
   );
   gpc1_1 gpc1927 (
      {stage0_55[152]},
      {stage1_55[88]}
   );
   gpc1_1 gpc1928 (
      {stage0_55[153]},
      {stage1_55[89]}
   );
   gpc1_1 gpc1929 (
      {stage0_55[154]},
      {stage1_55[90]}
   );
   gpc1_1 gpc1930 (
      {stage0_55[155]},
      {stage1_55[91]}
   );
   gpc1_1 gpc1931 (
      {stage0_55[156]},
      {stage1_55[92]}
   );
   gpc1_1 gpc1932 (
      {stage0_55[157]},
      {stage1_55[93]}
   );
   gpc1_1 gpc1933 (
      {stage0_55[158]},
      {stage1_55[94]}
   );
   gpc1_1 gpc1934 (
      {stage0_55[159]},
      {stage1_55[95]}
   );
   gpc1_1 gpc1935 (
      {stage0_55[160]},
      {stage1_55[96]}
   );
   gpc1_1 gpc1936 (
      {stage0_55[161]},
      {stage1_55[97]}
   );
   gpc1_1 gpc1937 (
      {stage0_56[148]},
      {stage1_56[66]}
   );
   gpc1_1 gpc1938 (
      {stage0_56[149]},
      {stage1_56[67]}
   );
   gpc1_1 gpc1939 (
      {stage0_56[150]},
      {stage1_56[68]}
   );
   gpc1_1 gpc1940 (
      {stage0_56[151]},
      {stage1_56[69]}
   );
   gpc1_1 gpc1941 (
      {stage0_56[152]},
      {stage1_56[70]}
   );
   gpc1_1 gpc1942 (
      {stage0_56[153]},
      {stage1_56[71]}
   );
   gpc1_1 gpc1943 (
      {stage0_56[154]},
      {stage1_56[72]}
   );
   gpc1_1 gpc1944 (
      {stage0_56[155]},
      {stage1_56[73]}
   );
   gpc1_1 gpc1945 (
      {stage0_56[156]},
      {stage1_56[74]}
   );
   gpc1_1 gpc1946 (
      {stage0_56[157]},
      {stage1_56[75]}
   );
   gpc1_1 gpc1947 (
      {stage0_56[158]},
      {stage1_56[76]}
   );
   gpc1_1 gpc1948 (
      {stage0_56[159]},
      {stage1_56[77]}
   );
   gpc1_1 gpc1949 (
      {stage0_56[160]},
      {stage1_56[78]}
   );
   gpc1_1 gpc1950 (
      {stage0_56[161]},
      {stage1_56[79]}
   );
   gpc1_1 gpc1951 (
      {stage0_57[156]},
      {stage1_57[66]}
   );
   gpc1_1 gpc1952 (
      {stage0_57[157]},
      {stage1_57[67]}
   );
   gpc1_1 gpc1953 (
      {stage0_57[158]},
      {stage1_57[68]}
   );
   gpc1_1 gpc1954 (
      {stage0_57[159]},
      {stage1_57[69]}
   );
   gpc1_1 gpc1955 (
      {stage0_57[160]},
      {stage1_57[70]}
   );
   gpc1_1 gpc1956 (
      {stage0_57[161]},
      {stage1_57[71]}
   );
   gpc1_1 gpc1957 (
      {stage0_58[144]},
      {stage1_58[56]}
   );
   gpc1_1 gpc1958 (
      {stage0_58[145]},
      {stage1_58[57]}
   );
   gpc1_1 gpc1959 (
      {stage0_58[146]},
      {stage1_58[58]}
   );
   gpc1_1 gpc1960 (
      {stage0_58[147]},
      {stage1_58[59]}
   );
   gpc1_1 gpc1961 (
      {stage0_58[148]},
      {stage1_58[60]}
   );
   gpc1_1 gpc1962 (
      {stage0_58[149]},
      {stage1_58[61]}
   );
   gpc1_1 gpc1963 (
      {stage0_58[150]},
      {stage1_58[62]}
   );
   gpc1_1 gpc1964 (
      {stage0_58[151]},
      {stage1_58[63]}
   );
   gpc1_1 gpc1965 (
      {stage0_58[152]},
      {stage1_58[64]}
   );
   gpc1_1 gpc1966 (
      {stage0_58[153]},
      {stage1_58[65]}
   );
   gpc1_1 gpc1967 (
      {stage0_58[154]},
      {stage1_58[66]}
   );
   gpc1_1 gpc1968 (
      {stage0_58[155]},
      {stage1_58[67]}
   );
   gpc1_1 gpc1969 (
      {stage0_58[156]},
      {stage1_58[68]}
   );
   gpc1_1 gpc1970 (
      {stage0_58[157]},
      {stage1_58[69]}
   );
   gpc1_1 gpc1971 (
      {stage0_58[158]},
      {stage1_58[70]}
   );
   gpc1_1 gpc1972 (
      {stage0_58[159]},
      {stage1_58[71]}
   );
   gpc1_1 gpc1973 (
      {stage0_58[160]},
      {stage1_58[72]}
   );
   gpc1_1 gpc1974 (
      {stage0_58[161]},
      {stage1_58[73]}
   );
   gpc1_1 gpc1975 (
      {stage0_59[132]},
      {stage1_59[50]}
   );
   gpc1_1 gpc1976 (
      {stage0_59[133]},
      {stage1_59[51]}
   );
   gpc1_1 gpc1977 (
      {stage0_59[134]},
      {stage1_59[52]}
   );
   gpc1_1 gpc1978 (
      {stage0_59[135]},
      {stage1_59[53]}
   );
   gpc1_1 gpc1979 (
      {stage0_59[136]},
      {stage1_59[54]}
   );
   gpc1_1 gpc1980 (
      {stage0_59[137]},
      {stage1_59[55]}
   );
   gpc1_1 gpc1981 (
      {stage0_59[138]},
      {stage1_59[56]}
   );
   gpc1_1 gpc1982 (
      {stage0_59[139]},
      {stage1_59[57]}
   );
   gpc1_1 gpc1983 (
      {stage0_59[140]},
      {stage1_59[58]}
   );
   gpc1_1 gpc1984 (
      {stage0_59[141]},
      {stage1_59[59]}
   );
   gpc1_1 gpc1985 (
      {stage0_59[142]},
      {stage1_59[60]}
   );
   gpc1_1 gpc1986 (
      {stage0_59[143]},
      {stage1_59[61]}
   );
   gpc1_1 gpc1987 (
      {stage0_59[144]},
      {stage1_59[62]}
   );
   gpc1_1 gpc1988 (
      {stage0_59[145]},
      {stage1_59[63]}
   );
   gpc1_1 gpc1989 (
      {stage0_59[146]},
      {stage1_59[64]}
   );
   gpc1_1 gpc1990 (
      {stage0_59[147]},
      {stage1_59[65]}
   );
   gpc1_1 gpc1991 (
      {stage0_59[148]},
      {stage1_59[66]}
   );
   gpc1_1 gpc1992 (
      {stage0_59[149]},
      {stage1_59[67]}
   );
   gpc1_1 gpc1993 (
      {stage0_59[150]},
      {stage1_59[68]}
   );
   gpc1_1 gpc1994 (
      {stage0_59[151]},
      {stage1_59[69]}
   );
   gpc1_1 gpc1995 (
      {stage0_59[152]},
      {stage1_59[70]}
   );
   gpc1_1 gpc1996 (
      {stage0_59[153]},
      {stage1_59[71]}
   );
   gpc1_1 gpc1997 (
      {stage0_59[154]},
      {stage1_59[72]}
   );
   gpc1_1 gpc1998 (
      {stage0_59[155]},
      {stage1_59[73]}
   );
   gpc1_1 gpc1999 (
      {stage0_59[156]},
      {stage1_59[74]}
   );
   gpc1_1 gpc2000 (
      {stage0_59[157]},
      {stage1_59[75]}
   );
   gpc1_1 gpc2001 (
      {stage0_59[158]},
      {stage1_59[76]}
   );
   gpc1_1 gpc2002 (
      {stage0_59[159]},
      {stage1_59[77]}
   );
   gpc1_1 gpc2003 (
      {stage0_59[160]},
      {stage1_59[78]}
   );
   gpc1_1 gpc2004 (
      {stage0_59[161]},
      {stage1_59[79]}
   );
   gpc1_1 gpc2005 (
      {stage0_61[144]},
      {stage1_61[73]}
   );
   gpc1_1 gpc2006 (
      {stage0_61[145]},
      {stage1_61[74]}
   );
   gpc1_1 gpc2007 (
      {stage0_61[146]},
      {stage1_61[75]}
   );
   gpc1_1 gpc2008 (
      {stage0_61[147]},
      {stage1_61[76]}
   );
   gpc1_1 gpc2009 (
      {stage0_61[148]},
      {stage1_61[77]}
   );
   gpc1_1 gpc2010 (
      {stage0_61[149]},
      {stage1_61[78]}
   );
   gpc1_1 gpc2011 (
      {stage0_61[150]},
      {stage1_61[79]}
   );
   gpc1_1 gpc2012 (
      {stage0_61[151]},
      {stage1_61[80]}
   );
   gpc1_1 gpc2013 (
      {stage0_61[152]},
      {stage1_61[81]}
   );
   gpc1_1 gpc2014 (
      {stage0_61[153]},
      {stage1_61[82]}
   );
   gpc1_1 gpc2015 (
      {stage0_61[154]},
      {stage1_61[83]}
   );
   gpc1_1 gpc2016 (
      {stage0_61[155]},
      {stage1_61[84]}
   );
   gpc1_1 gpc2017 (
      {stage0_61[156]},
      {stage1_61[85]}
   );
   gpc1_1 gpc2018 (
      {stage0_61[157]},
      {stage1_61[86]}
   );
   gpc1_1 gpc2019 (
      {stage0_61[158]},
      {stage1_61[87]}
   );
   gpc1_1 gpc2020 (
      {stage0_61[159]},
      {stage1_61[88]}
   );
   gpc1_1 gpc2021 (
      {stage0_61[160]},
      {stage1_61[89]}
   );
   gpc1_1 gpc2022 (
      {stage0_61[161]},
      {stage1_61[90]}
   );
   gpc1_1 gpc2023 (
      {stage0_62[126]},
      {stage1_62[51]}
   );
   gpc1_1 gpc2024 (
      {stage0_62[127]},
      {stage1_62[52]}
   );
   gpc1_1 gpc2025 (
      {stage0_62[128]},
      {stage1_62[53]}
   );
   gpc1_1 gpc2026 (
      {stage0_62[129]},
      {stage1_62[54]}
   );
   gpc1_1 gpc2027 (
      {stage0_62[130]},
      {stage1_62[55]}
   );
   gpc1_1 gpc2028 (
      {stage0_62[131]},
      {stage1_62[56]}
   );
   gpc1_1 gpc2029 (
      {stage0_62[132]},
      {stage1_62[57]}
   );
   gpc1_1 gpc2030 (
      {stage0_62[133]},
      {stage1_62[58]}
   );
   gpc1_1 gpc2031 (
      {stage0_62[134]},
      {stage1_62[59]}
   );
   gpc1_1 gpc2032 (
      {stage0_62[135]},
      {stage1_62[60]}
   );
   gpc1_1 gpc2033 (
      {stage0_62[136]},
      {stage1_62[61]}
   );
   gpc1_1 gpc2034 (
      {stage0_62[137]},
      {stage1_62[62]}
   );
   gpc1_1 gpc2035 (
      {stage0_62[138]},
      {stage1_62[63]}
   );
   gpc1_1 gpc2036 (
      {stage0_62[139]},
      {stage1_62[64]}
   );
   gpc1_1 gpc2037 (
      {stage0_62[140]},
      {stage1_62[65]}
   );
   gpc1_1 gpc2038 (
      {stage0_62[141]},
      {stage1_62[66]}
   );
   gpc1_1 gpc2039 (
      {stage0_62[142]},
      {stage1_62[67]}
   );
   gpc1_1 gpc2040 (
      {stage0_62[143]},
      {stage1_62[68]}
   );
   gpc1_1 gpc2041 (
      {stage0_62[144]},
      {stage1_62[69]}
   );
   gpc1_1 gpc2042 (
      {stage0_62[145]},
      {stage1_62[70]}
   );
   gpc1_1 gpc2043 (
      {stage0_62[146]},
      {stage1_62[71]}
   );
   gpc1_1 gpc2044 (
      {stage0_62[147]},
      {stage1_62[72]}
   );
   gpc1_1 gpc2045 (
      {stage0_62[148]},
      {stage1_62[73]}
   );
   gpc1_1 gpc2046 (
      {stage0_62[149]},
      {stage1_62[74]}
   );
   gpc1_1 gpc2047 (
      {stage0_62[150]},
      {stage1_62[75]}
   );
   gpc1_1 gpc2048 (
      {stage0_62[151]},
      {stage1_62[76]}
   );
   gpc1_1 gpc2049 (
      {stage0_62[152]},
      {stage1_62[77]}
   );
   gpc1_1 gpc2050 (
      {stage0_62[153]},
      {stage1_62[78]}
   );
   gpc1_1 gpc2051 (
      {stage0_62[154]},
      {stage1_62[79]}
   );
   gpc1_1 gpc2052 (
      {stage0_62[155]},
      {stage1_62[80]}
   );
   gpc1_1 gpc2053 (
      {stage0_62[156]},
      {stage1_62[81]}
   );
   gpc1_1 gpc2054 (
      {stage0_62[157]},
      {stage1_62[82]}
   );
   gpc1_1 gpc2055 (
      {stage0_62[158]},
      {stage1_62[83]}
   );
   gpc1_1 gpc2056 (
      {stage0_62[159]},
      {stage1_62[84]}
   );
   gpc1_1 gpc2057 (
      {stage0_62[160]},
      {stage1_62[85]}
   );
   gpc1_1 gpc2058 (
      {stage0_62[161]},
      {stage1_62[86]}
   );
   gpc1_1 gpc2059 (
      {stage0_63[144]},
      {stage1_63[45]}
   );
   gpc1_1 gpc2060 (
      {stage0_63[145]},
      {stage1_63[46]}
   );
   gpc1_1 gpc2061 (
      {stage0_63[146]},
      {stage1_63[47]}
   );
   gpc1_1 gpc2062 (
      {stage0_63[147]},
      {stage1_63[48]}
   );
   gpc1_1 gpc2063 (
      {stage0_63[148]},
      {stage1_63[49]}
   );
   gpc1_1 gpc2064 (
      {stage0_63[149]},
      {stage1_63[50]}
   );
   gpc1_1 gpc2065 (
      {stage0_63[150]},
      {stage1_63[51]}
   );
   gpc1_1 gpc2066 (
      {stage0_63[151]},
      {stage1_63[52]}
   );
   gpc1_1 gpc2067 (
      {stage0_63[152]},
      {stage1_63[53]}
   );
   gpc1_1 gpc2068 (
      {stage0_63[153]},
      {stage1_63[54]}
   );
   gpc1_1 gpc2069 (
      {stage0_63[154]},
      {stage1_63[55]}
   );
   gpc1_1 gpc2070 (
      {stage0_63[155]},
      {stage1_63[56]}
   );
   gpc1_1 gpc2071 (
      {stage0_63[156]},
      {stage1_63[57]}
   );
   gpc1_1 gpc2072 (
      {stage0_63[157]},
      {stage1_63[58]}
   );
   gpc1_1 gpc2073 (
      {stage0_63[158]},
      {stage1_63[59]}
   );
   gpc1_1 gpc2074 (
      {stage0_63[159]},
      {stage1_63[60]}
   );
   gpc1_1 gpc2075 (
      {stage0_63[160]},
      {stage1_63[61]}
   );
   gpc1_1 gpc2076 (
      {stage0_63[161]},
      {stage1_63[62]}
   );
   gpc1163_5 gpc2077 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc2078 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc2079 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc2080 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc2081 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc2082 (
      {stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25]},
      {stage1_1[18]},
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc2083 (
      {stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29], stage1_0[30]},
      {stage1_1[19]},
      {stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc2084 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8]},
      {stage2_5[0],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc2085 (
      {stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31]},
      {stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage2_5[1],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc606_5 gpc2086 (
      {stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37]},
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20]},
      {stage2_5[2],stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9]}
   );
   gpc1163_5 gpc2087 (
      {stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_5[0]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[0],stage2_5[3],stage2_4[10],stage2_3[10]}
   );
   gpc615_5 gpc2088 (
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28]},
      {stage1_4[6]},
      {stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5], stage1_5[6]},
      {stage2_7[1],stage2_6[1],stage2_5[4],stage2_4[11],stage2_3[11]}
   );
   gpc615_5 gpc2089 (
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_4[7]},
      {stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12]},
      {stage2_7[2],stage2_6[2],stage2_5[5],stage2_4[12],stage2_3[12]}
   );
   gpc615_5 gpc2090 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[8]},
      {stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17], stage1_5[18]},
      {stage2_7[3],stage2_6[3],stage2_5[6],stage2_4[13],stage2_3[13]}
   );
   gpc615_5 gpc2091 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[9]},
      {stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23], stage1_5[24]},
      {stage2_7[4],stage2_6[4],stage2_5[7],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc2092 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[10]},
      {stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage2_7[5],stage2_6[5],stage2_5[8],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc2093 (
      {stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage1_4[11]},
      {stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage2_7[6],stage2_6[6],stage2_5[9],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc2094 (
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58]},
      {stage1_4[12]},
      {stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42]},
      {stage2_7[7],stage2_6[7],stage2_5[10],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc2095 (
      {stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63]},
      {stage1_4[13]},
      {stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48]},
      {stage2_7[8],stage2_6[8],stage2_5[11],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc2096 (
      {stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67], stage1_3[68]},
      {stage1_4[14]},
      {stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53], stage1_5[54]},
      {stage2_7[9],stage2_6[9],stage2_5[12],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc2097 (
      {stage1_3[69], stage1_3[70], stage1_3[71], stage1_3[72], stage1_3[73]},
      {stage1_4[15]},
      {stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59], stage1_5[60]},
      {stage2_7[10],stage2_6[10],stage2_5[13],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc2098 (
      {stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77], stage1_3[78]},
      {stage1_4[16]},
      {stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66]},
      {stage2_7[11],stage2_6[11],stage2_5[14],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc2099 (
      {stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage1_4[17]},
      {stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71], stage1_5[72]},
      {stage2_7[12],stage2_6[12],stage2_5[15],stage2_4[22],stage2_3[22]}
   );
   gpc606_5 gpc2100 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[0],stage2_7[13],stage2_6[13],stage2_5[16],stage2_4[23]}
   );
   gpc606_5 gpc2101 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[1],stage2_7[14],stage2_6[14],stage2_5[17],stage2_4[24]}
   );
   gpc606_5 gpc2102 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[2],stage2_7[15],stage2_6[15],stage2_5[18],stage2_4[25]}
   );
   gpc606_5 gpc2103 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[3],stage2_7[16],stage2_6[16],stage2_5[19],stage2_4[26]}
   );
   gpc606_5 gpc2104 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[4],stage2_7[17],stage2_6[17],stage2_5[20],stage2_4[27]}
   );
   gpc606_5 gpc2105 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[5],stage2_7[18],stage2_6[18],stage2_5[21],stage2_4[28]}
   );
   gpc606_5 gpc2106 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[6],stage2_7[19],stage2_6[19],stage2_5[22],stage2_4[29]}
   );
   gpc606_5 gpc2107 (
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[7],stage2_7[20],stage2_6[20],stage2_5[23],stage2_4[30]}
   );
   gpc606_5 gpc2108 (
      {stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[8],stage2_7[21],stage2_6[21],stage2_5[24]}
   );
   gpc606_5 gpc2109 (
      {stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[9],stage2_7[22],stage2_6[22],stage2_5[25]}
   );
   gpc606_5 gpc2110 (
      {stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[10],stage2_7[23],stage2_6[23],stage2_5[26]}
   );
   gpc606_5 gpc2111 (
      {stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[11],stage2_7[24],stage2_6[24],stage2_5[27]}
   );
   gpc606_5 gpc2112 (
      {stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[12],stage2_7[25],stage2_6[25],stage2_5[28]}
   );
   gpc606_5 gpc2113 (
      {stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107], stage1_5[108]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[13],stage2_7[26],stage2_6[26],stage2_5[29]}
   );
   gpc615_5 gpc2114 (
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage1_7[36]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[6],stage2_8[14],stage2_7[27],stage2_6[27]}
   );
   gpc615_5 gpc2115 (
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], 1'b0},
      {stage1_7[37]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[7],stage2_8[15],stage2_7[28],stage2_6[28]}
   );
   gpc606_5 gpc2116 (
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[8],stage2_8[16],stage2_7[29]}
   );
   gpc615_5 gpc2117 (
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage1_8[12]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[3],stage2_9[9],stage2_8[17],stage2_7[30]}
   );
   gpc615_5 gpc2118 (
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_8[13]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[4],stage2_9[10],stage2_8[18],stage2_7[31]}
   );
   gpc615_5 gpc2119 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58]},
      {stage1_8[14]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[5],stage2_9[11],stage2_8[19],stage2_7[32]}
   );
   gpc615_5 gpc2120 (
      {stage1_7[59], stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63]},
      {stage1_8[15]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[6],stage2_9[12],stage2_8[20],stage2_7[33]}
   );
   gpc606_5 gpc2121 (
      {stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[5],stage2_10[7],stage2_9[13],stage2_8[21]}
   );
   gpc606_5 gpc2122 (
      {stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[6],stage2_10[8],stage2_9[14],stage2_8[22]}
   );
   gpc606_5 gpc2123 (
      {stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[7],stage2_10[9],stage2_9[15],stage2_8[23]}
   );
   gpc606_5 gpc2124 (
      {stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[8],stage2_10[10],stage2_9[16],stage2_8[24]}
   );
   gpc606_5 gpc2125 (
      {stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[9],stage2_10[11],stage2_9[17],stage2_8[25]}
   );
   gpc606_5 gpc2126 (
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[5],stage2_11[10],stage2_10[12],stage2_9[18]}
   );
   gpc606_5 gpc2127 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[6],stage2_11[11],stage2_10[13],stage2_9[19]}
   );
   gpc606_5 gpc2128 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[7],stage2_11[12],stage2_10[14],stage2_9[20]}
   );
   gpc606_5 gpc2129 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[8],stage2_11[13],stage2_10[15],stage2_9[21]}
   );
   gpc606_5 gpc2130 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[4],stage2_12[9],stage2_11[14],stage2_10[16]}
   );
   gpc606_5 gpc2131 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[5],stage2_12[10],stage2_11[15],stage2_10[17]}
   );
   gpc606_5 gpc2132 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[6],stage2_12[11],stage2_11[16],stage2_10[18]}
   );
   gpc606_5 gpc2133 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[7],stage2_12[12],stage2_11[17],stage2_10[19]}
   );
   gpc615_5 gpc2134 (
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58]},
      {stage1_11[24]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[8],stage2_12[13],stage2_11[18],stage2_10[20]}
   );
   gpc615_5 gpc2135 (
      {stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63]},
      {stage1_11[25]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[9],stage2_12[14],stage2_11[19],stage2_10[21]}
   );
   gpc615_5 gpc2136 (
      {stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68]},
      {stage1_11[26]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[10],stage2_12[15],stage2_11[20],stage2_10[22]}
   );
   gpc615_5 gpc2137 (
      {stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72], stage1_10[73]},
      {stage1_11[27]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[11],stage2_12[16],stage2_11[21],stage2_10[23]}
   );
   gpc615_5 gpc2138 (
      {stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78]},
      {stage1_11[28]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[12],stage2_12[17],stage2_11[22],stage2_10[24]}
   );
   gpc615_5 gpc2139 (
      {stage1_11[29], stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33]},
      {stage1_12[54]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[9],stage2_13[13],stage2_12[18],stage2_11[23]}
   );
   gpc615_5 gpc2140 (
      {stage1_11[34], stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38]},
      {stage1_12[55]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[10],stage2_13[14],stage2_12[19],stage2_11[24]}
   );
   gpc615_5 gpc2141 (
      {stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43]},
      {stage1_12[56]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[11],stage2_13[15],stage2_12[20],stage2_11[25]}
   );
   gpc615_5 gpc2142 (
      {stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_12[57]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[12],stage2_13[16],stage2_12[21],stage2_11[26]}
   );
   gpc615_5 gpc2143 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[58]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[13],stage2_13[17],stage2_12[22],stage2_11[27]}
   );
   gpc615_5 gpc2144 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58]},
      {stage1_12[59]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[14],stage2_13[18],stage2_12[23],stage2_11[28]}
   );
   gpc615_5 gpc2145 (
      {stage1_11[59], stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63]},
      {stage1_12[60]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[15],stage2_13[19],stage2_12[24],stage2_11[29]}
   );
   gpc615_5 gpc2146 (
      {stage1_11[64], stage1_11[65], stage1_11[66], stage1_11[67], stage1_11[68]},
      {stage1_12[61]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[16],stage2_13[20],stage2_12[25],stage2_11[30]}
   );
   gpc615_5 gpc2147 (
      {stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72], stage1_11[73]},
      {stage1_12[62]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[17],stage2_13[21],stage2_12[26],stage2_11[31]}
   );
   gpc606_5 gpc2148 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[9],stage2_14[18],stage2_13[22]}
   );
   gpc606_5 gpc2149 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[1],stage2_15[10],stage2_14[19],stage2_13[23]}
   );
   gpc615_5 gpc2150 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4]},
      {stage1_15[12]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[2],stage2_15[11],stage2_14[20]}
   );
   gpc615_5 gpc2151 (
      {stage1_14[5], stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9]},
      {stage1_15[13]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[3],stage2_15[12],stage2_14[21]}
   );
   gpc606_5 gpc2152 (
      {stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[4],stage2_15[13]}
   );
   gpc606_5 gpc2153 (
      {stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[5],stage2_15[14]}
   );
   gpc606_5 gpc2154 (
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[4],stage2_17[6],stage2_16[6],stage2_15[15]}
   );
   gpc606_5 gpc2155 (
      {stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[5],stage2_17[7],stage2_16[7],stage2_15[16]}
   );
   gpc606_5 gpc2156 (
      {stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[6],stage2_17[8],stage2_16[8],stage2_15[17]}
   );
   gpc606_5 gpc2157 (
      {stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48], stage1_15[49]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[7],stage2_17[9],stage2_16[9],stage2_15[18]}
   );
   gpc606_5 gpc2158 (
      {stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[8],stage2_17[10],stage2_16[10],stage2_15[19]}
   );
   gpc606_5 gpc2159 (
      {stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[9],stage2_17[11],stage2_16[11],stage2_15[20]}
   );
   gpc606_5 gpc2160 (
      {stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[10],stage2_17[12],stage2_16[12],stage2_15[21]}
   );
   gpc606_5 gpc2161 (
      {stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72], stage1_15[73]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[11],stage2_17[13],stage2_16[13],stage2_15[22]}
   );
   gpc606_5 gpc2162 (
      {stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77], stage1_15[78], stage1_15[79]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[12],stage2_17[14],stage2_16[14],stage2_15[23]}
   );
   gpc606_5 gpc2163 (
      {stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83], stage1_15[84], stage1_15[85]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[13],stage2_17[15],stage2_16[15],stage2_15[24]}
   );
   gpc606_5 gpc2164 (
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[12],stage2_18[14],stage2_17[16],stage2_16[16]}
   );
   gpc606_5 gpc2165 (
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[13],stage2_18[15],stage2_17[17],stage2_16[17]}
   );
   gpc606_5 gpc2166 (
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[14],stage2_18[16],stage2_17[18],stage2_16[18]}
   );
   gpc606_5 gpc2167 (
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[15],stage2_18[17],stage2_17[19],stage2_16[19]}
   );
   gpc606_5 gpc2168 (
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[16],stage2_18[18],stage2_17[20],stage2_16[20]}
   );
   gpc606_5 gpc2169 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[5],stage2_19[17],stage2_18[19],stage2_17[21]}
   );
   gpc606_5 gpc2170 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[6],stage2_19[18],stage2_18[20],stage2_17[22]}
   );
   gpc606_5 gpc2171 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[7],stage2_19[19],stage2_18[21],stage2_17[23]}
   );
   gpc615_5 gpc2172 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94]},
      {stage1_18[30]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[8],stage2_19[20],stage2_18[22],stage2_17[24]}
   );
   gpc615_5 gpc2173 (
      {stage1_17[95], stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99]},
      {stage1_18[31]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[9],stage2_19[21],stage2_18[23],stage2_17[25]}
   );
   gpc615_5 gpc2174 (
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36]},
      {stage1_19[30]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[5],stage2_20[10],stage2_19[22],stage2_18[24]}
   );
   gpc615_5 gpc2175 (
      {stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage1_19[31]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[6],stage2_20[11],stage2_19[23],stage2_18[25]}
   );
   gpc615_5 gpc2176 (
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46]},
      {stage1_19[32]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[7],stage2_20[12],stage2_19[24],stage2_18[26]}
   );
   gpc615_5 gpc2177 (
      {stage1_19[33], stage1_19[34], stage1_19[35], stage1_19[36], stage1_19[37]},
      {stage1_20[18]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[8],stage2_20[13],stage2_19[25]}
   );
   gpc615_5 gpc2178 (
      {stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41], stage1_19[42]},
      {stage1_20[19]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[4],stage2_21[9],stage2_20[14],stage2_19[26]}
   );
   gpc615_5 gpc2179 (
      {stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage1_20[20]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[5],stage2_21[10],stage2_20[15],stage2_19[27]}
   );
   gpc606_5 gpc2180 (
      {stage1_20[21], stage1_20[22], stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[3],stage2_22[6],stage2_21[11],stage2_20[16]}
   );
   gpc606_5 gpc2181 (
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[1],stage2_23[4],stage2_22[7],stage2_21[12]}
   );
   gpc606_5 gpc2182 (
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[2],stage2_23[5],stage2_22[8],stage2_21[13]}
   );
   gpc606_5 gpc2183 (
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[3],stage2_23[6],stage2_22[9],stage2_21[14]}
   );
   gpc606_5 gpc2184 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[4],stage2_23[7],stage2_22[10],stage2_21[15]}
   );
   gpc606_5 gpc2185 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[5],stage2_23[8],stage2_22[11],stage2_21[16]}
   );
   gpc1163_5 gpc2186 (
      {stage1_22[6], stage1_22[7], stage1_22[8]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage1_24[0]},
      {stage1_25[0]},
      {stage2_26[0],stage2_25[5],stage2_24[6],stage2_23[9],stage2_22[12]}
   );
   gpc1163_5 gpc2187 (
      {stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage1_24[1]},
      {stage1_25[1]},
      {stage2_26[1],stage2_25[6],stage2_24[7],stage2_23[10],stage2_22[13]}
   );
   gpc1163_5 gpc2188 (
      {stage1_22[12], stage1_22[13], stage1_22[14]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage1_24[2]},
      {stage1_25[2]},
      {stage2_26[2],stage2_25[7],stage2_24[8],stage2_23[11],stage2_22[14]}
   );
   gpc1163_5 gpc2189 (
      {stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage1_24[3]},
      {stage1_25[3]},
      {stage2_26[3],stage2_25[8],stage2_24[9],stage2_23[12],stage2_22[15]}
   );
   gpc1163_5 gpc2190 (
      {stage1_22[18], stage1_22[19], stage1_22[20]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage1_24[4]},
      {stage1_25[4]},
      {stage2_26[4],stage2_25[9],stage2_24[10],stage2_23[13],stage2_22[16]}
   );
   gpc1163_5 gpc2191 (
      {stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage1_24[5]},
      {stage1_25[5]},
      {stage2_26[5],stage2_25[10],stage2_24[11],stage2_23[14],stage2_22[17]}
   );
   gpc1163_5 gpc2192 (
      {stage1_22[24], stage1_22[25], stage1_22[26]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage1_24[6]},
      {stage1_25[6]},
      {stage2_26[6],stage2_25[11],stage2_24[12],stage2_23[15],stage2_22[18]}
   );
   gpc615_5 gpc2193 (
      {stage1_22[27], stage1_22[28], stage1_22[29], stage1_22[30], stage1_22[31]},
      {stage1_23[72]},
      {stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12]},
      {stage2_26[7],stage2_25[12],stage2_24[13],stage2_23[16],stage2_22[19]}
   );
   gpc615_5 gpc2194 (
      {stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35], stage1_22[36]},
      {stage1_23[73]},
      {stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18]},
      {stage2_26[8],stage2_25[13],stage2_24[14],stage2_23[17],stage2_22[20]}
   );
   gpc615_5 gpc2195 (
      {stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_23[74]},
      {stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24]},
      {stage2_26[9],stage2_25[14],stage2_24[15],stage2_23[18],stage2_22[21]}
   );
   gpc615_5 gpc2196 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46]},
      {stage1_23[75]},
      {stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29], stage1_24[30]},
      {stage2_26[10],stage2_25[15],stage2_24[16],stage2_23[19],stage2_22[22]}
   );
   gpc615_5 gpc2197 (
      {stage1_22[47], stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51]},
      {stage1_23[76]},
      {stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35], stage1_24[36]},
      {stage2_26[11],stage2_25[16],stage2_24[17],stage2_23[20],stage2_22[23]}
   );
   gpc615_5 gpc2198 (
      {stage1_22[52], stage1_22[53], stage1_22[54], stage1_22[55], stage1_22[56]},
      {stage1_23[77]},
      {stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41], stage1_24[42]},
      {stage2_26[12],stage2_25[17],stage2_24[18],stage2_23[21],stage2_22[24]}
   );
   gpc615_5 gpc2199 (
      {stage1_22[57], stage1_22[58], stage1_22[59], stage1_22[60], stage1_22[61]},
      {stage1_23[78]},
      {stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47], stage1_24[48]},
      {stage2_26[13],stage2_25[18],stage2_24[19],stage2_23[22],stage2_22[25]}
   );
   gpc606_5 gpc2200 (
      {stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82], stage1_23[83], stage1_23[84]},
      {stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12]},
      {stage2_27[0],stage2_26[14],stage2_25[19],stage2_24[20],stage2_23[23]}
   );
   gpc606_5 gpc2201 (
      {stage1_23[85], stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89], stage1_23[90]},
      {stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18]},
      {stage2_27[1],stage2_26[15],stage2_25[20],stage2_24[21],stage2_23[24]}
   );
   gpc606_5 gpc2202 (
      {stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95], stage1_23[96]},
      {stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23], stage1_25[24]},
      {stage2_27[2],stage2_26[16],stage2_25[21],stage2_24[22],stage2_23[25]}
   );
   gpc606_5 gpc2203 (
      {stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101], stage1_23[102]},
      {stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29], stage1_25[30]},
      {stage2_27[3],stage2_26[17],stage2_25[22],stage2_24[23],stage2_23[26]}
   );
   gpc606_5 gpc2204 (
      {stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107], stage1_23[108]},
      {stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35], stage1_25[36]},
      {stage2_27[4],stage2_26[18],stage2_25[23],stage2_24[24],stage2_23[27]}
   );
   gpc606_5 gpc2205 (
      {stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112], stage1_23[113], stage1_23[114]},
      {stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41], stage1_25[42]},
      {stage2_27[5],stage2_26[19],stage2_25[24],stage2_24[25],stage2_23[28]}
   );
   gpc606_5 gpc2206 (
      {stage1_23[115], stage1_23[116], stage1_23[117], stage1_23[118], stage1_23[119], stage1_23[120]},
      {stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47], stage1_25[48]},
      {stage2_27[6],stage2_26[20],stage2_25[25],stage2_24[26],stage2_23[29]}
   );
   gpc606_5 gpc2207 (
      {stage1_23[121], stage1_23[122], stage1_23[123], stage1_23[124], stage1_23[125], stage1_23[126]},
      {stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53], stage1_25[54]},
      {stage2_27[7],stage2_26[21],stage2_25[26],stage2_24[27],stage2_23[30]}
   );
   gpc615_5 gpc2208 (
      {stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage1_25[55]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[8],stage2_26[22],stage2_25[27],stage2_24[28]}
   );
   gpc615_5 gpc2209 (
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58]},
      {stage1_25[56]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[9],stage2_26[23],stage2_25[28],stage2_24[29]}
   );
   gpc615_5 gpc2210 (
      {stage1_24[59], stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63]},
      {stage1_25[57]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[10],stage2_26[24],stage2_25[29],stage2_24[30]}
   );
   gpc615_5 gpc2211 (
      {stage1_24[64], stage1_24[65], stage1_24[66], stage1_24[67], stage1_24[68]},
      {stage1_25[58]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[11],stage2_26[25],stage2_25[30],stage2_24[31]}
   );
   gpc606_5 gpc2212 (
      {stage1_25[59], stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[4],stage2_27[12],stage2_26[26],stage2_25[31]}
   );
   gpc606_5 gpc2213 (
      {stage1_25[65], stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[5],stage2_27[13],stage2_26[27],stage2_25[32]}
   );
   gpc606_5 gpc2214 (
      {stage1_25[71], stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[6],stage2_27[14],stage2_26[28],stage2_25[33]}
   );
   gpc606_5 gpc2215 (
      {stage1_25[77], stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[7],stage2_27[15],stage2_26[29],stage2_25[34]}
   );
   gpc2116_5 gpc2216 (
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage1_27[24]},
      {stage1_28[0]},
      {stage1_29[0], stage1_29[1]},
      {stage2_30[0],stage2_29[4],stage2_28[8],stage2_27[16],stage2_26[30]}
   );
   gpc2116_5 gpc2217 (
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage1_27[25]},
      {stage1_28[1]},
      {stage1_29[2], stage1_29[3]},
      {stage2_30[1],stage2_29[5],stage2_28[9],stage2_27[17],stage2_26[31]}
   );
   gpc2116_5 gpc2218 (
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage1_27[26]},
      {stage1_28[2]},
      {stage1_29[4], stage1_29[5]},
      {stage2_30[2],stage2_29[6],stage2_28[10],stage2_27[18],stage2_26[32]}
   );
   gpc2116_5 gpc2219 (
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage1_27[27]},
      {stage1_28[3]},
      {stage1_29[6], stage1_29[7]},
      {stage2_30[3],stage2_29[7],stage2_28[11],stage2_27[19],stage2_26[33]}
   );
   gpc2116_5 gpc2220 (
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage1_27[28]},
      {stage1_28[4]},
      {stage1_29[8], stage1_29[9]},
      {stage2_30[4],stage2_29[8],stage2_28[12],stage2_27[20],stage2_26[34]}
   );
   gpc615_5 gpc2221 (
      {stage1_27[29], stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33]},
      {stage1_28[5]},
      {stage1_29[10], stage1_29[11], stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15]},
      {stage2_31[0],stage2_30[5],stage2_29[9],stage2_28[13],stage2_27[21]}
   );
   gpc615_5 gpc2222 (
      {stage1_27[34], stage1_27[35], stage1_27[36], stage1_27[37], stage1_27[38]},
      {stage1_28[6]},
      {stage1_29[16], stage1_29[17], stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21]},
      {stage2_31[1],stage2_30[6],stage2_29[10],stage2_28[14],stage2_27[22]}
   );
   gpc615_5 gpc2223 (
      {stage1_27[39], stage1_27[40], stage1_27[41], stage1_27[42], stage1_27[43]},
      {stage1_28[7]},
      {stage1_29[22], stage1_29[23], stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27]},
      {stage2_31[2],stage2_30[7],stage2_29[11],stage2_28[15],stage2_27[23]}
   );
   gpc615_5 gpc2224 (
      {stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47], stage1_27[48]},
      {stage1_28[8]},
      {stage1_29[28], stage1_29[29], stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33]},
      {stage2_31[3],stage2_30[8],stage2_29[12],stage2_28[16],stage2_27[24]}
   );
   gpc606_5 gpc2225 (
      {stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12], stage1_28[13], stage1_28[14]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[4],stage2_30[9],stage2_29[13],stage2_28[17]}
   );
   gpc606_5 gpc2226 (
      {stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18], stage1_28[19], stage1_28[20]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[5],stage2_30[10],stage2_29[14],stage2_28[18]}
   );
   gpc606_5 gpc2227 (
      {stage1_28[21], stage1_28[22], stage1_28[23], stage1_28[24], stage1_28[25], stage1_28[26]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[6],stage2_30[11],stage2_29[15],stage2_28[19]}
   );
   gpc606_5 gpc2228 (
      {stage1_28[27], stage1_28[28], stage1_28[29], stage1_28[30], stage1_28[31], stage1_28[32]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[7],stage2_30[12],stage2_29[16],stage2_28[20]}
   );
   gpc606_5 gpc2229 (
      {stage1_28[33], stage1_28[34], stage1_28[35], stage1_28[36], stage1_28[37], stage1_28[38]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[8],stage2_30[13],stage2_29[17],stage2_28[21]}
   );
   gpc606_5 gpc2230 (
      {stage1_28[39], stage1_28[40], stage1_28[41], stage1_28[42], stage1_28[43], stage1_28[44]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[9],stage2_30[14],stage2_29[18],stage2_28[22]}
   );
   gpc606_5 gpc2231 (
      {stage1_28[45], stage1_28[46], stage1_28[47], stage1_28[48], stage1_28[49], stage1_28[50]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[10],stage2_30[15],stage2_29[19],stage2_28[23]}
   );
   gpc606_5 gpc2232 (
      {stage1_28[51], stage1_28[52], stage1_28[53], stage1_28[54], stage1_28[55], stage1_28[56]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[11],stage2_30[16],stage2_29[20],stage2_28[24]}
   );
   gpc606_5 gpc2233 (
      {stage1_28[57], stage1_28[58], stage1_28[59], stage1_28[60], stage1_28[61], stage1_28[62]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[12],stage2_30[17],stage2_29[21],stage2_28[25]}
   );
   gpc606_5 gpc2234 (
      {stage1_28[63], stage1_28[64], stage1_28[65], stage1_28[66], stage1_28[67], stage1_28[68]},
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage2_32[9],stage2_31[13],stage2_30[18],stage2_29[22],stage2_28[26]}
   );
   gpc606_5 gpc2235 (
      {stage1_29[34], stage1_29[35], stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[10],stage2_31[14],stage2_30[19],stage2_29[23]}
   );
   gpc606_5 gpc2236 (
      {stage1_29[40], stage1_29[41], stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[11],stage2_31[15],stage2_30[20],stage2_29[24]}
   );
   gpc606_5 gpc2237 (
      {stage1_29[46], stage1_29[47], stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[12],stage2_31[16],stage2_30[21],stage2_29[25]}
   );
   gpc606_5 gpc2238 (
      {stage1_29[52], stage1_29[53], stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[13],stage2_31[17],stage2_30[22],stage2_29[26]}
   );
   gpc606_5 gpc2239 (
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[4],stage2_32[14],stage2_31[18],stage2_30[23]}
   );
   gpc606_5 gpc2240 (
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[5],stage2_32[15],stage2_31[19],stage2_30[24]}
   );
   gpc606_5 gpc2241 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[6],stage2_32[16],stage2_31[20],stage2_30[25]}
   );
   gpc606_5 gpc2242 (
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[7],stage2_32[17],stage2_31[21],stage2_30[26]}
   );
   gpc615_5 gpc2243 (
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28]},
      {stage1_32[24]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[4],stage2_33[8],stage2_32[18],stage2_31[22]}
   );
   gpc615_5 gpc2244 (
      {stage1_31[29], stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33]},
      {stage1_32[25]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[5],stage2_33[9],stage2_32[19],stage2_31[23]}
   );
   gpc615_5 gpc2245 (
      {stage1_31[34], stage1_31[35], stage1_31[36], stage1_31[37], stage1_31[38]},
      {stage1_32[26]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[6],stage2_33[10],stage2_32[20],stage2_31[24]}
   );
   gpc615_5 gpc2246 (
      {stage1_31[39], stage1_31[40], stage1_31[41], stage1_31[42], stage1_31[43]},
      {stage1_32[27]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[7],stage2_33[11],stage2_32[21],stage2_31[25]}
   );
   gpc615_5 gpc2247 (
      {stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48]},
      {stage1_32[28]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[8],stage2_33[12],stage2_32[22],stage2_31[26]}
   );
   gpc615_5 gpc2248 (
      {stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage1_32[29]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[9],stage2_33[13],stage2_32[23],stage2_31[27]}
   );
   gpc615_5 gpc2249 (
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58]},
      {stage1_32[30]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[10],stage2_33[14],stage2_32[24],stage2_31[28]}
   );
   gpc615_5 gpc2250 (
      {stage1_31[59], stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63]},
      {stage1_32[31]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[11],stage2_33[15],stage2_32[25],stage2_31[29]}
   );
   gpc615_5 gpc2251 (
      {stage1_31[64], stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68]},
      {stage1_32[32]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[12],stage2_33[16],stage2_32[26],stage2_31[30]}
   );
   gpc615_5 gpc2252 (
      {stage1_31[69], stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73]},
      {stage1_32[33]},
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage2_35[9],stage2_34[13],stage2_33[17],stage2_32[27],stage2_31[31]}
   );
   gpc615_5 gpc2253 (
      {stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78]},
      {stage1_32[34]},
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage2_35[10],stage2_34[14],stage2_33[18],stage2_32[28],stage2_31[32]}
   );
   gpc615_5 gpc2254 (
      {stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage1_32[35]},
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71]},
      {stage2_35[11],stage2_34[15],stage2_33[19],stage2_32[29],stage2_31[33]}
   );
   gpc615_5 gpc2255 (
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88]},
      {stage1_32[36]},
      {stage1_33[72], stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77]},
      {stage2_35[12],stage2_34[16],stage2_33[20],stage2_32[30],stage2_31[34]}
   );
   gpc615_5 gpc2256 (
      {stage1_31[89], stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93]},
      {stage1_32[37]},
      {stage1_33[78], stage1_33[79], stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83]},
      {stage2_35[13],stage2_34[17],stage2_33[21],stage2_32[31],stage2_31[35]}
   );
   gpc606_5 gpc2257 (
      {stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[14],stage2_34[18],stage2_33[22],stage2_32[32]}
   );
   gpc606_5 gpc2258 (
      {stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[15],stage2_34[19],stage2_33[23],stage2_32[33]}
   );
   gpc606_5 gpc2259 (
      {stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[16],stage2_34[20],stage2_33[24],stage2_32[34]}
   );
   gpc606_5 gpc2260 (
      {stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[17],stage2_34[21],stage2_33[25],stage2_32[35]}
   );
   gpc606_5 gpc2261 (
      {stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[18],stage2_34[22],stage2_33[26],stage2_32[36]}
   );
   gpc606_5 gpc2262 (
      {stage1_33[84], stage1_33[85], stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[5],stage2_35[19],stage2_34[23],stage2_33[27]}
   );
   gpc606_5 gpc2263 (
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[1],stage2_36[6],stage2_35[20],stage2_34[24]}
   );
   gpc606_5 gpc2264 (
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[2],stage2_36[7],stage2_35[21],stage2_34[25]}
   );
   gpc606_5 gpc2265 (
      {stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[3],stage2_36[8],stage2_35[22],stage2_34[26]}
   );
   gpc615_5 gpc2266 (
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10]},
      {stage1_36[18]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[3],stage2_37[4],stage2_36[9],stage2_35[23]}
   );
   gpc615_5 gpc2267 (
      {stage1_35[11], stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15]},
      {stage1_36[19]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[4],stage2_37[5],stage2_36[10],stage2_35[24]}
   );
   gpc615_5 gpc2268 (
      {stage1_35[16], stage1_35[17], stage1_35[18], stage1_35[19], stage1_35[20]},
      {stage1_36[20]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[5],stage2_37[6],stage2_36[11],stage2_35[25]}
   );
   gpc615_5 gpc2269 (
      {stage1_35[21], stage1_35[22], stage1_35[23], stage1_35[24], stage1_35[25]},
      {stage1_36[21]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[6],stage2_37[7],stage2_36[12],stage2_35[26]}
   );
   gpc615_5 gpc2270 (
      {stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29], stage1_35[30]},
      {stage1_36[22]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[7],stage2_37[8],stage2_36[13],stage2_35[27]}
   );
   gpc615_5 gpc2271 (
      {stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage1_36[23]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[8],stage2_37[9],stage2_36[14],stage2_35[28]}
   );
   gpc615_5 gpc2272 (
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40]},
      {stage1_36[24]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[9],stage2_37[10],stage2_36[15],stage2_35[29]}
   );
   gpc615_5 gpc2273 (
      {stage1_35[41], stage1_35[42], stage1_35[43], stage1_35[44], stage1_35[45]},
      {stage1_36[25]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[10],stage2_37[11],stage2_36[16],stage2_35[30]}
   );
   gpc1343_5 gpc2274 (
      {stage1_36[26], stage1_36[27], stage1_36[28]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51]},
      {stage1_38[0], stage1_38[1], stage1_38[2]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[8],stage2_38[11],stage2_37[12],stage2_36[17]}
   );
   gpc606_5 gpc2275 (
      {stage1_36[29], stage1_36[30], stage1_36[31], stage1_36[32], stage1_36[33], stage1_36[34]},
      {stage1_38[3], stage1_38[4], stage1_38[5], stage1_38[6], stage1_38[7], stage1_38[8]},
      {stage2_40[1],stage2_39[9],stage2_38[12],stage2_37[13],stage2_36[18]}
   );
   gpc606_5 gpc2276 (
      {stage1_36[35], stage1_36[36], stage1_36[37], stage1_36[38], stage1_36[39], stage1_36[40]},
      {stage1_38[9], stage1_38[10], stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14]},
      {stage2_40[2],stage2_39[10],stage2_38[13],stage2_37[14],stage2_36[19]}
   );
   gpc606_5 gpc2277 (
      {stage1_36[41], stage1_36[42], stage1_36[43], stage1_36[44], stage1_36[45], stage1_36[46]},
      {stage1_38[15], stage1_38[16], stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20]},
      {stage2_40[3],stage2_39[11],stage2_38[14],stage2_37[15],stage2_36[20]}
   );
   gpc615_5 gpc2278 (
      {stage1_36[47], stage1_36[48], stage1_36[49], stage1_36[50], stage1_36[51]},
      {stage1_37[52]},
      {stage1_38[21], stage1_38[22], stage1_38[23], stage1_38[24], stage1_38[25], stage1_38[26]},
      {stage2_40[4],stage2_39[12],stage2_38[15],stage2_37[16],stage2_36[21]}
   );
   gpc615_5 gpc2279 (
      {stage1_36[52], stage1_36[53], stage1_36[54], stage1_36[55], stage1_36[56]},
      {stage1_37[53]},
      {stage1_38[27], stage1_38[28], stage1_38[29], stage1_38[30], stage1_38[31], stage1_38[32]},
      {stage2_40[5],stage2_39[13],stage2_38[16],stage2_37[17],stage2_36[22]}
   );
   gpc615_5 gpc2280 (
      {stage1_36[57], stage1_36[58], stage1_36[59], stage1_36[60], stage1_36[61]},
      {stage1_37[54]},
      {stage1_38[33], stage1_38[34], stage1_38[35], stage1_38[36], stage1_38[37], stage1_38[38]},
      {stage2_40[6],stage2_39[14],stage2_38[17],stage2_37[18],stage2_36[23]}
   );
   gpc615_5 gpc2281 (
      {stage1_36[62], stage1_36[63], stage1_36[64], stage1_36[65], stage1_36[66]},
      {stage1_37[55]},
      {stage1_38[39], stage1_38[40], stage1_38[41], stage1_38[42], stage1_38[43], stage1_38[44]},
      {stage2_40[7],stage2_39[15],stage2_38[18],stage2_37[19],stage2_36[24]}
   );
   gpc615_5 gpc2282 (
      {stage1_36[67], stage1_36[68], stage1_36[69], stage1_36[70], stage1_36[71]},
      {stage1_37[56]},
      {stage1_38[45], stage1_38[46], stage1_38[47], stage1_38[48], stage1_38[49], stage1_38[50]},
      {stage2_40[8],stage2_39[16],stage2_38[19],stage2_37[20],stage2_36[25]}
   );
   gpc606_5 gpc2283 (
      {stage1_37[57], stage1_37[58], stage1_37[59], stage1_37[60], stage1_37[61], stage1_37[62]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[9],stage2_39[17],stage2_38[20],stage2_37[21]}
   );
   gpc606_5 gpc2284 (
      {stage1_37[63], stage1_37[64], stage1_37[65], stage1_37[66], stage1_37[67], stage1_37[68]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[10],stage2_39[18],stage2_38[21],stage2_37[22]}
   );
   gpc606_5 gpc2285 (
      {stage1_37[69], stage1_37[70], stage1_37[71], stage1_37[72], stage1_37[73], stage1_37[74]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[11],stage2_39[19],stage2_38[22],stage2_37[23]}
   );
   gpc606_5 gpc2286 (
      {stage1_37[75], stage1_37[76], stage1_37[77], stage1_37[78], stage1_37[79], stage1_37[80]},
      {stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24]},
      {stage2_41[3],stage2_40[12],stage2_39[20],stage2_38[23],stage2_37[24]}
   );
   gpc606_5 gpc2287 (
      {stage1_37[81], stage1_37[82], stage1_37[83], stage1_37[84], stage1_37[85], stage1_37[86]},
      {stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30]},
      {stage2_41[4],stage2_40[13],stage2_39[21],stage2_38[24],stage2_37[25]}
   );
   gpc606_5 gpc2288 (
      {stage1_37[87], stage1_37[88], stage1_37[89], stage1_37[90], stage1_37[91], stage1_37[92]},
      {stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36]},
      {stage2_41[5],stage2_40[14],stage2_39[22],stage2_38[25],stage2_37[26]}
   );
   gpc606_5 gpc2289 (
      {stage1_37[93], stage1_37[94], stage1_37[95], stage1_37[96], stage1_37[97], stage1_37[98]},
      {stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42]},
      {stage2_41[6],stage2_40[15],stage2_39[23],stage2_38[26],stage2_37[27]}
   );
   gpc606_5 gpc2290 (
      {stage1_37[99], stage1_37[100], stage1_37[101], stage1_37[102], stage1_37[103], stage1_37[104]},
      {stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48]},
      {stage2_41[7],stage2_40[16],stage2_39[24],stage2_38[27],stage2_37[28]}
   );
   gpc606_5 gpc2291 (
      {stage1_37[105], stage1_37[106], stage1_37[107], stage1_37[108], stage1_37[109], stage1_37[110]},
      {stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54]},
      {stage2_41[8],stage2_40[17],stage2_39[25],stage2_38[28],stage2_37[29]}
   );
   gpc606_5 gpc2292 (
      {stage1_37[111], stage1_37[112], stage1_37[113], stage1_37[114], stage1_37[115], stage1_37[116]},
      {stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60]},
      {stage2_41[9],stage2_40[18],stage2_39[26],stage2_38[29],stage2_37[30]}
   );
   gpc615_5 gpc2293 (
      {stage1_38[51], stage1_38[52], stage1_38[53], stage1_38[54], stage1_38[55]},
      {stage1_39[61]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[10],stage2_40[19],stage2_39[27],stage2_38[30]}
   );
   gpc615_5 gpc2294 (
      {stage1_38[56], stage1_38[57], stage1_38[58], stage1_38[59], stage1_38[60]},
      {stage1_39[62]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[11],stage2_40[20],stage2_39[28],stage2_38[31]}
   );
   gpc615_5 gpc2295 (
      {stage1_38[61], stage1_38[62], stage1_38[63], stage1_38[64], stage1_38[65]},
      {stage1_39[63]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[12],stage2_40[21],stage2_39[29],stage2_38[32]}
   );
   gpc606_5 gpc2296 (
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[3],stage2_41[13],stage2_40[22]}
   );
   gpc606_5 gpc2297 (
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[1],stage2_42[4],stage2_41[14],stage2_40[23]}
   );
   gpc606_5 gpc2298 (
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[2],stage2_42[5],stage2_41[15],stage2_40[24]}
   );
   gpc606_5 gpc2299 (
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[3],stage2_42[6],stage2_41[16],stage2_40[25]}
   );
   gpc606_5 gpc2300 (
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[4],stage2_42[7],stage2_41[17],stage2_40[26]}
   );
   gpc606_5 gpc2301 (
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[5],stage2_42[8],stage2_41[18],stage2_40[27]}
   );
   gpc606_5 gpc2302 (
      {stage1_40[54], stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58], stage1_40[59]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[6],stage2_42[9],stage2_41[19],stage2_40[28]}
   );
   gpc606_5 gpc2303 (
      {stage1_40[60], stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64], stage1_40[65]},
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage2_44[7],stage2_43[7],stage2_42[10],stage2_41[20],stage2_40[29]}
   );
   gpc606_5 gpc2304 (
      {stage1_40[66], stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70], stage1_40[71]},
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage2_44[8],stage2_43[8],stage2_42[11],stage2_41[21],stage2_40[30]}
   );
   gpc606_5 gpc2305 (
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[9],stage2_43[9],stage2_42[12],stage2_41[22]}
   );
   gpc606_5 gpc2306 (
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[10],stage2_43[10],stage2_42[13],stage2_41[23]}
   );
   gpc606_5 gpc2307 (
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[11],stage2_43[11],stage2_42[14],stage2_41[24]}
   );
   gpc606_5 gpc2308 (
      {stage1_41[18], stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[12],stage2_43[12],stage2_42[15],stage2_41[25]}
   );
   gpc606_5 gpc2309 (
      {stage1_41[24], stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[13],stage2_43[13],stage2_42[16],stage2_41[26]}
   );
   gpc606_5 gpc2310 (
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[14],stage2_43[14],stage2_42[17],stage2_41[27]}
   );
   gpc606_5 gpc2311 (
      {stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[15],stage2_43[15],stage2_42[18],stage2_41[28]}
   );
   gpc606_5 gpc2312 (
      {stage1_41[42], stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[16],stage2_43[16],stage2_42[19],stage2_41[29]}
   );
   gpc606_5 gpc2313 (
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[8],stage2_44[17],stage2_43[17]}
   );
   gpc606_5 gpc2314 (
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[9],stage2_44[18],stage2_43[18]}
   );
   gpc606_5 gpc2315 (
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[2],stage2_45[10],stage2_44[19],stage2_43[19]}
   );
   gpc606_5 gpc2316 (
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[3],stage2_45[11],stage2_44[20],stage2_43[20]}
   );
   gpc606_5 gpc2317 (
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[4],stage2_45[12],stage2_44[21],stage2_43[21]}
   );
   gpc606_5 gpc2318 (
      {stage1_43[78], stage1_43[79], stage1_43[80], stage1_43[81], stage1_43[82], stage1_43[83]},
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage2_47[5],stage2_46[5],stage2_45[13],stage2_44[22],stage2_43[22]}
   );
   gpc606_5 gpc2319 (
      {stage1_43[84], stage1_43[85], stage1_43[86], stage1_43[87], stage1_43[88], stage1_43[89]},
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage2_47[6],stage2_46[6],stage2_45[14],stage2_44[23],stage2_43[23]}
   );
   gpc606_5 gpc2320 (
      {stage1_43[90], stage1_43[91], stage1_43[92], stage1_43[93], stage1_43[94], stage1_43[95]},
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage2_47[7],stage2_46[7],stage2_45[15],stage2_44[24],stage2_43[24]}
   );
   gpc606_5 gpc2321 (
      {stage1_43[96], stage1_43[97], stage1_43[98], stage1_43[99], stage1_43[100], stage1_43[101]},
      {stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51], stage1_45[52], stage1_45[53]},
      {stage2_47[8],stage2_46[8],stage2_45[16],stage2_44[25],stage2_43[25]}
   );
   gpc606_5 gpc2322 (
      {stage1_43[102], stage1_43[103], stage1_43[104], stage1_43[105], stage1_43[106], stage1_43[107]},
      {stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57], stage1_45[58], stage1_45[59]},
      {stage2_47[9],stage2_46[9],stage2_45[17],stage2_44[26],stage2_43[26]}
   );
   gpc606_5 gpc2323 (
      {stage1_43[108], stage1_43[109], stage1_43[110], stage1_43[111], stage1_43[112], stage1_43[113]},
      {stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63], stage1_45[64], stage1_45[65]},
      {stage2_47[10],stage2_46[10],stage2_45[18],stage2_44[27],stage2_43[27]}
   );
   gpc615_5 gpc2324 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4]},
      {stage1_45[66]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[11],stage2_46[11],stage2_45[19],stage2_44[28]}
   );
   gpc615_5 gpc2325 (
      {stage1_44[5], stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9]},
      {stage1_45[67]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[12],stage2_46[12],stage2_45[20],stage2_44[29]}
   );
   gpc606_5 gpc2326 (
      {stage1_45[68], stage1_45[69], stage1_45[70], stage1_45[71], stage1_45[72], stage1_45[73]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[2],stage2_47[13],stage2_46[13],stage2_45[21]}
   );
   gpc606_5 gpc2327 (
      {stage1_45[74], stage1_45[75], stage1_45[76], stage1_45[77], stage1_45[78], stage1_45[79]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[3],stage2_47[14],stage2_46[14],stage2_45[22]}
   );
   gpc606_5 gpc2328 (
      {stage1_45[80], stage1_45[81], stage1_45[82], stage1_45[83], stage1_45[84], stage1_45[85]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[4],stage2_47[15],stage2_46[15],stage2_45[23]}
   );
   gpc606_5 gpc2329 (
      {stage1_45[86], stage1_45[87], stage1_45[88], stage1_45[89], stage1_45[90], stage1_45[91]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[5],stage2_47[16],stage2_46[16],stage2_45[24]}
   );
   gpc615_5 gpc2330 (
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16]},
      {stage1_47[24]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[4],stage2_48[6],stage2_47[17],stage2_46[17]}
   );
   gpc615_5 gpc2331 (
      {stage1_46[17], stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21]},
      {stage1_47[25]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[5],stage2_48[7],stage2_47[18],stage2_46[18]}
   );
   gpc615_5 gpc2332 (
      {stage1_46[22], stage1_46[23], stage1_46[24], stage1_46[25], stage1_46[26]},
      {stage1_47[26]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[6],stage2_48[8],stage2_47[19],stage2_46[19]}
   );
   gpc615_5 gpc2333 (
      {stage1_46[27], stage1_46[28], stage1_46[29], stage1_46[30], stage1_46[31]},
      {stage1_47[27]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[7],stage2_48[9],stage2_47[20],stage2_46[20]}
   );
   gpc615_5 gpc2334 (
      {stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35], stage1_46[36]},
      {stage1_47[28]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[8],stage2_48[10],stage2_47[21],stage2_46[21]}
   );
   gpc615_5 gpc2335 (
      {stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage1_47[29]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[9],stage2_48[11],stage2_47[22],stage2_46[22]}
   );
   gpc615_5 gpc2336 (
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46]},
      {stage1_47[30]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[10],stage2_48[12],stage2_47[23],stage2_46[23]}
   );
   gpc615_5 gpc2337 (
      {stage1_46[47], stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51]},
      {stage1_47[31]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[11],stage2_48[13],stage2_47[24],stage2_46[24]}
   );
   gpc615_5 gpc2338 (
      {stage1_46[52], stage1_46[53], stage1_46[54], stage1_46[55], stage1_46[56]},
      {stage1_47[32]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[12],stage2_48[14],stage2_47[25],stage2_46[25]}
   );
   gpc606_5 gpc2339 (
      {stage1_47[33], stage1_47[34], stage1_47[35], stage1_47[36], stage1_47[37], stage1_47[38]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[9],stage2_49[13],stage2_48[15],stage2_47[26]}
   );
   gpc606_5 gpc2340 (
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[1],stage2_50[10],stage2_49[14],stage2_48[16]}
   );
   gpc606_5 gpc2341 (
      {stage1_48[60], stage1_48[61], stage1_48[62], stage1_48[63], stage1_48[64], stage1_48[65]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[2],stage2_50[11],stage2_49[15],stage2_48[17]}
   );
   gpc606_5 gpc2342 (
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[2],stage2_51[3],stage2_50[12],stage2_49[16]}
   );
   gpc606_5 gpc2343 (
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[3],stage2_51[4],stage2_50[13],stage2_49[17]}
   );
   gpc606_5 gpc2344 (
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[4],stage2_51[5],stage2_50[14],stage2_49[18]}
   );
   gpc606_5 gpc2345 (
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage2_53[3],stage2_52[5],stage2_51[6],stage2_50[15],stage2_49[19]}
   );
   gpc606_5 gpc2346 (
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage2_53[4],stage2_52[6],stage2_51[7],stage2_50[16],stage2_49[20]}
   );
   gpc606_5 gpc2347 (
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage2_53[5],stage2_52[7],stage2_51[8],stage2_50[17],stage2_49[21]}
   );
   gpc606_5 gpc2348 (
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39], stage1_51[40], stage1_51[41]},
      {stage2_53[6],stage2_52[8],stage2_51[9],stage2_50[18],stage2_49[22]}
   );
   gpc606_5 gpc2349 (
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45], stage1_51[46], stage1_51[47]},
      {stage2_53[7],stage2_52[9],stage2_51[10],stage2_50[19],stage2_49[23]}
   );
   gpc606_5 gpc2350 (
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage1_51[48], stage1_51[49], stage1_51[50], stage1_51[51], stage1_51[52], stage1_51[53]},
      {stage2_53[8],stage2_52[10],stage2_51[11],stage2_50[20],stage2_49[24]}
   );
   gpc606_5 gpc2351 (
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage1_51[54], stage1_51[55], stage1_51[56], stage1_51[57], stage1_51[58], stage1_51[59]},
      {stage2_53[9],stage2_52[11],stage2_51[12],stage2_50[21],stage2_49[25]}
   );
   gpc606_5 gpc2352 (
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage1_51[60], stage1_51[61], stage1_51[62], stage1_51[63], stage1_51[64], stage1_51[65]},
      {stage2_53[10],stage2_52[12],stage2_51[13],stage2_50[22],stage2_49[26]}
   );
   gpc606_5 gpc2353 (
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage1_51[66], stage1_51[67], stage1_51[68], stage1_51[69], stage1_51[70], stage1_51[71]},
      {stage2_53[11],stage2_52[13],stage2_51[14],stage2_50[23],stage2_49[27]}
   );
   gpc117_4 gpc2354 (
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17], stage1_50[18]},
      {stage1_51[72]},
      {stage1_52[0]},
      {stage2_53[12],stage2_52[14],stage2_51[15],stage2_50[24]}
   );
   gpc606_5 gpc2355 (
      {stage1_50[19], stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23], stage1_50[24]},
      {stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5], stage1_52[6]},
      {stage2_54[0],stage2_53[13],stage2_52[15],stage2_51[16],stage2_50[25]}
   );
   gpc606_5 gpc2356 (
      {stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29], stage1_50[30]},
      {stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11], stage1_52[12]},
      {stage2_54[1],stage2_53[14],stage2_52[16],stage2_51[17],stage2_50[26]}
   );
   gpc606_5 gpc2357 (
      {stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35], stage1_50[36]},
      {stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17], stage1_52[18]},
      {stage2_54[2],stage2_53[15],stage2_52[17],stage2_51[18],stage2_50[27]}
   );
   gpc615_5 gpc2358 (
      {stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage1_51[73]},
      {stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23], stage1_52[24]},
      {stage2_54[3],stage2_53[16],stage2_52[18],stage2_51[19],stage2_50[28]}
   );
   gpc615_5 gpc2359 (
      {stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45], stage1_50[46]},
      {stage1_51[74]},
      {stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28], stage1_52[29], stage1_52[30]},
      {stage2_54[4],stage2_53[17],stage2_52[19],stage2_51[20],stage2_50[29]}
   );
   gpc606_5 gpc2360 (
      {stage1_51[75], stage1_51[76], stage1_51[77], stage1_51[78], stage1_51[79], stage1_51[80]},
      {stage1_53[0], stage1_53[1], stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5]},
      {stage2_55[0],stage2_54[5],stage2_53[18],stage2_52[20],stage2_51[21]}
   );
   gpc606_5 gpc2361 (
      {stage1_51[81], stage1_51[82], stage1_51[83], stage1_51[84], stage1_51[85], stage1_51[86]},
      {stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11]},
      {stage2_55[1],stage2_54[6],stage2_53[19],stage2_52[21],stage2_51[22]}
   );
   gpc606_5 gpc2362 (
      {stage1_51[87], stage1_51[88], stage1_51[89], stage1_51[90], stage1_51[91], stage1_51[92]},
      {stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15], stage1_53[16], stage1_53[17]},
      {stage2_55[2],stage2_54[7],stage2_53[20],stage2_52[22],stage2_51[23]}
   );
   gpc606_5 gpc2363 (
      {stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34], stage1_52[35], stage1_52[36]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[3],stage2_54[8],stage2_53[21],stage2_52[23]}
   );
   gpc606_5 gpc2364 (
      {stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41], stage1_52[42]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[4],stage2_54[9],stage2_53[22],stage2_52[24]}
   );
   gpc606_5 gpc2365 (
      {stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47], stage1_52[48]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[5],stage2_54[10],stage2_53[23],stage2_52[25]}
   );
   gpc606_5 gpc2366 (
      {stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53], stage1_52[54]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[6],stage2_54[11],stage2_53[24],stage2_52[26]}
   );
   gpc606_5 gpc2367 (
      {stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59], stage1_52[60]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[7],stage2_54[12],stage2_53[25],stage2_52[27]}
   );
   gpc606_5 gpc2368 (
      {stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64], stage1_52[65], stage1_52[66]},
      {stage1_54[30], stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage2_56[5],stage2_55[8],stage2_54[13],stage2_53[26],stage2_52[28]}
   );
   gpc606_5 gpc2369 (
      {stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70], stage1_52[71], stage1_52[72]},
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40], stage1_54[41]},
      {stage2_56[6],stage2_55[9],stage2_54[14],stage2_53[27],stage2_52[29]}
   );
   gpc606_5 gpc2370 (
      {stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21], stage1_53[22], stage1_53[23]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[7],stage2_55[10],stage2_54[15],stage2_53[28]}
   );
   gpc606_5 gpc2371 (
      {stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[8],stage2_55[11],stage2_54[16],stage2_53[29]}
   );
   gpc606_5 gpc2372 (
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34], stage1_53[35]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[9],stage2_55[12],stage2_54[17],stage2_53[30]}
   );
   gpc606_5 gpc2373 (
      {stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39], stage1_53[40], stage1_53[41]},
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23]},
      {stage2_57[3],stage2_56[10],stage2_55[13],stage2_54[18],stage2_53[31]}
   );
   gpc606_5 gpc2374 (
      {stage1_53[42], stage1_53[43], stage1_53[44], stage1_53[45], stage1_53[46], stage1_53[47]},
      {stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29]},
      {stage2_57[4],stage2_56[11],stage2_55[14],stage2_54[19],stage2_53[32]}
   );
   gpc615_5 gpc2375 (
      {stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46]},
      {stage1_55[30]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[5],stage2_56[12],stage2_55[15],stage2_54[20]}
   );
   gpc615_5 gpc2376 (
      {stage1_54[47], stage1_54[48], stage1_54[49], stage1_54[50], stage1_54[51]},
      {stage1_55[31]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[6],stage2_56[13],stage2_55[16],stage2_54[21]}
   );
   gpc606_5 gpc2377 (
      {stage1_55[32], stage1_55[33], stage1_55[34], stage1_55[35], stage1_55[36], stage1_55[37]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[2],stage2_57[7],stage2_56[14],stage2_55[17]}
   );
   gpc615_5 gpc2378 (
      {stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41], stage1_55[42]},
      {stage1_56[12]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[3],stage2_57[8],stage2_56[15],stage2_55[18]}
   );
   gpc615_5 gpc2379 (
      {stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage1_56[13]},
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage2_59[2],stage2_58[4],stage2_57[9],stage2_56[16],stage2_55[19]}
   );
   gpc615_5 gpc2380 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[14]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[3],stage2_58[5],stage2_57[10],stage2_56[17],stage2_55[20]}
   );
   gpc615_5 gpc2381 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[15]},
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage2_59[4],stage2_58[6],stage2_57[11],stage2_56[18],stage2_55[21]}
   );
   gpc615_5 gpc2382 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[16]},
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage2_59[5],stage2_58[7],stage2_57[12],stage2_56[19],stage2_55[22]}
   );
   gpc615_5 gpc2383 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[17]},
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage2_59[6],stage2_58[8],stage2_57[13],stage2_56[20],stage2_55[23]}
   );
   gpc615_5 gpc2384 (
      {stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71], stage1_55[72]},
      {stage1_56[18]},
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage2_59[7],stage2_58[9],stage2_57[14],stage2_56[21],stage2_55[24]}
   );
   gpc615_5 gpc2385 (
      {stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage1_56[19]},
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage2_59[8],stage2_58[10],stage2_57[15],stage2_56[22],stage2_55[25]}
   );
   gpc615_5 gpc2386 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82]},
      {stage1_56[20]},
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage2_59[9],stage2_58[11],stage2_57[16],stage2_56[23],stage2_55[26]}
   );
   gpc615_5 gpc2387 (
      {stage1_55[83], stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87]},
      {stage1_56[21]},
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage2_59[10],stage2_58[12],stage2_57[17],stage2_56[24],stage2_55[27]}
   );
   gpc606_5 gpc2388 (
      {stage1_56[22], stage1_56[23], stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[11],stage2_58[13],stage2_57[18],stage2_56[25]}
   );
   gpc606_5 gpc2389 (
      {stage1_56[28], stage1_56[29], stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[12],stage2_58[14],stage2_57[19],stage2_56[26]}
   );
   gpc606_5 gpc2390 (
      {stage1_56[34], stage1_56[35], stage1_56[36], stage1_56[37], stage1_56[38], stage1_56[39]},
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage2_60[2],stage2_59[13],stage2_58[15],stage2_57[20],stage2_56[27]}
   );
   gpc606_5 gpc2391 (
      {stage1_56[40], stage1_56[41], stage1_56[42], stage1_56[43], stage1_56[44], stage1_56[45]},
      {stage1_58[18], stage1_58[19], stage1_58[20], stage1_58[21], stage1_58[22], stage1_58[23]},
      {stage2_60[3],stage2_59[14],stage2_58[16],stage2_57[21],stage2_56[28]}
   );
   gpc606_5 gpc2392 (
      {stage1_56[46], stage1_56[47], stage1_56[48], stage1_56[49], stage1_56[50], stage1_56[51]},
      {stage1_58[24], stage1_58[25], stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29]},
      {stage2_60[4],stage2_59[15],stage2_58[17],stage2_57[22],stage2_56[29]}
   );
   gpc606_5 gpc2393 (
      {stage1_56[52], stage1_56[53], stage1_56[54], stage1_56[55], stage1_56[56], stage1_56[57]},
      {stage1_58[30], stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage2_60[5],stage2_59[16],stage2_58[18],stage2_57[23],stage2_56[30]}
   );
   gpc606_5 gpc2394 (
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[0],stage2_60[6],stage2_59[17],stage2_58[19]}
   );
   gpc606_5 gpc2395 (
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[1],stage2_60[7],stage2_59[18],stage2_58[20]}
   );
   gpc606_5 gpc2396 (
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[2],stage2_60[8],stage2_59[19],stage2_58[21]}
   );
   gpc606_5 gpc2397 (
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage2_62[3],stage2_61[3],stage2_60[9],stage2_59[20],stage2_58[22]}
   );
   gpc615_5 gpc2398 (
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64]},
      {stage1_59[0]},
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage2_62[4],stage2_61[4],stage2_60[10],stage2_59[21],stage2_58[23]}
   );
   gpc606_5 gpc2399 (
      {stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5], stage1_59[6]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[5],stage2_61[5],stage2_60[11],stage2_59[22]}
   );
   gpc606_5 gpc2400 (
      {stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11], stage1_59[12]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[6],stage2_61[6],stage2_60[12],stage2_59[23]}
   );
   gpc606_5 gpc2401 (
      {stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17], stage1_59[18]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[7],stage2_61[7],stage2_60[13],stage2_59[24]}
   );
   gpc606_5 gpc2402 (
      {stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23], stage1_59[24]},
      {stage1_61[18], stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage2_63[3],stage2_62[8],stage2_61[8],stage2_60[14],stage2_59[25]}
   );
   gpc606_5 gpc2403 (
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[4],stage2_62[9],stage2_61[9],stage2_60[15]}
   );
   gpc606_5 gpc2404 (
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage2_64[1],stage2_63[5],stage2_62[10],stage2_61[10],stage2_60[16]}
   );
   gpc606_5 gpc2405 (
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage2_64[2],stage2_63[6],stage2_62[11],stage2_61[11],stage2_60[17]}
   );
   gpc606_5 gpc2406 (
      {stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51], stage1_60[52], stage1_60[53]},
      {stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage2_64[3],stage2_63[7],stage2_62[12],stage2_61[12],stage2_60[18]}
   );
   gpc606_5 gpc2407 (
      {stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57], stage1_60[58], stage1_60[59]},
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage2_64[4],stage2_63[8],stage2_62[13],stage2_61[13],stage2_60[19]}
   );
   gpc606_5 gpc2408 (
      {stage1_60[60], stage1_60[61], stage1_60[62], stage1_60[63], stage1_60[64], stage1_60[65]},
      {stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35]},
      {stage2_64[5],stage2_63[9],stage2_62[14],stage2_61[14],stage2_60[20]}
   );
   gpc606_5 gpc2409 (
      {stage1_61[24], stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[6],stage2_63[10],stage2_62[15],stage2_61[15]}
   );
   gpc606_5 gpc2410 (
      {stage1_61[30], stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage2_65[1],stage2_64[7],stage2_63[11],stage2_62[16],stage2_61[16]}
   );
   gpc606_5 gpc2411 (
      {stage1_61[36], stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage2_65[2],stage2_64[8],stage2_63[12],stage2_62[17],stage2_61[17]}
   );
   gpc2135_5 gpc2412 (
      {stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39], stage1_62[40]},
      {stage1_63[18], stage1_63[19], stage1_63[20]},
      {stage1_64[0]},
      {stage1_65[0], stage1_65[1]},
      {stage2_66[0],stage2_65[3],stage2_64[9],stage2_63[13],stage2_62[18]}
   );
   gpc2135_5 gpc2413 (
      {stage1_62[41], stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45]},
      {stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage1_64[1]},
      {stage1_65[2], stage1_65[3]},
      {stage2_66[1],stage2_65[4],stage2_64[10],stage2_63[14],stage2_62[19]}
   );
   gpc2135_5 gpc2414 (
      {stage1_62[46], stage1_62[47], stage1_62[48], stage1_62[49], stage1_62[50]},
      {stage1_63[24], stage1_63[25], stage1_63[26]},
      {stage1_64[2]},
      {stage1_65[4], stage1_65[5]},
      {stage2_66[2],stage2_65[5],stage2_64[11],stage2_63[15],stage2_62[20]}
   );
   gpc2135_5 gpc2415 (
      {stage1_62[51], stage1_62[52], stage1_62[53], stage1_62[54], stage1_62[55]},
      {stage1_63[27], stage1_63[28], stage1_63[29]},
      {stage1_64[3]},
      {stage1_65[6], stage1_65[7]},
      {stage2_66[3],stage2_65[6],stage2_64[12],stage2_63[16],stage2_62[21]}
   );
   gpc2135_5 gpc2416 (
      {stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59], stage1_62[60]},
      {stage1_63[30], stage1_63[31], stage1_63[32]},
      {stage1_64[4]},
      {stage1_65[8], stage1_65[9]},
      {stage2_66[4],stage2_65[7],stage2_64[13],stage2_63[17],stage2_62[22]}
   );
   gpc2135_5 gpc2417 (
      {stage1_62[61], stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65]},
      {stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage1_64[5]},
      {stage1_65[10], stage1_65[11]},
      {stage2_66[5],stage2_65[8],stage2_64[14],stage2_63[18],stage2_62[23]}
   );
   gpc606_5 gpc2418 (
      {stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69], stage1_62[70], stage1_62[71]},
      {stage1_64[6], stage1_64[7], stage1_64[8], stage1_64[9], stage1_64[10], stage1_64[11]},
      {stage2_66[6],stage2_65[9],stage2_64[15],stage2_63[19],stage2_62[24]}
   );
   gpc606_5 gpc2419 (
      {stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75], stage1_62[76], stage1_62[77]},
      {stage1_64[12], stage1_64[13], stage1_64[14], stage1_64[15], stage1_64[16], stage1_64[17]},
      {stage2_66[7],stage2_65[10],stage2_64[16],stage2_63[20],stage2_62[25]}
   );
   gpc606_5 gpc2420 (
      {stage1_63[36], stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41]},
      {stage1_65[12], stage1_65[13], stage1_65[14], stage1_65[15], stage1_65[16], stage1_65[17]},
      {stage2_67[0],stage2_66[8],stage2_65[11],stage2_64[17],stage2_63[21]}
   );
   gpc606_5 gpc2421 (
      {stage1_63[42], stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47]},
      {stage1_65[18], stage1_65[19], stage1_65[20], stage1_65[21], stage1_65[22], stage1_65[23]},
      {stage2_67[1],stage2_66[9],stage2_65[12],stage2_64[18],stage2_63[22]}
   );
   gpc1_1 gpc2422 (
      {stage1_0[31]},
      {stage2_0[7]}
   );
   gpc1_1 gpc2423 (
      {stage1_0[32]},
      {stage2_0[8]}
   );
   gpc1_1 gpc2424 (
      {stage1_0[33]},
      {stage2_0[9]}
   );
   gpc1_1 gpc2425 (
      {stage1_1[38]},
      {stage2_1[10]}
   );
   gpc1_1 gpc2426 (
      {stage1_1[39]},
      {stage2_1[11]}
   );
   gpc1_1 gpc2427 (
      {stage1_1[40]},
      {stage2_1[12]}
   );
   gpc1_1 gpc2428 (
      {stage1_1[41]},
      {stage2_1[13]}
   );
   gpc1_1 gpc2429 (
      {stage1_1[42]},
      {stage2_1[14]}
   );
   gpc1_1 gpc2430 (
      {stage1_1[43]},
      {stage2_1[15]}
   );
   gpc1_1 gpc2431 (
      {stage1_1[44]},
      {stage2_1[16]}
   );
   gpc1_1 gpc2432 (
      {stage1_1[45]},
      {stage2_1[17]}
   );
   gpc1_1 gpc2433 (
      {stage1_1[46]},
      {stage2_1[18]}
   );
   gpc1_1 gpc2434 (
      {stage1_2[27]},
      {stage2_2[10]}
   );
   gpc1_1 gpc2435 (
      {stage1_2[28]},
      {stage2_2[11]}
   );
   gpc1_1 gpc2436 (
      {stage1_2[29]},
      {stage2_2[12]}
   );
   gpc1_1 gpc2437 (
      {stage1_2[30]},
      {stage2_2[13]}
   );
   gpc1_1 gpc2438 (
      {stage1_2[31]},
      {stage2_2[14]}
   );
   gpc1_1 gpc2439 (
      {stage1_2[32]},
      {stage2_2[15]}
   );
   gpc1_1 gpc2440 (
      {stage1_2[33]},
      {stage2_2[16]}
   );
   gpc1_1 gpc2441 (
      {stage1_2[34]},
      {stage2_2[17]}
   );
   gpc1_1 gpc2442 (
      {stage1_2[35]},
      {stage2_2[18]}
   );
   gpc1_1 gpc2443 (
      {stage1_2[36]},
      {stage2_2[19]}
   );
   gpc1_1 gpc2444 (
      {stage1_2[37]},
      {stage2_2[20]}
   );
   gpc1_1 gpc2445 (
      {stage1_2[38]},
      {stage2_2[21]}
   );
   gpc1_1 gpc2446 (
      {stage1_2[39]},
      {stage2_2[22]}
   );
   gpc1_1 gpc2447 (
      {stage1_2[40]},
      {stage2_2[23]}
   );
   gpc1_1 gpc2448 (
      {stage1_2[41]},
      {stage2_2[24]}
   );
   gpc1_1 gpc2449 (
      {stage1_2[42]},
      {stage2_2[25]}
   );
   gpc1_1 gpc2450 (
      {stage1_2[43]},
      {stage2_2[26]}
   );
   gpc1_1 gpc2451 (
      {stage1_2[44]},
      {stage2_2[27]}
   );
   gpc1_1 gpc2452 (
      {stage1_2[45]},
      {stage2_2[28]}
   );
   gpc1_1 gpc2453 (
      {stage1_2[46]},
      {stage2_2[29]}
   );
   gpc1_1 gpc2454 (
      {stage1_2[47]},
      {stage2_2[30]}
   );
   gpc1_1 gpc2455 (
      {stage1_2[48]},
      {stage2_2[31]}
   );
   gpc1_1 gpc2456 (
      {stage1_2[49]},
      {stage2_2[32]}
   );
   gpc1_1 gpc2457 (
      {stage1_2[50]},
      {stage2_2[33]}
   );
   gpc1_1 gpc2458 (
      {stage1_2[51]},
      {stage2_2[34]}
   );
   gpc1_1 gpc2459 (
      {stage1_2[52]},
      {stage2_2[35]}
   );
   gpc1_1 gpc2460 (
      {stage1_2[53]},
      {stage2_2[36]}
   );
   gpc1_1 gpc2461 (
      {stage1_2[54]},
      {stage2_2[37]}
   );
   gpc1_1 gpc2462 (
      {stage1_4[66]},
      {stage2_4[31]}
   );
   gpc1_1 gpc2463 (
      {stage1_4[67]},
      {stage2_4[32]}
   );
   gpc1_1 gpc2464 (
      {stage1_4[68]},
      {stage2_4[33]}
   );
   gpc1_1 gpc2465 (
      {stage1_4[69]},
      {stage2_4[34]}
   );
   gpc1_1 gpc2466 (
      {stage1_4[70]},
      {stage2_4[35]}
   );
   gpc1_1 gpc2467 (
      {stage1_4[71]},
      {stage2_4[36]}
   );
   gpc1_1 gpc2468 (
      {stage1_4[72]},
      {stage2_4[37]}
   );
   gpc1_1 gpc2469 (
      {stage1_4[73]},
      {stage2_4[38]}
   );
   gpc1_1 gpc2470 (
      {stage1_4[74]},
      {stage2_4[39]}
   );
   gpc1_1 gpc2471 (
      {stage1_4[75]},
      {stage2_4[40]}
   );
   gpc1_1 gpc2472 (
      {stage1_4[76]},
      {stage2_4[41]}
   );
   gpc1_1 gpc2473 (
      {stage1_4[77]},
      {stage2_4[42]}
   );
   gpc1_1 gpc2474 (
      {stage1_4[78]},
      {stage2_4[43]}
   );
   gpc1_1 gpc2475 (
      {stage1_4[79]},
      {stage2_4[44]}
   );
   gpc1_1 gpc2476 (
      {stage1_4[80]},
      {stage2_4[45]}
   );
   gpc1_1 gpc2477 (
      {stage1_4[81]},
      {stage2_4[46]}
   );
   gpc1_1 gpc2478 (
      {stage1_4[82]},
      {stage2_4[47]}
   );
   gpc1_1 gpc2479 (
      {stage1_5[109]},
      {stage2_5[30]}
   );
   gpc1_1 gpc2480 (
      {stage1_5[110]},
      {stage2_5[31]}
   );
   gpc1_1 gpc2481 (
      {stage1_5[111]},
      {stage2_5[32]}
   );
   gpc1_1 gpc2482 (
      {stage1_5[112]},
      {stage2_5[33]}
   );
   gpc1_1 gpc2483 (
      {stage1_5[113]},
      {stage2_5[34]}
   );
   gpc1_1 gpc2484 (
      {stage1_5[114]},
      {stage2_5[35]}
   );
   gpc1_1 gpc2485 (
      {stage1_7[64]},
      {stage2_7[34]}
   );
   gpc1_1 gpc2486 (
      {stage1_7[65]},
      {stage2_7[35]}
   );
   gpc1_1 gpc2487 (
      {stage1_7[66]},
      {stage2_7[36]}
   );
   gpc1_1 gpc2488 (
      {stage1_7[67]},
      {stage2_7[37]}
   );
   gpc1_1 gpc2489 (
      {stage1_7[68]},
      {stage2_7[38]}
   );
   gpc1_1 gpc2490 (
      {stage1_7[69]},
      {stage2_7[39]}
   );
   gpc1_1 gpc2491 (
      {stage1_7[70]},
      {stage2_7[40]}
   );
   gpc1_1 gpc2492 (
      {stage1_8[46]},
      {stage2_8[26]}
   );
   gpc1_1 gpc2493 (
      {stage1_8[47]},
      {stage2_8[27]}
   );
   gpc1_1 gpc2494 (
      {stage1_8[48]},
      {stage2_8[28]}
   );
   gpc1_1 gpc2495 (
      {stage1_8[49]},
      {stage2_8[29]}
   );
   gpc1_1 gpc2496 (
      {stage1_8[50]},
      {stage2_8[30]}
   );
   gpc1_1 gpc2497 (
      {stage1_8[51]},
      {stage2_8[31]}
   );
   gpc1_1 gpc2498 (
      {stage1_8[52]},
      {stage2_8[32]}
   );
   gpc1_1 gpc2499 (
      {stage1_8[53]},
      {stage2_8[33]}
   );
   gpc1_1 gpc2500 (
      {stage1_8[54]},
      {stage2_8[34]}
   );
   gpc1_1 gpc2501 (
      {stage1_8[55]},
      {stage2_8[35]}
   );
   gpc1_1 gpc2502 (
      {stage1_8[56]},
      {stage2_8[36]}
   );
   gpc1_1 gpc2503 (
      {stage1_8[57]},
      {stage2_8[37]}
   );
   gpc1_1 gpc2504 (
      {stage1_8[58]},
      {stage2_8[38]}
   );
   gpc1_1 gpc2505 (
      {stage1_8[59]},
      {stage2_8[39]}
   );
   gpc1_1 gpc2506 (
      {stage1_8[60]},
      {stage2_8[40]}
   );
   gpc1_1 gpc2507 (
      {stage1_8[61]},
      {stage2_8[41]}
   );
   gpc1_1 gpc2508 (
      {stage1_8[62]},
      {stage2_8[42]}
   );
   gpc1_1 gpc2509 (
      {stage1_8[63]},
      {stage2_8[43]}
   );
   gpc1_1 gpc2510 (
      {stage1_8[64]},
      {stage2_8[44]}
   );
   gpc1_1 gpc2511 (
      {stage1_8[65]},
      {stage2_8[45]}
   );
   gpc1_1 gpc2512 (
      {stage1_8[66]},
      {stage2_8[46]}
   );
   gpc1_1 gpc2513 (
      {stage1_8[67]},
      {stage2_8[47]}
   );
   gpc1_1 gpc2514 (
      {stage1_8[68]},
      {stage2_8[48]}
   );
   gpc1_1 gpc2515 (
      {stage1_8[69]},
      {stage2_8[49]}
   );
   gpc1_1 gpc2516 (
      {stage1_8[70]},
      {stage2_8[50]}
   );
   gpc1_1 gpc2517 (
      {stage1_8[71]},
      {stage2_8[51]}
   );
   gpc1_1 gpc2518 (
      {stage1_8[72]},
      {stage2_8[52]}
   );
   gpc1_1 gpc2519 (
      {stage1_8[73]},
      {stage2_8[53]}
   );
   gpc1_1 gpc2520 (
      {stage1_8[74]},
      {stage2_8[54]}
   );
   gpc1_1 gpc2521 (
      {stage1_8[75]},
      {stage2_8[55]}
   );
   gpc1_1 gpc2522 (
      {stage1_8[76]},
      {stage2_8[56]}
   );
   gpc1_1 gpc2523 (
      {stage1_8[77]},
      {stage2_8[57]}
   );
   gpc1_1 gpc2524 (
      {stage1_8[78]},
      {stage2_8[58]}
   );
   gpc1_1 gpc2525 (
      {stage1_8[79]},
      {stage2_8[59]}
   );
   gpc1_1 gpc2526 (
      {stage1_8[80]},
      {stage2_8[60]}
   );
   gpc1_1 gpc2527 (
      {stage1_9[54]},
      {stage2_9[22]}
   );
   gpc1_1 gpc2528 (
      {stage1_9[55]},
      {stage2_9[23]}
   );
   gpc1_1 gpc2529 (
      {stage1_9[56]},
      {stage2_9[24]}
   );
   gpc1_1 gpc2530 (
      {stage1_9[57]},
      {stage2_9[25]}
   );
   gpc1_1 gpc2531 (
      {stage1_10[79]},
      {stage2_10[25]}
   );
   gpc1_1 gpc2532 (
      {stage1_10[80]},
      {stage2_10[26]}
   );
   gpc1_1 gpc2533 (
      {stage1_10[81]},
      {stage2_10[27]}
   );
   gpc1_1 gpc2534 (
      {stage1_10[82]},
      {stage2_10[28]}
   );
   gpc1_1 gpc2535 (
      {stage1_10[83]},
      {stage2_10[29]}
   );
   gpc1_1 gpc2536 (
      {stage1_10[84]},
      {stage2_10[30]}
   );
   gpc1_1 gpc2537 (
      {stage1_10[85]},
      {stage2_10[31]}
   );
   gpc1_1 gpc2538 (
      {stage1_10[86]},
      {stage2_10[32]}
   );
   gpc1_1 gpc2539 (
      {stage1_10[87]},
      {stage2_10[33]}
   );
   gpc1_1 gpc2540 (
      {stage1_10[88]},
      {stage2_10[34]}
   );
   gpc1_1 gpc2541 (
      {stage1_10[89]},
      {stage2_10[35]}
   );
   gpc1_1 gpc2542 (
      {stage1_10[90]},
      {stage2_10[36]}
   );
   gpc1_1 gpc2543 (
      {stage1_10[91]},
      {stage2_10[37]}
   );
   gpc1_1 gpc2544 (
      {stage1_10[92]},
      {stage2_10[38]}
   );
   gpc1_1 gpc2545 (
      {stage1_10[93]},
      {stage2_10[39]}
   );
   gpc1_1 gpc2546 (
      {stage1_10[94]},
      {stage2_10[40]}
   );
   gpc1_1 gpc2547 (
      {stage1_11[74]},
      {stage2_11[32]}
   );
   gpc1_1 gpc2548 (
      {stage1_11[75]},
      {stage2_11[33]}
   );
   gpc1_1 gpc2549 (
      {stage1_11[76]},
      {stage2_11[34]}
   );
   gpc1_1 gpc2550 (
      {stage1_11[77]},
      {stage2_11[35]}
   );
   gpc1_1 gpc2551 (
      {stage1_11[78]},
      {stage2_11[36]}
   );
   gpc1_1 gpc2552 (
      {stage1_11[79]},
      {stage2_11[37]}
   );
   gpc1_1 gpc2553 (
      {stage1_11[80]},
      {stage2_11[38]}
   );
   gpc1_1 gpc2554 (
      {stage1_12[63]},
      {stage2_12[27]}
   );
   gpc1_1 gpc2555 (
      {stage1_12[64]},
      {stage2_12[28]}
   );
   gpc1_1 gpc2556 (
      {stage1_12[65]},
      {stage2_12[29]}
   );
   gpc1_1 gpc2557 (
      {stage1_12[66]},
      {stage2_12[30]}
   );
   gpc1_1 gpc2558 (
      {stage1_13[66]},
      {stage2_13[24]}
   );
   gpc1_1 gpc2559 (
      {stage1_13[67]},
      {stage2_13[25]}
   );
   gpc1_1 gpc2560 (
      {stage1_13[68]},
      {stage2_13[26]}
   );
   gpc1_1 gpc2561 (
      {stage1_13[69]},
      {stage2_13[27]}
   );
   gpc1_1 gpc2562 (
      {stage1_13[70]},
      {stage2_13[28]}
   );
   gpc1_1 gpc2563 (
      {stage1_13[71]},
      {stage2_13[29]}
   );
   gpc1_1 gpc2564 (
      {stage1_13[72]},
      {stage2_13[30]}
   );
   gpc1_1 gpc2565 (
      {stage1_13[73]},
      {stage2_13[31]}
   );
   gpc1_1 gpc2566 (
      {stage1_13[74]},
      {stage2_13[32]}
   );
   gpc1_1 gpc2567 (
      {stage1_13[75]},
      {stage2_13[33]}
   );
   gpc1_1 gpc2568 (
      {stage1_13[76]},
      {stage2_13[34]}
   );
   gpc1_1 gpc2569 (
      {stage1_13[77]},
      {stage2_13[35]}
   );
   gpc1_1 gpc2570 (
      {stage1_13[78]},
      {stage2_13[36]}
   );
   gpc1_1 gpc2571 (
      {stage1_13[79]},
      {stage2_13[37]}
   );
   gpc1_1 gpc2572 (
      {stage1_13[80]},
      {stage2_13[38]}
   );
   gpc1_1 gpc2573 (
      {stage1_13[81]},
      {stage2_13[39]}
   );
   gpc1_1 gpc2574 (
      {stage1_13[82]},
      {stage2_13[40]}
   );
   gpc1_1 gpc2575 (
      {stage1_13[83]},
      {stage2_13[41]}
   );
   gpc1_1 gpc2576 (
      {stage1_13[84]},
      {stage2_13[42]}
   );
   gpc1_1 gpc2577 (
      {stage1_13[85]},
      {stage2_13[43]}
   );
   gpc1_1 gpc2578 (
      {stage1_13[86]},
      {stage2_13[44]}
   );
   gpc1_1 gpc2579 (
      {stage1_14[10]},
      {stage2_14[22]}
   );
   gpc1_1 gpc2580 (
      {stage1_14[11]},
      {stage2_14[23]}
   );
   gpc1_1 gpc2581 (
      {stage1_14[12]},
      {stage2_14[24]}
   );
   gpc1_1 gpc2582 (
      {stage1_14[13]},
      {stage2_14[25]}
   );
   gpc1_1 gpc2583 (
      {stage1_14[14]},
      {stage2_14[26]}
   );
   gpc1_1 gpc2584 (
      {stage1_14[15]},
      {stage2_14[27]}
   );
   gpc1_1 gpc2585 (
      {stage1_14[16]},
      {stage2_14[28]}
   );
   gpc1_1 gpc2586 (
      {stage1_14[17]},
      {stage2_14[29]}
   );
   gpc1_1 gpc2587 (
      {stage1_14[18]},
      {stage2_14[30]}
   );
   gpc1_1 gpc2588 (
      {stage1_14[19]},
      {stage2_14[31]}
   );
   gpc1_1 gpc2589 (
      {stage1_14[20]},
      {stage2_14[32]}
   );
   gpc1_1 gpc2590 (
      {stage1_14[21]},
      {stage2_14[33]}
   );
   gpc1_1 gpc2591 (
      {stage1_14[22]},
      {stage2_14[34]}
   );
   gpc1_1 gpc2592 (
      {stage1_14[23]},
      {stage2_14[35]}
   );
   gpc1_1 gpc2593 (
      {stage1_14[24]},
      {stage2_14[36]}
   );
   gpc1_1 gpc2594 (
      {stage1_14[25]},
      {stage2_14[37]}
   );
   gpc1_1 gpc2595 (
      {stage1_14[26]},
      {stage2_14[38]}
   );
   gpc1_1 gpc2596 (
      {stage1_14[27]},
      {stage2_14[39]}
   );
   gpc1_1 gpc2597 (
      {stage1_14[28]},
      {stage2_14[40]}
   );
   gpc1_1 gpc2598 (
      {stage1_14[29]},
      {stage2_14[41]}
   );
   gpc1_1 gpc2599 (
      {stage1_14[30]},
      {stage2_14[42]}
   );
   gpc1_1 gpc2600 (
      {stage1_14[31]},
      {stage2_14[43]}
   );
   gpc1_1 gpc2601 (
      {stage1_14[32]},
      {stage2_14[44]}
   );
   gpc1_1 gpc2602 (
      {stage1_14[33]},
      {stage2_14[45]}
   );
   gpc1_1 gpc2603 (
      {stage1_14[34]},
      {stage2_14[46]}
   );
   gpc1_1 gpc2604 (
      {stage1_14[35]},
      {stage2_14[47]}
   );
   gpc1_1 gpc2605 (
      {stage1_14[36]},
      {stage2_14[48]}
   );
   gpc1_1 gpc2606 (
      {stage1_14[37]},
      {stage2_14[49]}
   );
   gpc1_1 gpc2607 (
      {stage1_14[38]},
      {stage2_14[50]}
   );
   gpc1_1 gpc2608 (
      {stage1_14[39]},
      {stage2_14[51]}
   );
   gpc1_1 gpc2609 (
      {stage1_14[40]},
      {stage2_14[52]}
   );
   gpc1_1 gpc2610 (
      {stage1_14[41]},
      {stage2_14[53]}
   );
   gpc1_1 gpc2611 (
      {stage1_14[42]},
      {stage2_14[54]}
   );
   gpc1_1 gpc2612 (
      {stage1_14[43]},
      {stage2_14[55]}
   );
   gpc1_1 gpc2613 (
      {stage1_14[44]},
      {stage2_14[56]}
   );
   gpc1_1 gpc2614 (
      {stage1_14[45]},
      {stage2_14[57]}
   );
   gpc1_1 gpc2615 (
      {stage1_14[46]},
      {stage2_14[58]}
   );
   gpc1_1 gpc2616 (
      {stage1_14[47]},
      {stage2_14[59]}
   );
   gpc1_1 gpc2617 (
      {stage1_14[48]},
      {stage2_14[60]}
   );
   gpc1_1 gpc2618 (
      {stage1_14[49]},
      {stage2_14[61]}
   );
   gpc1_1 gpc2619 (
      {stage1_14[50]},
      {stage2_14[62]}
   );
   gpc1_1 gpc2620 (
      {stage1_14[51]},
      {stage2_14[63]}
   );
   gpc1_1 gpc2621 (
      {stage1_14[52]},
      {stage2_14[64]}
   );
   gpc1_1 gpc2622 (
      {stage1_14[53]},
      {stage2_14[65]}
   );
   gpc1_1 gpc2623 (
      {stage1_14[54]},
      {stage2_14[66]}
   );
   gpc1_1 gpc2624 (
      {stage1_14[55]},
      {stage2_14[67]}
   );
   gpc1_1 gpc2625 (
      {stage1_14[56]},
      {stage2_14[68]}
   );
   gpc1_1 gpc2626 (
      {stage1_14[57]},
      {stage2_14[69]}
   );
   gpc1_1 gpc2627 (
      {stage1_14[58]},
      {stage2_14[70]}
   );
   gpc1_1 gpc2628 (
      {stage1_14[59]},
      {stage2_14[71]}
   );
   gpc1_1 gpc2629 (
      {stage1_14[60]},
      {stage2_14[72]}
   );
   gpc1_1 gpc2630 (
      {stage1_14[61]},
      {stage2_14[73]}
   );
   gpc1_1 gpc2631 (
      {stage1_15[86]},
      {stage2_15[25]}
   );
   gpc1_1 gpc2632 (
      {stage1_15[87]},
      {stage2_15[26]}
   );
   gpc1_1 gpc2633 (
      {stage1_15[88]},
      {stage2_15[27]}
   );
   gpc1_1 gpc2634 (
      {stage1_15[89]},
      {stage2_15[28]}
   );
   gpc1_1 gpc2635 (
      {stage1_15[90]},
      {stage2_15[29]}
   );
   gpc1_1 gpc2636 (
      {stage1_15[91]},
      {stage2_15[30]}
   );
   gpc1_1 gpc2637 (
      {stage1_15[92]},
      {stage2_15[31]}
   );
   gpc1_1 gpc2638 (
      {stage1_15[93]},
      {stage2_15[32]}
   );
   gpc1_1 gpc2639 (
      {stage1_15[94]},
      {stage2_15[33]}
   );
   gpc1_1 gpc2640 (
      {stage1_15[95]},
      {stage2_15[34]}
   );
   gpc1_1 gpc2641 (
      {stage1_15[96]},
      {stage2_15[35]}
   );
   gpc1_1 gpc2642 (
      {stage1_15[97]},
      {stage2_15[36]}
   );
   gpc1_1 gpc2643 (
      {stage1_16[42]},
      {stage2_16[21]}
   );
   gpc1_1 gpc2644 (
      {stage1_16[43]},
      {stage2_16[22]}
   );
   gpc1_1 gpc2645 (
      {stage1_16[44]},
      {stage2_16[23]}
   );
   gpc1_1 gpc2646 (
      {stage1_16[45]},
      {stage2_16[24]}
   );
   gpc1_1 gpc2647 (
      {stage1_16[46]},
      {stage2_16[25]}
   );
   gpc1_1 gpc2648 (
      {stage1_16[47]},
      {stage2_16[26]}
   );
   gpc1_1 gpc2649 (
      {stage1_16[48]},
      {stage2_16[27]}
   );
   gpc1_1 gpc2650 (
      {stage1_16[49]},
      {stage2_16[28]}
   );
   gpc1_1 gpc2651 (
      {stage1_16[50]},
      {stage2_16[29]}
   );
   gpc1_1 gpc2652 (
      {stage1_16[51]},
      {stage2_16[30]}
   );
   gpc1_1 gpc2653 (
      {stage1_16[52]},
      {stage2_16[31]}
   );
   gpc1_1 gpc2654 (
      {stage1_16[53]},
      {stage2_16[32]}
   );
   gpc1_1 gpc2655 (
      {stage1_16[54]},
      {stage2_16[33]}
   );
   gpc1_1 gpc2656 (
      {stage1_16[55]},
      {stage2_16[34]}
   );
   gpc1_1 gpc2657 (
      {stage1_16[56]},
      {stage2_16[35]}
   );
   gpc1_1 gpc2658 (
      {stage1_16[57]},
      {stage2_16[36]}
   );
   gpc1_1 gpc2659 (
      {stage1_16[58]},
      {stage2_16[37]}
   );
   gpc1_1 gpc2660 (
      {stage1_16[59]},
      {stage2_16[38]}
   );
   gpc1_1 gpc2661 (
      {stage1_16[60]},
      {stage2_16[39]}
   );
   gpc1_1 gpc2662 (
      {stage1_16[61]},
      {stage2_16[40]}
   );
   gpc1_1 gpc2663 (
      {stage1_16[62]},
      {stage2_16[41]}
   );
   gpc1_1 gpc2664 (
      {stage1_16[63]},
      {stage2_16[42]}
   );
   gpc1_1 gpc2665 (
      {stage1_16[64]},
      {stage2_16[43]}
   );
   gpc1_1 gpc2666 (
      {stage1_16[65]},
      {stage2_16[44]}
   );
   gpc1_1 gpc2667 (
      {stage1_16[66]},
      {stage2_16[45]}
   );
   gpc1_1 gpc2668 (
      {stage1_16[67]},
      {stage2_16[46]}
   );
   gpc1_1 gpc2669 (
      {stage1_17[100]},
      {stage2_17[26]}
   );
   gpc1_1 gpc2670 (
      {stage1_17[101]},
      {stage2_17[27]}
   );
   gpc1_1 gpc2671 (
      {stage1_17[102]},
      {stage2_17[28]}
   );
   gpc1_1 gpc2672 (
      {stage1_17[103]},
      {stage2_17[29]}
   );
   gpc1_1 gpc2673 (
      {stage1_17[104]},
      {stage2_17[30]}
   );
   gpc1_1 gpc2674 (
      {stage1_17[105]},
      {stage2_17[31]}
   );
   gpc1_1 gpc2675 (
      {stage1_17[106]},
      {stage2_17[32]}
   );
   gpc1_1 gpc2676 (
      {stage1_17[107]},
      {stage2_17[33]}
   );
   gpc1_1 gpc2677 (
      {stage1_17[108]},
      {stage2_17[34]}
   );
   gpc1_1 gpc2678 (
      {stage1_17[109]},
      {stage2_17[35]}
   );
   gpc1_1 gpc2679 (
      {stage1_17[110]},
      {stage2_17[36]}
   );
   gpc1_1 gpc2680 (
      {stage1_17[111]},
      {stage2_17[37]}
   );
   gpc1_1 gpc2681 (
      {stage1_17[112]},
      {stage2_17[38]}
   );
   gpc1_1 gpc2682 (
      {stage1_17[113]},
      {stage2_17[39]}
   );
   gpc1_1 gpc2683 (
      {stage1_18[47]},
      {stage2_18[27]}
   );
   gpc1_1 gpc2684 (
      {stage1_18[48]},
      {stage2_18[28]}
   );
   gpc1_1 gpc2685 (
      {stage1_18[49]},
      {stage2_18[29]}
   );
   gpc1_1 gpc2686 (
      {stage1_18[50]},
      {stage2_18[30]}
   );
   gpc1_1 gpc2687 (
      {stage1_18[51]},
      {stage2_18[31]}
   );
   gpc1_1 gpc2688 (
      {stage1_18[52]},
      {stage2_18[32]}
   );
   gpc1_1 gpc2689 (
      {stage1_18[53]},
      {stage2_18[33]}
   );
   gpc1_1 gpc2690 (
      {stage1_18[54]},
      {stage2_18[34]}
   );
   gpc1_1 gpc2691 (
      {stage1_18[55]},
      {stage2_18[35]}
   );
   gpc1_1 gpc2692 (
      {stage1_18[56]},
      {stage2_18[36]}
   );
   gpc1_1 gpc2693 (
      {stage1_18[57]},
      {stage2_18[37]}
   );
   gpc1_1 gpc2694 (
      {stage1_18[58]},
      {stage2_18[38]}
   );
   gpc1_1 gpc2695 (
      {stage1_18[59]},
      {stage2_18[39]}
   );
   gpc1_1 gpc2696 (
      {stage1_18[60]},
      {stage2_18[40]}
   );
   gpc1_1 gpc2697 (
      {stage1_18[61]},
      {stage2_18[41]}
   );
   gpc1_1 gpc2698 (
      {stage1_18[62]},
      {stage2_18[42]}
   );
   gpc1_1 gpc2699 (
      {stage1_19[48]},
      {stage2_19[28]}
   );
   gpc1_1 gpc2700 (
      {stage1_19[49]},
      {stage2_19[29]}
   );
   gpc1_1 gpc2701 (
      {stage1_19[50]},
      {stage2_19[30]}
   );
   gpc1_1 gpc2702 (
      {stage1_19[51]},
      {stage2_19[31]}
   );
   gpc1_1 gpc2703 (
      {stage1_19[52]},
      {stage2_19[32]}
   );
   gpc1_1 gpc2704 (
      {stage1_19[53]},
      {stage2_19[33]}
   );
   gpc1_1 gpc2705 (
      {stage1_19[54]},
      {stage2_19[34]}
   );
   gpc1_1 gpc2706 (
      {stage1_19[55]},
      {stage2_19[35]}
   );
   gpc1_1 gpc2707 (
      {stage1_19[56]},
      {stage2_19[36]}
   );
   gpc1_1 gpc2708 (
      {stage1_19[57]},
      {stage2_19[37]}
   );
   gpc1_1 gpc2709 (
      {stage1_19[58]},
      {stage2_19[38]}
   );
   gpc1_1 gpc2710 (
      {stage1_19[59]},
      {stage2_19[39]}
   );
   gpc1_1 gpc2711 (
      {stage1_19[60]},
      {stage2_19[40]}
   );
   gpc1_1 gpc2712 (
      {stage1_19[61]},
      {stage2_19[41]}
   );
   gpc1_1 gpc2713 (
      {stage1_19[62]},
      {stage2_19[42]}
   );
   gpc1_1 gpc2714 (
      {stage1_19[63]},
      {stage2_19[43]}
   );
   gpc1_1 gpc2715 (
      {stage1_19[64]},
      {stage2_19[44]}
   );
   gpc1_1 gpc2716 (
      {stage1_19[65]},
      {stage2_19[45]}
   );
   gpc1_1 gpc2717 (
      {stage1_19[66]},
      {stage2_19[46]}
   );
   gpc1_1 gpc2718 (
      {stage1_19[67]},
      {stage2_19[47]}
   );
   gpc1_1 gpc2719 (
      {stage1_19[68]},
      {stage2_19[48]}
   );
   gpc1_1 gpc2720 (
      {stage1_19[69]},
      {stage2_19[49]}
   );
   gpc1_1 gpc2721 (
      {stage1_19[70]},
      {stage2_19[50]}
   );
   gpc1_1 gpc2722 (
      {stage1_20[27]},
      {stage2_20[17]}
   );
   gpc1_1 gpc2723 (
      {stage1_20[28]},
      {stage2_20[18]}
   );
   gpc1_1 gpc2724 (
      {stage1_20[29]},
      {stage2_20[19]}
   );
   gpc1_1 gpc2725 (
      {stage1_20[30]},
      {stage2_20[20]}
   );
   gpc1_1 gpc2726 (
      {stage1_20[31]},
      {stage2_20[21]}
   );
   gpc1_1 gpc2727 (
      {stage1_20[32]},
      {stage2_20[22]}
   );
   gpc1_1 gpc2728 (
      {stage1_20[33]},
      {stage2_20[23]}
   );
   gpc1_1 gpc2729 (
      {stage1_20[34]},
      {stage2_20[24]}
   );
   gpc1_1 gpc2730 (
      {stage1_20[35]},
      {stage2_20[25]}
   );
   gpc1_1 gpc2731 (
      {stage1_20[36]},
      {stage2_20[26]}
   );
   gpc1_1 gpc2732 (
      {stage1_20[37]},
      {stage2_20[27]}
   );
   gpc1_1 gpc2733 (
      {stage1_20[38]},
      {stage2_20[28]}
   );
   gpc1_1 gpc2734 (
      {stage1_20[39]},
      {stage2_20[29]}
   );
   gpc1_1 gpc2735 (
      {stage1_20[40]},
      {stage2_20[30]}
   );
   gpc1_1 gpc2736 (
      {stage1_20[41]},
      {stage2_20[31]}
   );
   gpc1_1 gpc2737 (
      {stage1_20[42]},
      {stage2_20[32]}
   );
   gpc1_1 gpc2738 (
      {stage1_20[43]},
      {stage2_20[33]}
   );
   gpc1_1 gpc2739 (
      {stage1_20[44]},
      {stage2_20[34]}
   );
   gpc1_1 gpc2740 (
      {stage1_20[45]},
      {stage2_20[35]}
   );
   gpc1_1 gpc2741 (
      {stage1_20[46]},
      {stage2_20[36]}
   );
   gpc1_1 gpc2742 (
      {stage1_20[47]},
      {stage2_20[37]}
   );
   gpc1_1 gpc2743 (
      {stage1_20[48]},
      {stage2_20[38]}
   );
   gpc1_1 gpc2744 (
      {stage1_20[49]},
      {stage2_20[39]}
   );
   gpc1_1 gpc2745 (
      {stage1_20[50]},
      {stage2_20[40]}
   );
   gpc1_1 gpc2746 (
      {stage1_20[51]},
      {stage2_20[41]}
   );
   gpc1_1 gpc2747 (
      {stage1_20[52]},
      {stage2_20[42]}
   );
   gpc1_1 gpc2748 (
      {stage1_20[53]},
      {stage2_20[43]}
   );
   gpc1_1 gpc2749 (
      {stage1_20[54]},
      {stage2_20[44]}
   );
   gpc1_1 gpc2750 (
      {stage1_20[55]},
      {stage2_20[45]}
   );
   gpc1_1 gpc2751 (
      {stage1_20[56]},
      {stage2_20[46]}
   );
   gpc1_1 gpc2752 (
      {stage1_20[57]},
      {stage2_20[47]}
   );
   gpc1_1 gpc2753 (
      {stage1_20[58]},
      {stage2_20[48]}
   );
   gpc1_1 gpc2754 (
      {stage1_20[59]},
      {stage2_20[49]}
   );
   gpc1_1 gpc2755 (
      {stage1_20[60]},
      {stage2_20[50]}
   );
   gpc1_1 gpc2756 (
      {stage1_20[61]},
      {stage2_20[51]}
   );
   gpc1_1 gpc2757 (
      {stage1_20[62]},
      {stage2_20[52]}
   );
   gpc1_1 gpc2758 (
      {stage1_20[63]},
      {stage2_20[53]}
   );
   gpc1_1 gpc2759 (
      {stage1_20[64]},
      {stage2_20[54]}
   );
   gpc1_1 gpc2760 (
      {stage1_20[65]},
      {stage2_20[55]}
   );
   gpc1_1 gpc2761 (
      {stage1_20[66]},
      {stage2_20[56]}
   );
   gpc1_1 gpc2762 (
      {stage1_20[67]},
      {stage2_20[57]}
   );
   gpc1_1 gpc2763 (
      {stage1_21[48]},
      {stage2_21[17]}
   );
   gpc1_1 gpc2764 (
      {stage1_21[49]},
      {stage2_21[18]}
   );
   gpc1_1 gpc2765 (
      {stage1_21[50]},
      {stage2_21[19]}
   );
   gpc1_1 gpc2766 (
      {stage1_21[51]},
      {stage2_21[20]}
   );
   gpc1_1 gpc2767 (
      {stage1_21[52]},
      {stage2_21[21]}
   );
   gpc1_1 gpc2768 (
      {stage1_21[53]},
      {stage2_21[22]}
   );
   gpc1_1 gpc2769 (
      {stage1_21[54]},
      {stage2_21[23]}
   );
   gpc1_1 gpc2770 (
      {stage1_21[55]},
      {stage2_21[24]}
   );
   gpc1_1 gpc2771 (
      {stage1_21[56]},
      {stage2_21[25]}
   );
   gpc1_1 gpc2772 (
      {stage1_21[57]},
      {stage2_21[26]}
   );
   gpc1_1 gpc2773 (
      {stage1_21[58]},
      {stage2_21[27]}
   );
   gpc1_1 gpc2774 (
      {stage1_21[59]},
      {stage2_21[28]}
   );
   gpc1_1 gpc2775 (
      {stage1_21[60]},
      {stage2_21[29]}
   );
   gpc1_1 gpc2776 (
      {stage1_21[61]},
      {stage2_21[30]}
   );
   gpc1_1 gpc2777 (
      {stage1_21[62]},
      {stage2_21[31]}
   );
   gpc1_1 gpc2778 (
      {stage1_21[63]},
      {stage2_21[32]}
   );
   gpc1_1 gpc2779 (
      {stage1_21[64]},
      {stage2_21[33]}
   );
   gpc1_1 gpc2780 (
      {stage1_21[65]},
      {stage2_21[34]}
   );
   gpc1_1 gpc2781 (
      {stage1_21[66]},
      {stage2_21[35]}
   );
   gpc1_1 gpc2782 (
      {stage1_21[67]},
      {stage2_21[36]}
   );
   gpc1_1 gpc2783 (
      {stage1_21[68]},
      {stage2_21[37]}
   );
   gpc1_1 gpc2784 (
      {stage1_21[69]},
      {stage2_21[38]}
   );
   gpc1_1 gpc2785 (
      {stage1_21[70]},
      {stage2_21[39]}
   );
   gpc1_1 gpc2786 (
      {stage1_22[62]},
      {stage2_22[26]}
   );
   gpc1_1 gpc2787 (
      {stage1_22[63]},
      {stage2_22[27]}
   );
   gpc1_1 gpc2788 (
      {stage1_22[64]},
      {stage2_22[28]}
   );
   gpc1_1 gpc2789 (
      {stage1_22[65]},
      {stage2_22[29]}
   );
   gpc1_1 gpc2790 (
      {stage1_22[66]},
      {stage2_22[30]}
   );
   gpc1_1 gpc2791 (
      {stage1_23[127]},
      {stage2_23[31]}
   );
   gpc1_1 gpc2792 (
      {stage1_23[128]},
      {stage2_23[32]}
   );
   gpc1_1 gpc2793 (
      {stage1_23[129]},
      {stage2_23[33]}
   );
   gpc1_1 gpc2794 (
      {stage1_23[130]},
      {stage2_23[34]}
   );
   gpc1_1 gpc2795 (
      {stage1_23[131]},
      {stage2_23[35]}
   );
   gpc1_1 gpc2796 (
      {stage1_23[132]},
      {stage2_23[36]}
   );
   gpc1_1 gpc2797 (
      {stage1_23[133]},
      {stage2_23[37]}
   );
   gpc1_1 gpc2798 (
      {stage1_23[134]},
      {stage2_23[38]}
   );
   gpc1_1 gpc2799 (
      {stage1_23[135]},
      {stage2_23[39]}
   );
   gpc1_1 gpc2800 (
      {stage1_23[136]},
      {stage2_23[40]}
   );
   gpc1_1 gpc2801 (
      {stage1_23[137]},
      {stage2_23[41]}
   );
   gpc1_1 gpc2802 (
      {stage1_23[138]},
      {stage2_23[42]}
   );
   gpc1_1 gpc2803 (
      {stage1_23[139]},
      {stage2_23[43]}
   );
   gpc1_1 gpc2804 (
      {stage1_23[140]},
      {stage2_23[44]}
   );
   gpc1_1 gpc2805 (
      {stage1_23[141]},
      {stage2_23[45]}
   );
   gpc1_1 gpc2806 (
      {stage1_23[142]},
      {stage2_23[46]}
   );
   gpc1_1 gpc2807 (
      {stage1_24[69]},
      {stage2_24[32]}
   );
   gpc1_1 gpc2808 (
      {stage1_24[70]},
      {stage2_24[33]}
   );
   gpc1_1 gpc2809 (
      {stage1_24[71]},
      {stage2_24[34]}
   );
   gpc1_1 gpc2810 (
      {stage1_24[72]},
      {stage2_24[35]}
   );
   gpc1_1 gpc2811 (
      {stage1_24[73]},
      {stage2_24[36]}
   );
   gpc1_1 gpc2812 (
      {stage1_24[74]},
      {stage2_24[37]}
   );
   gpc1_1 gpc2813 (
      {stage1_24[75]},
      {stage2_24[38]}
   );
   gpc1_1 gpc2814 (
      {stage1_24[76]},
      {stage2_24[39]}
   );
   gpc1_1 gpc2815 (
      {stage1_24[77]},
      {stage2_24[40]}
   );
   gpc1_1 gpc2816 (
      {stage1_24[78]},
      {stage2_24[41]}
   );
   gpc1_1 gpc2817 (
      {stage1_24[79]},
      {stage2_24[42]}
   );
   gpc1_1 gpc2818 (
      {stage1_24[80]},
      {stage2_24[43]}
   );
   gpc1_1 gpc2819 (
      {stage1_24[81]},
      {stage2_24[44]}
   );
   gpc1_1 gpc2820 (
      {stage1_24[82]},
      {stage2_24[45]}
   );
   gpc1_1 gpc2821 (
      {stage1_25[83]},
      {stage2_25[35]}
   );
   gpc1_1 gpc2822 (
      {stage1_25[84]},
      {stage2_25[36]}
   );
   gpc1_1 gpc2823 (
      {stage1_26[54]},
      {stage2_26[35]}
   );
   gpc1_1 gpc2824 (
      {stage1_26[55]},
      {stage2_26[36]}
   );
   gpc1_1 gpc2825 (
      {stage1_26[56]},
      {stage2_26[37]}
   );
   gpc1_1 gpc2826 (
      {stage1_26[57]},
      {stage2_26[38]}
   );
   gpc1_1 gpc2827 (
      {stage1_26[58]},
      {stage2_26[39]}
   );
   gpc1_1 gpc2828 (
      {stage1_26[59]},
      {stage2_26[40]}
   );
   gpc1_1 gpc2829 (
      {stage1_26[60]},
      {stage2_26[41]}
   );
   gpc1_1 gpc2830 (
      {stage1_26[61]},
      {stage2_26[42]}
   );
   gpc1_1 gpc2831 (
      {stage1_26[62]},
      {stage2_26[43]}
   );
   gpc1_1 gpc2832 (
      {stage1_26[63]},
      {stage2_26[44]}
   );
   gpc1_1 gpc2833 (
      {stage1_26[64]},
      {stage2_26[45]}
   );
   gpc1_1 gpc2834 (
      {stage1_26[65]},
      {stage2_26[46]}
   );
   gpc1_1 gpc2835 (
      {stage1_26[66]},
      {stage2_26[47]}
   );
   gpc1_1 gpc2836 (
      {stage1_26[67]},
      {stage2_26[48]}
   );
   gpc1_1 gpc2837 (
      {stage1_26[68]},
      {stage2_26[49]}
   );
   gpc1_1 gpc2838 (
      {stage1_26[69]},
      {stage2_26[50]}
   );
   gpc1_1 gpc2839 (
      {stage1_26[70]},
      {stage2_26[51]}
   );
   gpc1_1 gpc2840 (
      {stage1_26[71]},
      {stage2_26[52]}
   );
   gpc1_1 gpc2841 (
      {stage1_27[49]},
      {stage2_27[25]}
   );
   gpc1_1 gpc2842 (
      {stage1_27[50]},
      {stage2_27[26]}
   );
   gpc1_1 gpc2843 (
      {stage1_27[51]},
      {stage2_27[27]}
   );
   gpc1_1 gpc2844 (
      {stage1_27[52]},
      {stage2_27[28]}
   );
   gpc1_1 gpc2845 (
      {stage1_27[53]},
      {stage2_27[29]}
   );
   gpc1_1 gpc2846 (
      {stage1_27[54]},
      {stage2_27[30]}
   );
   gpc1_1 gpc2847 (
      {stage1_27[55]},
      {stage2_27[31]}
   );
   gpc1_1 gpc2848 (
      {stage1_27[56]},
      {stage2_27[32]}
   );
   gpc1_1 gpc2849 (
      {stage1_27[57]},
      {stage2_27[33]}
   );
   gpc1_1 gpc2850 (
      {stage1_27[58]},
      {stage2_27[34]}
   );
   gpc1_1 gpc2851 (
      {stage1_27[59]},
      {stage2_27[35]}
   );
   gpc1_1 gpc2852 (
      {stage1_27[60]},
      {stage2_27[36]}
   );
   gpc1_1 gpc2853 (
      {stage1_27[61]},
      {stage2_27[37]}
   );
   gpc1_1 gpc2854 (
      {stage1_27[62]},
      {stage2_27[38]}
   );
   gpc1_1 gpc2855 (
      {stage1_27[63]},
      {stage2_27[39]}
   );
   gpc1_1 gpc2856 (
      {stage1_27[64]},
      {stage2_27[40]}
   );
   gpc1_1 gpc2857 (
      {stage1_27[65]},
      {stage2_27[41]}
   );
   gpc1_1 gpc2858 (
      {stage1_27[66]},
      {stage2_27[42]}
   );
   gpc1_1 gpc2859 (
      {stage1_27[67]},
      {stage2_27[43]}
   );
   gpc1_1 gpc2860 (
      {stage1_27[68]},
      {stage2_27[44]}
   );
   gpc1_1 gpc2861 (
      {stage1_27[69]},
      {stage2_27[45]}
   );
   gpc1_1 gpc2862 (
      {stage1_27[70]},
      {stage2_27[46]}
   );
   gpc1_1 gpc2863 (
      {stage1_27[71]},
      {stage2_27[47]}
   );
   gpc1_1 gpc2864 (
      {stage1_27[72]},
      {stage2_27[48]}
   );
   gpc1_1 gpc2865 (
      {stage1_27[73]},
      {stage2_27[49]}
   );
   gpc1_1 gpc2866 (
      {stage1_28[69]},
      {stage2_28[27]}
   );
   gpc1_1 gpc2867 (
      {stage1_28[70]},
      {stage2_28[28]}
   );
   gpc1_1 gpc2868 (
      {stage1_28[71]},
      {stage2_28[29]}
   );
   gpc1_1 gpc2869 (
      {stage1_28[72]},
      {stage2_28[30]}
   );
   gpc1_1 gpc2870 (
      {stage1_28[73]},
      {stage2_28[31]}
   );
   gpc1_1 gpc2871 (
      {stage1_28[74]},
      {stage2_28[32]}
   );
   gpc1_1 gpc2872 (
      {stage1_28[75]},
      {stage2_28[33]}
   );
   gpc1_1 gpc2873 (
      {stage1_28[76]},
      {stage2_28[34]}
   );
   gpc1_1 gpc2874 (
      {stage1_29[58]},
      {stage2_29[27]}
   );
   gpc1_1 gpc2875 (
      {stage1_29[59]},
      {stage2_29[28]}
   );
   gpc1_1 gpc2876 (
      {stage1_29[60]},
      {stage2_29[29]}
   );
   gpc1_1 gpc2877 (
      {stage1_29[61]},
      {stage2_29[30]}
   );
   gpc1_1 gpc2878 (
      {stage1_29[62]},
      {stage2_29[31]}
   );
   gpc1_1 gpc2879 (
      {stage1_29[63]},
      {stage2_29[32]}
   );
   gpc1_1 gpc2880 (
      {stage1_29[64]},
      {stage2_29[33]}
   );
   gpc1_1 gpc2881 (
      {stage1_29[65]},
      {stage2_29[34]}
   );
   gpc1_1 gpc2882 (
      {stage1_29[66]},
      {stage2_29[35]}
   );
   gpc1_1 gpc2883 (
      {stage1_29[67]},
      {stage2_29[36]}
   );
   gpc1_1 gpc2884 (
      {stage1_29[68]},
      {stage2_29[37]}
   );
   gpc1_1 gpc2885 (
      {stage1_29[69]},
      {stage2_29[38]}
   );
   gpc1_1 gpc2886 (
      {stage1_29[70]},
      {stage2_29[39]}
   );
   gpc1_1 gpc2887 (
      {stage1_29[71]},
      {stage2_29[40]}
   );
   gpc1_1 gpc2888 (
      {stage1_29[72]},
      {stage2_29[41]}
   );
   gpc1_1 gpc2889 (
      {stage1_29[73]},
      {stage2_29[42]}
   );
   gpc1_1 gpc2890 (
      {stage1_29[74]},
      {stage2_29[43]}
   );
   gpc1_1 gpc2891 (
      {stage1_29[75]},
      {stage2_29[44]}
   );
   gpc1_1 gpc2892 (
      {stage1_29[76]},
      {stage2_29[45]}
   );
   gpc1_1 gpc2893 (
      {stage1_29[77]},
      {stage2_29[46]}
   );
   gpc1_1 gpc2894 (
      {stage1_29[78]},
      {stage2_29[47]}
   );
   gpc1_1 gpc2895 (
      {stage1_29[79]},
      {stage2_29[48]}
   );
   gpc1_1 gpc2896 (
      {stage1_29[80]},
      {stage2_29[49]}
   );
   gpc1_1 gpc2897 (
      {stage1_30[84]},
      {stage2_30[27]}
   );
   gpc1_1 gpc2898 (
      {stage1_30[85]},
      {stage2_30[28]}
   );
   gpc1_1 gpc2899 (
      {stage1_30[86]},
      {stage2_30[29]}
   );
   gpc1_1 gpc2900 (
      {stage1_30[87]},
      {stage2_30[30]}
   );
   gpc1_1 gpc2901 (
      {stage1_30[88]},
      {stage2_30[31]}
   );
   gpc1_1 gpc2902 (
      {stage1_30[89]},
      {stage2_30[32]}
   );
   gpc1_1 gpc2903 (
      {stage1_30[90]},
      {stage2_30[33]}
   );
   gpc1_1 gpc2904 (
      {stage1_30[91]},
      {stage2_30[34]}
   );
   gpc1_1 gpc2905 (
      {stage1_30[92]},
      {stage2_30[35]}
   );
   gpc1_1 gpc2906 (
      {stage1_30[93]},
      {stage2_30[36]}
   );
   gpc1_1 gpc2907 (
      {stage1_30[94]},
      {stage2_30[37]}
   );
   gpc1_1 gpc2908 (
      {stage1_30[95]},
      {stage2_30[38]}
   );
   gpc1_1 gpc2909 (
      {stage1_30[96]},
      {stage2_30[39]}
   );
   gpc1_1 gpc2910 (
      {stage1_30[97]},
      {stage2_30[40]}
   );
   gpc1_1 gpc2911 (
      {stage1_30[98]},
      {stage2_30[41]}
   );
   gpc1_1 gpc2912 (
      {stage1_30[99]},
      {stage2_30[42]}
   );
   gpc1_1 gpc2913 (
      {stage1_30[100]},
      {stage2_30[43]}
   );
   gpc1_1 gpc2914 (
      {stage1_30[101]},
      {stage2_30[44]}
   );
   gpc1_1 gpc2915 (
      {stage1_30[102]},
      {stage2_30[45]}
   );
   gpc1_1 gpc2916 (
      {stage1_30[103]},
      {stage2_30[46]}
   );
   gpc1_1 gpc2917 (
      {stage1_30[104]},
      {stage2_30[47]}
   );
   gpc1_1 gpc2918 (
      {stage1_30[105]},
      {stage2_30[48]}
   );
   gpc1_1 gpc2919 (
      {stage1_30[106]},
      {stage2_30[49]}
   );
   gpc1_1 gpc2920 (
      {stage1_31[94]},
      {stage2_31[36]}
   );
   gpc1_1 gpc2921 (
      {stage1_31[95]},
      {stage2_31[37]}
   );
   gpc1_1 gpc2922 (
      {stage1_31[96]},
      {stage2_31[38]}
   );
   gpc1_1 gpc2923 (
      {stage1_32[68]},
      {stage2_32[37]}
   );
   gpc1_1 gpc2924 (
      {stage1_32[69]},
      {stage2_32[38]}
   );
   gpc1_1 gpc2925 (
      {stage1_32[70]},
      {stage2_32[39]}
   );
   gpc1_1 gpc2926 (
      {stage1_32[71]},
      {stage2_32[40]}
   );
   gpc1_1 gpc2927 (
      {stage1_32[72]},
      {stage2_32[41]}
   );
   gpc1_1 gpc2928 (
      {stage1_32[73]},
      {stage2_32[42]}
   );
   gpc1_1 gpc2929 (
      {stage1_32[74]},
      {stage2_32[43]}
   );
   gpc1_1 gpc2930 (
      {stage1_32[75]},
      {stage2_32[44]}
   );
   gpc1_1 gpc2931 (
      {stage1_32[76]},
      {stage2_32[45]}
   );
   gpc1_1 gpc2932 (
      {stage1_32[77]},
      {stage2_32[46]}
   );
   gpc1_1 gpc2933 (
      {stage1_32[78]},
      {stage2_32[47]}
   );
   gpc1_1 gpc2934 (
      {stage1_32[79]},
      {stage2_32[48]}
   );
   gpc1_1 gpc2935 (
      {stage1_32[80]},
      {stage2_32[49]}
   );
   gpc1_1 gpc2936 (
      {stage1_32[81]},
      {stage2_32[50]}
   );
   gpc1_1 gpc2937 (
      {stage1_32[82]},
      {stage2_32[51]}
   );
   gpc1_1 gpc2938 (
      {stage1_32[83]},
      {stage2_32[52]}
   );
   gpc1_1 gpc2939 (
      {stage1_32[84]},
      {stage2_32[53]}
   );
   gpc1_1 gpc2940 (
      {stage1_32[85]},
      {stage2_32[54]}
   );
   gpc1_1 gpc2941 (
      {stage1_32[86]},
      {stage2_32[55]}
   );
   gpc1_1 gpc2942 (
      {stage1_34[48]},
      {stage2_34[27]}
   );
   gpc1_1 gpc2943 (
      {stage1_34[49]},
      {stage2_34[28]}
   );
   gpc1_1 gpc2944 (
      {stage1_34[50]},
      {stage2_34[29]}
   );
   gpc1_1 gpc2945 (
      {stage1_34[51]},
      {stage2_34[30]}
   );
   gpc1_1 gpc2946 (
      {stage1_34[52]},
      {stage2_34[31]}
   );
   gpc1_1 gpc2947 (
      {stage1_34[53]},
      {stage2_34[32]}
   );
   gpc1_1 gpc2948 (
      {stage1_34[54]},
      {stage2_34[33]}
   );
   gpc1_1 gpc2949 (
      {stage1_34[55]},
      {stage2_34[34]}
   );
   gpc1_1 gpc2950 (
      {stage1_35[46]},
      {stage2_35[31]}
   );
   gpc1_1 gpc2951 (
      {stage1_35[47]},
      {stage2_35[32]}
   );
   gpc1_1 gpc2952 (
      {stage1_35[48]},
      {stage2_35[33]}
   );
   gpc1_1 gpc2953 (
      {stage1_35[49]},
      {stage2_35[34]}
   );
   gpc1_1 gpc2954 (
      {stage1_35[50]},
      {stage2_35[35]}
   );
   gpc1_1 gpc2955 (
      {stage1_35[51]},
      {stage2_35[36]}
   );
   gpc1_1 gpc2956 (
      {stage1_35[52]},
      {stage2_35[37]}
   );
   gpc1_1 gpc2957 (
      {stage1_35[53]},
      {stage2_35[38]}
   );
   gpc1_1 gpc2958 (
      {stage1_35[54]},
      {stage2_35[39]}
   );
   gpc1_1 gpc2959 (
      {stage1_35[55]},
      {stage2_35[40]}
   );
   gpc1_1 gpc2960 (
      {stage1_35[56]},
      {stage2_35[41]}
   );
   gpc1_1 gpc2961 (
      {stage1_35[57]},
      {stage2_35[42]}
   );
   gpc1_1 gpc2962 (
      {stage1_35[58]},
      {stage2_35[43]}
   );
   gpc1_1 gpc2963 (
      {stage1_35[59]},
      {stage2_35[44]}
   );
   gpc1_1 gpc2964 (
      {stage1_36[72]},
      {stage2_36[26]}
   );
   gpc1_1 gpc2965 (
      {stage1_36[73]},
      {stage2_36[27]}
   );
   gpc1_1 gpc2966 (
      {stage1_36[74]},
      {stage2_36[28]}
   );
   gpc1_1 gpc2967 (
      {stage1_36[75]},
      {stage2_36[29]}
   );
   gpc1_1 gpc2968 (
      {stage1_36[76]},
      {stage2_36[30]}
   );
   gpc1_1 gpc2969 (
      {stage1_36[77]},
      {stage2_36[31]}
   );
   gpc1_1 gpc2970 (
      {stage1_36[78]},
      {stage2_36[32]}
   );
   gpc1_1 gpc2971 (
      {stage1_36[79]},
      {stage2_36[33]}
   );
   gpc1_1 gpc2972 (
      {stage1_36[80]},
      {stage2_36[34]}
   );
   gpc1_1 gpc2973 (
      {stage1_36[81]},
      {stage2_36[35]}
   );
   gpc1_1 gpc2974 (
      {stage1_36[82]},
      {stage2_36[36]}
   );
   gpc1_1 gpc2975 (
      {stage1_37[117]},
      {stage2_37[31]}
   );
   gpc1_1 gpc2976 (
      {stage1_37[118]},
      {stage2_37[32]}
   );
   gpc1_1 gpc2977 (
      {stage1_37[119]},
      {stage2_37[33]}
   );
   gpc1_1 gpc2978 (
      {stage1_37[120]},
      {stage2_37[34]}
   );
   gpc1_1 gpc2979 (
      {stage1_37[121]},
      {stage2_37[35]}
   );
   gpc1_1 gpc2980 (
      {stage1_37[122]},
      {stage2_37[36]}
   );
   gpc1_1 gpc2981 (
      {stage1_37[123]},
      {stage2_37[37]}
   );
   gpc1_1 gpc2982 (
      {stage1_37[124]},
      {stage2_37[38]}
   );
   gpc1_1 gpc2983 (
      {stage1_37[125]},
      {stage2_37[39]}
   );
   gpc1_1 gpc2984 (
      {stage1_37[126]},
      {stage2_37[40]}
   );
   gpc1_1 gpc2985 (
      {stage1_37[127]},
      {stage2_37[41]}
   );
   gpc1_1 gpc2986 (
      {stage1_39[64]},
      {stage2_39[30]}
   );
   gpc1_1 gpc2987 (
      {stage1_39[65]},
      {stage2_39[31]}
   );
   gpc1_1 gpc2988 (
      {stage1_39[66]},
      {stage2_39[32]}
   );
   gpc1_1 gpc2989 (
      {stage1_39[67]},
      {stage2_39[33]}
   );
   gpc1_1 gpc2990 (
      {stage1_40[72]},
      {stage2_40[31]}
   );
   gpc1_1 gpc2991 (
      {stage1_40[73]},
      {stage2_40[32]}
   );
   gpc1_1 gpc2992 (
      {stage1_40[74]},
      {stage2_40[33]}
   );
   gpc1_1 gpc2993 (
      {stage1_40[75]},
      {stage2_40[34]}
   );
   gpc1_1 gpc2994 (
      {stage1_40[76]},
      {stage2_40[35]}
   );
   gpc1_1 gpc2995 (
      {stage1_40[77]},
      {stage2_40[36]}
   );
   gpc1_1 gpc2996 (
      {stage1_40[78]},
      {stage2_40[37]}
   );
   gpc1_1 gpc2997 (
      {stage1_40[79]},
      {stage2_40[38]}
   );
   gpc1_1 gpc2998 (
      {stage1_40[80]},
      {stage2_40[39]}
   );
   gpc1_1 gpc2999 (
      {stage1_40[81]},
      {stage2_40[40]}
   );
   gpc1_1 gpc3000 (
      {stage1_41[48]},
      {stage2_41[30]}
   );
   gpc1_1 gpc3001 (
      {stage1_41[49]},
      {stage2_41[31]}
   );
   gpc1_1 gpc3002 (
      {stage1_41[50]},
      {stage2_41[32]}
   );
   gpc1_1 gpc3003 (
      {stage1_41[51]},
      {stage2_41[33]}
   );
   gpc1_1 gpc3004 (
      {stage1_41[52]},
      {stage2_41[34]}
   );
   gpc1_1 gpc3005 (
      {stage1_41[53]},
      {stage2_41[35]}
   );
   gpc1_1 gpc3006 (
      {stage1_41[54]},
      {stage2_41[36]}
   );
   gpc1_1 gpc3007 (
      {stage1_41[55]},
      {stage2_41[37]}
   );
   gpc1_1 gpc3008 (
      {stage1_41[56]},
      {stage2_41[38]}
   );
   gpc1_1 gpc3009 (
      {stage1_41[57]},
      {stage2_41[39]}
   );
   gpc1_1 gpc3010 (
      {stage1_41[58]},
      {stage2_41[40]}
   );
   gpc1_1 gpc3011 (
      {stage1_41[59]},
      {stage2_41[41]}
   );
   gpc1_1 gpc3012 (
      {stage1_41[60]},
      {stage2_41[42]}
   );
   gpc1_1 gpc3013 (
      {stage1_41[61]},
      {stage2_41[43]}
   );
   gpc1_1 gpc3014 (
      {stage1_41[62]},
      {stage2_41[44]}
   );
   gpc1_1 gpc3015 (
      {stage1_41[63]},
      {stage2_41[45]}
   );
   gpc1_1 gpc3016 (
      {stage1_41[64]},
      {stage2_41[46]}
   );
   gpc1_1 gpc3017 (
      {stage1_41[65]},
      {stage2_41[47]}
   );
   gpc1_1 gpc3018 (
      {stage1_41[66]},
      {stage2_41[48]}
   );
   gpc1_1 gpc3019 (
      {stage1_41[67]},
      {stage2_41[49]}
   );
   gpc1_1 gpc3020 (
      {stage1_41[68]},
      {stage2_41[50]}
   );
   gpc1_1 gpc3021 (
      {stage1_41[69]},
      {stage2_41[51]}
   );
   gpc1_1 gpc3022 (
      {stage1_41[70]},
      {stage2_41[52]}
   );
   gpc1_1 gpc3023 (
      {stage1_41[71]},
      {stage2_41[53]}
   );
   gpc1_1 gpc3024 (
      {stage1_41[72]},
      {stage2_41[54]}
   );
   gpc1_1 gpc3025 (
      {stage1_41[73]},
      {stage2_41[55]}
   );
   gpc1_1 gpc3026 (
      {stage1_42[54]},
      {stage2_42[20]}
   );
   gpc1_1 gpc3027 (
      {stage1_42[55]},
      {stage2_42[21]}
   );
   gpc1_1 gpc3028 (
      {stage1_42[56]},
      {stage2_42[22]}
   );
   gpc1_1 gpc3029 (
      {stage1_42[57]},
      {stage2_42[23]}
   );
   gpc1_1 gpc3030 (
      {stage1_42[58]},
      {stage2_42[24]}
   );
   gpc1_1 gpc3031 (
      {stage1_42[59]},
      {stage2_42[25]}
   );
   gpc1_1 gpc3032 (
      {stage1_42[60]},
      {stage2_42[26]}
   );
   gpc1_1 gpc3033 (
      {stage1_42[61]},
      {stage2_42[27]}
   );
   gpc1_1 gpc3034 (
      {stage1_42[62]},
      {stage2_42[28]}
   );
   gpc1_1 gpc3035 (
      {stage1_42[63]},
      {stage2_42[29]}
   );
   gpc1_1 gpc3036 (
      {stage1_42[64]},
      {stage2_42[30]}
   );
   gpc1_1 gpc3037 (
      {stage1_42[65]},
      {stage2_42[31]}
   );
   gpc1_1 gpc3038 (
      {stage1_42[66]},
      {stage2_42[32]}
   );
   gpc1_1 gpc3039 (
      {stage1_42[67]},
      {stage2_42[33]}
   );
   gpc1_1 gpc3040 (
      {stage1_42[68]},
      {stage2_42[34]}
   );
   gpc1_1 gpc3041 (
      {stage1_42[69]},
      {stage2_42[35]}
   );
   gpc1_1 gpc3042 (
      {stage1_42[70]},
      {stage2_42[36]}
   );
   gpc1_1 gpc3043 (
      {stage1_42[71]},
      {stage2_42[37]}
   );
   gpc1_1 gpc3044 (
      {stage1_42[72]},
      {stage2_42[38]}
   );
   gpc1_1 gpc3045 (
      {stage1_42[73]},
      {stage2_42[39]}
   );
   gpc1_1 gpc3046 (
      {stage1_42[74]},
      {stage2_42[40]}
   );
   gpc1_1 gpc3047 (
      {stage1_42[75]},
      {stage2_42[41]}
   );
   gpc1_1 gpc3048 (
      {stage1_42[76]},
      {stage2_42[42]}
   );
   gpc1_1 gpc3049 (
      {stage1_42[77]},
      {stage2_42[43]}
   );
   gpc1_1 gpc3050 (
      {stage1_42[78]},
      {stage2_42[44]}
   );
   gpc1_1 gpc3051 (
      {stage1_42[79]},
      {stage2_42[45]}
   );
   gpc1_1 gpc3052 (
      {stage1_42[80]},
      {stage2_42[46]}
   );
   gpc1_1 gpc3053 (
      {stage1_42[81]},
      {stage2_42[47]}
   );
   gpc1_1 gpc3054 (
      {stage1_42[82]},
      {stage2_42[48]}
   );
   gpc1_1 gpc3055 (
      {stage1_42[83]},
      {stage2_42[49]}
   );
   gpc1_1 gpc3056 (
      {stage1_42[84]},
      {stage2_42[50]}
   );
   gpc1_1 gpc3057 (
      {stage1_42[85]},
      {stage2_42[51]}
   );
   gpc1_1 gpc3058 (
      {stage1_42[86]},
      {stage2_42[52]}
   );
   gpc1_1 gpc3059 (
      {stage1_42[87]},
      {stage2_42[53]}
   );
   gpc1_1 gpc3060 (
      {stage1_42[88]},
      {stage2_42[54]}
   );
   gpc1_1 gpc3061 (
      {stage1_42[89]},
      {stage2_42[55]}
   );
   gpc1_1 gpc3062 (
      {stage1_42[90]},
      {stage2_42[56]}
   );
   gpc1_1 gpc3063 (
      {stage1_42[91]},
      {stage2_42[57]}
   );
   gpc1_1 gpc3064 (
      {stage1_42[92]},
      {stage2_42[58]}
   );
   gpc1_1 gpc3065 (
      {stage1_42[93]},
      {stage2_42[59]}
   );
   gpc1_1 gpc3066 (
      {stage1_42[94]},
      {stage2_42[60]}
   );
   gpc1_1 gpc3067 (
      {stage1_42[95]},
      {stage2_42[61]}
   );
   gpc1_1 gpc3068 (
      {stage1_43[114]},
      {stage2_43[28]}
   );
   gpc1_1 gpc3069 (
      {stage1_43[115]},
      {stage2_43[29]}
   );
   gpc1_1 gpc3070 (
      {stage1_43[116]},
      {stage2_43[30]}
   );
   gpc1_1 gpc3071 (
      {stage1_43[117]},
      {stage2_43[31]}
   );
   gpc1_1 gpc3072 (
      {stage1_43[118]},
      {stage2_43[32]}
   );
   gpc1_1 gpc3073 (
      {stage1_43[119]},
      {stage2_43[33]}
   );
   gpc1_1 gpc3074 (
      {stage1_43[120]},
      {stage2_43[34]}
   );
   gpc1_1 gpc3075 (
      {stage1_43[121]},
      {stage2_43[35]}
   );
   gpc1_1 gpc3076 (
      {stage1_43[122]},
      {stage2_43[36]}
   );
   gpc1_1 gpc3077 (
      {stage1_43[123]},
      {stage2_43[37]}
   );
   gpc1_1 gpc3078 (
      {stage1_43[124]},
      {stage2_43[38]}
   );
   gpc1_1 gpc3079 (
      {stage1_43[125]},
      {stage2_43[39]}
   );
   gpc1_1 gpc3080 (
      {stage1_43[126]},
      {stage2_43[40]}
   );
   gpc1_1 gpc3081 (
      {stage1_43[127]},
      {stage2_43[41]}
   );
   gpc1_1 gpc3082 (
      {stage1_43[128]},
      {stage2_43[42]}
   );
   gpc1_1 gpc3083 (
      {stage1_43[129]},
      {stage2_43[43]}
   );
   gpc1_1 gpc3084 (
      {stage1_43[130]},
      {stage2_43[44]}
   );
   gpc1_1 gpc3085 (
      {stage1_43[131]},
      {stage2_43[45]}
   );
   gpc1_1 gpc3086 (
      {stage1_43[132]},
      {stage2_43[46]}
   );
   gpc1_1 gpc3087 (
      {stage1_43[133]},
      {stage2_43[47]}
   );
   gpc1_1 gpc3088 (
      {stage1_43[134]},
      {stage2_43[48]}
   );
   gpc1_1 gpc3089 (
      {stage1_43[135]},
      {stage2_43[49]}
   );
   gpc1_1 gpc3090 (
      {stage1_43[136]},
      {stage2_43[50]}
   );
   gpc1_1 gpc3091 (
      {stage1_43[137]},
      {stage2_43[51]}
   );
   gpc1_1 gpc3092 (
      {stage1_44[10]},
      {stage2_44[30]}
   );
   gpc1_1 gpc3093 (
      {stage1_44[11]},
      {stage2_44[31]}
   );
   gpc1_1 gpc3094 (
      {stage1_44[12]},
      {stage2_44[32]}
   );
   gpc1_1 gpc3095 (
      {stage1_44[13]},
      {stage2_44[33]}
   );
   gpc1_1 gpc3096 (
      {stage1_44[14]},
      {stage2_44[34]}
   );
   gpc1_1 gpc3097 (
      {stage1_44[15]},
      {stage2_44[35]}
   );
   gpc1_1 gpc3098 (
      {stage1_44[16]},
      {stage2_44[36]}
   );
   gpc1_1 gpc3099 (
      {stage1_44[17]},
      {stage2_44[37]}
   );
   gpc1_1 gpc3100 (
      {stage1_44[18]},
      {stage2_44[38]}
   );
   gpc1_1 gpc3101 (
      {stage1_44[19]},
      {stage2_44[39]}
   );
   gpc1_1 gpc3102 (
      {stage1_44[20]},
      {stage2_44[40]}
   );
   gpc1_1 gpc3103 (
      {stage1_44[21]},
      {stage2_44[41]}
   );
   gpc1_1 gpc3104 (
      {stage1_44[22]},
      {stage2_44[42]}
   );
   gpc1_1 gpc3105 (
      {stage1_44[23]},
      {stage2_44[43]}
   );
   gpc1_1 gpc3106 (
      {stage1_44[24]},
      {stage2_44[44]}
   );
   gpc1_1 gpc3107 (
      {stage1_44[25]},
      {stage2_44[45]}
   );
   gpc1_1 gpc3108 (
      {stage1_44[26]},
      {stage2_44[46]}
   );
   gpc1_1 gpc3109 (
      {stage1_44[27]},
      {stage2_44[47]}
   );
   gpc1_1 gpc3110 (
      {stage1_44[28]},
      {stage2_44[48]}
   );
   gpc1_1 gpc3111 (
      {stage1_44[29]},
      {stage2_44[49]}
   );
   gpc1_1 gpc3112 (
      {stage1_44[30]},
      {stage2_44[50]}
   );
   gpc1_1 gpc3113 (
      {stage1_44[31]},
      {stage2_44[51]}
   );
   gpc1_1 gpc3114 (
      {stage1_44[32]},
      {stage2_44[52]}
   );
   gpc1_1 gpc3115 (
      {stage1_44[33]},
      {stage2_44[53]}
   );
   gpc1_1 gpc3116 (
      {stage1_44[34]},
      {stage2_44[54]}
   );
   gpc1_1 gpc3117 (
      {stage1_44[35]},
      {stage2_44[55]}
   );
   gpc1_1 gpc3118 (
      {stage1_44[36]},
      {stage2_44[56]}
   );
   gpc1_1 gpc3119 (
      {stage1_44[37]},
      {stage2_44[57]}
   );
   gpc1_1 gpc3120 (
      {stage1_44[38]},
      {stage2_44[58]}
   );
   gpc1_1 gpc3121 (
      {stage1_44[39]},
      {stage2_44[59]}
   );
   gpc1_1 gpc3122 (
      {stage1_44[40]},
      {stage2_44[60]}
   );
   gpc1_1 gpc3123 (
      {stage1_44[41]},
      {stage2_44[61]}
   );
   gpc1_1 gpc3124 (
      {stage1_44[42]},
      {stage2_44[62]}
   );
   gpc1_1 gpc3125 (
      {stage1_44[43]},
      {stage2_44[63]}
   );
   gpc1_1 gpc3126 (
      {stage1_44[44]},
      {stage2_44[64]}
   );
   gpc1_1 gpc3127 (
      {stage1_44[45]},
      {stage2_44[65]}
   );
   gpc1_1 gpc3128 (
      {stage1_45[92]},
      {stage2_45[25]}
   );
   gpc1_1 gpc3129 (
      {stage1_46[57]},
      {stage2_46[26]}
   );
   gpc1_1 gpc3130 (
      {stage1_46[58]},
      {stage2_46[27]}
   );
   gpc1_1 gpc3131 (
      {stage1_46[59]},
      {stage2_46[28]}
   );
   gpc1_1 gpc3132 (
      {stage1_46[60]},
      {stage2_46[29]}
   );
   gpc1_1 gpc3133 (
      {stage1_46[61]},
      {stage2_46[30]}
   );
   gpc1_1 gpc3134 (
      {stage1_46[62]},
      {stage2_46[31]}
   );
   gpc1_1 gpc3135 (
      {stage1_46[63]},
      {stage2_46[32]}
   );
   gpc1_1 gpc3136 (
      {stage1_47[39]},
      {stage2_47[27]}
   );
   gpc1_1 gpc3137 (
      {stage1_47[40]},
      {stage2_47[28]}
   );
   gpc1_1 gpc3138 (
      {stage1_47[41]},
      {stage2_47[29]}
   );
   gpc1_1 gpc3139 (
      {stage1_47[42]},
      {stage2_47[30]}
   );
   gpc1_1 gpc3140 (
      {stage1_47[43]},
      {stage2_47[31]}
   );
   gpc1_1 gpc3141 (
      {stage1_47[44]},
      {stage2_47[32]}
   );
   gpc1_1 gpc3142 (
      {stage1_47[45]},
      {stage2_47[33]}
   );
   gpc1_1 gpc3143 (
      {stage1_47[46]},
      {stage2_47[34]}
   );
   gpc1_1 gpc3144 (
      {stage1_47[47]},
      {stage2_47[35]}
   );
   gpc1_1 gpc3145 (
      {stage1_47[48]},
      {stage2_47[36]}
   );
   gpc1_1 gpc3146 (
      {stage1_47[49]},
      {stage2_47[37]}
   );
   gpc1_1 gpc3147 (
      {stage1_47[50]},
      {stage2_47[38]}
   );
   gpc1_1 gpc3148 (
      {stage1_47[51]},
      {stage2_47[39]}
   );
   gpc1_1 gpc3149 (
      {stage1_47[52]},
      {stage2_47[40]}
   );
   gpc1_1 gpc3150 (
      {stage1_47[53]},
      {stage2_47[41]}
   );
   gpc1_1 gpc3151 (
      {stage1_47[54]},
      {stage2_47[42]}
   );
   gpc1_1 gpc3152 (
      {stage1_47[55]},
      {stage2_47[43]}
   );
   gpc1_1 gpc3153 (
      {stage1_47[56]},
      {stage2_47[44]}
   );
   gpc1_1 gpc3154 (
      {stage1_47[57]},
      {stage2_47[45]}
   );
   gpc1_1 gpc3155 (
      {stage1_48[66]},
      {stage2_48[18]}
   );
   gpc1_1 gpc3156 (
      {stage1_48[67]},
      {stage2_48[19]}
   );
   gpc1_1 gpc3157 (
      {stage1_48[68]},
      {stage2_48[20]}
   );
   gpc1_1 gpc3158 (
      {stage1_48[69]},
      {stage2_48[21]}
   );
   gpc1_1 gpc3159 (
      {stage1_48[70]},
      {stage2_48[22]}
   );
   gpc1_1 gpc3160 (
      {stage1_48[71]},
      {stage2_48[23]}
   );
   gpc1_1 gpc3161 (
      {stage1_49[78]},
      {stage2_49[28]}
   );
   gpc1_1 gpc3162 (
      {stage1_49[79]},
      {stage2_49[29]}
   );
   gpc1_1 gpc3163 (
      {stage1_49[80]},
      {stage2_49[30]}
   );
   gpc1_1 gpc3164 (
      {stage1_49[81]},
      {stage2_49[31]}
   );
   gpc1_1 gpc3165 (
      {stage1_49[82]},
      {stage2_49[32]}
   );
   gpc1_1 gpc3166 (
      {stage1_49[83]},
      {stage2_49[33]}
   );
   gpc1_1 gpc3167 (
      {stage1_49[84]},
      {stage2_49[34]}
   );
   gpc1_1 gpc3168 (
      {stage1_49[85]},
      {stage2_49[35]}
   );
   gpc1_1 gpc3169 (
      {stage1_49[86]},
      {stage2_49[36]}
   );
   gpc1_1 gpc3170 (
      {stage1_50[47]},
      {stage2_50[30]}
   );
   gpc1_1 gpc3171 (
      {stage1_50[48]},
      {stage2_50[31]}
   );
   gpc1_1 gpc3172 (
      {stage1_50[49]},
      {stage2_50[32]}
   );
   gpc1_1 gpc3173 (
      {stage1_50[50]},
      {stage2_50[33]}
   );
   gpc1_1 gpc3174 (
      {stage1_50[51]},
      {stage2_50[34]}
   );
   gpc1_1 gpc3175 (
      {stage1_50[52]},
      {stage2_50[35]}
   );
   gpc1_1 gpc3176 (
      {stage1_50[53]},
      {stage2_50[36]}
   );
   gpc1_1 gpc3177 (
      {stage1_50[54]},
      {stage2_50[37]}
   );
   gpc1_1 gpc3178 (
      {stage1_50[55]},
      {stage2_50[38]}
   );
   gpc1_1 gpc3179 (
      {stage1_50[56]},
      {stage2_50[39]}
   );
   gpc1_1 gpc3180 (
      {stage1_50[57]},
      {stage2_50[40]}
   );
   gpc1_1 gpc3181 (
      {stage1_51[93]},
      {stage2_51[24]}
   );
   gpc1_1 gpc3182 (
      {stage1_52[73]},
      {stage2_52[30]}
   );
   gpc1_1 gpc3183 (
      {stage1_52[74]},
      {stage2_52[31]}
   );
   gpc1_1 gpc3184 (
      {stage1_52[75]},
      {stage2_52[32]}
   );
   gpc1_1 gpc3185 (
      {stage1_52[76]},
      {stage2_52[33]}
   );
   gpc1_1 gpc3186 (
      {stage1_53[48]},
      {stage2_53[33]}
   );
   gpc1_1 gpc3187 (
      {stage1_53[49]},
      {stage2_53[34]}
   );
   gpc1_1 gpc3188 (
      {stage1_53[50]},
      {stage2_53[35]}
   );
   gpc1_1 gpc3189 (
      {stage1_53[51]},
      {stage2_53[36]}
   );
   gpc1_1 gpc3190 (
      {stage1_53[52]},
      {stage2_53[37]}
   );
   gpc1_1 gpc3191 (
      {stage1_53[53]},
      {stage2_53[38]}
   );
   gpc1_1 gpc3192 (
      {stage1_53[54]},
      {stage2_53[39]}
   );
   gpc1_1 gpc3193 (
      {stage1_53[55]},
      {stage2_53[40]}
   );
   gpc1_1 gpc3194 (
      {stage1_53[56]},
      {stage2_53[41]}
   );
   gpc1_1 gpc3195 (
      {stage1_53[57]},
      {stage2_53[42]}
   );
   gpc1_1 gpc3196 (
      {stage1_53[58]},
      {stage2_53[43]}
   );
   gpc1_1 gpc3197 (
      {stage1_53[59]},
      {stage2_53[44]}
   );
   gpc1_1 gpc3198 (
      {stage1_53[60]},
      {stage2_53[45]}
   );
   gpc1_1 gpc3199 (
      {stage1_53[61]},
      {stage2_53[46]}
   );
   gpc1_1 gpc3200 (
      {stage1_53[62]},
      {stage2_53[47]}
   );
   gpc1_1 gpc3201 (
      {stage1_53[63]},
      {stage2_53[48]}
   );
   gpc1_1 gpc3202 (
      {stage1_53[64]},
      {stage2_53[49]}
   );
   gpc1_1 gpc3203 (
      {stage1_53[65]},
      {stage2_53[50]}
   );
   gpc1_1 gpc3204 (
      {stage1_54[52]},
      {stage2_54[22]}
   );
   gpc1_1 gpc3205 (
      {stage1_54[53]},
      {stage2_54[23]}
   );
   gpc1_1 gpc3206 (
      {stage1_54[54]},
      {stage2_54[24]}
   );
   gpc1_1 gpc3207 (
      {stage1_54[55]},
      {stage2_54[25]}
   );
   gpc1_1 gpc3208 (
      {stage1_54[56]},
      {stage2_54[26]}
   );
   gpc1_1 gpc3209 (
      {stage1_54[57]},
      {stage2_54[27]}
   );
   gpc1_1 gpc3210 (
      {stage1_55[88]},
      {stage2_55[28]}
   );
   gpc1_1 gpc3211 (
      {stage1_55[89]},
      {stage2_55[29]}
   );
   gpc1_1 gpc3212 (
      {stage1_55[90]},
      {stage2_55[30]}
   );
   gpc1_1 gpc3213 (
      {stage1_55[91]},
      {stage2_55[31]}
   );
   gpc1_1 gpc3214 (
      {stage1_55[92]},
      {stage2_55[32]}
   );
   gpc1_1 gpc3215 (
      {stage1_55[93]},
      {stage2_55[33]}
   );
   gpc1_1 gpc3216 (
      {stage1_55[94]},
      {stage2_55[34]}
   );
   gpc1_1 gpc3217 (
      {stage1_55[95]},
      {stage2_55[35]}
   );
   gpc1_1 gpc3218 (
      {stage1_55[96]},
      {stage2_55[36]}
   );
   gpc1_1 gpc3219 (
      {stage1_55[97]},
      {stage2_55[37]}
   );
   gpc1_1 gpc3220 (
      {stage1_56[58]},
      {stage2_56[31]}
   );
   gpc1_1 gpc3221 (
      {stage1_56[59]},
      {stage2_56[32]}
   );
   gpc1_1 gpc3222 (
      {stage1_56[60]},
      {stage2_56[33]}
   );
   gpc1_1 gpc3223 (
      {stage1_56[61]},
      {stage2_56[34]}
   );
   gpc1_1 gpc3224 (
      {stage1_56[62]},
      {stage2_56[35]}
   );
   gpc1_1 gpc3225 (
      {stage1_56[63]},
      {stage2_56[36]}
   );
   gpc1_1 gpc3226 (
      {stage1_56[64]},
      {stage2_56[37]}
   );
   gpc1_1 gpc3227 (
      {stage1_56[65]},
      {stage2_56[38]}
   );
   gpc1_1 gpc3228 (
      {stage1_56[66]},
      {stage2_56[39]}
   );
   gpc1_1 gpc3229 (
      {stage1_56[67]},
      {stage2_56[40]}
   );
   gpc1_1 gpc3230 (
      {stage1_56[68]},
      {stage2_56[41]}
   );
   gpc1_1 gpc3231 (
      {stage1_56[69]},
      {stage2_56[42]}
   );
   gpc1_1 gpc3232 (
      {stage1_56[70]},
      {stage2_56[43]}
   );
   gpc1_1 gpc3233 (
      {stage1_56[71]},
      {stage2_56[44]}
   );
   gpc1_1 gpc3234 (
      {stage1_56[72]},
      {stage2_56[45]}
   );
   gpc1_1 gpc3235 (
      {stage1_56[73]},
      {stage2_56[46]}
   );
   gpc1_1 gpc3236 (
      {stage1_56[74]},
      {stage2_56[47]}
   );
   gpc1_1 gpc3237 (
      {stage1_56[75]},
      {stage2_56[48]}
   );
   gpc1_1 gpc3238 (
      {stage1_56[76]},
      {stage2_56[49]}
   );
   gpc1_1 gpc3239 (
      {stage1_56[77]},
      {stage2_56[50]}
   );
   gpc1_1 gpc3240 (
      {stage1_56[78]},
      {stage2_56[51]}
   );
   gpc1_1 gpc3241 (
      {stage1_56[79]},
      {stage2_56[52]}
   );
   gpc1_1 gpc3242 (
      {stage1_57[66]},
      {stage2_57[24]}
   );
   gpc1_1 gpc3243 (
      {stage1_57[67]},
      {stage2_57[25]}
   );
   gpc1_1 gpc3244 (
      {stage1_57[68]},
      {stage2_57[26]}
   );
   gpc1_1 gpc3245 (
      {stage1_57[69]},
      {stage2_57[27]}
   );
   gpc1_1 gpc3246 (
      {stage1_57[70]},
      {stage2_57[28]}
   );
   gpc1_1 gpc3247 (
      {stage1_57[71]},
      {stage2_57[29]}
   );
   gpc1_1 gpc3248 (
      {stage1_58[65]},
      {stage2_58[24]}
   );
   gpc1_1 gpc3249 (
      {stage1_58[66]},
      {stage2_58[25]}
   );
   gpc1_1 gpc3250 (
      {stage1_58[67]},
      {stage2_58[26]}
   );
   gpc1_1 gpc3251 (
      {stage1_58[68]},
      {stage2_58[27]}
   );
   gpc1_1 gpc3252 (
      {stage1_58[69]},
      {stage2_58[28]}
   );
   gpc1_1 gpc3253 (
      {stage1_58[70]},
      {stage2_58[29]}
   );
   gpc1_1 gpc3254 (
      {stage1_58[71]},
      {stage2_58[30]}
   );
   gpc1_1 gpc3255 (
      {stage1_58[72]},
      {stage2_58[31]}
   );
   gpc1_1 gpc3256 (
      {stage1_58[73]},
      {stage2_58[32]}
   );
   gpc1_1 gpc3257 (
      {stage1_59[25]},
      {stage2_59[26]}
   );
   gpc1_1 gpc3258 (
      {stage1_59[26]},
      {stage2_59[27]}
   );
   gpc1_1 gpc3259 (
      {stage1_59[27]},
      {stage2_59[28]}
   );
   gpc1_1 gpc3260 (
      {stage1_59[28]},
      {stage2_59[29]}
   );
   gpc1_1 gpc3261 (
      {stage1_59[29]},
      {stage2_59[30]}
   );
   gpc1_1 gpc3262 (
      {stage1_59[30]},
      {stage2_59[31]}
   );
   gpc1_1 gpc3263 (
      {stage1_59[31]},
      {stage2_59[32]}
   );
   gpc1_1 gpc3264 (
      {stage1_59[32]},
      {stage2_59[33]}
   );
   gpc1_1 gpc3265 (
      {stage1_59[33]},
      {stage2_59[34]}
   );
   gpc1_1 gpc3266 (
      {stage1_59[34]},
      {stage2_59[35]}
   );
   gpc1_1 gpc3267 (
      {stage1_59[35]},
      {stage2_59[36]}
   );
   gpc1_1 gpc3268 (
      {stage1_59[36]},
      {stage2_59[37]}
   );
   gpc1_1 gpc3269 (
      {stage1_59[37]},
      {stage2_59[38]}
   );
   gpc1_1 gpc3270 (
      {stage1_59[38]},
      {stage2_59[39]}
   );
   gpc1_1 gpc3271 (
      {stage1_59[39]},
      {stage2_59[40]}
   );
   gpc1_1 gpc3272 (
      {stage1_59[40]},
      {stage2_59[41]}
   );
   gpc1_1 gpc3273 (
      {stage1_59[41]},
      {stage2_59[42]}
   );
   gpc1_1 gpc3274 (
      {stage1_59[42]},
      {stage2_59[43]}
   );
   gpc1_1 gpc3275 (
      {stage1_59[43]},
      {stage2_59[44]}
   );
   gpc1_1 gpc3276 (
      {stage1_59[44]},
      {stage2_59[45]}
   );
   gpc1_1 gpc3277 (
      {stage1_59[45]},
      {stage2_59[46]}
   );
   gpc1_1 gpc3278 (
      {stage1_59[46]},
      {stage2_59[47]}
   );
   gpc1_1 gpc3279 (
      {stage1_59[47]},
      {stage2_59[48]}
   );
   gpc1_1 gpc3280 (
      {stage1_59[48]},
      {stage2_59[49]}
   );
   gpc1_1 gpc3281 (
      {stage1_59[49]},
      {stage2_59[50]}
   );
   gpc1_1 gpc3282 (
      {stage1_59[50]},
      {stage2_59[51]}
   );
   gpc1_1 gpc3283 (
      {stage1_59[51]},
      {stage2_59[52]}
   );
   gpc1_1 gpc3284 (
      {stage1_59[52]},
      {stage2_59[53]}
   );
   gpc1_1 gpc3285 (
      {stage1_59[53]},
      {stage2_59[54]}
   );
   gpc1_1 gpc3286 (
      {stage1_59[54]},
      {stage2_59[55]}
   );
   gpc1_1 gpc3287 (
      {stage1_59[55]},
      {stage2_59[56]}
   );
   gpc1_1 gpc3288 (
      {stage1_59[56]},
      {stage2_59[57]}
   );
   gpc1_1 gpc3289 (
      {stage1_59[57]},
      {stage2_59[58]}
   );
   gpc1_1 gpc3290 (
      {stage1_59[58]},
      {stage2_59[59]}
   );
   gpc1_1 gpc3291 (
      {stage1_59[59]},
      {stage2_59[60]}
   );
   gpc1_1 gpc3292 (
      {stage1_59[60]},
      {stage2_59[61]}
   );
   gpc1_1 gpc3293 (
      {stage1_59[61]},
      {stage2_59[62]}
   );
   gpc1_1 gpc3294 (
      {stage1_59[62]},
      {stage2_59[63]}
   );
   gpc1_1 gpc3295 (
      {stage1_59[63]},
      {stage2_59[64]}
   );
   gpc1_1 gpc3296 (
      {stage1_59[64]},
      {stage2_59[65]}
   );
   gpc1_1 gpc3297 (
      {stage1_59[65]},
      {stage2_59[66]}
   );
   gpc1_1 gpc3298 (
      {stage1_59[66]},
      {stage2_59[67]}
   );
   gpc1_1 gpc3299 (
      {stage1_59[67]},
      {stage2_59[68]}
   );
   gpc1_1 gpc3300 (
      {stage1_59[68]},
      {stage2_59[69]}
   );
   gpc1_1 gpc3301 (
      {stage1_59[69]},
      {stage2_59[70]}
   );
   gpc1_1 gpc3302 (
      {stage1_59[70]},
      {stage2_59[71]}
   );
   gpc1_1 gpc3303 (
      {stage1_59[71]},
      {stage2_59[72]}
   );
   gpc1_1 gpc3304 (
      {stage1_59[72]},
      {stage2_59[73]}
   );
   gpc1_1 gpc3305 (
      {stage1_59[73]},
      {stage2_59[74]}
   );
   gpc1_1 gpc3306 (
      {stage1_59[74]},
      {stage2_59[75]}
   );
   gpc1_1 gpc3307 (
      {stage1_59[75]},
      {stage2_59[76]}
   );
   gpc1_1 gpc3308 (
      {stage1_59[76]},
      {stage2_59[77]}
   );
   gpc1_1 gpc3309 (
      {stage1_59[77]},
      {stage2_59[78]}
   );
   gpc1_1 gpc3310 (
      {stage1_59[78]},
      {stage2_59[79]}
   );
   gpc1_1 gpc3311 (
      {stage1_59[79]},
      {stage2_59[80]}
   );
   gpc1_1 gpc3312 (
      {stage1_60[66]},
      {stage2_60[21]}
   );
   gpc1_1 gpc3313 (
      {stage1_61[42]},
      {stage2_61[18]}
   );
   gpc1_1 gpc3314 (
      {stage1_61[43]},
      {stage2_61[19]}
   );
   gpc1_1 gpc3315 (
      {stage1_61[44]},
      {stage2_61[20]}
   );
   gpc1_1 gpc3316 (
      {stage1_61[45]},
      {stage2_61[21]}
   );
   gpc1_1 gpc3317 (
      {stage1_61[46]},
      {stage2_61[22]}
   );
   gpc1_1 gpc3318 (
      {stage1_61[47]},
      {stage2_61[23]}
   );
   gpc1_1 gpc3319 (
      {stage1_61[48]},
      {stage2_61[24]}
   );
   gpc1_1 gpc3320 (
      {stage1_61[49]},
      {stage2_61[25]}
   );
   gpc1_1 gpc3321 (
      {stage1_61[50]},
      {stage2_61[26]}
   );
   gpc1_1 gpc3322 (
      {stage1_61[51]},
      {stage2_61[27]}
   );
   gpc1_1 gpc3323 (
      {stage1_61[52]},
      {stage2_61[28]}
   );
   gpc1_1 gpc3324 (
      {stage1_61[53]},
      {stage2_61[29]}
   );
   gpc1_1 gpc3325 (
      {stage1_61[54]},
      {stage2_61[30]}
   );
   gpc1_1 gpc3326 (
      {stage1_61[55]},
      {stage2_61[31]}
   );
   gpc1_1 gpc3327 (
      {stage1_61[56]},
      {stage2_61[32]}
   );
   gpc1_1 gpc3328 (
      {stage1_61[57]},
      {stage2_61[33]}
   );
   gpc1_1 gpc3329 (
      {stage1_61[58]},
      {stage2_61[34]}
   );
   gpc1_1 gpc3330 (
      {stage1_61[59]},
      {stage2_61[35]}
   );
   gpc1_1 gpc3331 (
      {stage1_61[60]},
      {stage2_61[36]}
   );
   gpc1_1 gpc3332 (
      {stage1_61[61]},
      {stage2_61[37]}
   );
   gpc1_1 gpc3333 (
      {stage1_61[62]},
      {stage2_61[38]}
   );
   gpc1_1 gpc3334 (
      {stage1_61[63]},
      {stage2_61[39]}
   );
   gpc1_1 gpc3335 (
      {stage1_61[64]},
      {stage2_61[40]}
   );
   gpc1_1 gpc3336 (
      {stage1_61[65]},
      {stage2_61[41]}
   );
   gpc1_1 gpc3337 (
      {stage1_61[66]},
      {stage2_61[42]}
   );
   gpc1_1 gpc3338 (
      {stage1_61[67]},
      {stage2_61[43]}
   );
   gpc1_1 gpc3339 (
      {stage1_61[68]},
      {stage2_61[44]}
   );
   gpc1_1 gpc3340 (
      {stage1_61[69]},
      {stage2_61[45]}
   );
   gpc1_1 gpc3341 (
      {stage1_61[70]},
      {stage2_61[46]}
   );
   gpc1_1 gpc3342 (
      {stage1_61[71]},
      {stage2_61[47]}
   );
   gpc1_1 gpc3343 (
      {stage1_61[72]},
      {stage2_61[48]}
   );
   gpc1_1 gpc3344 (
      {stage1_61[73]},
      {stage2_61[49]}
   );
   gpc1_1 gpc3345 (
      {stage1_61[74]},
      {stage2_61[50]}
   );
   gpc1_1 gpc3346 (
      {stage1_61[75]},
      {stage2_61[51]}
   );
   gpc1_1 gpc3347 (
      {stage1_61[76]},
      {stage2_61[52]}
   );
   gpc1_1 gpc3348 (
      {stage1_61[77]},
      {stage2_61[53]}
   );
   gpc1_1 gpc3349 (
      {stage1_61[78]},
      {stage2_61[54]}
   );
   gpc1_1 gpc3350 (
      {stage1_61[79]},
      {stage2_61[55]}
   );
   gpc1_1 gpc3351 (
      {stage1_61[80]},
      {stage2_61[56]}
   );
   gpc1_1 gpc3352 (
      {stage1_61[81]},
      {stage2_61[57]}
   );
   gpc1_1 gpc3353 (
      {stage1_61[82]},
      {stage2_61[58]}
   );
   gpc1_1 gpc3354 (
      {stage1_61[83]},
      {stage2_61[59]}
   );
   gpc1_1 gpc3355 (
      {stage1_61[84]},
      {stage2_61[60]}
   );
   gpc1_1 gpc3356 (
      {stage1_61[85]},
      {stage2_61[61]}
   );
   gpc1_1 gpc3357 (
      {stage1_61[86]},
      {stage2_61[62]}
   );
   gpc1_1 gpc3358 (
      {stage1_61[87]},
      {stage2_61[63]}
   );
   gpc1_1 gpc3359 (
      {stage1_61[88]},
      {stage2_61[64]}
   );
   gpc1_1 gpc3360 (
      {stage1_61[89]},
      {stage2_61[65]}
   );
   gpc1_1 gpc3361 (
      {stage1_61[90]},
      {stage2_61[66]}
   );
   gpc1_1 gpc3362 (
      {stage1_62[78]},
      {stage2_62[26]}
   );
   gpc1_1 gpc3363 (
      {stage1_62[79]},
      {stage2_62[27]}
   );
   gpc1_1 gpc3364 (
      {stage1_62[80]},
      {stage2_62[28]}
   );
   gpc1_1 gpc3365 (
      {stage1_62[81]},
      {stage2_62[29]}
   );
   gpc1_1 gpc3366 (
      {stage1_62[82]},
      {stage2_62[30]}
   );
   gpc1_1 gpc3367 (
      {stage1_62[83]},
      {stage2_62[31]}
   );
   gpc1_1 gpc3368 (
      {stage1_62[84]},
      {stage2_62[32]}
   );
   gpc1_1 gpc3369 (
      {stage1_62[85]},
      {stage2_62[33]}
   );
   gpc1_1 gpc3370 (
      {stage1_62[86]},
      {stage2_62[34]}
   );
   gpc1_1 gpc3371 (
      {stage1_63[48]},
      {stage2_63[23]}
   );
   gpc1_1 gpc3372 (
      {stage1_63[49]},
      {stage2_63[24]}
   );
   gpc1_1 gpc3373 (
      {stage1_63[50]},
      {stage2_63[25]}
   );
   gpc1_1 gpc3374 (
      {stage1_63[51]},
      {stage2_63[26]}
   );
   gpc1_1 gpc3375 (
      {stage1_63[52]},
      {stage2_63[27]}
   );
   gpc1_1 gpc3376 (
      {stage1_63[53]},
      {stage2_63[28]}
   );
   gpc1_1 gpc3377 (
      {stage1_63[54]},
      {stage2_63[29]}
   );
   gpc1_1 gpc3378 (
      {stage1_63[55]},
      {stage2_63[30]}
   );
   gpc1_1 gpc3379 (
      {stage1_63[56]},
      {stage2_63[31]}
   );
   gpc1_1 gpc3380 (
      {stage1_63[57]},
      {stage2_63[32]}
   );
   gpc1_1 gpc3381 (
      {stage1_63[58]},
      {stage2_63[33]}
   );
   gpc1_1 gpc3382 (
      {stage1_63[59]},
      {stage2_63[34]}
   );
   gpc1_1 gpc3383 (
      {stage1_63[60]},
      {stage2_63[35]}
   );
   gpc1_1 gpc3384 (
      {stage1_63[61]},
      {stage2_63[36]}
   );
   gpc1_1 gpc3385 (
      {stage1_63[62]},
      {stage2_63[37]}
   );
   gpc1_1 gpc3386 (
      {stage1_64[18]},
      {stage2_64[19]}
   );
   gpc1_1 gpc3387 (
      {stage1_64[19]},
      {stage2_64[20]}
   );
   gpc1_1 gpc3388 (
      {stage1_64[20]},
      {stage2_64[21]}
   );
   gpc1_1 gpc3389 (
      {stage1_64[21]},
      {stage2_64[22]}
   );
   gpc1_1 gpc3390 (
      {stage1_64[22]},
      {stage2_64[23]}
   );
   gpc1_1 gpc3391 (
      {stage1_64[23]},
      {stage2_64[24]}
   );
   gpc1_1 gpc3392 (
      {stage1_64[24]},
      {stage2_64[25]}
   );
   gpc1_1 gpc3393 (
      {stage1_64[25]},
      {stage2_64[26]}
   );
   gpc1_1 gpc3394 (
      {stage1_64[26]},
      {stage2_64[27]}
   );
   gpc1_1 gpc3395 (
      {stage1_64[27]},
      {stage2_64[28]}
   );
   gpc1_1 gpc3396 (
      {stage1_64[28]},
      {stage2_64[29]}
   );
   gpc1_1 gpc3397 (
      {stage1_64[29]},
      {stage2_64[30]}
   );
   gpc1_1 gpc3398 (
      {stage1_64[30]},
      {stage2_64[31]}
   );
   gpc1_1 gpc3399 (
      {stage1_64[31]},
      {stage2_64[32]}
   );
   gpc1_1 gpc3400 (
      {stage1_64[32]},
      {stage2_64[33]}
   );
   gpc1_1 gpc3401 (
      {stage1_64[33]},
      {stage2_64[34]}
   );
   gpc1_1 gpc3402 (
      {stage1_64[34]},
      {stage2_64[35]}
   );
   gpc1_1 gpc3403 (
      {stage1_64[35]},
      {stage2_64[36]}
   );
   gpc1_1 gpc3404 (
      {stage1_64[36]},
      {stage2_64[37]}
   );
   gpc1_1 gpc3405 (
      {stage1_64[37]},
      {stage2_64[38]}
   );
   gpc1_1 gpc3406 (
      {stage1_64[38]},
      {stage2_64[39]}
   );
   gpc1_1 gpc3407 (
      {stage1_64[39]},
      {stage2_64[40]}
   );
   gpc1_1 gpc3408 (
      {stage1_64[40]},
      {stage2_64[41]}
   );
   gpc1_1 gpc3409 (
      {stage1_64[41]},
      {stage2_64[42]}
   );
   gpc1_1 gpc3410 (
      {stage1_64[42]},
      {stage2_64[43]}
   );
   gpc1_1 gpc3411 (
      {stage1_64[43]},
      {stage2_64[44]}
   );
   gpc1_1 gpc3412 (
      {stage1_64[44]},
      {stage2_64[45]}
   );
   gpc1163_5 gpc3413 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc3414 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc3415 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc606_5 gpc3416 (
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[2],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc3417 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage2_3[1]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[3],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc3418 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[2]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[4],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc615_5 gpc3419 (
      {stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_3[3]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[5],stage3_4[6],stage3_3[6],stage3_2[6]}
   );
   gpc615_5 gpc3420 (
      {stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8]},
      {stage2_4[36]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[6],stage3_5[6],stage3_4[7],stage3_3[7]}
   );
   gpc615_5 gpc3421 (
      {stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[37]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[7],stage3_5[7],stage3_4[8],stage3_3[8]}
   );
   gpc615_5 gpc3422 (
      {stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage2_4[38]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[8],stage3_5[8],stage3_4[9],stage3_3[9]}
   );
   gpc606_5 gpc3423 (
      {stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42], stage2_4[43], stage2_4[44]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[9],stage3_5[9],stage3_4[10]}
   );
   gpc606_5 gpc3424 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[1],stage3_7[4],stage3_6[10],stage3_5[10]}
   );
   gpc606_5 gpc3425 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[2],stage3_7[5],stage3_6[11],stage3_5[11]}
   );
   gpc606_5 gpc3426 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[2],stage3_8[3],stage3_7[6],stage3_6[12]}
   );
   gpc606_5 gpc3427 (
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[3],stage3_8[4],stage3_7[7],stage3_6[13]}
   );
   gpc606_5 gpc3428 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[4],stage3_8[5],stage3_7[8],stage3_6[14]}
   );
   gpc207_4 gpc3429 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18]},
      {stage2_9[0], stage2_9[1]},
      {stage3_10[3],stage3_9[5],stage3_8[6],stage3_7[9]}
   );
   gpc207_4 gpc3430 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25]},
      {stage2_9[2], stage2_9[3]},
      {stage3_10[4],stage3_9[6],stage3_8[7],stage3_7[10]}
   );
   gpc606_5 gpc3431 (
      {stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage2_9[4], stage2_9[5], stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9]},
      {stage3_11[0],stage3_10[5],stage3_9[7],stage3_8[8],stage3_7[11]}
   );
   gpc615_5 gpc3432 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[18]},
      {stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15]},
      {stage3_11[1],stage3_10[6],stage3_9[8],stage3_8[9],stage3_7[12]}
   );
   gpc606_5 gpc3433 (
      {stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[7],stage3_9[9],stage3_8[10]}
   );
   gpc606_5 gpc3434 (
      {stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[3],stage3_10[8],stage3_9[10],stage3_8[11]}
   );
   gpc606_5 gpc3435 (
      {stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[4],stage3_10[9],stage3_9[11],stage3_8[12]}
   );
   gpc606_5 gpc3436 (
      {stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[5],stage3_10[10],stage3_9[12],stage3_8[13]}
   );
   gpc606_5 gpc3437 (
      {stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47], stage2_8[48]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[6],stage3_10[11],stage3_9[13],stage3_8[14]}
   );
   gpc606_5 gpc3438 (
      {stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[7],stage3_10[12],stage3_9[14],stage3_8[15]}
   );
   gpc606_5 gpc3439 (
      {stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59], stage2_8[60]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], 1'b0},
      {stage3_12[6],stage3_11[8],stage3_10[13],stage3_9[15],stage3_8[16]}
   );
   gpc606_5 gpc3440 (
      {stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[7],stage3_11[9],stage3_10[14],stage3_9[16]}
   );
   gpc606_5 gpc3441 (
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[1],stage3_12[8],stage3_11[10]}
   );
   gpc606_5 gpc3442 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[2],stage3_12[9],stage3_11[11]}
   );
   gpc606_5 gpc3443 (
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[3],stage3_12[10],stage3_11[12]}
   );
   gpc606_5 gpc3444 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[3],stage3_13[4],stage3_12[11],stage3_11[13]}
   );
   gpc606_5 gpc3445 (
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[4],stage3_13[5],stage3_12[12],stage3_11[14]}
   );
   gpc606_5 gpc3446 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[5],stage3_14[5],stage3_13[6],stage3_12[13]}
   );
   gpc606_5 gpc3447 (
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[6],stage3_14[6],stage3_13[7],stage3_12[14]}
   );
   gpc606_5 gpc3448 (
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[7],stage3_14[7],stage3_13[8],stage3_12[15]}
   );
   gpc606_5 gpc3449 (
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[8],stage3_14[8],stage3_13[9],stage3_12[16]}
   );
   gpc606_5 gpc3450 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[9],stage3_14[9],stage3_13[10]}
   );
   gpc615_5 gpc3451 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28]},
      {stage2_15[6]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[1],stage3_16[5],stage3_15[10],stage3_14[10]}
   );
   gpc615_5 gpc3452 (
      {stage2_14[29], stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33]},
      {stage2_15[7]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[2],stage3_16[6],stage3_15[11],stage3_14[11]}
   );
   gpc615_5 gpc3453 (
      {stage2_14[34], stage2_14[35], stage2_14[36], stage2_14[37], stage2_14[38]},
      {stage2_15[8]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[3],stage3_16[7],stage3_15[12],stage3_14[12]}
   );
   gpc615_5 gpc3454 (
      {stage2_14[39], stage2_14[40], stage2_14[41], stage2_14[42], stage2_14[43]},
      {stage2_15[9]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[4],stage3_16[8],stage3_15[13],stage3_14[13]}
   );
   gpc615_5 gpc3455 (
      {stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47], stage2_14[48]},
      {stage2_15[10]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[5],stage3_16[9],stage3_15[14],stage3_14[14]}
   );
   gpc615_5 gpc3456 (
      {stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage2_15[11]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[6],stage3_16[10],stage3_15[15],stage3_14[15]}
   );
   gpc615_5 gpc3457 (
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16]},
      {stage2_16[36]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[6],stage3_17[7],stage3_16[11],stage3_15[16]}
   );
   gpc606_5 gpc3458 (
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[1],stage3_18[7],stage3_17[8]}
   );
   gpc606_5 gpc3459 (
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[1],stage3_19[2],stage3_18[8],stage3_17[9]}
   );
   gpc606_5 gpc3460 (
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[2],stage3_19[3],stage3_18[9],stage3_17[10]}
   );
   gpc606_5 gpc3461 (
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage3_21[3],stage3_20[3],stage3_19[4],stage3_18[10],stage3_17[11]}
   );
   gpc606_5 gpc3462 (
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage2_19[24], stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage3_21[4],stage3_20[4],stage3_19[5],stage3_18[11],stage3_17[12]}
   );
   gpc615_5 gpc3463 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4]},
      {stage2_19[30]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[5],stage3_20[5],stage3_19[6],stage3_18[12]}
   );
   gpc615_5 gpc3464 (
      {stage2_18[5], stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9]},
      {stage2_19[31]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[6],stage3_20[6],stage3_19[7],stage3_18[13]}
   );
   gpc615_5 gpc3465 (
      {stage2_18[10], stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14]},
      {stage2_19[32]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[7],stage3_20[7],stage3_19[8],stage3_18[14]}
   );
   gpc615_5 gpc3466 (
      {stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19]},
      {stage2_19[33]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[8],stage3_20[8],stage3_19[9],stage3_18[15]}
   );
   gpc615_5 gpc3467 (
      {stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24]},
      {stage2_19[34]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[9],stage3_20[9],stage3_19[10],stage3_18[16]}
   );
   gpc615_5 gpc3468 (
      {stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage2_19[35]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[10],stage3_20[10],stage3_19[11],stage3_18[17]}
   );
   gpc615_5 gpc3469 (
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34]},
      {stage2_19[36]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[11],stage3_20[11],stage3_19[12],stage3_18[18]}
   );
   gpc615_5 gpc3470 (
      {stage2_18[35], stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39]},
      {stage2_19[37]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[12],stage3_20[12],stage3_19[13],stage3_18[19]}
   );
   gpc615_5 gpc3471 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4]},
      {stage2_22[0]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[8],stage3_21[13]}
   );
   gpc615_5 gpc3472 (
      {stage2_21[5], stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9]},
      {stage2_22[1]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[9],stage3_21[14]}
   );
   gpc615_5 gpc3473 (
      {stage2_21[10], stage2_21[11], stage2_21[12], stage2_21[13], stage2_21[14]},
      {stage2_22[2]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[10],stage3_21[15]}
   );
   gpc615_5 gpc3474 (
      {stage2_21[15], stage2_21[16], stage2_21[17], stage2_21[18], stage2_21[19]},
      {stage2_22[3]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[11],stage3_21[16]}
   );
   gpc615_5 gpc3475 (
      {stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23], stage2_21[24]},
      {stage2_22[4]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[12],stage3_21[17]}
   );
   gpc615_5 gpc3476 (
      {stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage2_22[5]},
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage3_25[5],stage3_24[5],stage3_23[5],stage3_22[13],stage3_21[18]}
   );
   gpc615_5 gpc3477 (
      {stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33], stage2_21[34]},
      {stage2_22[6]},
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage3_25[6],stage3_24[6],stage3_23[6],stage3_22[14],stage3_21[19]}
   );
   gpc615_5 gpc3478 (
      {stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage2_23[42]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[7],stage3_24[7],stage3_23[7],stage3_22[15]}
   );
   gpc615_5 gpc3479 (
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16]},
      {stage2_23[43]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[8],stage3_24[8],stage3_23[8],stage3_22[16]}
   );
   gpc615_5 gpc3480 (
      {stage2_22[17], stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21]},
      {stage2_23[44]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[9],stage3_24[9],stage3_23[9],stage3_22[17]}
   );
   gpc615_5 gpc3481 (
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[3],stage3_25[10],stage3_24[10]}
   );
   gpc615_5 gpc3482 (
      {stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27]},
      {stage2_25[1]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[1],stage3_26[4],stage3_25[11],stage3_24[11]}
   );
   gpc615_5 gpc3483 (
      {stage2_24[28], stage2_24[29], stage2_24[30], stage2_24[31], stage2_24[32]},
      {stage2_25[2]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[2],stage3_26[5],stage3_25[12],stage3_24[12]}
   );
   gpc606_5 gpc3484 (
      {stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6], stage2_25[7], stage2_25[8]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[3],stage3_27[3],stage3_26[6],stage3_25[13]}
   );
   gpc606_5 gpc3485 (
      {stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12], stage2_25[13], stage2_25[14]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[4],stage3_27[4],stage3_26[7],stage3_25[14]}
   );
   gpc606_5 gpc3486 (
      {stage2_25[15], stage2_25[16], stage2_25[17], stage2_25[18], stage2_25[19], stage2_25[20]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[5],stage3_27[5],stage3_26[8],stage3_25[15]}
   );
   gpc606_5 gpc3487 (
      {stage2_25[21], stage2_25[22], stage2_25[23], stage2_25[24], stage2_25[25], stage2_25[26]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[6],stage3_27[6],stage3_26[9],stage3_25[16]}
   );
   gpc606_5 gpc3488 (
      {stage2_25[27], stage2_25[28], stage2_25[29], stage2_25[30], stage2_25[31], stage2_25[32]},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[7],stage3_27[7],stage3_26[10],stage3_25[17]}
   );
   gpc207_4 gpc3489 (
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24]},
      {stage2_28[0], stage2_28[1]},
      {stage3_29[5],stage3_28[8],stage3_27[8],stage3_26[11]}
   );
   gpc207_4 gpc3490 (
      {stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31]},
      {stage2_28[2], stage2_28[3]},
      {stage3_29[6],stage3_28[9],stage3_27[9],stage3_26[12]}
   );
   gpc207_4 gpc3491 (
      {stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38]},
      {stage2_28[4], stage2_28[5]},
      {stage3_29[7],stage3_28[10],stage3_27[10],stage3_26[13]}
   );
   gpc207_4 gpc3492 (
      {stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45]},
      {stage2_28[6], stage2_28[7]},
      {stage3_29[8],stage3_28[11],stage3_27[11],stage3_26[14]}
   );
   gpc207_4 gpc3493 (
      {stage2_26[46], stage2_26[47], stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52]},
      {stage2_28[8], stage2_28[9]},
      {stage3_29[9],stage3_28[12],stage3_27[12],stage3_26[15]}
   );
   gpc606_5 gpc3494 (
      {stage2_27[30], stage2_27[31], stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[0],stage3_29[10],stage3_28[13],stage3_27[13]}
   );
   gpc606_5 gpc3495 (
      {stage2_27[36], stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[1],stage3_29[11],stage3_28[14],stage3_27[14]}
   );
   gpc615_5 gpc3496 (
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46]},
      {stage2_28[10]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[2],stage3_29[12],stage3_28[15],stage3_27[15]}
   );
   gpc606_5 gpc3497 (
      {stage2_28[11], stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[3],stage3_30[3],stage3_29[13],stage3_28[16]}
   );
   gpc606_5 gpc3498 (
      {stage2_28[17], stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[4],stage3_30[4],stage3_29[14],stage3_28[17]}
   );
   gpc606_5 gpc3499 (
      {stage2_28[23], stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[5],stage3_30[5],stage3_29[15],stage3_28[18]}
   );
   gpc606_5 gpc3500 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[6],stage3_30[6],stage3_29[16],stage3_28[19]}
   );
   gpc606_5 gpc3501 (
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[4],stage3_31[7],stage3_30[7],stage3_29[17]}
   );
   gpc606_5 gpc3502 (
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[5],stage3_31[8],stage3_30[8],stage3_29[18]}
   );
   gpc606_5 gpc3503 (
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[6],stage3_31[9],stage3_30[9],stage3_29[19]}
   );
   gpc606_5 gpc3504 (
      {stage2_29[36], stage2_29[37], stage2_29[38], stage2_29[39], stage2_29[40], stage2_29[41]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[3],stage3_32[7],stage3_31[10],stage3_30[10],stage3_29[20]}
   );
   gpc606_5 gpc3505 (
      {stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[4],stage3_32[8],stage3_31[11],stage3_30[11],stage3_29[21]}
   );
   gpc615_5 gpc3506 (
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28]},
      {stage2_31[30]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[5],stage3_32[9],stage3_31[12],stage3_30[12]}
   );
   gpc615_5 gpc3507 (
      {stage2_30[29], stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33]},
      {stage2_31[31]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[6],stage3_32[10],stage3_31[13],stage3_30[13]}
   );
   gpc615_5 gpc3508 (
      {stage2_30[34], stage2_30[35], stage2_30[36], stage2_30[37], stage2_30[38]},
      {stage2_31[32]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[7],stage3_32[11],stage3_31[14],stage3_30[14]}
   );
   gpc606_5 gpc3509 (
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[0],stage3_34[3],stage3_33[8],stage3_32[12]}
   );
   gpc606_5 gpc3510 (
      {stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[1],stage3_34[4],stage3_33[9],stage3_32[13]}
   );
   gpc606_5 gpc3511 (
      {stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[2],stage3_34[5],stage3_33[10],stage3_32[14]}
   );
   gpc7_3 gpc3512 (
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5], stage2_33[6]},
      {stage3_35[3],stage3_34[6],stage3_33[11]}
   );
   gpc7_3 gpc3513 (
      {stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11], stage2_33[12], stage2_33[13]},
      {stage3_35[4],stage3_34[7],stage3_33[12]}
   );
   gpc7_3 gpc3514 (
      {stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17], stage2_33[18], stage2_33[19], stage2_33[20]},
      {stage3_35[5],stage3_34[8],stage3_33[13]}
   );
   gpc7_3 gpc3515 (
      {stage2_33[21], stage2_33[22], stage2_33[23], stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27]},
      {stage3_35[6],stage3_34[9],stage3_33[14]}
   );
   gpc615_5 gpc3516 (
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22]},
      {stage2_35[0]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[0],stage3_36[3],stage3_35[7],stage3_34[10]}
   );
   gpc606_5 gpc3517 (
      {stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5], stage2_35[6]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[1],stage3_37[1],stage3_36[4],stage3_35[8]}
   );
   gpc606_5 gpc3518 (
      {stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11], stage2_35[12]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage3_39[1],stage3_38[2],stage3_37[2],stage3_36[5],stage3_35[9]}
   );
   gpc615_5 gpc3519 (
      {stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16], stage2_35[17]},
      {stage2_36[6]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage3_39[2],stage3_38[3],stage3_37[3],stage3_36[6],stage3_35[10]}
   );
   gpc615_5 gpc3520 (
      {stage2_35[18], stage2_35[19], stage2_35[20], stage2_35[21], stage2_35[22]},
      {stage2_36[7]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[3],stage3_38[4],stage3_37[4],stage3_36[7],stage3_35[11]}
   );
   gpc615_5 gpc3521 (
      {stage2_35[23], stage2_35[24], stage2_35[25], stage2_35[26], stage2_35[27]},
      {stage2_36[8]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[4],stage3_38[5],stage3_37[5],stage3_36[8],stage3_35[12]}
   );
   gpc615_5 gpc3522 (
      {stage2_35[28], stage2_35[29], stage2_35[30], stage2_35[31], stage2_35[32]},
      {stage2_36[9]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[5],stage3_38[6],stage3_37[6],stage3_36[9],stage3_35[13]}
   );
   gpc606_5 gpc3523 (
      {stage2_36[10], stage2_36[11], stage2_36[12], stage2_36[13], stage2_36[14], stage2_36[15]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[6],stage3_38[7],stage3_37[7],stage3_36[10]}
   );
   gpc606_5 gpc3524 (
      {stage2_36[16], stage2_36[17], stage2_36[18], stage2_36[19], stage2_36[20], stage2_36[21]},
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11]},
      {stage3_40[1],stage3_39[7],stage3_38[8],stage3_37[8],stage3_36[11]}
   );
   gpc606_5 gpc3525 (
      {stage2_36[22], stage2_36[23], stage2_36[24], stage2_36[25], stage2_36[26], stage2_36[27]},
      {stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17]},
      {stage3_40[2],stage3_39[8],stage3_38[9],stage3_37[9],stage3_36[12]}
   );
   gpc606_5 gpc3526 (
      {stage2_36[28], stage2_36[29], stage2_36[30], stage2_36[31], stage2_36[32], stage2_36[33]},
      {stage2_38[18], stage2_38[19], stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23]},
      {stage3_40[3],stage3_39[9],stage3_38[10],stage3_37[10],stage3_36[13]}
   );
   gpc606_5 gpc3527 (
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[4],stage3_39[10],stage3_38[11],stage3_37[11]}
   );
   gpc615_5 gpc3528 (
      {stage2_38[24], stage2_38[25], stage2_38[26], stage2_38[27], stage2_38[28]},
      {stage2_39[6]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[1],stage3_40[5],stage3_39[11],stage3_38[12]}
   );
   gpc615_5 gpc3529 (
      {stage2_38[29], stage2_38[30], stage2_38[31], stage2_38[32], 1'b0},
      {stage2_39[7]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[2],stage3_40[6],stage3_39[12],stage3_38[13]}
   );
   gpc606_5 gpc3530 (
      {stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11], stage2_39[12], stage2_39[13]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[2],stage3_41[3],stage3_40[7],stage3_39[13]}
   );
   gpc606_5 gpc3531 (
      {stage2_39[14], stage2_39[15], stage2_39[16], stage2_39[17], stage2_39[18], stage2_39[19]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[3],stage3_41[4],stage3_40[8],stage3_39[14]}
   );
   gpc606_5 gpc3532 (
      {stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23], stage2_39[24], stage2_39[25]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[4],stage3_41[5],stage3_40[9],stage3_39[15]}
   );
   gpc606_5 gpc3533 (
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[3],stage3_42[5],stage3_41[6],stage3_40[10]}
   );
   gpc606_5 gpc3534 (
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[4],stage3_42[6],stage3_41[7],stage3_40[11]}
   );
   gpc606_5 gpc3535 (
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage2_42[12], stage2_42[13], stage2_42[14], stage2_42[15], stage2_42[16], stage2_42[17]},
      {stage3_44[2],stage3_43[5],stage3_42[7],stage3_41[8],stage3_40[12]}
   );
   gpc606_5 gpc3536 (
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage2_43[0], stage2_43[1], stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5]},
      {stage3_45[0],stage3_44[3],stage3_43[6],stage3_42[8],stage3_41[9]}
   );
   gpc606_5 gpc3537 (
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage2_43[6], stage2_43[7], stage2_43[8], stage2_43[9], stage2_43[10], stage2_43[11]},
      {stage3_45[1],stage3_44[4],stage3_43[7],stage3_42[9],stage3_41[10]}
   );
   gpc615_5 gpc3538 (
      {stage2_41[30], stage2_41[31], stage2_41[32], stage2_41[33], stage2_41[34]},
      {stage2_42[18]},
      {stage2_43[12], stage2_43[13], stage2_43[14], stage2_43[15], stage2_43[16], stage2_43[17]},
      {stage3_45[2],stage3_44[5],stage3_43[8],stage3_42[10],stage3_41[11]}
   );
   gpc615_5 gpc3539 (
      {stage2_41[35], stage2_41[36], stage2_41[37], stage2_41[38], stage2_41[39]},
      {stage2_42[19]},
      {stage2_43[18], stage2_43[19], stage2_43[20], stage2_43[21], stage2_43[22], stage2_43[23]},
      {stage3_45[3],stage3_44[6],stage3_43[9],stage3_42[11],stage3_41[12]}
   );
   gpc615_5 gpc3540 (
      {stage2_41[40], stage2_41[41], stage2_41[42], stage2_41[43], stage2_41[44]},
      {stage2_42[20]},
      {stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27], stage2_43[28], stage2_43[29]},
      {stage3_45[4],stage3_44[7],stage3_43[10],stage3_42[12],stage3_41[13]}
   );
   gpc615_5 gpc3541 (
      {stage2_42[21], stage2_42[22], stage2_42[23], stage2_42[24], stage2_42[25]},
      {stage2_43[30]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[5],stage3_44[8],stage3_43[11],stage3_42[13]}
   );
   gpc615_5 gpc3542 (
      {stage2_42[26], stage2_42[27], stage2_42[28], stage2_42[29], stage2_42[30]},
      {stage2_43[31]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[6],stage3_44[9],stage3_43[12],stage3_42[14]}
   );
   gpc615_5 gpc3543 (
      {stage2_42[31], stage2_42[32], stage2_42[33], stage2_42[34], stage2_42[35]},
      {stage2_43[32]},
      {stage2_44[12], stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17]},
      {stage3_46[2],stage3_45[7],stage3_44[10],stage3_43[13],stage3_42[15]}
   );
   gpc615_5 gpc3544 (
      {stage2_42[36], stage2_42[37], stage2_42[38], stage2_42[39], stage2_42[40]},
      {stage2_43[33]},
      {stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23]},
      {stage3_46[3],stage3_45[8],stage3_44[11],stage3_43[14],stage3_42[16]}
   );
   gpc615_5 gpc3545 (
      {stage2_42[41], stage2_42[42], stage2_42[43], stage2_42[44], stage2_42[45]},
      {stage2_43[34]},
      {stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage3_46[4],stage3_45[9],stage3_44[12],stage3_43[15],stage3_42[17]}
   );
   gpc615_5 gpc3546 (
      {stage2_42[46], stage2_42[47], stage2_42[48], stage2_42[49], stage2_42[50]},
      {stage2_43[35]},
      {stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33], stage2_44[34], stage2_44[35]},
      {stage3_46[5],stage3_45[10],stage3_44[13],stage3_43[16],stage3_42[18]}
   );
   gpc615_5 gpc3547 (
      {stage2_42[51], stage2_42[52], stage2_42[53], stage2_42[54], stage2_42[55]},
      {stage2_43[36]},
      {stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39], stage2_44[40], stage2_44[41]},
      {stage3_46[6],stage3_45[11],stage3_44[14],stage3_43[17],stage3_42[19]}
   );
   gpc615_5 gpc3548 (
      {stage2_43[37], stage2_43[38], stage2_43[39], stage2_43[40], stage2_43[41]},
      {stage2_44[42]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[7],stage3_45[12],stage3_44[15],stage3_43[18]}
   );
   gpc615_5 gpc3549 (
      {stage2_43[42], stage2_43[43], stage2_43[44], stage2_43[45], stage2_43[46]},
      {stage2_44[43]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[8],stage3_45[13],stage3_44[16],stage3_43[19]}
   );
   gpc615_5 gpc3550 (
      {stage2_43[47], stage2_43[48], stage2_43[49], stage2_43[50], stage2_43[51]},
      {stage2_44[44]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[9],stage3_45[14],stage3_44[17],stage3_43[20]}
   );
   gpc615_5 gpc3551 (
      {stage2_44[45], stage2_44[46], stage2_44[47], stage2_44[48], stage2_44[49]},
      {stage2_45[18]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[3],stage3_46[10],stage3_45[15],stage3_44[18]}
   );
   gpc615_5 gpc3552 (
      {stage2_44[50], stage2_44[51], stage2_44[52], stage2_44[53], stage2_44[54]},
      {stage2_45[19]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[4],stage3_46[11],stage3_45[16],stage3_44[19]}
   );
   gpc606_5 gpc3553 (
      {stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23], stage2_45[24], stage2_45[25]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[2],stage3_47[5],stage3_46[12],stage3_45[17]}
   );
   gpc606_5 gpc3554 (
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[1],stage3_48[3],stage3_47[6],stage3_46[13]}
   );
   gpc1325_5 gpc3555 (
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22]},
      {stage2_47[6], stage2_47[7]},
      {stage2_48[6], stage2_48[7], stage2_48[8]},
      {stage2_49[0]},
      {stage3_50[1],stage3_49[2],stage3_48[4],stage3_47[7],stage3_46[14]}
   );
   gpc1325_5 gpc3556 (
      {stage2_46[23], stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27]},
      {stage2_47[8], stage2_47[9]},
      {stage2_48[9], stage2_48[10], stage2_48[11]},
      {stage2_49[1]},
      {stage3_50[2],stage3_49[3],stage3_48[5],stage3_47[8],stage3_46[15]}
   );
   gpc1325_5 gpc3557 (
      {stage2_46[28], stage2_46[29], stage2_46[30], stage2_46[31], stage2_46[32]},
      {stage2_47[10], stage2_47[11]},
      {stage2_48[12], stage2_48[13], stage2_48[14]},
      {stage2_49[2]},
      {stage3_50[3],stage3_49[4],stage3_48[6],stage3_47[9],stage3_46[16]}
   );
   gpc615_5 gpc3558 (
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16]},
      {stage2_48[15]},
      {stage2_49[3], stage2_49[4], stage2_49[5], stage2_49[6], stage2_49[7], stage2_49[8]},
      {stage3_51[0],stage3_50[4],stage3_49[5],stage3_48[7],stage3_47[10]}
   );
   gpc615_5 gpc3559 (
      {stage2_47[17], stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21]},
      {stage2_48[16]},
      {stage2_49[9], stage2_49[10], stage2_49[11], stage2_49[12], stage2_49[13], stage2_49[14]},
      {stage3_51[1],stage3_50[5],stage3_49[6],stage3_48[8],stage3_47[11]}
   );
   gpc615_5 gpc3560 (
      {stage2_47[22], stage2_47[23], stage2_47[24], stage2_47[25], stage2_47[26]},
      {stage2_48[17]},
      {stage2_49[15], stage2_49[16], stage2_49[17], stage2_49[18], stage2_49[19], stage2_49[20]},
      {stage3_51[2],stage3_50[6],stage3_49[7],stage3_48[9],stage3_47[12]}
   );
   gpc615_5 gpc3561 (
      {stage2_47[27], stage2_47[28], stage2_47[29], stage2_47[30], stage2_47[31]},
      {stage2_48[18]},
      {stage2_49[21], stage2_49[22], stage2_49[23], stage2_49[24], stage2_49[25], stage2_49[26]},
      {stage3_51[3],stage3_50[7],stage3_49[8],stage3_48[10],stage3_47[13]}
   );
   gpc615_5 gpc3562 (
      {stage2_47[32], stage2_47[33], stage2_47[34], stage2_47[35], stage2_47[36]},
      {stage2_48[19]},
      {stage2_49[27], stage2_49[28], stage2_49[29], stage2_49[30], stage2_49[31], stage2_49[32]},
      {stage3_51[4],stage3_50[8],stage3_49[9],stage3_48[11],stage3_47[14]}
   );
   gpc2116_5 gpc3563 (
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage2_51[0]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1]},
      {stage3_54[0],stage3_53[0],stage3_52[0],stage3_51[5],stage3_50[9]}
   );
   gpc2116_5 gpc3564 (
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage2_51[1]},
      {stage2_52[1]},
      {stage2_53[2], stage2_53[3]},
      {stage3_54[1],stage3_53[1],stage3_52[1],stage3_51[6],stage3_50[10]}
   );
   gpc615_5 gpc3565 (
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16]},
      {stage2_51[2]},
      {stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5], stage2_52[6], stage2_52[7]},
      {stage3_54[2],stage3_53[2],stage3_52[2],stage3_51[7],stage3_50[11]}
   );
   gpc615_5 gpc3566 (
      {stage2_50[17], stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21]},
      {stage2_51[3]},
      {stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11], stage2_52[12], stage2_52[13]},
      {stage3_54[3],stage3_53[3],stage3_52[3],stage3_51[8],stage3_50[12]}
   );
   gpc615_5 gpc3567 (
      {stage2_51[4], stage2_51[5], stage2_51[6], stage2_51[7], stage2_51[8]},
      {stage2_52[14]},
      {stage2_53[4], stage2_53[5], stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9]},
      {stage3_55[0],stage3_54[4],stage3_53[4],stage3_52[4],stage3_51[9]}
   );
   gpc615_5 gpc3568 (
      {stage2_51[9], stage2_51[10], stage2_51[11], stage2_51[12], stage2_51[13]},
      {stage2_52[15]},
      {stage2_53[10], stage2_53[11], stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15]},
      {stage3_55[1],stage3_54[5],stage3_53[5],stage3_52[5],stage3_51[10]}
   );
   gpc615_5 gpc3569 (
      {stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17], stage2_51[18]},
      {stage2_52[16]},
      {stage2_53[16], stage2_53[17], stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21]},
      {stage3_55[2],stage3_54[6],stage3_53[6],stage3_52[6],stage3_51[11]}
   );
   gpc615_5 gpc3570 (
      {stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23]},
      {stage2_52[17]},
      {stage2_53[22], stage2_53[23], stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27]},
      {stage3_55[3],stage3_54[7],stage3_53[7],stage3_52[7],stage3_51[12]}
   );
   gpc606_5 gpc3571 (
      {stage2_53[28], stage2_53[29], stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[0],stage3_55[4],stage3_54[8],stage3_53[8]}
   );
   gpc606_5 gpc3572 (
      {stage2_53[34], stage2_53[35], stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[1],stage3_55[5],stage3_54[9],stage3_53[9]}
   );
   gpc606_5 gpc3573 (
      {stage2_53[40], stage2_53[41], stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage3_57[2],stage3_56[2],stage3_55[6],stage3_54[10],stage3_53[10]}
   );
   gpc606_5 gpc3574 (
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[3],stage3_56[3],stage3_55[7],stage3_54[11]}
   );
   gpc606_5 gpc3575 (
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[4],stage3_56[4],stage3_55[8],stage3_54[12]}
   );
   gpc606_5 gpc3576 (
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[5],stage3_56[5],stage3_55[9],stage3_54[13]}
   );
   gpc615_5 gpc3577 (
      {stage2_54[18], stage2_54[19], stage2_54[20], stage2_54[21], stage2_54[22]},
      {stage2_55[18]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[6],stage3_56[6],stage3_55[10],stage3_54[14]}
   );
   gpc615_5 gpc3578 (
      {stage2_54[23], stage2_54[24], stage2_54[25], stage2_54[26], stage2_54[27]},
      {stage2_55[19]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[7],stage3_56[7],stage3_55[11],stage3_54[15]}
   );
   gpc615_5 gpc3579 (
      {stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23], stage2_55[24]},
      {stage2_56[30]},
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5]},
      {stage3_59[0],stage3_58[5],stage3_57[8],stage3_56[8],stage3_55[12]}
   );
   gpc615_5 gpc3580 (
      {stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage2_56[31]},
      {stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage3_59[1],stage3_58[6],stage3_57[9],stage3_56[9],stage3_55[13]}
   );
   gpc615_5 gpc3581 (
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34]},
      {stage2_56[32]},
      {stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16], stage2_57[17]},
      {stage3_59[2],stage3_58[7],stage3_57[10],stage3_56[10],stage3_55[14]}
   );
   gpc606_5 gpc3582 (
      {stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22], stage2_57[23]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[0],stage3_59[3],stage3_58[8],stage3_57[11]}
   );
   gpc606_5 gpc3583 (
      {stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28], stage2_57[29]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[1],stage3_59[4],stage3_58[9],stage3_57[12]}
   );
   gpc1163_5 gpc3584 (
      {stage2_58[0], stage2_58[1], stage2_58[2]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage2_60[0]},
      {stage2_61[0]},
      {stage3_62[0],stage3_61[2],stage3_60[2],stage3_59[5],stage3_58[10]}
   );
   gpc615_5 gpc3585 (
      {stage2_58[3], stage2_58[4], stage2_58[5], stage2_58[6], stage2_58[7]},
      {stage2_59[18]},
      {stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5], stage2_60[6]},
      {stage3_62[1],stage3_61[3],stage3_60[3],stage3_59[6],stage3_58[11]}
   );
   gpc615_5 gpc3586 (
      {stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11], stage2_58[12]},
      {stage2_59[19]},
      {stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11], stage2_60[12]},
      {stage3_62[2],stage3_61[4],stage3_60[4],stage3_59[7],stage3_58[12]}
   );
   gpc135_4 gpc3587 (
      {stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23], stage2_59[24]},
      {stage2_60[13], stage2_60[14], stage2_60[15]},
      {stage2_61[1]},
      {stage3_62[3],stage3_61[5],stage3_60[5],stage3_59[8]}
   );
   gpc606_5 gpc3588 (
      {stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29], stage2_59[30]},
      {stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5], stage2_61[6], stage2_61[7]},
      {stage3_63[0],stage3_62[4],stage3_61[6],stage3_60[6],stage3_59[9]}
   );
   gpc606_5 gpc3589 (
      {stage2_59[31], stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35], stage2_59[36]},
      {stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11], stage2_61[12], stage2_61[13]},
      {stage3_63[1],stage3_62[5],stage3_61[7],stage3_60[7],stage3_59[10]}
   );
   gpc606_5 gpc3590 (
      {stage2_59[37], stage2_59[38], stage2_59[39], stage2_59[40], stage2_59[41], stage2_59[42]},
      {stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17], stage2_61[18], stage2_61[19]},
      {stage3_63[2],stage3_62[6],stage3_61[8],stage3_60[8],stage3_59[11]}
   );
   gpc606_5 gpc3591 (
      {stage2_59[43], stage2_59[44], stage2_59[45], stage2_59[46], stage2_59[47], stage2_59[48]},
      {stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23], stage2_61[24], stage2_61[25]},
      {stage3_63[3],stage3_62[7],stage3_61[9],stage3_60[9],stage3_59[12]}
   );
   gpc606_5 gpc3592 (
      {stage2_59[49], stage2_59[50], stage2_59[51], stage2_59[52], stage2_59[53], stage2_59[54]},
      {stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29], stage2_61[30], stage2_61[31]},
      {stage3_63[4],stage3_62[8],stage3_61[10],stage3_60[10],stage3_59[13]}
   );
   gpc615_5 gpc3593 (
      {stage2_59[55], stage2_59[56], stage2_59[57], stage2_59[58], stage2_59[59]},
      {stage2_60[16]},
      {stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35], stage2_61[36], stage2_61[37]},
      {stage3_63[5],stage3_62[9],stage3_61[11],stage3_60[11],stage3_59[14]}
   );
   gpc615_5 gpc3594 (
      {stage2_59[60], stage2_59[61], stage2_59[62], stage2_59[63], stage2_59[64]},
      {stage2_60[17]},
      {stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41], stage2_61[42], stage2_61[43]},
      {stage3_63[6],stage3_62[10],stage3_61[12],stage3_60[12],stage3_59[15]}
   );
   gpc615_5 gpc3595 (
      {stage2_59[65], stage2_59[66], stage2_59[67], stage2_59[68], stage2_59[69]},
      {stage2_60[18]},
      {stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47], stage2_61[48], stage2_61[49]},
      {stage3_63[7],stage3_62[11],stage3_61[13],stage3_60[13],stage3_59[16]}
   );
   gpc606_5 gpc3596 (
      {stage2_60[19], stage2_60[20], stage2_60[21], 1'b0, 1'b0, 1'b0},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[8],stage3_62[12],stage3_61[14],stage3_60[14]}
   );
   gpc1163_5 gpc3597 (
      {stage2_61[50], stage2_61[51], stage2_61[52]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage2_63[0]},
      {stage2_64[0]},
      {stage3_65[0],stage3_64[1],stage3_63[9],stage3_62[13],stage3_61[15]}
   );
   gpc606_5 gpc3598 (
      {stage2_61[53], stage2_61[54], stage2_61[55], stage2_61[56], stage2_61[57], stage2_61[58]},
      {stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5], stage2_63[6]},
      {stage3_65[1],stage3_64[2],stage3_63[10],stage3_62[14],stage3_61[16]}
   );
   gpc1163_5 gpc3599 (
      {stage2_62[12], stage2_62[13], stage2_62[14]},
      {stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11], stage2_63[12]},
      {stage2_64[1]},
      {stage2_65[0]},
      {stage3_66[0],stage3_65[2],stage3_64[3],stage3_63[11],stage3_62[15]}
   );
   gpc1163_5 gpc3600 (
      {stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage2_63[13], stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17], stage2_63[18]},
      {stage2_64[2]},
      {stage2_65[1]},
      {stage3_66[1],stage3_65[3],stage3_64[4],stage3_63[12],stage3_62[16]}
   );
   gpc1163_5 gpc3601 (
      {stage2_62[18], stage2_62[19], stage2_62[20]},
      {stage2_63[19], stage2_63[20], stage2_63[21], stage2_63[22], stage2_63[23], stage2_63[24]},
      {stage2_64[3]},
      {stage2_65[2]},
      {stage3_66[2],stage3_65[4],stage3_64[5],stage3_63[13],stage3_62[17]}
   );
   gpc1163_5 gpc3602 (
      {stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage2_63[25], stage2_63[26], stage2_63[27], stage2_63[28], stage2_63[29], stage2_63[30]},
      {stage2_64[4]},
      {stage2_65[3]},
      {stage3_66[3],stage3_65[5],stage3_64[6],stage3_63[14],stage3_62[18]}
   );
   gpc606_5 gpc3603 (
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage2_64[5], stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10]},
      {stage3_66[4],stage3_65[6],stage3_64[7],stage3_63[15],stage3_62[19]}
   );
   gpc615_5 gpc3604 (
      {stage2_62[30], stage2_62[31], stage2_62[32], stage2_62[33], stage2_62[34]},
      {stage2_63[31]},
      {stage2_64[11], stage2_64[12], stage2_64[13], stage2_64[14], stage2_64[15], stage2_64[16]},
      {stage3_66[5],stage3_65[7],stage3_64[8],stage3_63[16],stage3_62[20]}
   );
   gpc606_5 gpc3605 (
      {stage2_63[32], stage2_63[33], stage2_63[34], stage2_63[35], stage2_63[36], stage2_63[37]},
      {stage2_65[4], stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8], stage2_65[9]},
      {stage3_67[0],stage3_66[6],stage3_65[8],stage3_64[9],stage3_63[17]}
   );
   gpc606_5 gpc3606 (
      {stage2_64[17], stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21], stage2_64[22]},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3], stage2_66[4], stage2_66[5]},
      {stage3_68[0],stage3_67[1],stage3_66[7],stage3_65[9],stage3_64[10]}
   );
   gpc606_5 gpc3607 (
      {stage2_64[23], stage2_64[24], stage2_64[25], stage2_64[26], stage2_64[27], stage2_64[28]},
      {stage2_66[6], stage2_66[7], stage2_66[8], stage2_66[9], 1'b0, 1'b0},
      {stage3_68[1],stage3_67[2],stage3_66[8],stage3_65[10],stage3_64[11]}
   );
   gpc1_1 gpc3608 (
      {stage2_0[3]},
      {stage3_0[1]}
   );
   gpc1_1 gpc3609 (
      {stage2_0[4]},
      {stage3_0[2]}
   );
   gpc1_1 gpc3610 (
      {stage2_0[5]},
      {stage3_0[3]}
   );
   gpc1_1 gpc3611 (
      {stage2_0[6]},
      {stage3_0[4]}
   );
   gpc1_1 gpc3612 (
      {stage2_0[7]},
      {stage3_0[5]}
   );
   gpc1_1 gpc3613 (
      {stage2_0[8]},
      {stage3_0[6]}
   );
   gpc1_1 gpc3614 (
      {stage2_0[9]},
      {stage3_0[7]}
   );
   gpc1_1 gpc3615 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc3616 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc3617 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc3618 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc3619 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc3620 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc3621 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc3622 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc3623 (
      {stage2_1[14]},
      {stage3_1[9]}
   );
   gpc1_1 gpc3624 (
      {stage2_1[15]},
      {stage3_1[10]}
   );
   gpc1_1 gpc3625 (
      {stage2_1[16]},
      {stage3_1[11]}
   );
   gpc1_1 gpc3626 (
      {stage2_1[17]},
      {stage3_1[12]}
   );
   gpc1_1 gpc3627 (
      {stage2_1[18]},
      {stage3_1[13]}
   );
   gpc1_1 gpc3628 (
      {stage2_2[34]},
      {stage3_2[7]}
   );
   gpc1_1 gpc3629 (
      {stage2_2[35]},
      {stage3_2[8]}
   );
   gpc1_1 gpc3630 (
      {stage2_2[36]},
      {stage3_2[9]}
   );
   gpc1_1 gpc3631 (
      {stage2_2[37]},
      {stage3_2[10]}
   );
   gpc1_1 gpc3632 (
      {stage2_3[19]},
      {stage3_3[10]}
   );
   gpc1_1 gpc3633 (
      {stage2_3[20]},
      {stage3_3[11]}
   );
   gpc1_1 gpc3634 (
      {stage2_3[21]},
      {stage3_3[12]}
   );
   gpc1_1 gpc3635 (
      {stage2_3[22]},
      {stage3_3[13]}
   );
   gpc1_1 gpc3636 (
      {stage2_4[45]},
      {stage3_4[11]}
   );
   gpc1_1 gpc3637 (
      {stage2_4[46]},
      {stage3_4[12]}
   );
   gpc1_1 gpc3638 (
      {stage2_4[47]},
      {stage3_4[13]}
   );
   gpc1_1 gpc3639 (
      {stage2_5[30]},
      {stage3_5[12]}
   );
   gpc1_1 gpc3640 (
      {stage2_5[31]},
      {stage3_5[13]}
   );
   gpc1_1 gpc3641 (
      {stage2_5[32]},
      {stage3_5[14]}
   );
   gpc1_1 gpc3642 (
      {stage2_5[33]},
      {stage3_5[15]}
   );
   gpc1_1 gpc3643 (
      {stage2_5[34]},
      {stage3_5[16]}
   );
   gpc1_1 gpc3644 (
      {stage2_5[35]},
      {stage3_5[17]}
   );
   gpc1_1 gpc3645 (
      {stage2_6[24]},
      {stage3_6[15]}
   );
   gpc1_1 gpc3646 (
      {stage2_6[25]},
      {stage3_6[16]}
   );
   gpc1_1 gpc3647 (
      {stage2_6[26]},
      {stage3_6[17]}
   );
   gpc1_1 gpc3648 (
      {stage2_6[27]},
      {stage3_6[18]}
   );
   gpc1_1 gpc3649 (
      {stage2_6[28]},
      {stage3_6[19]}
   );
   gpc1_1 gpc3650 (
      {stage2_7[37]},
      {stage3_7[13]}
   );
   gpc1_1 gpc3651 (
      {stage2_7[38]},
      {stage3_7[14]}
   );
   gpc1_1 gpc3652 (
      {stage2_7[39]},
      {stage3_7[15]}
   );
   gpc1_1 gpc3653 (
      {stage2_7[40]},
      {stage3_7[16]}
   );
   gpc1_1 gpc3654 (
      {stage2_9[22]},
      {stage3_9[17]}
   );
   gpc1_1 gpc3655 (
      {stage2_9[23]},
      {stage3_9[18]}
   );
   gpc1_1 gpc3656 (
      {stage2_9[24]},
      {stage3_9[19]}
   );
   gpc1_1 gpc3657 (
      {stage2_9[25]},
      {stage3_9[20]}
   );
   gpc1_1 gpc3658 (
      {stage2_11[36]},
      {stage3_11[15]}
   );
   gpc1_1 gpc3659 (
      {stage2_11[37]},
      {stage3_11[16]}
   );
   gpc1_1 gpc3660 (
      {stage2_11[38]},
      {stage3_11[17]}
   );
   gpc1_1 gpc3661 (
      {stage2_12[24]},
      {stage3_12[17]}
   );
   gpc1_1 gpc3662 (
      {stage2_12[25]},
      {stage3_12[18]}
   );
   gpc1_1 gpc3663 (
      {stage2_12[26]},
      {stage3_12[19]}
   );
   gpc1_1 gpc3664 (
      {stage2_12[27]},
      {stage3_12[20]}
   );
   gpc1_1 gpc3665 (
      {stage2_12[28]},
      {stage3_12[21]}
   );
   gpc1_1 gpc3666 (
      {stage2_12[29]},
      {stage3_12[22]}
   );
   gpc1_1 gpc3667 (
      {stage2_12[30]},
      {stage3_12[23]}
   );
   gpc1_1 gpc3668 (
      {stage2_13[36]},
      {stage3_13[11]}
   );
   gpc1_1 gpc3669 (
      {stage2_13[37]},
      {stage3_13[12]}
   );
   gpc1_1 gpc3670 (
      {stage2_13[38]},
      {stage3_13[13]}
   );
   gpc1_1 gpc3671 (
      {stage2_13[39]},
      {stage3_13[14]}
   );
   gpc1_1 gpc3672 (
      {stage2_13[40]},
      {stage3_13[15]}
   );
   gpc1_1 gpc3673 (
      {stage2_13[41]},
      {stage3_13[16]}
   );
   gpc1_1 gpc3674 (
      {stage2_13[42]},
      {stage3_13[17]}
   );
   gpc1_1 gpc3675 (
      {stage2_13[43]},
      {stage3_13[18]}
   );
   gpc1_1 gpc3676 (
      {stage2_13[44]},
      {stage3_13[19]}
   );
   gpc1_1 gpc3677 (
      {stage2_14[54]},
      {stage3_14[16]}
   );
   gpc1_1 gpc3678 (
      {stage2_14[55]},
      {stage3_14[17]}
   );
   gpc1_1 gpc3679 (
      {stage2_14[56]},
      {stage3_14[18]}
   );
   gpc1_1 gpc3680 (
      {stage2_14[57]},
      {stage3_14[19]}
   );
   gpc1_1 gpc3681 (
      {stage2_14[58]},
      {stage3_14[20]}
   );
   gpc1_1 gpc3682 (
      {stage2_14[59]},
      {stage3_14[21]}
   );
   gpc1_1 gpc3683 (
      {stage2_14[60]},
      {stage3_14[22]}
   );
   gpc1_1 gpc3684 (
      {stage2_14[61]},
      {stage3_14[23]}
   );
   gpc1_1 gpc3685 (
      {stage2_14[62]},
      {stage3_14[24]}
   );
   gpc1_1 gpc3686 (
      {stage2_14[63]},
      {stage3_14[25]}
   );
   gpc1_1 gpc3687 (
      {stage2_14[64]},
      {stage3_14[26]}
   );
   gpc1_1 gpc3688 (
      {stage2_14[65]},
      {stage3_14[27]}
   );
   gpc1_1 gpc3689 (
      {stage2_14[66]},
      {stage3_14[28]}
   );
   gpc1_1 gpc3690 (
      {stage2_14[67]},
      {stage3_14[29]}
   );
   gpc1_1 gpc3691 (
      {stage2_14[68]},
      {stage3_14[30]}
   );
   gpc1_1 gpc3692 (
      {stage2_14[69]},
      {stage3_14[31]}
   );
   gpc1_1 gpc3693 (
      {stage2_14[70]},
      {stage3_14[32]}
   );
   gpc1_1 gpc3694 (
      {stage2_14[71]},
      {stage3_14[33]}
   );
   gpc1_1 gpc3695 (
      {stage2_14[72]},
      {stage3_14[34]}
   );
   gpc1_1 gpc3696 (
      {stage2_14[73]},
      {stage3_14[35]}
   );
   gpc1_1 gpc3697 (
      {stage2_15[17]},
      {stage3_15[17]}
   );
   gpc1_1 gpc3698 (
      {stage2_15[18]},
      {stage3_15[18]}
   );
   gpc1_1 gpc3699 (
      {stage2_15[19]},
      {stage3_15[19]}
   );
   gpc1_1 gpc3700 (
      {stage2_15[20]},
      {stage3_15[20]}
   );
   gpc1_1 gpc3701 (
      {stage2_15[21]},
      {stage3_15[21]}
   );
   gpc1_1 gpc3702 (
      {stage2_15[22]},
      {stage3_15[22]}
   );
   gpc1_1 gpc3703 (
      {stage2_15[23]},
      {stage3_15[23]}
   );
   gpc1_1 gpc3704 (
      {stage2_15[24]},
      {stage3_15[24]}
   );
   gpc1_1 gpc3705 (
      {stage2_15[25]},
      {stage3_15[25]}
   );
   gpc1_1 gpc3706 (
      {stage2_15[26]},
      {stage3_15[26]}
   );
   gpc1_1 gpc3707 (
      {stage2_15[27]},
      {stage3_15[27]}
   );
   gpc1_1 gpc3708 (
      {stage2_15[28]},
      {stage3_15[28]}
   );
   gpc1_1 gpc3709 (
      {stage2_15[29]},
      {stage3_15[29]}
   );
   gpc1_1 gpc3710 (
      {stage2_15[30]},
      {stage3_15[30]}
   );
   gpc1_1 gpc3711 (
      {stage2_15[31]},
      {stage3_15[31]}
   );
   gpc1_1 gpc3712 (
      {stage2_15[32]},
      {stage3_15[32]}
   );
   gpc1_1 gpc3713 (
      {stage2_15[33]},
      {stage3_15[33]}
   );
   gpc1_1 gpc3714 (
      {stage2_15[34]},
      {stage3_15[34]}
   );
   gpc1_1 gpc3715 (
      {stage2_15[35]},
      {stage3_15[35]}
   );
   gpc1_1 gpc3716 (
      {stage2_15[36]},
      {stage3_15[36]}
   );
   gpc1_1 gpc3717 (
      {stage2_16[37]},
      {stage3_16[12]}
   );
   gpc1_1 gpc3718 (
      {stage2_16[38]},
      {stage3_16[13]}
   );
   gpc1_1 gpc3719 (
      {stage2_16[39]},
      {stage3_16[14]}
   );
   gpc1_1 gpc3720 (
      {stage2_16[40]},
      {stage3_16[15]}
   );
   gpc1_1 gpc3721 (
      {stage2_16[41]},
      {stage3_16[16]}
   );
   gpc1_1 gpc3722 (
      {stage2_16[42]},
      {stage3_16[17]}
   );
   gpc1_1 gpc3723 (
      {stage2_16[43]},
      {stage3_16[18]}
   );
   gpc1_1 gpc3724 (
      {stage2_16[44]},
      {stage3_16[19]}
   );
   gpc1_1 gpc3725 (
      {stage2_16[45]},
      {stage3_16[20]}
   );
   gpc1_1 gpc3726 (
      {stage2_16[46]},
      {stage3_16[21]}
   );
   gpc1_1 gpc3727 (
      {stage2_17[36]},
      {stage3_17[13]}
   );
   gpc1_1 gpc3728 (
      {stage2_17[37]},
      {stage3_17[14]}
   );
   gpc1_1 gpc3729 (
      {stage2_17[38]},
      {stage3_17[15]}
   );
   gpc1_1 gpc3730 (
      {stage2_17[39]},
      {stage3_17[16]}
   );
   gpc1_1 gpc3731 (
      {stage2_18[40]},
      {stage3_18[20]}
   );
   gpc1_1 gpc3732 (
      {stage2_18[41]},
      {stage3_18[21]}
   );
   gpc1_1 gpc3733 (
      {stage2_18[42]},
      {stage3_18[22]}
   );
   gpc1_1 gpc3734 (
      {stage2_19[38]},
      {stage3_19[14]}
   );
   gpc1_1 gpc3735 (
      {stage2_19[39]},
      {stage3_19[15]}
   );
   gpc1_1 gpc3736 (
      {stage2_19[40]},
      {stage3_19[16]}
   );
   gpc1_1 gpc3737 (
      {stage2_19[41]},
      {stage3_19[17]}
   );
   gpc1_1 gpc3738 (
      {stage2_19[42]},
      {stage3_19[18]}
   );
   gpc1_1 gpc3739 (
      {stage2_19[43]},
      {stage3_19[19]}
   );
   gpc1_1 gpc3740 (
      {stage2_19[44]},
      {stage3_19[20]}
   );
   gpc1_1 gpc3741 (
      {stage2_19[45]},
      {stage3_19[21]}
   );
   gpc1_1 gpc3742 (
      {stage2_19[46]},
      {stage3_19[22]}
   );
   gpc1_1 gpc3743 (
      {stage2_19[47]},
      {stage3_19[23]}
   );
   gpc1_1 gpc3744 (
      {stage2_19[48]},
      {stage3_19[24]}
   );
   gpc1_1 gpc3745 (
      {stage2_19[49]},
      {stage3_19[25]}
   );
   gpc1_1 gpc3746 (
      {stage2_19[50]},
      {stage3_19[26]}
   );
   gpc1_1 gpc3747 (
      {stage2_20[48]},
      {stage3_20[13]}
   );
   gpc1_1 gpc3748 (
      {stage2_20[49]},
      {stage3_20[14]}
   );
   gpc1_1 gpc3749 (
      {stage2_20[50]},
      {stage3_20[15]}
   );
   gpc1_1 gpc3750 (
      {stage2_20[51]},
      {stage3_20[16]}
   );
   gpc1_1 gpc3751 (
      {stage2_20[52]},
      {stage3_20[17]}
   );
   gpc1_1 gpc3752 (
      {stage2_20[53]},
      {stage3_20[18]}
   );
   gpc1_1 gpc3753 (
      {stage2_20[54]},
      {stage3_20[19]}
   );
   gpc1_1 gpc3754 (
      {stage2_20[55]},
      {stage3_20[20]}
   );
   gpc1_1 gpc3755 (
      {stage2_20[56]},
      {stage3_20[21]}
   );
   gpc1_1 gpc3756 (
      {stage2_20[57]},
      {stage3_20[22]}
   );
   gpc1_1 gpc3757 (
      {stage2_21[35]},
      {stage3_21[20]}
   );
   gpc1_1 gpc3758 (
      {stage2_21[36]},
      {stage3_21[21]}
   );
   gpc1_1 gpc3759 (
      {stage2_21[37]},
      {stage3_21[22]}
   );
   gpc1_1 gpc3760 (
      {stage2_21[38]},
      {stage3_21[23]}
   );
   gpc1_1 gpc3761 (
      {stage2_21[39]},
      {stage3_21[24]}
   );
   gpc1_1 gpc3762 (
      {stage2_22[22]},
      {stage3_22[18]}
   );
   gpc1_1 gpc3763 (
      {stage2_22[23]},
      {stage3_22[19]}
   );
   gpc1_1 gpc3764 (
      {stage2_22[24]},
      {stage3_22[20]}
   );
   gpc1_1 gpc3765 (
      {stage2_22[25]},
      {stage3_22[21]}
   );
   gpc1_1 gpc3766 (
      {stage2_22[26]},
      {stage3_22[22]}
   );
   gpc1_1 gpc3767 (
      {stage2_22[27]},
      {stage3_22[23]}
   );
   gpc1_1 gpc3768 (
      {stage2_22[28]},
      {stage3_22[24]}
   );
   gpc1_1 gpc3769 (
      {stage2_22[29]},
      {stage3_22[25]}
   );
   gpc1_1 gpc3770 (
      {stage2_22[30]},
      {stage3_22[26]}
   );
   gpc1_1 gpc3771 (
      {stage2_23[45]},
      {stage3_23[10]}
   );
   gpc1_1 gpc3772 (
      {stage2_23[46]},
      {stage3_23[11]}
   );
   gpc1_1 gpc3773 (
      {stage2_24[33]},
      {stage3_24[13]}
   );
   gpc1_1 gpc3774 (
      {stage2_24[34]},
      {stage3_24[14]}
   );
   gpc1_1 gpc3775 (
      {stage2_24[35]},
      {stage3_24[15]}
   );
   gpc1_1 gpc3776 (
      {stage2_24[36]},
      {stage3_24[16]}
   );
   gpc1_1 gpc3777 (
      {stage2_24[37]},
      {stage3_24[17]}
   );
   gpc1_1 gpc3778 (
      {stage2_24[38]},
      {stage3_24[18]}
   );
   gpc1_1 gpc3779 (
      {stage2_24[39]},
      {stage3_24[19]}
   );
   gpc1_1 gpc3780 (
      {stage2_24[40]},
      {stage3_24[20]}
   );
   gpc1_1 gpc3781 (
      {stage2_24[41]},
      {stage3_24[21]}
   );
   gpc1_1 gpc3782 (
      {stage2_24[42]},
      {stage3_24[22]}
   );
   gpc1_1 gpc3783 (
      {stage2_24[43]},
      {stage3_24[23]}
   );
   gpc1_1 gpc3784 (
      {stage2_24[44]},
      {stage3_24[24]}
   );
   gpc1_1 gpc3785 (
      {stage2_24[45]},
      {stage3_24[25]}
   );
   gpc1_1 gpc3786 (
      {stage2_25[33]},
      {stage3_25[18]}
   );
   gpc1_1 gpc3787 (
      {stage2_25[34]},
      {stage3_25[19]}
   );
   gpc1_1 gpc3788 (
      {stage2_25[35]},
      {stage3_25[20]}
   );
   gpc1_1 gpc3789 (
      {stage2_25[36]},
      {stage3_25[21]}
   );
   gpc1_1 gpc3790 (
      {stage2_27[47]},
      {stage3_27[16]}
   );
   gpc1_1 gpc3791 (
      {stage2_27[48]},
      {stage3_27[17]}
   );
   gpc1_1 gpc3792 (
      {stage2_27[49]},
      {stage3_27[18]}
   );
   gpc1_1 gpc3793 (
      {stage2_29[48]},
      {stage3_29[22]}
   );
   gpc1_1 gpc3794 (
      {stage2_29[49]},
      {stage3_29[23]}
   );
   gpc1_1 gpc3795 (
      {stage2_30[39]},
      {stage3_30[15]}
   );
   gpc1_1 gpc3796 (
      {stage2_30[40]},
      {stage3_30[16]}
   );
   gpc1_1 gpc3797 (
      {stage2_30[41]},
      {stage3_30[17]}
   );
   gpc1_1 gpc3798 (
      {stage2_30[42]},
      {stage3_30[18]}
   );
   gpc1_1 gpc3799 (
      {stage2_30[43]},
      {stage3_30[19]}
   );
   gpc1_1 gpc3800 (
      {stage2_30[44]},
      {stage3_30[20]}
   );
   gpc1_1 gpc3801 (
      {stage2_30[45]},
      {stage3_30[21]}
   );
   gpc1_1 gpc3802 (
      {stage2_30[46]},
      {stage3_30[22]}
   );
   gpc1_1 gpc3803 (
      {stage2_30[47]},
      {stage3_30[23]}
   );
   gpc1_1 gpc3804 (
      {stage2_30[48]},
      {stage3_30[24]}
   );
   gpc1_1 gpc3805 (
      {stage2_30[49]},
      {stage3_30[25]}
   );
   gpc1_1 gpc3806 (
      {stage2_31[33]},
      {stage3_31[15]}
   );
   gpc1_1 gpc3807 (
      {stage2_31[34]},
      {stage3_31[16]}
   );
   gpc1_1 gpc3808 (
      {stage2_31[35]},
      {stage3_31[17]}
   );
   gpc1_1 gpc3809 (
      {stage2_31[36]},
      {stage3_31[18]}
   );
   gpc1_1 gpc3810 (
      {stage2_31[37]},
      {stage3_31[19]}
   );
   gpc1_1 gpc3811 (
      {stage2_31[38]},
      {stage3_31[20]}
   );
   gpc1_1 gpc3812 (
      {stage2_32[36]},
      {stage3_32[15]}
   );
   gpc1_1 gpc3813 (
      {stage2_32[37]},
      {stage3_32[16]}
   );
   gpc1_1 gpc3814 (
      {stage2_32[38]},
      {stage3_32[17]}
   );
   gpc1_1 gpc3815 (
      {stage2_32[39]},
      {stage3_32[18]}
   );
   gpc1_1 gpc3816 (
      {stage2_32[40]},
      {stage3_32[19]}
   );
   gpc1_1 gpc3817 (
      {stage2_32[41]},
      {stage3_32[20]}
   );
   gpc1_1 gpc3818 (
      {stage2_32[42]},
      {stage3_32[21]}
   );
   gpc1_1 gpc3819 (
      {stage2_32[43]},
      {stage3_32[22]}
   );
   gpc1_1 gpc3820 (
      {stage2_32[44]},
      {stage3_32[23]}
   );
   gpc1_1 gpc3821 (
      {stage2_32[45]},
      {stage3_32[24]}
   );
   gpc1_1 gpc3822 (
      {stage2_32[46]},
      {stage3_32[25]}
   );
   gpc1_1 gpc3823 (
      {stage2_32[47]},
      {stage3_32[26]}
   );
   gpc1_1 gpc3824 (
      {stage2_32[48]},
      {stage3_32[27]}
   );
   gpc1_1 gpc3825 (
      {stage2_32[49]},
      {stage3_32[28]}
   );
   gpc1_1 gpc3826 (
      {stage2_32[50]},
      {stage3_32[29]}
   );
   gpc1_1 gpc3827 (
      {stage2_32[51]},
      {stage3_32[30]}
   );
   gpc1_1 gpc3828 (
      {stage2_32[52]},
      {stage3_32[31]}
   );
   gpc1_1 gpc3829 (
      {stage2_32[53]},
      {stage3_32[32]}
   );
   gpc1_1 gpc3830 (
      {stage2_32[54]},
      {stage3_32[33]}
   );
   gpc1_1 gpc3831 (
      {stage2_32[55]},
      {stage3_32[34]}
   );
   gpc1_1 gpc3832 (
      {stage2_34[23]},
      {stage3_34[11]}
   );
   gpc1_1 gpc3833 (
      {stage2_34[24]},
      {stage3_34[12]}
   );
   gpc1_1 gpc3834 (
      {stage2_34[25]},
      {stage3_34[13]}
   );
   gpc1_1 gpc3835 (
      {stage2_34[26]},
      {stage3_34[14]}
   );
   gpc1_1 gpc3836 (
      {stage2_34[27]},
      {stage3_34[15]}
   );
   gpc1_1 gpc3837 (
      {stage2_34[28]},
      {stage3_34[16]}
   );
   gpc1_1 gpc3838 (
      {stage2_34[29]},
      {stage3_34[17]}
   );
   gpc1_1 gpc3839 (
      {stage2_34[30]},
      {stage3_34[18]}
   );
   gpc1_1 gpc3840 (
      {stage2_34[31]},
      {stage3_34[19]}
   );
   gpc1_1 gpc3841 (
      {stage2_34[32]},
      {stage3_34[20]}
   );
   gpc1_1 gpc3842 (
      {stage2_34[33]},
      {stage3_34[21]}
   );
   gpc1_1 gpc3843 (
      {stage2_34[34]},
      {stage3_34[22]}
   );
   gpc1_1 gpc3844 (
      {stage2_35[33]},
      {stage3_35[14]}
   );
   gpc1_1 gpc3845 (
      {stage2_35[34]},
      {stage3_35[15]}
   );
   gpc1_1 gpc3846 (
      {stage2_35[35]},
      {stage3_35[16]}
   );
   gpc1_1 gpc3847 (
      {stage2_35[36]},
      {stage3_35[17]}
   );
   gpc1_1 gpc3848 (
      {stage2_35[37]},
      {stage3_35[18]}
   );
   gpc1_1 gpc3849 (
      {stage2_35[38]},
      {stage3_35[19]}
   );
   gpc1_1 gpc3850 (
      {stage2_35[39]},
      {stage3_35[20]}
   );
   gpc1_1 gpc3851 (
      {stage2_35[40]},
      {stage3_35[21]}
   );
   gpc1_1 gpc3852 (
      {stage2_35[41]},
      {stage3_35[22]}
   );
   gpc1_1 gpc3853 (
      {stage2_35[42]},
      {stage3_35[23]}
   );
   gpc1_1 gpc3854 (
      {stage2_35[43]},
      {stage3_35[24]}
   );
   gpc1_1 gpc3855 (
      {stage2_35[44]},
      {stage3_35[25]}
   );
   gpc1_1 gpc3856 (
      {stage2_36[34]},
      {stage3_36[14]}
   );
   gpc1_1 gpc3857 (
      {stage2_36[35]},
      {stage3_36[15]}
   );
   gpc1_1 gpc3858 (
      {stage2_36[36]},
      {stage3_36[16]}
   );
   gpc1_1 gpc3859 (
      {stage2_39[26]},
      {stage3_39[16]}
   );
   gpc1_1 gpc3860 (
      {stage2_39[27]},
      {stage3_39[17]}
   );
   gpc1_1 gpc3861 (
      {stage2_39[28]},
      {stage3_39[18]}
   );
   gpc1_1 gpc3862 (
      {stage2_39[29]},
      {stage3_39[19]}
   );
   gpc1_1 gpc3863 (
      {stage2_39[30]},
      {stage3_39[20]}
   );
   gpc1_1 gpc3864 (
      {stage2_39[31]},
      {stage3_39[21]}
   );
   gpc1_1 gpc3865 (
      {stage2_39[32]},
      {stage3_39[22]}
   );
   gpc1_1 gpc3866 (
      {stage2_39[33]},
      {stage3_39[23]}
   );
   gpc1_1 gpc3867 (
      {stage2_40[30]},
      {stage3_40[13]}
   );
   gpc1_1 gpc3868 (
      {stage2_40[31]},
      {stage3_40[14]}
   );
   gpc1_1 gpc3869 (
      {stage2_40[32]},
      {stage3_40[15]}
   );
   gpc1_1 gpc3870 (
      {stage2_40[33]},
      {stage3_40[16]}
   );
   gpc1_1 gpc3871 (
      {stage2_40[34]},
      {stage3_40[17]}
   );
   gpc1_1 gpc3872 (
      {stage2_40[35]},
      {stage3_40[18]}
   );
   gpc1_1 gpc3873 (
      {stage2_40[36]},
      {stage3_40[19]}
   );
   gpc1_1 gpc3874 (
      {stage2_40[37]},
      {stage3_40[20]}
   );
   gpc1_1 gpc3875 (
      {stage2_40[38]},
      {stage3_40[21]}
   );
   gpc1_1 gpc3876 (
      {stage2_40[39]},
      {stage3_40[22]}
   );
   gpc1_1 gpc3877 (
      {stage2_40[40]},
      {stage3_40[23]}
   );
   gpc1_1 gpc3878 (
      {stage2_41[45]},
      {stage3_41[14]}
   );
   gpc1_1 gpc3879 (
      {stage2_41[46]},
      {stage3_41[15]}
   );
   gpc1_1 gpc3880 (
      {stage2_41[47]},
      {stage3_41[16]}
   );
   gpc1_1 gpc3881 (
      {stage2_41[48]},
      {stage3_41[17]}
   );
   gpc1_1 gpc3882 (
      {stage2_41[49]},
      {stage3_41[18]}
   );
   gpc1_1 gpc3883 (
      {stage2_41[50]},
      {stage3_41[19]}
   );
   gpc1_1 gpc3884 (
      {stage2_41[51]},
      {stage3_41[20]}
   );
   gpc1_1 gpc3885 (
      {stage2_41[52]},
      {stage3_41[21]}
   );
   gpc1_1 gpc3886 (
      {stage2_41[53]},
      {stage3_41[22]}
   );
   gpc1_1 gpc3887 (
      {stage2_41[54]},
      {stage3_41[23]}
   );
   gpc1_1 gpc3888 (
      {stage2_41[55]},
      {stage3_41[24]}
   );
   gpc1_1 gpc3889 (
      {stage2_42[56]},
      {stage3_42[20]}
   );
   gpc1_1 gpc3890 (
      {stage2_42[57]},
      {stage3_42[21]}
   );
   gpc1_1 gpc3891 (
      {stage2_42[58]},
      {stage3_42[22]}
   );
   gpc1_1 gpc3892 (
      {stage2_42[59]},
      {stage3_42[23]}
   );
   gpc1_1 gpc3893 (
      {stage2_42[60]},
      {stage3_42[24]}
   );
   gpc1_1 gpc3894 (
      {stage2_42[61]},
      {stage3_42[25]}
   );
   gpc1_1 gpc3895 (
      {stage2_44[55]},
      {stage3_44[20]}
   );
   gpc1_1 gpc3896 (
      {stage2_44[56]},
      {stage3_44[21]}
   );
   gpc1_1 gpc3897 (
      {stage2_44[57]},
      {stage3_44[22]}
   );
   gpc1_1 gpc3898 (
      {stage2_44[58]},
      {stage3_44[23]}
   );
   gpc1_1 gpc3899 (
      {stage2_44[59]},
      {stage3_44[24]}
   );
   gpc1_1 gpc3900 (
      {stage2_44[60]},
      {stage3_44[25]}
   );
   gpc1_1 gpc3901 (
      {stage2_44[61]},
      {stage3_44[26]}
   );
   gpc1_1 gpc3902 (
      {stage2_44[62]},
      {stage3_44[27]}
   );
   gpc1_1 gpc3903 (
      {stage2_44[63]},
      {stage3_44[28]}
   );
   gpc1_1 gpc3904 (
      {stage2_44[64]},
      {stage3_44[29]}
   );
   gpc1_1 gpc3905 (
      {stage2_44[65]},
      {stage3_44[30]}
   );
   gpc1_1 gpc3906 (
      {stage2_47[37]},
      {stage3_47[15]}
   );
   gpc1_1 gpc3907 (
      {stage2_47[38]},
      {stage3_47[16]}
   );
   gpc1_1 gpc3908 (
      {stage2_47[39]},
      {stage3_47[17]}
   );
   gpc1_1 gpc3909 (
      {stage2_47[40]},
      {stage3_47[18]}
   );
   gpc1_1 gpc3910 (
      {stage2_47[41]},
      {stage3_47[19]}
   );
   gpc1_1 gpc3911 (
      {stage2_47[42]},
      {stage3_47[20]}
   );
   gpc1_1 gpc3912 (
      {stage2_47[43]},
      {stage3_47[21]}
   );
   gpc1_1 gpc3913 (
      {stage2_47[44]},
      {stage3_47[22]}
   );
   gpc1_1 gpc3914 (
      {stage2_47[45]},
      {stage3_47[23]}
   );
   gpc1_1 gpc3915 (
      {stage2_48[20]},
      {stage3_48[12]}
   );
   gpc1_1 gpc3916 (
      {stage2_48[21]},
      {stage3_48[13]}
   );
   gpc1_1 gpc3917 (
      {stage2_48[22]},
      {stage3_48[14]}
   );
   gpc1_1 gpc3918 (
      {stage2_48[23]},
      {stage3_48[15]}
   );
   gpc1_1 gpc3919 (
      {stage2_49[33]},
      {stage3_49[10]}
   );
   gpc1_1 gpc3920 (
      {stage2_49[34]},
      {stage3_49[11]}
   );
   gpc1_1 gpc3921 (
      {stage2_49[35]},
      {stage3_49[12]}
   );
   gpc1_1 gpc3922 (
      {stage2_49[36]},
      {stage3_49[13]}
   );
   gpc1_1 gpc3923 (
      {stage2_50[22]},
      {stage3_50[13]}
   );
   gpc1_1 gpc3924 (
      {stage2_50[23]},
      {stage3_50[14]}
   );
   gpc1_1 gpc3925 (
      {stage2_50[24]},
      {stage3_50[15]}
   );
   gpc1_1 gpc3926 (
      {stage2_50[25]},
      {stage3_50[16]}
   );
   gpc1_1 gpc3927 (
      {stage2_50[26]},
      {stage3_50[17]}
   );
   gpc1_1 gpc3928 (
      {stage2_50[27]},
      {stage3_50[18]}
   );
   gpc1_1 gpc3929 (
      {stage2_50[28]},
      {stage3_50[19]}
   );
   gpc1_1 gpc3930 (
      {stage2_50[29]},
      {stage3_50[20]}
   );
   gpc1_1 gpc3931 (
      {stage2_50[30]},
      {stage3_50[21]}
   );
   gpc1_1 gpc3932 (
      {stage2_50[31]},
      {stage3_50[22]}
   );
   gpc1_1 gpc3933 (
      {stage2_50[32]},
      {stage3_50[23]}
   );
   gpc1_1 gpc3934 (
      {stage2_50[33]},
      {stage3_50[24]}
   );
   gpc1_1 gpc3935 (
      {stage2_50[34]},
      {stage3_50[25]}
   );
   gpc1_1 gpc3936 (
      {stage2_50[35]},
      {stage3_50[26]}
   );
   gpc1_1 gpc3937 (
      {stage2_50[36]},
      {stage3_50[27]}
   );
   gpc1_1 gpc3938 (
      {stage2_50[37]},
      {stage3_50[28]}
   );
   gpc1_1 gpc3939 (
      {stage2_50[38]},
      {stage3_50[29]}
   );
   gpc1_1 gpc3940 (
      {stage2_50[39]},
      {stage3_50[30]}
   );
   gpc1_1 gpc3941 (
      {stage2_50[40]},
      {stage3_50[31]}
   );
   gpc1_1 gpc3942 (
      {stage2_51[24]},
      {stage3_51[13]}
   );
   gpc1_1 gpc3943 (
      {stage2_52[18]},
      {stage3_52[8]}
   );
   gpc1_1 gpc3944 (
      {stage2_52[19]},
      {stage3_52[9]}
   );
   gpc1_1 gpc3945 (
      {stage2_52[20]},
      {stage3_52[10]}
   );
   gpc1_1 gpc3946 (
      {stage2_52[21]},
      {stage3_52[11]}
   );
   gpc1_1 gpc3947 (
      {stage2_52[22]},
      {stage3_52[12]}
   );
   gpc1_1 gpc3948 (
      {stage2_52[23]},
      {stage3_52[13]}
   );
   gpc1_1 gpc3949 (
      {stage2_52[24]},
      {stage3_52[14]}
   );
   gpc1_1 gpc3950 (
      {stage2_52[25]},
      {stage3_52[15]}
   );
   gpc1_1 gpc3951 (
      {stage2_52[26]},
      {stage3_52[16]}
   );
   gpc1_1 gpc3952 (
      {stage2_52[27]},
      {stage3_52[17]}
   );
   gpc1_1 gpc3953 (
      {stage2_52[28]},
      {stage3_52[18]}
   );
   gpc1_1 gpc3954 (
      {stage2_52[29]},
      {stage3_52[19]}
   );
   gpc1_1 gpc3955 (
      {stage2_52[30]},
      {stage3_52[20]}
   );
   gpc1_1 gpc3956 (
      {stage2_52[31]},
      {stage3_52[21]}
   );
   gpc1_1 gpc3957 (
      {stage2_52[32]},
      {stage3_52[22]}
   );
   gpc1_1 gpc3958 (
      {stage2_52[33]},
      {stage3_52[23]}
   );
   gpc1_1 gpc3959 (
      {stage2_53[46]},
      {stage3_53[11]}
   );
   gpc1_1 gpc3960 (
      {stage2_53[47]},
      {stage3_53[12]}
   );
   gpc1_1 gpc3961 (
      {stage2_53[48]},
      {stage3_53[13]}
   );
   gpc1_1 gpc3962 (
      {stage2_53[49]},
      {stage3_53[14]}
   );
   gpc1_1 gpc3963 (
      {stage2_53[50]},
      {stage3_53[15]}
   );
   gpc1_1 gpc3964 (
      {stage2_55[35]},
      {stage3_55[15]}
   );
   gpc1_1 gpc3965 (
      {stage2_55[36]},
      {stage3_55[16]}
   );
   gpc1_1 gpc3966 (
      {stage2_55[37]},
      {stage3_55[17]}
   );
   gpc1_1 gpc3967 (
      {stage2_56[33]},
      {stage3_56[11]}
   );
   gpc1_1 gpc3968 (
      {stage2_56[34]},
      {stage3_56[12]}
   );
   gpc1_1 gpc3969 (
      {stage2_56[35]},
      {stage3_56[13]}
   );
   gpc1_1 gpc3970 (
      {stage2_56[36]},
      {stage3_56[14]}
   );
   gpc1_1 gpc3971 (
      {stage2_56[37]},
      {stage3_56[15]}
   );
   gpc1_1 gpc3972 (
      {stage2_56[38]},
      {stage3_56[16]}
   );
   gpc1_1 gpc3973 (
      {stage2_56[39]},
      {stage3_56[17]}
   );
   gpc1_1 gpc3974 (
      {stage2_56[40]},
      {stage3_56[18]}
   );
   gpc1_1 gpc3975 (
      {stage2_56[41]},
      {stage3_56[19]}
   );
   gpc1_1 gpc3976 (
      {stage2_56[42]},
      {stage3_56[20]}
   );
   gpc1_1 gpc3977 (
      {stage2_56[43]},
      {stage3_56[21]}
   );
   gpc1_1 gpc3978 (
      {stage2_56[44]},
      {stage3_56[22]}
   );
   gpc1_1 gpc3979 (
      {stage2_56[45]},
      {stage3_56[23]}
   );
   gpc1_1 gpc3980 (
      {stage2_56[46]},
      {stage3_56[24]}
   );
   gpc1_1 gpc3981 (
      {stage2_56[47]},
      {stage3_56[25]}
   );
   gpc1_1 gpc3982 (
      {stage2_56[48]},
      {stage3_56[26]}
   );
   gpc1_1 gpc3983 (
      {stage2_56[49]},
      {stage3_56[27]}
   );
   gpc1_1 gpc3984 (
      {stage2_56[50]},
      {stage3_56[28]}
   );
   gpc1_1 gpc3985 (
      {stage2_56[51]},
      {stage3_56[29]}
   );
   gpc1_1 gpc3986 (
      {stage2_56[52]},
      {stage3_56[30]}
   );
   gpc1_1 gpc3987 (
      {stage2_58[13]},
      {stage3_58[13]}
   );
   gpc1_1 gpc3988 (
      {stage2_58[14]},
      {stage3_58[14]}
   );
   gpc1_1 gpc3989 (
      {stage2_58[15]},
      {stage3_58[15]}
   );
   gpc1_1 gpc3990 (
      {stage2_58[16]},
      {stage3_58[16]}
   );
   gpc1_1 gpc3991 (
      {stage2_58[17]},
      {stage3_58[17]}
   );
   gpc1_1 gpc3992 (
      {stage2_58[18]},
      {stage3_58[18]}
   );
   gpc1_1 gpc3993 (
      {stage2_58[19]},
      {stage3_58[19]}
   );
   gpc1_1 gpc3994 (
      {stage2_58[20]},
      {stage3_58[20]}
   );
   gpc1_1 gpc3995 (
      {stage2_58[21]},
      {stage3_58[21]}
   );
   gpc1_1 gpc3996 (
      {stage2_58[22]},
      {stage3_58[22]}
   );
   gpc1_1 gpc3997 (
      {stage2_58[23]},
      {stage3_58[23]}
   );
   gpc1_1 gpc3998 (
      {stage2_58[24]},
      {stage3_58[24]}
   );
   gpc1_1 gpc3999 (
      {stage2_58[25]},
      {stage3_58[25]}
   );
   gpc1_1 gpc4000 (
      {stage2_58[26]},
      {stage3_58[26]}
   );
   gpc1_1 gpc4001 (
      {stage2_58[27]},
      {stage3_58[27]}
   );
   gpc1_1 gpc4002 (
      {stage2_58[28]},
      {stage3_58[28]}
   );
   gpc1_1 gpc4003 (
      {stage2_58[29]},
      {stage3_58[29]}
   );
   gpc1_1 gpc4004 (
      {stage2_58[30]},
      {stage3_58[30]}
   );
   gpc1_1 gpc4005 (
      {stage2_58[31]},
      {stage3_58[31]}
   );
   gpc1_1 gpc4006 (
      {stage2_58[32]},
      {stage3_58[32]}
   );
   gpc1_1 gpc4007 (
      {stage2_59[70]},
      {stage3_59[17]}
   );
   gpc1_1 gpc4008 (
      {stage2_59[71]},
      {stage3_59[18]}
   );
   gpc1_1 gpc4009 (
      {stage2_59[72]},
      {stage3_59[19]}
   );
   gpc1_1 gpc4010 (
      {stage2_59[73]},
      {stage3_59[20]}
   );
   gpc1_1 gpc4011 (
      {stage2_59[74]},
      {stage3_59[21]}
   );
   gpc1_1 gpc4012 (
      {stage2_59[75]},
      {stage3_59[22]}
   );
   gpc1_1 gpc4013 (
      {stage2_59[76]},
      {stage3_59[23]}
   );
   gpc1_1 gpc4014 (
      {stage2_59[77]},
      {stage3_59[24]}
   );
   gpc1_1 gpc4015 (
      {stage2_59[78]},
      {stage3_59[25]}
   );
   gpc1_1 gpc4016 (
      {stage2_59[79]},
      {stage3_59[26]}
   );
   gpc1_1 gpc4017 (
      {stage2_59[80]},
      {stage3_59[27]}
   );
   gpc1_1 gpc4018 (
      {stage2_61[59]},
      {stage3_61[17]}
   );
   gpc1_1 gpc4019 (
      {stage2_61[60]},
      {stage3_61[18]}
   );
   gpc1_1 gpc4020 (
      {stage2_61[61]},
      {stage3_61[19]}
   );
   gpc1_1 gpc4021 (
      {stage2_61[62]},
      {stage3_61[20]}
   );
   gpc1_1 gpc4022 (
      {stage2_61[63]},
      {stage3_61[21]}
   );
   gpc1_1 gpc4023 (
      {stage2_61[64]},
      {stage3_61[22]}
   );
   gpc1_1 gpc4024 (
      {stage2_61[65]},
      {stage3_61[23]}
   );
   gpc1_1 gpc4025 (
      {stage2_61[66]},
      {stage3_61[24]}
   );
   gpc1_1 gpc4026 (
      {stage2_64[29]},
      {stage3_64[12]}
   );
   gpc1_1 gpc4027 (
      {stage2_64[30]},
      {stage3_64[13]}
   );
   gpc1_1 gpc4028 (
      {stage2_64[31]},
      {stage3_64[14]}
   );
   gpc1_1 gpc4029 (
      {stage2_64[32]},
      {stage3_64[15]}
   );
   gpc1_1 gpc4030 (
      {stage2_64[33]},
      {stage3_64[16]}
   );
   gpc1_1 gpc4031 (
      {stage2_64[34]},
      {stage3_64[17]}
   );
   gpc1_1 gpc4032 (
      {stage2_64[35]},
      {stage3_64[18]}
   );
   gpc1_1 gpc4033 (
      {stage2_64[36]},
      {stage3_64[19]}
   );
   gpc1_1 gpc4034 (
      {stage2_64[37]},
      {stage3_64[20]}
   );
   gpc1_1 gpc4035 (
      {stage2_64[38]},
      {stage3_64[21]}
   );
   gpc1_1 gpc4036 (
      {stage2_64[39]},
      {stage3_64[22]}
   );
   gpc1_1 gpc4037 (
      {stage2_64[40]},
      {stage3_64[23]}
   );
   gpc1_1 gpc4038 (
      {stage2_64[41]},
      {stage3_64[24]}
   );
   gpc1_1 gpc4039 (
      {stage2_64[42]},
      {stage3_64[25]}
   );
   gpc1_1 gpc4040 (
      {stage2_64[43]},
      {stage3_64[26]}
   );
   gpc1_1 gpc4041 (
      {stage2_64[44]},
      {stage3_64[27]}
   );
   gpc1_1 gpc4042 (
      {stage2_64[45]},
      {stage3_64[28]}
   );
   gpc1_1 gpc4043 (
      {stage2_65[10]},
      {stage3_65[11]}
   );
   gpc1_1 gpc4044 (
      {stage2_65[11]},
      {stage3_65[12]}
   );
   gpc1_1 gpc4045 (
      {stage2_65[12]},
      {stage3_65[13]}
   );
   gpc1_1 gpc4046 (
      {stage2_67[0]},
      {stage3_67[3]}
   );
   gpc1_1 gpc4047 (
      {stage2_67[1]},
      {stage3_67[4]}
   );
   gpc1163_5 gpc4048 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[0]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1163_5 gpc4049 (
      {stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_2[1]},
      {stage3_3[1]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc615_5 gpc4050 (
      {stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5], stage3_2[6]},
      {stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc606_5 gpc4051 (
      {stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6], stage3_3[7], stage3_3[8]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[3],stage4_3[3]}
   );
   gpc606_5 gpc4052 (
      {stage3_3[9], stage3_3[10], stage3_3[11], stage3_3[12], stage3_3[13], 1'b0},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[4],stage4_3[4]}
   );
   gpc615_5 gpc4053 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_5[12]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[2],stage4_6[3],stage4_5[3],stage4_4[5]}
   );
   gpc615_5 gpc4054 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[4]}
   );
   gpc207_4 gpc4055 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_9[0], stage3_9[1]},
      {stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[4]}
   );
   gpc207_4 gpc4056 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14]},
      {stage3_9[2], stage3_9[3]},
      {stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc4057 (
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[3],stage4_9[3],stage4_8[4]}
   );
   gpc2135_5 gpc4058 (
      {stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7], stage3_9[8]},
      {stage3_10[6], stage3_10[7], stage3_10[8]},
      {stage3_11[0]},
      {stage3_12[0], stage3_12[1]},
      {stage4_13[0],stage4_12[1],stage4_11[1],stage4_10[4],stage4_9[4]}
   );
   gpc606_5 gpc4059 (
      {stage3_9[9], stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14]},
      {stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5], stage3_11[6]},
      {stage4_13[1],stage4_12[2],stage4_11[2],stage4_10[5],stage4_9[5]}
   );
   gpc606_5 gpc4060 (
      {stage3_9[15], stage3_9[16], stage3_9[17], stage3_9[18], stage3_9[19], stage3_9[20]},
      {stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11], stage3_11[12]},
      {stage4_13[2],stage4_12[3],stage4_11[3],stage4_10[6],stage4_9[6]}
   );
   gpc2135_5 gpc4061 (
      {stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage3_11[13], stage3_11[14], stage3_11[15]},
      {stage3_12[2]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[0],stage4_13[3],stage4_12[4],stage4_11[4],stage4_10[7]}
   );
   gpc207_4 gpc4062 (
      {stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage3_14[0], stage3_14[1]},
      {stage4_15[0],stage4_14[1],stage4_13[4],stage4_12[5]}
   );
   gpc207_4 gpc4063 (
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16]},
      {stage3_14[2], stage3_14[3]},
      {stage4_15[1],stage4_14[2],stage4_13[5],stage4_12[6]}
   );
   gpc606_5 gpc4064 (
      {stage3_12[17], stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22]},
      {stage3_14[4], stage3_14[5], stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9]},
      {stage4_16[0],stage4_15[2],stage4_14[3],stage4_13[6],stage4_12[7]}
   );
   gpc606_5 gpc4065 (
      {stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[3],stage4_14[4],stage4_13[7]}
   );
   gpc606_5 gpc4066 (
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[4],stage4_14[5],stage4_13[8]}
   );
   gpc606_5 gpc4067 (
      {stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[3],stage4_15[5],stage4_14[6],stage4_13[9]}
   );
   gpc117_4 gpc4068 (
      {stage3_14[10], stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[18]},
      {stage3_16[0]},
      {stage4_17[3],stage4_16[4],stage4_15[6],stage4_14[7]}
   );
   gpc117_4 gpc4069 (
      {stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage3_15[19]},
      {stage3_16[1]},
      {stage4_17[4],stage4_16[5],stage4_15[7],stage4_14[8]}
   );
   gpc117_4 gpc4070 (
      {stage3_14[24], stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage3_15[20]},
      {stage3_16[2]},
      {stage4_17[5],stage4_16[6],stage4_15[8],stage4_14[9]}
   );
   gpc117_4 gpc4071 (
      {stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35], 1'b0, 1'b0},
      {stage3_15[21]},
      {stage3_16[3]},
      {stage4_17[6],stage4_16[7],stage4_15[9],stage4_14[10]}
   );
   gpc615_5 gpc4072 (
      {stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25], stage3_15[26]},
      {stage3_16[4]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[0],stage4_17[7],stage4_16[8],stage4_15[10]}
   );
   gpc615_5 gpc4073 (
      {stage3_15[27], stage3_15[28], stage3_15[29], stage3_15[30], stage3_15[31]},
      {stage3_16[5]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[1],stage4_17[8],stage4_16[9],stage4_15[11]}
   );
   gpc606_5 gpc4074 (
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[2],stage4_18[2],stage4_17[9],stage4_16[10]}
   );
   gpc606_5 gpc4075 (
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[3],stage4_18[3],stage4_17[10],stage4_16[11]}
   );
   gpc606_5 gpc4076 (
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], 1'b0, 1'b0},
      {stage3_18[12], stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17]},
      {stage4_20[2],stage4_19[4],stage4_18[4],stage4_17[11],stage4_16[12]}
   );
   gpc615_5 gpc4077 (
      {stage3_18[18], stage3_18[19], stage3_18[20], stage3_18[21], stage3_18[22]},
      {stage3_19[0]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[3],stage4_19[5],stage4_18[5]}
   );
   gpc615_5 gpc4078 (
      {stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage3_20[6]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[1],stage4_21[1],stage4_20[4],stage4_19[6]}
   );
   gpc615_5 gpc4079 (
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10]},
      {stage3_20[7]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[2],stage4_21[2],stage4_20[5],stage4_19[7]}
   );
   gpc615_5 gpc4080 (
      {stage3_19[11], stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15]},
      {stage3_20[8]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[3],stage4_21[3],stage4_20[6],stage4_19[8]}
   );
   gpc615_5 gpc4081 (
      {stage3_19[16], stage3_19[17], stage3_19[18], stage3_19[19], stage3_19[20]},
      {stage3_20[9]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[4],stage4_21[4],stage4_20[7],stage4_19[9]}
   );
   gpc606_5 gpc4082 (
      {stage3_20[10], stage3_20[11], stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[4],stage4_22[5],stage4_21[5],stage4_20[8]}
   );
   gpc606_5 gpc4083 (
      {stage3_20[16], stage3_20[17], stage3_20[18], stage3_20[19], stage3_20[20], stage3_20[21]},
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11]},
      {stage4_24[1],stage4_23[5],stage4_22[6],stage4_21[6],stage4_20[9]}
   );
   gpc615_5 gpc4084 (
      {stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16]},
      {stage3_23[0]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[0],stage4_24[2],stage4_23[6],stage4_22[7]}
   );
   gpc615_5 gpc4085 (
      {stage3_22[17], stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21]},
      {stage3_23[1]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[1],stage4_24[3],stage4_23[7],stage4_22[8]}
   );
   gpc615_5 gpc4086 (
      {stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage3_24[12]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[2],stage4_25[2],stage4_24[4],stage4_23[8]}
   );
   gpc615_5 gpc4087 (
      {stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage3_24[13]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[3],stage4_25[3],stage4_24[5],stage4_23[9]}
   );
   gpc615_5 gpc4088 (
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16]},
      {stage3_26[0]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[2],stage4_26[4],stage4_25[4]}
   );
   gpc615_5 gpc4089 (
      {stage3_25[17], stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21]},
      {stage3_26[1]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[1],stage4_27[3],stage4_26[5],stage4_25[5]}
   );
   gpc117_4 gpc4090 (
      {stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5], stage3_26[6], stage3_26[7], stage3_26[8]},
      {stage3_27[12]},
      {stage3_28[0]},
      {stage4_29[2],stage4_28[2],stage4_27[4],stage4_26[6]}
   );
   gpc207_4 gpc4091 (
      {stage3_26[9], stage3_26[10], stage3_26[11], stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15]},
      {stage3_28[1], stage3_28[2]},
      {stage4_29[3],stage4_28[3],stage4_27[5],stage4_26[7]}
   );
   gpc606_5 gpc4092 (
      {stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17], stage3_27[18]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[0],stage4_29[4],stage4_28[4],stage4_27[6]}
   );
   gpc606_5 gpc4093 (
      {stage3_28[3], stage3_28[4], stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[5],stage4_28[5]}
   );
   gpc606_5 gpc4094 (
      {stage3_28[9], stage3_28[10], stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[2],stage4_30[2],stage4_29[6],stage4_28[6]}
   );
   gpc606_5 gpc4095 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[2],stage4_31[3],stage4_30[3],stage4_29[7]}
   );
   gpc606_5 gpc4096 (
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[3],stage4_31[4],stage4_30[4],stage4_29[8]}
   );
   gpc606_5 gpc4097 (
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[4],stage4_31[5],stage4_30[5],stage4_29[9]}
   );
   gpc615_5 gpc4098 (
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16]},
      {stage3_31[18]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[3],stage4_32[5],stage4_31[6],stage4_30[6]}
   );
   gpc606_5 gpc4099 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[0],stage4_34[1],stage4_33[4],stage4_32[6]}
   );
   gpc606_5 gpc4100 (
      {stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[1],stage4_34[2],stage4_33[5],stage4_32[7]}
   );
   gpc606_5 gpc4101 (
      {stage3_32[18], stage3_32[19], stage3_32[20], stage3_32[21], stage3_32[22], stage3_32[23]},
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage4_36[2],stage4_35[2],stage4_34[3],stage4_33[6],stage4_32[8]}
   );
   gpc606_5 gpc4102 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[3],stage4_35[3],stage4_34[4],stage4_33[7]}
   );
   gpc606_5 gpc4103 (
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[1],stage4_36[4],stage4_35[4],stage4_34[5],stage4_33[8]}
   );
   gpc1343_5 gpc4104 (
      {stage3_35[12], stage3_35[13], stage3_35[14]},
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3]},
      {stage3_37[0], stage3_37[1], stage3_37[2]},
      {stage3_38[0]},
      {stage4_39[0],stage4_38[0],stage4_37[2],stage4_36[5],stage4_35[5]}
   );
   gpc1343_5 gpc4105 (
      {stage3_35[15], stage3_35[16], stage3_35[17]},
      {stage3_36[4], stage3_36[5], stage3_36[6], stage3_36[7]},
      {stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage3_38[1]},
      {stage4_39[1],stage4_38[1],stage4_37[3],stage4_36[6],stage4_35[6]}
   );
   gpc1343_5 gpc4106 (
      {stage3_35[18], stage3_35[19], stage3_35[20]},
      {stage3_36[8], stage3_36[9], stage3_36[10], stage3_36[11]},
      {stage3_37[6], stage3_37[7], stage3_37[8]},
      {stage3_38[2]},
      {stage4_39[2],stage4_38[2],stage4_37[4],stage4_36[7],stage4_35[7]}
   );
   gpc1343_5 gpc4107 (
      {stage3_35[21], stage3_35[22], stage3_35[23]},
      {stage3_36[12], stage3_36[13], stage3_36[14], stage3_36[15]},
      {stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage3_38[3]},
      {stage4_39[3],stage4_38[3],stage4_37[5],stage4_36[8],stage4_35[8]}
   );
   gpc615_5 gpc4108 (
      {stage3_38[4], stage3_38[5], stage3_38[6], stage3_38[7], stage3_38[8]},
      {stage3_39[0]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[0],stage4_40[0],stage4_39[4],stage4_38[4]}
   );
   gpc615_5 gpc4109 (
      {stage3_38[9], stage3_38[10], stage3_38[11], stage3_38[12], stage3_38[13]},
      {stage3_39[1]},
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage4_42[1],stage4_41[1],stage4_40[1],stage4_39[5],stage4_38[5]}
   );
   gpc117_4 gpc4110 (
      {stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5], stage3_39[6], stage3_39[7], stage3_39[8]},
      {stage3_40[12]},
      {stage3_41[0]},
      {stage4_42[2],stage4_41[2],stage4_40[2],stage4_39[6]}
   );
   gpc117_4 gpc4111 (
      {stage3_39[9], stage3_39[10], stage3_39[11], stage3_39[12], stage3_39[13], stage3_39[14], stage3_39[15]},
      {stage3_40[13]},
      {stage3_41[1]},
      {stage4_42[3],stage4_41[3],stage4_40[3],stage4_39[7]}
   );
   gpc117_4 gpc4112 (
      {stage3_39[16], stage3_39[17], stage3_39[18], stage3_39[19], stage3_39[20], stage3_39[21], stage3_39[22]},
      {stage3_40[14]},
      {stage3_41[2]},
      {stage4_42[4],stage4_41[4],stage4_40[4],stage4_39[8]}
   );
   gpc606_5 gpc4113 (
      {stage3_41[3], stage3_41[4], stage3_41[5], stage3_41[6], stage3_41[7], stage3_41[8]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[0],stage4_42[5],stage4_41[5]}
   );
   gpc606_5 gpc4114 (
      {stage3_41[9], stage3_41[10], stage3_41[11], stage3_41[12], stage3_41[13], stage3_41[14]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[1],stage4_43[1],stage4_42[6],stage4_41[6]}
   );
   gpc615_5 gpc4115 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4]},
      {stage3_43[12]},
      {stage3_44[0], stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage4_46[0],stage4_45[2],stage4_44[2],stage4_43[2],stage4_42[7]}
   );
   gpc615_5 gpc4116 (
      {stage3_42[5], stage3_42[6], stage3_42[7], stage3_42[8], stage3_42[9]},
      {stage3_43[13]},
      {stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9], stage3_44[10], stage3_44[11]},
      {stage4_46[1],stage4_45[3],stage4_44[3],stage4_43[3],stage4_42[8]}
   );
   gpc615_5 gpc4117 (
      {stage3_42[10], stage3_42[11], stage3_42[12], stage3_42[13], stage3_42[14]},
      {stage3_43[14]},
      {stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15], stage3_44[16], stage3_44[17]},
      {stage4_46[2],stage4_45[4],stage4_44[4],stage4_43[4],stage4_42[9]}
   );
   gpc615_5 gpc4118 (
      {stage3_42[15], stage3_42[16], stage3_42[17], stage3_42[18], stage3_42[19]},
      {stage3_43[15]},
      {stage3_44[18], stage3_44[19], stage3_44[20], stage3_44[21], stage3_44[22], stage3_44[23]},
      {stage4_46[3],stage4_45[5],stage4_44[5],stage4_43[5],stage4_42[10]}
   );
   gpc615_5 gpc4119 (
      {stage3_43[16], stage3_43[17], stage3_43[18], stage3_43[19], stage3_43[20]},
      {stage3_44[24]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[4],stage4_45[6],stage4_44[6],stage4_43[6]}
   );
   gpc606_5 gpc4120 (
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage3_47[0], stage3_47[1], stage3_47[2], stage3_47[3], stage3_47[4], stage3_47[5]},
      {stage4_49[0],stage4_48[0],stage4_47[1],stage4_46[5],stage4_45[7]}
   );
   gpc606_5 gpc4121 (
      {stage3_45[12], stage3_45[13], stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage3_47[6], stage3_47[7], stage3_47[8], stage3_47[9], stage3_47[10], stage3_47[11]},
      {stage4_49[1],stage4_48[1],stage4_47[2],stage4_46[6],stage4_45[8]}
   );
   gpc207_4 gpc4122 (
      {stage3_46[0], stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5], stage3_46[6]},
      {stage3_48[0], stage3_48[1]},
      {stage4_49[2],stage4_48[2],stage4_47[3],stage4_46[7]}
   );
   gpc606_5 gpc4123 (
      {stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5], stage3_48[6], stage3_48[7]},
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage4_52[0],stage4_51[0],stage4_50[0],stage4_49[3],stage4_48[3]}
   );
   gpc606_5 gpc4124 (
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[1],stage4_51[1],stage4_50[1],stage4_49[4]}
   );
   gpc7_3 gpc4125 (
      {stage3_50[6], stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12]},
      {stage4_52[2],stage4_51[2],stage4_50[2]}
   );
   gpc606_5 gpc4126 (
      {stage3_50[13], stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17], stage3_50[18]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[1],stage4_52[3],stage4_51[3],stage4_50[3]}
   );
   gpc606_5 gpc4127 (
      {stage3_50[19], stage3_50[20], stage3_50[21], stage3_50[22], stage3_50[23], stage3_50[24]},
      {stage3_52[6], stage3_52[7], stage3_52[8], stage3_52[9], stage3_52[10], stage3_52[11]},
      {stage4_54[1],stage4_53[2],stage4_52[4],stage4_51[4],stage4_50[4]}
   );
   gpc606_5 gpc4128 (
      {stage3_50[25], stage3_50[26], stage3_50[27], stage3_50[28], stage3_50[29], stage3_50[30]},
      {stage3_52[12], stage3_52[13], stage3_52[14], stage3_52[15], stage3_52[16], stage3_52[17]},
      {stage4_54[2],stage4_53[3],stage4_52[5],stage4_51[5],stage4_50[5]}
   );
   gpc606_5 gpc4129 (
      {stage3_51[6], stage3_51[7], stage3_51[8], stage3_51[9], stage3_51[10], stage3_51[11]},
      {stage3_53[0], stage3_53[1], stage3_53[2], stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage4_55[0],stage4_54[3],stage4_53[4],stage4_52[6],stage4_51[6]}
   );
   gpc615_5 gpc4130 (
      {stage3_52[18], stage3_52[19], stage3_52[20], stage3_52[21], stage3_52[22]},
      {stage3_53[6]},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage4_56[0],stage4_55[1],stage4_54[4],stage4_53[5],stage4_52[7]}
   );
   gpc606_5 gpc4131 (
      {stage3_54[6], stage3_54[7], stage3_54[8], stage3_54[9], stage3_54[10], stage3_54[11]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage4_58[0],stage4_57[0],stage4_56[1],stage4_55[2],stage4_54[5]}
   );
   gpc615_5 gpc4132 (
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4]},
      {stage3_56[6]},
      {stage3_57[0], stage3_57[1], stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage4_59[0],stage4_58[1],stage4_57[1],stage4_56[2],stage4_55[3]}
   );
   gpc606_5 gpc4133 (
      {stage3_56[7], stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11], stage3_56[12]},
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage4_60[0],stage4_59[1],stage4_58[2],stage4_57[2],stage4_56[3]}
   );
   gpc606_5 gpc4134 (
      {stage3_56[13], stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17], stage3_56[18]},
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11]},
      {stage4_60[1],stage4_59[2],stage4_58[3],stage4_57[3],stage4_56[4]}
   );
   gpc615_5 gpc4135 (
      {stage3_56[19], stage3_56[20], stage3_56[21], stage3_56[22], stage3_56[23]},
      {stage3_57[6]},
      {stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15], stage3_58[16], stage3_58[17]},
      {stage4_60[2],stage4_59[3],stage4_58[4],stage4_57[4],stage4_56[5]}
   );
   gpc606_5 gpc4136 (
      {stage3_57[7], stage3_57[8], stage3_57[9], stage3_57[10], stage3_57[11], stage3_57[12]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[3],stage4_59[4],stage4_58[5],stage4_57[5]}
   );
   gpc606_5 gpc4137 (
      {stage3_59[6], stage3_59[7], stage3_59[8], stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {stage4_63[0],stage4_62[0],stage4_61[1],stage4_60[4],stage4_59[5]}
   );
   gpc606_5 gpc4138 (
      {stage3_59[12], stage3_59[13], stage3_59[14], stage3_59[15], stage3_59[16], stage3_59[17]},
      {stage3_61[6], stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11]},
      {stage4_63[1],stage4_62[1],stage4_61[2],stage4_60[5],stage4_59[6]}
   );
   gpc606_5 gpc4139 (
      {stage3_60[0], stage3_60[1], stage3_60[2], stage3_60[3], stage3_60[4], stage3_60[5]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[2],stage4_62[2],stage4_61[3],stage4_60[6]}
   );
   gpc606_5 gpc4140 (
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage4_66[0],stage4_65[0],stage4_64[1],stage4_63[3],stage4_62[3]}
   );
   gpc606_5 gpc4141 (
      {stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15], stage3_62[16], stage3_62[17]},
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage4_66[1],stage4_65[1],stage4_64[2],stage4_63[4],stage4_62[4]}
   );
   gpc606_5 gpc4142 (
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[2],stage4_65[2],stage4_64[3],stage4_63[5]}
   );
   gpc606_5 gpc4143 (
      {stage3_63[6], stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11]},
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage4_67[1],stage4_66[3],stage4_65[3],stage4_64[4],stage4_63[6]}
   );
   gpc1_1 gpc4144 (
      {stage3_0[6]},
      {stage4_0[2]}
   );
   gpc1_1 gpc4145 (
      {stage3_0[7]},
      {stage4_0[3]}
   );
   gpc1_1 gpc4146 (
      {stage3_1[12]},
      {stage4_1[2]}
   );
   gpc1_1 gpc4147 (
      {stage3_1[13]},
      {stage4_1[3]}
   );
   gpc1_1 gpc4148 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc4149 (
      {stage3_2[8]},
      {stage4_2[4]}
   );
   gpc1_1 gpc4150 (
      {stage3_2[9]},
      {stage4_2[5]}
   );
   gpc1_1 gpc4151 (
      {stage3_2[10]},
      {stage4_2[6]}
   );
   gpc1_1 gpc4152 (
      {stage3_4[11]},
      {stage4_4[6]}
   );
   gpc1_1 gpc4153 (
      {stage3_4[12]},
      {stage4_4[7]}
   );
   gpc1_1 gpc4154 (
      {stage3_4[13]},
      {stage4_4[8]}
   );
   gpc1_1 gpc4155 (
      {stage3_5[13]},
      {stage4_5[4]}
   );
   gpc1_1 gpc4156 (
      {stage3_5[14]},
      {stage4_5[5]}
   );
   gpc1_1 gpc4157 (
      {stage3_5[15]},
      {stage4_5[6]}
   );
   gpc1_1 gpc4158 (
      {stage3_5[16]},
      {stage4_5[7]}
   );
   gpc1_1 gpc4159 (
      {stage3_5[17]},
      {stage4_5[8]}
   );
   gpc1_1 gpc4160 (
      {stage3_6[11]},
      {stage4_6[5]}
   );
   gpc1_1 gpc4161 (
      {stage3_6[12]},
      {stage4_6[6]}
   );
   gpc1_1 gpc4162 (
      {stage3_6[13]},
      {stage4_6[7]}
   );
   gpc1_1 gpc4163 (
      {stage3_6[14]},
      {stage4_6[8]}
   );
   gpc1_1 gpc4164 (
      {stage3_6[15]},
      {stage4_6[9]}
   );
   gpc1_1 gpc4165 (
      {stage3_6[16]},
      {stage4_6[10]}
   );
   gpc1_1 gpc4166 (
      {stage3_6[17]},
      {stage4_6[11]}
   );
   gpc1_1 gpc4167 (
      {stage3_6[18]},
      {stage4_6[12]}
   );
   gpc1_1 gpc4168 (
      {stage3_6[19]},
      {stage4_6[13]}
   );
   gpc1_1 gpc4169 (
      {stage3_7[15]},
      {stage4_7[6]}
   );
   gpc1_1 gpc4170 (
      {stage3_7[16]},
      {stage4_7[7]}
   );
   gpc1_1 gpc4171 (
      {stage3_8[12]},
      {stage4_8[5]}
   );
   gpc1_1 gpc4172 (
      {stage3_8[13]},
      {stage4_8[6]}
   );
   gpc1_1 gpc4173 (
      {stage3_8[14]},
      {stage4_8[7]}
   );
   gpc1_1 gpc4174 (
      {stage3_8[15]},
      {stage4_8[8]}
   );
   gpc1_1 gpc4175 (
      {stage3_8[16]},
      {stage4_8[9]}
   );
   gpc1_1 gpc4176 (
      {stage3_10[14]},
      {stage4_10[8]}
   );
   gpc1_1 gpc4177 (
      {stage3_11[16]},
      {stage4_11[5]}
   );
   gpc1_1 gpc4178 (
      {stage3_11[17]},
      {stage4_11[6]}
   );
   gpc1_1 gpc4179 (
      {stage3_12[23]},
      {stage4_12[8]}
   );
   gpc1_1 gpc4180 (
      {stage3_15[32]},
      {stage4_15[12]}
   );
   gpc1_1 gpc4181 (
      {stage3_15[33]},
      {stage4_15[13]}
   );
   gpc1_1 gpc4182 (
      {stage3_15[34]},
      {stage4_15[14]}
   );
   gpc1_1 gpc4183 (
      {stage3_15[35]},
      {stage4_15[15]}
   );
   gpc1_1 gpc4184 (
      {stage3_15[36]},
      {stage4_15[16]}
   );
   gpc1_1 gpc4185 (
      {stage3_17[12]},
      {stage4_17[12]}
   );
   gpc1_1 gpc4186 (
      {stage3_17[13]},
      {stage4_17[13]}
   );
   gpc1_1 gpc4187 (
      {stage3_17[14]},
      {stage4_17[14]}
   );
   gpc1_1 gpc4188 (
      {stage3_17[15]},
      {stage4_17[15]}
   );
   gpc1_1 gpc4189 (
      {stage3_17[16]},
      {stage4_17[16]}
   );
   gpc1_1 gpc4190 (
      {stage3_19[21]},
      {stage4_19[10]}
   );
   gpc1_1 gpc4191 (
      {stage3_19[22]},
      {stage4_19[11]}
   );
   gpc1_1 gpc4192 (
      {stage3_19[23]},
      {stage4_19[12]}
   );
   gpc1_1 gpc4193 (
      {stage3_19[24]},
      {stage4_19[13]}
   );
   gpc1_1 gpc4194 (
      {stage3_19[25]},
      {stage4_19[14]}
   );
   gpc1_1 gpc4195 (
      {stage3_19[26]},
      {stage4_19[15]}
   );
   gpc1_1 gpc4196 (
      {stage3_20[22]},
      {stage4_20[10]}
   );
   gpc1_1 gpc4197 (
      {stage3_21[24]},
      {stage4_21[7]}
   );
   gpc1_1 gpc4198 (
      {stage3_22[22]},
      {stage4_22[9]}
   );
   gpc1_1 gpc4199 (
      {stage3_22[23]},
      {stage4_22[10]}
   );
   gpc1_1 gpc4200 (
      {stage3_22[24]},
      {stage4_22[11]}
   );
   gpc1_1 gpc4201 (
      {stage3_22[25]},
      {stage4_22[12]}
   );
   gpc1_1 gpc4202 (
      {stage3_22[26]},
      {stage4_22[13]}
   );
   gpc1_1 gpc4203 (
      {stage3_24[14]},
      {stage4_24[6]}
   );
   gpc1_1 gpc4204 (
      {stage3_24[15]},
      {stage4_24[7]}
   );
   gpc1_1 gpc4205 (
      {stage3_24[16]},
      {stage4_24[8]}
   );
   gpc1_1 gpc4206 (
      {stage3_24[17]},
      {stage4_24[9]}
   );
   gpc1_1 gpc4207 (
      {stage3_24[18]},
      {stage4_24[10]}
   );
   gpc1_1 gpc4208 (
      {stage3_24[19]},
      {stage4_24[11]}
   );
   gpc1_1 gpc4209 (
      {stage3_24[20]},
      {stage4_24[12]}
   );
   gpc1_1 gpc4210 (
      {stage3_24[21]},
      {stage4_24[13]}
   );
   gpc1_1 gpc4211 (
      {stage3_24[22]},
      {stage4_24[14]}
   );
   gpc1_1 gpc4212 (
      {stage3_24[23]},
      {stage4_24[15]}
   );
   gpc1_1 gpc4213 (
      {stage3_24[24]},
      {stage4_24[16]}
   );
   gpc1_1 gpc4214 (
      {stage3_24[25]},
      {stage4_24[17]}
   );
   gpc1_1 gpc4215 (
      {stage3_28[15]},
      {stage4_28[7]}
   );
   gpc1_1 gpc4216 (
      {stage3_28[16]},
      {stage4_28[8]}
   );
   gpc1_1 gpc4217 (
      {stage3_28[17]},
      {stage4_28[9]}
   );
   gpc1_1 gpc4218 (
      {stage3_28[18]},
      {stage4_28[10]}
   );
   gpc1_1 gpc4219 (
      {stage3_28[19]},
      {stage4_28[11]}
   );
   gpc1_1 gpc4220 (
      {stage3_30[17]},
      {stage4_30[7]}
   );
   gpc1_1 gpc4221 (
      {stage3_30[18]},
      {stage4_30[8]}
   );
   gpc1_1 gpc4222 (
      {stage3_30[19]},
      {stage4_30[9]}
   );
   gpc1_1 gpc4223 (
      {stage3_30[20]},
      {stage4_30[10]}
   );
   gpc1_1 gpc4224 (
      {stage3_30[21]},
      {stage4_30[11]}
   );
   gpc1_1 gpc4225 (
      {stage3_30[22]},
      {stage4_30[12]}
   );
   gpc1_1 gpc4226 (
      {stage3_30[23]},
      {stage4_30[13]}
   );
   gpc1_1 gpc4227 (
      {stage3_30[24]},
      {stage4_30[14]}
   );
   gpc1_1 gpc4228 (
      {stage3_30[25]},
      {stage4_30[15]}
   );
   gpc1_1 gpc4229 (
      {stage3_31[19]},
      {stage4_31[7]}
   );
   gpc1_1 gpc4230 (
      {stage3_31[20]},
      {stage4_31[8]}
   );
   gpc1_1 gpc4231 (
      {stage3_32[24]},
      {stage4_32[9]}
   );
   gpc1_1 gpc4232 (
      {stage3_32[25]},
      {stage4_32[10]}
   );
   gpc1_1 gpc4233 (
      {stage3_32[26]},
      {stage4_32[11]}
   );
   gpc1_1 gpc4234 (
      {stage3_32[27]},
      {stage4_32[12]}
   );
   gpc1_1 gpc4235 (
      {stage3_32[28]},
      {stage4_32[13]}
   );
   gpc1_1 gpc4236 (
      {stage3_32[29]},
      {stage4_32[14]}
   );
   gpc1_1 gpc4237 (
      {stage3_32[30]},
      {stage4_32[15]}
   );
   gpc1_1 gpc4238 (
      {stage3_32[31]},
      {stage4_32[16]}
   );
   gpc1_1 gpc4239 (
      {stage3_32[32]},
      {stage4_32[17]}
   );
   gpc1_1 gpc4240 (
      {stage3_32[33]},
      {stage4_32[18]}
   );
   gpc1_1 gpc4241 (
      {stage3_32[34]},
      {stage4_32[19]}
   );
   gpc1_1 gpc4242 (
      {stage3_33[12]},
      {stage4_33[9]}
   );
   gpc1_1 gpc4243 (
      {stage3_33[13]},
      {stage4_33[10]}
   );
   gpc1_1 gpc4244 (
      {stage3_33[14]},
      {stage4_33[11]}
   );
   gpc1_1 gpc4245 (
      {stage3_34[18]},
      {stage4_34[6]}
   );
   gpc1_1 gpc4246 (
      {stage3_34[19]},
      {stage4_34[7]}
   );
   gpc1_1 gpc4247 (
      {stage3_34[20]},
      {stage4_34[8]}
   );
   gpc1_1 gpc4248 (
      {stage3_34[21]},
      {stage4_34[9]}
   );
   gpc1_1 gpc4249 (
      {stage3_34[22]},
      {stage4_34[10]}
   );
   gpc1_1 gpc4250 (
      {stage3_35[24]},
      {stage4_35[9]}
   );
   gpc1_1 gpc4251 (
      {stage3_35[25]},
      {stage4_35[10]}
   );
   gpc1_1 gpc4252 (
      {stage3_36[16]},
      {stage4_36[9]}
   );
   gpc1_1 gpc4253 (
      {stage3_39[23]},
      {stage4_39[9]}
   );
   gpc1_1 gpc4254 (
      {stage3_40[15]},
      {stage4_40[5]}
   );
   gpc1_1 gpc4255 (
      {stage3_40[16]},
      {stage4_40[6]}
   );
   gpc1_1 gpc4256 (
      {stage3_40[17]},
      {stage4_40[7]}
   );
   gpc1_1 gpc4257 (
      {stage3_40[18]},
      {stage4_40[8]}
   );
   gpc1_1 gpc4258 (
      {stage3_40[19]},
      {stage4_40[9]}
   );
   gpc1_1 gpc4259 (
      {stage3_40[20]},
      {stage4_40[10]}
   );
   gpc1_1 gpc4260 (
      {stage3_40[21]},
      {stage4_40[11]}
   );
   gpc1_1 gpc4261 (
      {stage3_40[22]},
      {stage4_40[12]}
   );
   gpc1_1 gpc4262 (
      {stage3_40[23]},
      {stage4_40[13]}
   );
   gpc1_1 gpc4263 (
      {stage3_41[15]},
      {stage4_41[7]}
   );
   gpc1_1 gpc4264 (
      {stage3_41[16]},
      {stage4_41[8]}
   );
   gpc1_1 gpc4265 (
      {stage3_41[17]},
      {stage4_41[9]}
   );
   gpc1_1 gpc4266 (
      {stage3_41[18]},
      {stage4_41[10]}
   );
   gpc1_1 gpc4267 (
      {stage3_41[19]},
      {stage4_41[11]}
   );
   gpc1_1 gpc4268 (
      {stage3_41[20]},
      {stage4_41[12]}
   );
   gpc1_1 gpc4269 (
      {stage3_41[21]},
      {stage4_41[13]}
   );
   gpc1_1 gpc4270 (
      {stage3_41[22]},
      {stage4_41[14]}
   );
   gpc1_1 gpc4271 (
      {stage3_41[23]},
      {stage4_41[15]}
   );
   gpc1_1 gpc4272 (
      {stage3_41[24]},
      {stage4_41[16]}
   );
   gpc1_1 gpc4273 (
      {stage3_42[20]},
      {stage4_42[11]}
   );
   gpc1_1 gpc4274 (
      {stage3_42[21]},
      {stage4_42[12]}
   );
   gpc1_1 gpc4275 (
      {stage3_42[22]},
      {stage4_42[13]}
   );
   gpc1_1 gpc4276 (
      {stage3_42[23]},
      {stage4_42[14]}
   );
   gpc1_1 gpc4277 (
      {stage3_42[24]},
      {stage4_42[15]}
   );
   gpc1_1 gpc4278 (
      {stage3_42[25]},
      {stage4_42[16]}
   );
   gpc1_1 gpc4279 (
      {stage3_44[25]},
      {stage4_44[7]}
   );
   gpc1_1 gpc4280 (
      {stage3_44[26]},
      {stage4_44[8]}
   );
   gpc1_1 gpc4281 (
      {stage3_44[27]},
      {stage4_44[9]}
   );
   gpc1_1 gpc4282 (
      {stage3_44[28]},
      {stage4_44[10]}
   );
   gpc1_1 gpc4283 (
      {stage3_44[29]},
      {stage4_44[11]}
   );
   gpc1_1 gpc4284 (
      {stage3_44[30]},
      {stage4_44[12]}
   );
   gpc1_1 gpc4285 (
      {stage3_46[7]},
      {stage4_46[8]}
   );
   gpc1_1 gpc4286 (
      {stage3_46[8]},
      {stage4_46[9]}
   );
   gpc1_1 gpc4287 (
      {stage3_46[9]},
      {stage4_46[10]}
   );
   gpc1_1 gpc4288 (
      {stage3_46[10]},
      {stage4_46[11]}
   );
   gpc1_1 gpc4289 (
      {stage3_46[11]},
      {stage4_46[12]}
   );
   gpc1_1 gpc4290 (
      {stage3_46[12]},
      {stage4_46[13]}
   );
   gpc1_1 gpc4291 (
      {stage3_46[13]},
      {stage4_46[14]}
   );
   gpc1_1 gpc4292 (
      {stage3_46[14]},
      {stage4_46[15]}
   );
   gpc1_1 gpc4293 (
      {stage3_46[15]},
      {stage4_46[16]}
   );
   gpc1_1 gpc4294 (
      {stage3_46[16]},
      {stage4_46[17]}
   );
   gpc1_1 gpc4295 (
      {stage3_47[12]},
      {stage4_47[4]}
   );
   gpc1_1 gpc4296 (
      {stage3_47[13]},
      {stage4_47[5]}
   );
   gpc1_1 gpc4297 (
      {stage3_47[14]},
      {stage4_47[6]}
   );
   gpc1_1 gpc4298 (
      {stage3_47[15]},
      {stage4_47[7]}
   );
   gpc1_1 gpc4299 (
      {stage3_47[16]},
      {stage4_47[8]}
   );
   gpc1_1 gpc4300 (
      {stage3_47[17]},
      {stage4_47[9]}
   );
   gpc1_1 gpc4301 (
      {stage3_47[18]},
      {stage4_47[10]}
   );
   gpc1_1 gpc4302 (
      {stage3_47[19]},
      {stage4_47[11]}
   );
   gpc1_1 gpc4303 (
      {stage3_47[20]},
      {stage4_47[12]}
   );
   gpc1_1 gpc4304 (
      {stage3_47[21]},
      {stage4_47[13]}
   );
   gpc1_1 gpc4305 (
      {stage3_47[22]},
      {stage4_47[14]}
   );
   gpc1_1 gpc4306 (
      {stage3_47[23]},
      {stage4_47[15]}
   );
   gpc1_1 gpc4307 (
      {stage3_48[8]},
      {stage4_48[4]}
   );
   gpc1_1 gpc4308 (
      {stage3_48[9]},
      {stage4_48[5]}
   );
   gpc1_1 gpc4309 (
      {stage3_48[10]},
      {stage4_48[6]}
   );
   gpc1_1 gpc4310 (
      {stage3_48[11]},
      {stage4_48[7]}
   );
   gpc1_1 gpc4311 (
      {stage3_48[12]},
      {stage4_48[8]}
   );
   gpc1_1 gpc4312 (
      {stage3_48[13]},
      {stage4_48[9]}
   );
   gpc1_1 gpc4313 (
      {stage3_48[14]},
      {stage4_48[10]}
   );
   gpc1_1 gpc4314 (
      {stage3_48[15]},
      {stage4_48[11]}
   );
   gpc1_1 gpc4315 (
      {stage3_49[6]},
      {stage4_49[5]}
   );
   gpc1_1 gpc4316 (
      {stage3_49[7]},
      {stage4_49[6]}
   );
   gpc1_1 gpc4317 (
      {stage3_49[8]},
      {stage4_49[7]}
   );
   gpc1_1 gpc4318 (
      {stage3_49[9]},
      {stage4_49[8]}
   );
   gpc1_1 gpc4319 (
      {stage3_49[10]},
      {stage4_49[9]}
   );
   gpc1_1 gpc4320 (
      {stage3_49[11]},
      {stage4_49[10]}
   );
   gpc1_1 gpc4321 (
      {stage3_49[12]},
      {stage4_49[11]}
   );
   gpc1_1 gpc4322 (
      {stage3_49[13]},
      {stage4_49[12]}
   );
   gpc1_1 gpc4323 (
      {stage3_50[31]},
      {stage4_50[6]}
   );
   gpc1_1 gpc4324 (
      {stage3_51[12]},
      {stage4_51[7]}
   );
   gpc1_1 gpc4325 (
      {stage3_51[13]},
      {stage4_51[8]}
   );
   gpc1_1 gpc4326 (
      {stage3_52[23]},
      {stage4_52[8]}
   );
   gpc1_1 gpc4327 (
      {stage3_53[7]},
      {stage4_53[6]}
   );
   gpc1_1 gpc4328 (
      {stage3_53[8]},
      {stage4_53[7]}
   );
   gpc1_1 gpc4329 (
      {stage3_53[9]},
      {stage4_53[8]}
   );
   gpc1_1 gpc4330 (
      {stage3_53[10]},
      {stage4_53[9]}
   );
   gpc1_1 gpc4331 (
      {stage3_53[11]},
      {stage4_53[10]}
   );
   gpc1_1 gpc4332 (
      {stage3_53[12]},
      {stage4_53[11]}
   );
   gpc1_1 gpc4333 (
      {stage3_53[13]},
      {stage4_53[12]}
   );
   gpc1_1 gpc4334 (
      {stage3_53[14]},
      {stage4_53[13]}
   );
   gpc1_1 gpc4335 (
      {stage3_53[15]},
      {stage4_53[14]}
   );
   gpc1_1 gpc4336 (
      {stage3_54[12]},
      {stage4_54[6]}
   );
   gpc1_1 gpc4337 (
      {stage3_54[13]},
      {stage4_54[7]}
   );
   gpc1_1 gpc4338 (
      {stage3_54[14]},
      {stage4_54[8]}
   );
   gpc1_1 gpc4339 (
      {stage3_54[15]},
      {stage4_54[9]}
   );
   gpc1_1 gpc4340 (
      {stage3_55[5]},
      {stage4_55[4]}
   );
   gpc1_1 gpc4341 (
      {stage3_55[6]},
      {stage4_55[5]}
   );
   gpc1_1 gpc4342 (
      {stage3_55[7]},
      {stage4_55[6]}
   );
   gpc1_1 gpc4343 (
      {stage3_55[8]},
      {stage4_55[7]}
   );
   gpc1_1 gpc4344 (
      {stage3_55[9]},
      {stage4_55[8]}
   );
   gpc1_1 gpc4345 (
      {stage3_55[10]},
      {stage4_55[9]}
   );
   gpc1_1 gpc4346 (
      {stage3_55[11]},
      {stage4_55[10]}
   );
   gpc1_1 gpc4347 (
      {stage3_55[12]},
      {stage4_55[11]}
   );
   gpc1_1 gpc4348 (
      {stage3_55[13]},
      {stage4_55[12]}
   );
   gpc1_1 gpc4349 (
      {stage3_55[14]},
      {stage4_55[13]}
   );
   gpc1_1 gpc4350 (
      {stage3_55[15]},
      {stage4_55[14]}
   );
   gpc1_1 gpc4351 (
      {stage3_55[16]},
      {stage4_55[15]}
   );
   gpc1_1 gpc4352 (
      {stage3_55[17]},
      {stage4_55[16]}
   );
   gpc1_1 gpc4353 (
      {stage3_56[24]},
      {stage4_56[6]}
   );
   gpc1_1 gpc4354 (
      {stage3_56[25]},
      {stage4_56[7]}
   );
   gpc1_1 gpc4355 (
      {stage3_56[26]},
      {stage4_56[8]}
   );
   gpc1_1 gpc4356 (
      {stage3_56[27]},
      {stage4_56[9]}
   );
   gpc1_1 gpc4357 (
      {stage3_56[28]},
      {stage4_56[10]}
   );
   gpc1_1 gpc4358 (
      {stage3_56[29]},
      {stage4_56[11]}
   );
   gpc1_1 gpc4359 (
      {stage3_56[30]},
      {stage4_56[12]}
   );
   gpc1_1 gpc4360 (
      {stage3_58[18]},
      {stage4_58[6]}
   );
   gpc1_1 gpc4361 (
      {stage3_58[19]},
      {stage4_58[7]}
   );
   gpc1_1 gpc4362 (
      {stage3_58[20]},
      {stage4_58[8]}
   );
   gpc1_1 gpc4363 (
      {stage3_58[21]},
      {stage4_58[9]}
   );
   gpc1_1 gpc4364 (
      {stage3_58[22]},
      {stage4_58[10]}
   );
   gpc1_1 gpc4365 (
      {stage3_58[23]},
      {stage4_58[11]}
   );
   gpc1_1 gpc4366 (
      {stage3_58[24]},
      {stage4_58[12]}
   );
   gpc1_1 gpc4367 (
      {stage3_58[25]},
      {stage4_58[13]}
   );
   gpc1_1 gpc4368 (
      {stage3_58[26]},
      {stage4_58[14]}
   );
   gpc1_1 gpc4369 (
      {stage3_58[27]},
      {stage4_58[15]}
   );
   gpc1_1 gpc4370 (
      {stage3_58[28]},
      {stage4_58[16]}
   );
   gpc1_1 gpc4371 (
      {stage3_58[29]},
      {stage4_58[17]}
   );
   gpc1_1 gpc4372 (
      {stage3_58[30]},
      {stage4_58[18]}
   );
   gpc1_1 gpc4373 (
      {stage3_58[31]},
      {stage4_58[19]}
   );
   gpc1_1 gpc4374 (
      {stage3_58[32]},
      {stage4_58[20]}
   );
   gpc1_1 gpc4375 (
      {stage3_59[18]},
      {stage4_59[7]}
   );
   gpc1_1 gpc4376 (
      {stage3_59[19]},
      {stage4_59[8]}
   );
   gpc1_1 gpc4377 (
      {stage3_59[20]},
      {stage4_59[9]}
   );
   gpc1_1 gpc4378 (
      {stage3_59[21]},
      {stage4_59[10]}
   );
   gpc1_1 gpc4379 (
      {stage3_59[22]},
      {stage4_59[11]}
   );
   gpc1_1 gpc4380 (
      {stage3_59[23]},
      {stage4_59[12]}
   );
   gpc1_1 gpc4381 (
      {stage3_59[24]},
      {stage4_59[13]}
   );
   gpc1_1 gpc4382 (
      {stage3_59[25]},
      {stage4_59[14]}
   );
   gpc1_1 gpc4383 (
      {stage3_59[26]},
      {stage4_59[15]}
   );
   gpc1_1 gpc4384 (
      {stage3_59[27]},
      {stage4_59[16]}
   );
   gpc1_1 gpc4385 (
      {stage3_60[6]},
      {stage4_60[7]}
   );
   gpc1_1 gpc4386 (
      {stage3_60[7]},
      {stage4_60[8]}
   );
   gpc1_1 gpc4387 (
      {stage3_60[8]},
      {stage4_60[9]}
   );
   gpc1_1 gpc4388 (
      {stage3_60[9]},
      {stage4_60[10]}
   );
   gpc1_1 gpc4389 (
      {stage3_60[10]},
      {stage4_60[11]}
   );
   gpc1_1 gpc4390 (
      {stage3_60[11]},
      {stage4_60[12]}
   );
   gpc1_1 gpc4391 (
      {stage3_60[12]},
      {stage4_60[13]}
   );
   gpc1_1 gpc4392 (
      {stage3_60[13]},
      {stage4_60[14]}
   );
   gpc1_1 gpc4393 (
      {stage3_60[14]},
      {stage4_60[15]}
   );
   gpc1_1 gpc4394 (
      {stage3_61[12]},
      {stage4_61[4]}
   );
   gpc1_1 gpc4395 (
      {stage3_61[13]},
      {stage4_61[5]}
   );
   gpc1_1 gpc4396 (
      {stage3_61[14]},
      {stage4_61[6]}
   );
   gpc1_1 gpc4397 (
      {stage3_61[15]},
      {stage4_61[7]}
   );
   gpc1_1 gpc4398 (
      {stage3_61[16]},
      {stage4_61[8]}
   );
   gpc1_1 gpc4399 (
      {stage3_61[17]},
      {stage4_61[9]}
   );
   gpc1_1 gpc4400 (
      {stage3_61[18]},
      {stage4_61[10]}
   );
   gpc1_1 gpc4401 (
      {stage3_61[19]},
      {stage4_61[11]}
   );
   gpc1_1 gpc4402 (
      {stage3_61[20]},
      {stage4_61[12]}
   );
   gpc1_1 gpc4403 (
      {stage3_61[21]},
      {stage4_61[13]}
   );
   gpc1_1 gpc4404 (
      {stage3_61[22]},
      {stage4_61[14]}
   );
   gpc1_1 gpc4405 (
      {stage3_61[23]},
      {stage4_61[15]}
   );
   gpc1_1 gpc4406 (
      {stage3_61[24]},
      {stage4_61[16]}
   );
   gpc1_1 gpc4407 (
      {stage3_62[18]},
      {stage4_62[5]}
   );
   gpc1_1 gpc4408 (
      {stage3_62[19]},
      {stage4_62[6]}
   );
   gpc1_1 gpc4409 (
      {stage3_62[20]},
      {stage4_62[7]}
   );
   gpc1_1 gpc4410 (
      {stage3_63[12]},
      {stage4_63[7]}
   );
   gpc1_1 gpc4411 (
      {stage3_63[13]},
      {stage4_63[8]}
   );
   gpc1_1 gpc4412 (
      {stage3_63[14]},
      {stage4_63[9]}
   );
   gpc1_1 gpc4413 (
      {stage3_63[15]},
      {stage4_63[10]}
   );
   gpc1_1 gpc4414 (
      {stage3_63[16]},
      {stage4_63[11]}
   );
   gpc1_1 gpc4415 (
      {stage3_63[17]},
      {stage4_63[12]}
   );
   gpc1_1 gpc4416 (
      {stage3_64[12]},
      {stage4_64[5]}
   );
   gpc1_1 gpc4417 (
      {stage3_64[13]},
      {stage4_64[6]}
   );
   gpc1_1 gpc4418 (
      {stage3_64[14]},
      {stage4_64[7]}
   );
   gpc1_1 gpc4419 (
      {stage3_64[15]},
      {stage4_64[8]}
   );
   gpc1_1 gpc4420 (
      {stage3_64[16]},
      {stage4_64[9]}
   );
   gpc1_1 gpc4421 (
      {stage3_64[17]},
      {stage4_64[10]}
   );
   gpc1_1 gpc4422 (
      {stage3_64[18]},
      {stage4_64[11]}
   );
   gpc1_1 gpc4423 (
      {stage3_64[19]},
      {stage4_64[12]}
   );
   gpc1_1 gpc4424 (
      {stage3_64[20]},
      {stage4_64[13]}
   );
   gpc1_1 gpc4425 (
      {stage3_64[21]},
      {stage4_64[14]}
   );
   gpc1_1 gpc4426 (
      {stage3_64[22]},
      {stage4_64[15]}
   );
   gpc1_1 gpc4427 (
      {stage3_64[23]},
      {stage4_64[16]}
   );
   gpc1_1 gpc4428 (
      {stage3_64[24]},
      {stage4_64[17]}
   );
   gpc1_1 gpc4429 (
      {stage3_64[25]},
      {stage4_64[18]}
   );
   gpc1_1 gpc4430 (
      {stage3_64[26]},
      {stage4_64[19]}
   );
   gpc1_1 gpc4431 (
      {stage3_64[27]},
      {stage4_64[20]}
   );
   gpc1_1 gpc4432 (
      {stage3_64[28]},
      {stage4_64[21]}
   );
   gpc1_1 gpc4433 (
      {stage3_65[12]},
      {stage4_65[4]}
   );
   gpc1_1 gpc4434 (
      {stage3_65[13]},
      {stage4_65[5]}
   );
   gpc1_1 gpc4435 (
      {stage3_66[0]},
      {stage4_66[4]}
   );
   gpc1_1 gpc4436 (
      {stage3_66[1]},
      {stage4_66[5]}
   );
   gpc1_1 gpc4437 (
      {stage3_66[2]},
      {stage4_66[6]}
   );
   gpc1_1 gpc4438 (
      {stage3_66[3]},
      {stage4_66[7]}
   );
   gpc1_1 gpc4439 (
      {stage3_66[4]},
      {stage4_66[8]}
   );
   gpc1_1 gpc4440 (
      {stage3_66[5]},
      {stage4_66[9]}
   );
   gpc1_1 gpc4441 (
      {stage3_66[6]},
      {stage4_66[10]}
   );
   gpc1_1 gpc4442 (
      {stage3_66[7]},
      {stage4_66[11]}
   );
   gpc1_1 gpc4443 (
      {stage3_66[8]},
      {stage4_66[12]}
   );
   gpc1_1 gpc4444 (
      {stage3_67[0]},
      {stage4_67[2]}
   );
   gpc1_1 gpc4445 (
      {stage3_67[1]},
      {stage4_67[3]}
   );
   gpc1_1 gpc4446 (
      {stage3_67[2]},
      {stage4_67[4]}
   );
   gpc1_1 gpc4447 (
      {stage3_67[3]},
      {stage4_67[5]}
   );
   gpc1_1 gpc4448 (
      {stage3_67[4]},
      {stage4_67[6]}
   );
   gpc1_1 gpc4449 (
      {stage3_68[0]},
      {stage4_68[0]}
   );
   gpc1_1 gpc4450 (
      {stage3_68[1]},
      {stage4_68[1]}
   );
   gpc1343_5 gpc4451 (
      {stage4_0[0], stage4_0[1], stage4_0[2]},
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3]},
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc4452 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[1]}
   );
   gpc606_5 gpc4453 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[1]}
   );
   gpc615_5 gpc4454 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[2]}
   );
   gpc606_5 gpc4455 (
      {stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[1],stage5_11[1],stage5_10[1],stage5_9[2]}
   );
   gpc606_5 gpc4456 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1]}
   );
   gpc615_5 gpc4457 (
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4]},
      {stage4_15[6]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[1]}
   );
   gpc615_5 gpc4458 (
      {stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage4_16[6]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[1],stage5_17[2],stage5_16[2],stage5_15[2]}
   );
   gpc606_5 gpc4459 (
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[1],stage5_18[2],stage5_17[3]}
   );
   gpc606_5 gpc4460 (
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], 1'b0},
      {stage4_19[6], stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage5_21[1],stage5_20[1],stage5_19[2],stage5_18[3],stage5_17[4]}
   );
   gpc615_5 gpc4461 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4]},
      {stage4_19[12]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[2],stage5_20[2],stage5_19[3],stage5_18[4]}
   );
   gpc606_5 gpc4462 (
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], 1'b0},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[0],stage5_22[1],stage5_21[3],stage5_20[3]}
   );
   gpc7_3 gpc4463 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5], stage4_21[6]},
      {stage5_23[1],stage5_22[2],stage5_21[4]}
   );
   gpc606_5 gpc4464 (
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[0],stage5_25[0],stage5_24[1],stage5_23[2]}
   );
   gpc1406_5 gpc4465 (
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3]},
      {stage4_27[0]},
      {stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[1],stage5_24[2]}
   );
   gpc1406_5 gpc4466 (
      {stage4_24[6], stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11]},
      {stage4_26[4], stage4_26[5], stage4_26[6], stage4_26[7]},
      {stage4_27[1]},
      {stage5_28[1],stage5_27[2],stage5_26[2],stage5_25[2],stage5_24[3]}
   );
   gpc615_5 gpc4467 (
      {stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5], stage4_27[6]},
      {stage4_28[0]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[0],stage5_29[0],stage5_28[2],stage5_27[3]}
   );
   gpc2135_5 gpc4468 (
      {stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage4_29[6], stage4_29[7], stage4_29[8]},
      {stage4_30[0]},
      {stage4_31[0], stage4_31[1]},
      {stage5_32[0],stage5_31[1],stage5_30[1],stage5_29[1],stage5_28[3]}
   );
   gpc606_5 gpc4469 (
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6]},
      {stage5_32[1],stage5_31[2],stage5_30[2],stage5_29[2],stage5_28[4]}
   );
   gpc615_5 gpc4470 (
      {stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage4_31[2]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[0],stage5_32[2],stage5_31[3],stage5_30[3]}
   );
   gpc615_5 gpc4471 (
      {stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15], 1'b0},
      {stage4_31[3]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[1],stage5_32[3],stage5_31[4],stage5_30[4]}
   );
   gpc615_5 gpc4472 (
      {stage4_31[4], stage4_31[5], stage4_31[6], stage4_31[7], stage4_31[8]},
      {stage4_32[12]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[2],stage5_33[2],stage5_32[4],stage5_31[5]}
   );
   gpc1343_5 gpc4473 (
      {stage4_33[6], stage4_33[7], stage4_33[8]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3]},
      {stage4_35[0], stage4_35[1], stage4_35[2]},
      {stage4_36[0]},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[3],stage5_33[3]}
   );
   gpc1343_5 gpc4474 (
      {stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_34[4], stage4_34[5], stage4_34[6], stage4_34[7]},
      {stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage4_36[1]},
      {stage5_37[1],stage5_36[1],stage5_35[2],stage5_34[4],stage5_33[4]}
   );
   gpc615_5 gpc4475 (
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10]},
      {stage4_36[2]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage5_39[0],stage5_38[0],stage5_37[2],stage5_36[2],stage5_35[3]}
   );
   gpc606_5 gpc4476 (
      {stage4_36[3], stage4_36[4], stage4_36[5], stage4_36[6], stage4_36[7], stage4_36[8]},
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5]},
      {stage5_40[0],stage5_39[1],stage5_38[1],stage5_37[3],stage5_36[3]}
   );
   gpc207_4 gpc4477 (
      {stage4_39[0], stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5], stage4_39[6]},
      {stage4_41[0], stage4_41[1]},
      {stage5_42[0],stage5_41[0],stage5_40[1],stage5_39[2]}
   );
   gpc606_5 gpc4478 (
      {stage4_40[0], stage4_40[1], stage4_40[2], stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[0],stage5_42[1],stage5_41[1],stage5_40[2]}
   );
   gpc606_5 gpc4479 (
      {stage4_40[6], stage4_40[7], stage4_40[8], stage4_40[9], stage4_40[10], stage4_40[11]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[1],stage5_42[2],stage5_41[2],stage5_40[3]}
   );
   gpc606_5 gpc4480 (
      {stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5], stage4_41[6], stage4_41[7]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[2],stage5_43[2],stage5_42[3],stage5_41[3]}
   );
   gpc615_5 gpc4481 (
      {stage4_42[12], stage4_42[13], stage4_42[14], stage4_42[15], stage4_42[16]},
      {stage4_43[6]},
      {stage4_44[0], stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage5_46[0],stage5_45[1],stage5_44[3],stage5_43[3],stage5_42[4]}
   );
   gpc606_5 gpc4482 (
      {stage4_44[6], stage4_44[7], stage4_44[8], stage4_44[9], stage4_44[10], stage4_44[11]},
      {stage4_46[0], stage4_46[1], stage4_46[2], stage4_46[3], stage4_46[4], stage4_46[5]},
      {stage5_48[0],stage5_47[0],stage5_46[1],stage5_45[2],stage5_44[4]}
   );
   gpc23_3 gpc4483 (
      {stage4_45[0], stage4_45[1], stage4_45[2]},
      {stage4_46[6], stage4_46[7]},
      {stage5_47[1],stage5_46[2],stage5_45[3]}
   );
   gpc606_5 gpc4484 (
      {stage4_45[3], stage4_45[4], stage4_45[5], stage4_45[6], stage4_45[7], stage4_45[8]},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4], stage4_47[5]},
      {stage5_49[0],stage5_48[1],stage5_47[2],stage5_46[3],stage5_45[4]}
   );
   gpc615_5 gpc4485 (
      {stage4_46[8], stage4_46[9], stage4_46[10], stage4_46[11], stage4_46[12]},
      {stage4_47[6]},
      {stage4_48[0], stage4_48[1], stage4_48[2], stage4_48[3], stage4_48[4], stage4_48[5]},
      {stage5_50[0],stage5_49[1],stage5_48[2],stage5_47[3],stage5_46[4]}
   );
   gpc615_5 gpc4486 (
      {stage4_46[13], stage4_46[14], stage4_46[15], stage4_46[16], stage4_46[17]},
      {stage4_47[7]},
      {stage4_48[6], stage4_48[7], stage4_48[8], stage4_48[9], stage4_48[10], stage4_48[11]},
      {stage5_50[1],stage5_49[2],stage5_48[3],stage5_47[4],stage5_46[5]}
   );
   gpc135_4 gpc4487 (
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4]},
      {stage4_50[0], stage4_50[1], stage4_50[2]},
      {stage4_51[0]},
      {stage5_52[0],stage5_51[0],stage5_50[2],stage5_49[3]}
   );
   gpc606_5 gpc4488 (
      {stage4_49[5], stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10]},
      {stage4_51[1], stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5], stage4_51[6]},
      {stage5_53[0],stage5_52[1],stage5_51[1],stage5_50[3],stage5_49[4]}
   );
   gpc615_5 gpc4489 (
      {stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6], 1'b0},
      {stage4_51[7]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[1],stage5_52[2],stage5_51[2],stage5_50[4]}
   );
   gpc606_5 gpc4490 (
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[0],stage5_55[0],stage5_54[1],stage5_53[2]}
   );
   gpc606_5 gpc4491 (
      {stage4_53[6], stage4_53[7], stage4_53[8], stage4_53[9], stage4_53[10], stage4_53[11]},
      {stage4_55[6], stage4_55[7], stage4_55[8], stage4_55[9], stage4_55[10], stage4_55[11]},
      {stage5_57[1],stage5_56[1],stage5_55[1],stage5_54[2],stage5_53[3]}
   );
   gpc615_5 gpc4492 (
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4]},
      {stage4_55[12]},
      {stage4_56[0], stage4_56[1], stage4_56[2], stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage5_58[0],stage5_57[2],stage5_56[2],stage5_55[2],stage5_54[3]}
   );
   gpc606_5 gpc4493 (
      {stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10], stage4_56[11]},
      {stage4_58[0], stage4_58[1], stage4_58[2], stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage5_60[0],stage5_59[0],stage5_58[1],stage5_57[3],stage5_56[3]}
   );
   gpc1343_5 gpc4494 (
      {stage4_57[0], stage4_57[1], stage4_57[2]},
      {stage4_58[6], stage4_58[7], stage4_58[8], stage4_58[9]},
      {stage4_59[0], stage4_59[1], stage4_59[2]},
      {stage4_60[0]},
      {stage5_61[0],stage5_60[1],stage5_59[1],stage5_58[2],stage5_57[4]}
   );
   gpc1343_5 gpc4495 (
      {stage4_57[3], stage4_57[4], stage4_57[5]},
      {stage4_58[10], stage4_58[11], stage4_58[12], stage4_58[13]},
      {stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_60[1]},
      {stage5_61[1],stage5_60[2],stage5_59[2],stage5_58[3],stage5_57[5]}
   );
   gpc606_5 gpc4496 (
      {stage4_58[14], stage4_58[15], stage4_58[16], stage4_58[17], stage4_58[18], stage4_58[19]},
      {stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5], stage4_60[6], stage4_60[7]},
      {stage5_62[0],stage5_61[2],stage5_60[3],stage5_59[3],stage5_58[4]}
   );
   gpc606_5 gpc4497 (
      {stage4_59[6], stage4_59[7], stage4_59[8], stage4_59[9], stage4_59[10], stage4_59[11]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[1],stage5_61[3],stage5_60[4],stage5_59[4]}
   );
   gpc606_5 gpc4498 (
      {stage4_59[12], stage4_59[13], stage4_59[14], stage4_59[15], stage4_59[16], 1'b0},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[2],stage5_61[4],stage5_60[5],stage5_59[5]}
   );
   gpc606_5 gpc4499 (
      {stage4_60[8], stage4_60[9], stage4_60[10], stage4_60[11], stage4_60[12], stage4_60[13]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[2],stage5_62[3],stage5_61[5],stage5_60[6]}
   );
   gpc135_4 gpc4500 (
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4]},
      {stage4_64[0], stage4_64[1], stage4_64[2]},
      {stage4_65[0]},
      {stage5_66[0],stage5_65[0],stage5_64[1],stage5_63[3]}
   );
   gpc606_5 gpc4501 (
      {stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6], stage4_64[7], stage4_64[8]},
      {stage4_66[0], stage4_66[1], stage4_66[2], stage4_66[3], stage4_66[4], stage4_66[5]},
      {stage5_68[0],stage5_67[0],stage5_66[1],stage5_65[1],stage5_64[2]}
   );
   gpc606_5 gpc4502 (
      {stage4_64[9], stage4_64[10], stage4_64[11], stage4_64[12], stage4_64[13], stage4_64[14]},
      {stage4_66[6], stage4_66[7], stage4_66[8], stage4_66[9], stage4_66[10], stage4_66[11]},
      {stage5_68[1],stage5_67[1],stage5_66[2],stage5_65[2],stage5_64[3]}
   );
   gpc606_5 gpc4503 (
      {stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5], 1'b0},
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], stage4_67[4], stage4_67[5]},
      {stage5_69[0],stage5_68[2],stage5_67[2],stage5_66[3],stage5_65[3]}
   );
   gpc1_1 gpc4504 (
      {stage4_0[3]},
      {stage5_0[1]}
   );
   gpc1_1 gpc4505 (
      {stage4_2[3]},
      {stage5_2[1]}
   );
   gpc1_1 gpc4506 (
      {stage4_2[4]},
      {stage5_2[2]}
   );
   gpc1_1 gpc4507 (
      {stage4_2[5]},
      {stage5_2[3]}
   );
   gpc1_1 gpc4508 (
      {stage4_2[6]},
      {stage5_2[4]}
   );
   gpc1_1 gpc4509 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc4510 (
      {stage4_3[2]},
      {stage5_3[2]}
   );
   gpc1_1 gpc4511 (
      {stage4_3[3]},
      {stage5_3[3]}
   );
   gpc1_1 gpc4512 (
      {stage4_3[4]},
      {stage5_3[4]}
   );
   gpc1_1 gpc4513 (
      {stage4_4[6]},
      {stage5_4[2]}
   );
   gpc1_1 gpc4514 (
      {stage4_4[7]},
      {stage5_4[3]}
   );
   gpc1_1 gpc4515 (
      {stage4_4[8]},
      {stage5_4[4]}
   );
   gpc1_1 gpc4516 (
      {stage4_5[6]},
      {stage5_5[2]}
   );
   gpc1_1 gpc4517 (
      {stage4_5[7]},
      {stage5_5[3]}
   );
   gpc1_1 gpc4518 (
      {stage4_5[8]},
      {stage5_5[4]}
   );
   gpc1_1 gpc4519 (
      {stage4_6[6]},
      {stage5_6[2]}
   );
   gpc1_1 gpc4520 (
      {stage4_6[7]},
      {stage5_6[3]}
   );
   gpc1_1 gpc4521 (
      {stage4_6[8]},
      {stage5_6[4]}
   );
   gpc1_1 gpc4522 (
      {stage4_6[9]},
      {stage5_6[5]}
   );
   gpc1_1 gpc4523 (
      {stage4_6[10]},
      {stage5_6[6]}
   );
   gpc1_1 gpc4524 (
      {stage4_6[11]},
      {stage5_6[7]}
   );
   gpc1_1 gpc4525 (
      {stage4_6[12]},
      {stage5_6[8]}
   );
   gpc1_1 gpc4526 (
      {stage4_6[13]},
      {stage5_6[9]}
   );
   gpc1_1 gpc4527 (
      {stage4_7[6]},
      {stage5_7[2]}
   );
   gpc1_1 gpc4528 (
      {stage4_7[7]},
      {stage5_7[3]}
   );
   gpc1_1 gpc4529 (
      {stage4_8[5]},
      {stage5_8[3]}
   );
   gpc1_1 gpc4530 (
      {stage4_8[6]},
      {stage5_8[4]}
   );
   gpc1_1 gpc4531 (
      {stage4_8[7]},
      {stage5_8[5]}
   );
   gpc1_1 gpc4532 (
      {stage4_8[8]},
      {stage5_8[6]}
   );
   gpc1_1 gpc4533 (
      {stage4_8[9]},
      {stage5_8[7]}
   );
   gpc1_1 gpc4534 (
      {stage4_10[6]},
      {stage5_10[2]}
   );
   gpc1_1 gpc4535 (
      {stage4_10[7]},
      {stage5_10[3]}
   );
   gpc1_1 gpc4536 (
      {stage4_10[8]},
      {stage5_10[4]}
   );
   gpc1_1 gpc4537 (
      {stage4_11[6]},
      {stage5_11[2]}
   );
   gpc1_1 gpc4538 (
      {stage4_12[0]},
      {stage5_12[2]}
   );
   gpc1_1 gpc4539 (
      {stage4_12[1]},
      {stage5_12[3]}
   );
   gpc1_1 gpc4540 (
      {stage4_12[2]},
      {stage5_12[4]}
   );
   gpc1_1 gpc4541 (
      {stage4_12[3]},
      {stage5_12[5]}
   );
   gpc1_1 gpc4542 (
      {stage4_12[4]},
      {stage5_12[6]}
   );
   gpc1_1 gpc4543 (
      {stage4_12[5]},
      {stage5_12[7]}
   );
   gpc1_1 gpc4544 (
      {stage4_12[6]},
      {stage5_12[8]}
   );
   gpc1_1 gpc4545 (
      {stage4_12[7]},
      {stage5_12[9]}
   );
   gpc1_1 gpc4546 (
      {stage4_12[8]},
      {stage5_12[10]}
   );
   gpc1_1 gpc4547 (
      {stage4_13[6]},
      {stage5_13[2]}
   );
   gpc1_1 gpc4548 (
      {stage4_13[7]},
      {stage5_13[3]}
   );
   gpc1_1 gpc4549 (
      {stage4_13[8]},
      {stage5_13[4]}
   );
   gpc1_1 gpc4550 (
      {stage4_13[9]},
      {stage5_13[5]}
   );
   gpc1_1 gpc4551 (
      {stage4_14[5]},
      {stage5_14[2]}
   );
   gpc1_1 gpc4552 (
      {stage4_14[6]},
      {stage5_14[3]}
   );
   gpc1_1 gpc4553 (
      {stage4_14[7]},
      {stage5_14[4]}
   );
   gpc1_1 gpc4554 (
      {stage4_14[8]},
      {stage5_14[5]}
   );
   gpc1_1 gpc4555 (
      {stage4_14[9]},
      {stage5_14[6]}
   );
   gpc1_1 gpc4556 (
      {stage4_14[10]},
      {stage5_14[7]}
   );
   gpc1_1 gpc4557 (
      {stage4_15[12]},
      {stage5_15[3]}
   );
   gpc1_1 gpc4558 (
      {stage4_15[13]},
      {stage5_15[4]}
   );
   gpc1_1 gpc4559 (
      {stage4_15[14]},
      {stage5_15[5]}
   );
   gpc1_1 gpc4560 (
      {stage4_15[15]},
      {stage5_15[6]}
   );
   gpc1_1 gpc4561 (
      {stage4_15[16]},
      {stage5_15[7]}
   );
   gpc1_1 gpc4562 (
      {stage4_16[7]},
      {stage5_16[3]}
   );
   gpc1_1 gpc4563 (
      {stage4_16[8]},
      {stage5_16[4]}
   );
   gpc1_1 gpc4564 (
      {stage4_16[9]},
      {stage5_16[5]}
   );
   gpc1_1 gpc4565 (
      {stage4_16[10]},
      {stage5_16[6]}
   );
   gpc1_1 gpc4566 (
      {stage4_16[11]},
      {stage5_16[7]}
   );
   gpc1_1 gpc4567 (
      {stage4_16[12]},
      {stage5_16[8]}
   );
   gpc1_1 gpc4568 (
      {stage4_18[5]},
      {stage5_18[5]}
   );
   gpc1_1 gpc4569 (
      {stage4_19[13]},
      {stage5_19[4]}
   );
   gpc1_1 gpc4570 (
      {stage4_19[14]},
      {stage5_19[5]}
   );
   gpc1_1 gpc4571 (
      {stage4_19[15]},
      {stage5_19[6]}
   );
   gpc1_1 gpc4572 (
      {stage4_21[7]},
      {stage5_21[5]}
   );
   gpc1_1 gpc4573 (
      {stage4_22[6]},
      {stage5_22[3]}
   );
   gpc1_1 gpc4574 (
      {stage4_22[7]},
      {stage5_22[4]}
   );
   gpc1_1 gpc4575 (
      {stage4_22[8]},
      {stage5_22[5]}
   );
   gpc1_1 gpc4576 (
      {stage4_22[9]},
      {stage5_22[6]}
   );
   gpc1_1 gpc4577 (
      {stage4_22[10]},
      {stage5_22[7]}
   );
   gpc1_1 gpc4578 (
      {stage4_22[11]},
      {stage5_22[8]}
   );
   gpc1_1 gpc4579 (
      {stage4_22[12]},
      {stage5_22[9]}
   );
   gpc1_1 gpc4580 (
      {stage4_22[13]},
      {stage5_22[10]}
   );
   gpc1_1 gpc4581 (
      {stage4_23[6]},
      {stage5_23[3]}
   );
   gpc1_1 gpc4582 (
      {stage4_23[7]},
      {stage5_23[4]}
   );
   gpc1_1 gpc4583 (
      {stage4_23[8]},
      {stage5_23[5]}
   );
   gpc1_1 gpc4584 (
      {stage4_23[9]},
      {stage5_23[6]}
   );
   gpc1_1 gpc4585 (
      {stage4_24[12]},
      {stage5_24[4]}
   );
   gpc1_1 gpc4586 (
      {stage4_24[13]},
      {stage5_24[5]}
   );
   gpc1_1 gpc4587 (
      {stage4_24[14]},
      {stage5_24[6]}
   );
   gpc1_1 gpc4588 (
      {stage4_24[15]},
      {stage5_24[7]}
   );
   gpc1_1 gpc4589 (
      {stage4_24[16]},
      {stage5_24[8]}
   );
   gpc1_1 gpc4590 (
      {stage4_24[17]},
      {stage5_24[9]}
   );
   gpc1_1 gpc4591 (
      {stage4_29[9]},
      {stage5_29[3]}
   );
   gpc1_1 gpc4592 (
      {stage4_32[13]},
      {stage5_32[5]}
   );
   gpc1_1 gpc4593 (
      {stage4_32[14]},
      {stage5_32[6]}
   );
   gpc1_1 gpc4594 (
      {stage4_32[15]},
      {stage5_32[7]}
   );
   gpc1_1 gpc4595 (
      {stage4_32[16]},
      {stage5_32[8]}
   );
   gpc1_1 gpc4596 (
      {stage4_32[17]},
      {stage5_32[9]}
   );
   gpc1_1 gpc4597 (
      {stage4_32[18]},
      {stage5_32[10]}
   );
   gpc1_1 gpc4598 (
      {stage4_32[19]},
      {stage5_32[11]}
   );
   gpc1_1 gpc4599 (
      {stage4_34[8]},
      {stage5_34[5]}
   );
   gpc1_1 gpc4600 (
      {stage4_34[9]},
      {stage5_34[6]}
   );
   gpc1_1 gpc4601 (
      {stage4_34[10]},
      {stage5_34[7]}
   );
   gpc1_1 gpc4602 (
      {stage4_36[9]},
      {stage5_36[4]}
   );
   gpc1_1 gpc4603 (
      {stage4_39[7]},
      {stage5_39[3]}
   );
   gpc1_1 gpc4604 (
      {stage4_39[8]},
      {stage5_39[4]}
   );
   gpc1_1 gpc4605 (
      {stage4_39[9]},
      {stage5_39[5]}
   );
   gpc1_1 gpc4606 (
      {stage4_40[12]},
      {stage5_40[4]}
   );
   gpc1_1 gpc4607 (
      {stage4_40[13]},
      {stage5_40[5]}
   );
   gpc1_1 gpc4608 (
      {stage4_41[8]},
      {stage5_41[4]}
   );
   gpc1_1 gpc4609 (
      {stage4_41[9]},
      {stage5_41[5]}
   );
   gpc1_1 gpc4610 (
      {stage4_41[10]},
      {stage5_41[6]}
   );
   gpc1_1 gpc4611 (
      {stage4_41[11]},
      {stage5_41[7]}
   );
   gpc1_1 gpc4612 (
      {stage4_41[12]},
      {stage5_41[8]}
   );
   gpc1_1 gpc4613 (
      {stage4_41[13]},
      {stage5_41[9]}
   );
   gpc1_1 gpc4614 (
      {stage4_41[14]},
      {stage5_41[10]}
   );
   gpc1_1 gpc4615 (
      {stage4_41[15]},
      {stage5_41[11]}
   );
   gpc1_1 gpc4616 (
      {stage4_41[16]},
      {stage5_41[12]}
   );
   gpc1_1 gpc4617 (
      {stage4_44[12]},
      {stage5_44[5]}
   );
   gpc1_1 gpc4618 (
      {stage4_47[8]},
      {stage5_47[5]}
   );
   gpc1_1 gpc4619 (
      {stage4_47[9]},
      {stage5_47[6]}
   );
   gpc1_1 gpc4620 (
      {stage4_47[10]},
      {stage5_47[7]}
   );
   gpc1_1 gpc4621 (
      {stage4_47[11]},
      {stage5_47[8]}
   );
   gpc1_1 gpc4622 (
      {stage4_47[12]},
      {stage5_47[9]}
   );
   gpc1_1 gpc4623 (
      {stage4_47[13]},
      {stage5_47[10]}
   );
   gpc1_1 gpc4624 (
      {stage4_47[14]},
      {stage5_47[11]}
   );
   gpc1_1 gpc4625 (
      {stage4_47[15]},
      {stage5_47[12]}
   );
   gpc1_1 gpc4626 (
      {stage4_49[11]},
      {stage5_49[5]}
   );
   gpc1_1 gpc4627 (
      {stage4_49[12]},
      {stage5_49[6]}
   );
   gpc1_1 gpc4628 (
      {stage4_51[8]},
      {stage5_51[3]}
   );
   gpc1_1 gpc4629 (
      {stage4_52[6]},
      {stage5_52[3]}
   );
   gpc1_1 gpc4630 (
      {stage4_52[7]},
      {stage5_52[4]}
   );
   gpc1_1 gpc4631 (
      {stage4_52[8]},
      {stage5_52[5]}
   );
   gpc1_1 gpc4632 (
      {stage4_53[12]},
      {stage5_53[4]}
   );
   gpc1_1 gpc4633 (
      {stage4_53[13]},
      {stage5_53[5]}
   );
   gpc1_1 gpc4634 (
      {stage4_53[14]},
      {stage5_53[6]}
   );
   gpc1_1 gpc4635 (
      {stage4_54[5]},
      {stage5_54[4]}
   );
   gpc1_1 gpc4636 (
      {stage4_54[6]},
      {stage5_54[5]}
   );
   gpc1_1 gpc4637 (
      {stage4_54[7]},
      {stage5_54[6]}
   );
   gpc1_1 gpc4638 (
      {stage4_54[8]},
      {stage5_54[7]}
   );
   gpc1_1 gpc4639 (
      {stage4_54[9]},
      {stage5_54[8]}
   );
   gpc1_1 gpc4640 (
      {stage4_55[13]},
      {stage5_55[3]}
   );
   gpc1_1 gpc4641 (
      {stage4_55[14]},
      {stage5_55[4]}
   );
   gpc1_1 gpc4642 (
      {stage4_55[15]},
      {stage5_55[5]}
   );
   gpc1_1 gpc4643 (
      {stage4_55[16]},
      {stage5_55[6]}
   );
   gpc1_1 gpc4644 (
      {stage4_56[12]},
      {stage5_56[4]}
   );
   gpc1_1 gpc4645 (
      {stage4_58[20]},
      {stage5_58[5]}
   );
   gpc1_1 gpc4646 (
      {stage4_60[14]},
      {stage5_60[7]}
   );
   gpc1_1 gpc4647 (
      {stage4_60[15]},
      {stage5_60[8]}
   );
   gpc1_1 gpc4648 (
      {stage4_61[12]},
      {stage5_61[6]}
   );
   gpc1_1 gpc4649 (
      {stage4_61[13]},
      {stage5_61[7]}
   );
   gpc1_1 gpc4650 (
      {stage4_61[14]},
      {stage5_61[8]}
   );
   gpc1_1 gpc4651 (
      {stage4_61[15]},
      {stage5_61[9]}
   );
   gpc1_1 gpc4652 (
      {stage4_61[16]},
      {stage5_61[10]}
   );
   gpc1_1 gpc4653 (
      {stage4_62[6]},
      {stage5_62[4]}
   );
   gpc1_1 gpc4654 (
      {stage4_62[7]},
      {stage5_62[5]}
   );
   gpc1_1 gpc4655 (
      {stage4_63[5]},
      {stage5_63[4]}
   );
   gpc1_1 gpc4656 (
      {stage4_63[6]},
      {stage5_63[5]}
   );
   gpc1_1 gpc4657 (
      {stage4_63[7]},
      {stage5_63[6]}
   );
   gpc1_1 gpc4658 (
      {stage4_63[8]},
      {stage5_63[7]}
   );
   gpc1_1 gpc4659 (
      {stage4_63[9]},
      {stage5_63[8]}
   );
   gpc1_1 gpc4660 (
      {stage4_63[10]},
      {stage5_63[9]}
   );
   gpc1_1 gpc4661 (
      {stage4_63[11]},
      {stage5_63[10]}
   );
   gpc1_1 gpc4662 (
      {stage4_63[12]},
      {stage5_63[11]}
   );
   gpc1_1 gpc4663 (
      {stage4_64[15]},
      {stage5_64[4]}
   );
   gpc1_1 gpc4664 (
      {stage4_64[16]},
      {stage5_64[5]}
   );
   gpc1_1 gpc4665 (
      {stage4_64[17]},
      {stage5_64[6]}
   );
   gpc1_1 gpc4666 (
      {stage4_64[18]},
      {stage5_64[7]}
   );
   gpc1_1 gpc4667 (
      {stage4_64[19]},
      {stage5_64[8]}
   );
   gpc1_1 gpc4668 (
      {stage4_64[20]},
      {stage5_64[9]}
   );
   gpc1_1 gpc4669 (
      {stage4_64[21]},
      {stage5_64[10]}
   );
   gpc1_1 gpc4670 (
      {stage4_66[12]},
      {stage5_66[4]}
   );
   gpc1_1 gpc4671 (
      {stage4_67[6]},
      {stage5_67[3]}
   );
   gpc1_1 gpc4672 (
      {stage4_68[0]},
      {stage5_68[3]}
   );
   gpc1_1 gpc4673 (
      {stage4_68[1]},
      {stage5_68[4]}
   );
   gpc615_5 gpc4674 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], 1'b0},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc1415_5 gpc4675 (
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc1415_5 gpc4676 (
      {stage5_6[5], stage5_6[6], stage5_6[7], stage5_6[8], stage5_6[9]},
      {stage5_7[1]},
      {stage5_8[4], stage5_8[5], stage5_8[6], stage5_8[7]},
      {stage5_9[1]},
      {stage6_10[1],stage6_9[1],stage6_8[1],stage6_7[2],stage6_6[2]}
   );
   gpc606_5 gpc4677 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[0]}
   );
   gpc606_5 gpc4678 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[1],stage6_13[1]}
   );
   gpc606_5 gpc4679 (
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5]},
      {stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[2]}
   );
   gpc2135_5 gpc4680 (
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4]},
      {stage5_20[0], stage5_20[1], stage5_20[2]},
      {stage5_21[0]},
      {stage5_22[0], stage5_22[1]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[1],stage6_19[1]}
   );
   gpc1163_5 gpc4681 (
      {stage5_22[2], stage5_22[3], stage5_22[4]},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5]},
      {stage5_24[0]},
      {stage5_25[0]},
      {stage6_26[0],stage6_25[0],stage6_24[0],stage6_23[1],stage6_22[1]}
   );
   gpc615_5 gpc4682 (
      {stage5_22[5], stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9]},
      {stage5_23[6]},
      {stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6]},
      {stage6_26[1],stage6_25[1],stage6_24[1],stage6_23[2],stage6_22[2]}
   );
   gpc1343_5 gpc4683 (
      {stage5_24[7], stage5_24[8], stage5_24[9]},
      {stage5_25[1], stage5_25[2], 1'b0, 1'b0},
      {stage5_26[0], stage5_26[1], stage5_26[2]},
      {stage5_27[0]},
      {stage6_28[0],stage6_27[0],stage6_26[2],stage6_25[2],stage6_24[2]}
   );
   gpc3_2 gpc4684 (
      {stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage6_28[1],stage6_27[1]}
   );
   gpc606_5 gpc4685 (
      {stage5_28[0], stage5_28[1], stage5_28[2], stage5_28[3], stage5_28[4], 1'b0},
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], 1'b0},
      {stage6_32[0],stage6_31[0],stage6_30[0],stage6_29[0],stage6_28[2]}
   );
   gpc606_5 gpc4686 (
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], 1'b0, 1'b0},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[1],stage6_31[1],stage6_30[1],stage6_29[1]}
   );
   gpc606_5 gpc4687 (
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[0],stage6_34[0],stage6_33[1],stage6_32[2]}
   );
   gpc615_5 gpc4688 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4]},
      {stage5_34[6]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], 1'b0, 1'b0},
      {stage6_37[0],stage6_36[1],stage6_35[1],stage6_34[1],stage6_33[2]}
   );
   gpc615_5 gpc4689 (
      {stage5_38[0], stage5_38[1], 1'b0, 1'b0, 1'b0},
      {stage5_39[0]},
      {stage5_40[0], stage5_40[1], stage5_40[2], stage5_40[3], stage5_40[4], stage5_40[5]},
      {stage6_42[0],stage6_41[0],stage6_40[0],stage6_39[0],stage6_38[0]}
   );
   gpc606_5 gpc4690 (
      {stage5_39[1], stage5_39[2], stage5_39[3], stage5_39[4], stage5_39[5], 1'b0},
      {stage5_41[0], stage5_41[1], stage5_41[2], stage5_41[3], stage5_41[4], stage5_41[5]},
      {stage6_43[0],stage6_42[1],stage6_41[1],stage6_40[1],stage6_39[1]}
   );
   gpc606_5 gpc4691 (
      {stage5_41[6], stage5_41[7], stage5_41[8], stage5_41[9], stage5_41[10], stage5_41[11]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3], 1'b0, 1'b0},
      {stage6_45[0],stage6_44[0],stage6_43[1],stage6_42[2],stage6_41[2]}
   );
   gpc606_5 gpc4692 (
      {stage5_44[0], stage5_44[1], stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5]},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage6_48[0],stage6_47[0],stage6_46[0],stage6_45[1],stage6_44[1]}
   );
   gpc606_5 gpc4693 (
      {stage5_45[0], stage5_45[1], stage5_45[2], stage5_45[3], stage5_45[4], 1'b0},
      {stage5_47[0], stage5_47[1], stage5_47[2], stage5_47[3], stage5_47[4], stage5_47[5]},
      {stage6_49[0],stage6_48[1],stage6_47[1],stage6_46[1],stage6_45[2]}
   );
   gpc615_5 gpc4694 (
      {stage5_47[6], stage5_47[7], stage5_47[8], stage5_47[9], stage5_47[10]},
      {stage5_48[0]},
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5]},
      {stage6_51[0],stage6_50[0],stage6_49[1],stage6_48[2],stage6_47[2]}
   );
   gpc1343_5 gpc4695 (
      {stage5_50[0], stage5_50[1], stage5_50[2]},
      {stage5_51[0], stage5_51[1], stage5_51[2], stage5_51[3]},
      {stage5_52[0], stage5_52[1], stage5_52[2]},
      {stage5_53[0]},
      {stage6_54[0],stage6_53[0],stage6_52[0],stage6_51[1],stage6_50[1]}
   );
   gpc223_4 gpc4696 (
      {stage5_53[1], stage5_53[2], stage5_53[3]},
      {stage5_54[0], stage5_54[1]},
      {stage5_55[0], stage5_55[1]},
      {stage6_56[0],stage6_55[0],stage6_54[1],stage6_53[1]}
   );
   gpc207_4 gpc4697 (
      {stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5], stage5_54[6], stage5_54[7], stage5_54[8]},
      {stage5_56[0], stage5_56[1]},
      {stage6_57[0],stage6_56[1],stage6_55[1],stage6_54[2]}
   );
   gpc615_5 gpc4698 (
      {stage5_55[2], stage5_55[3], stage5_55[4], stage5_55[5], stage5_55[6]},
      {stage5_56[2]},
      {stage5_57[0], stage5_57[1], stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5]},
      {stage6_59[0],stage6_58[0],stage6_57[1],stage6_56[2],stage6_55[2]}
   );
   gpc606_5 gpc4699 (
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4], stage5_58[5]},
      {stage5_60[0], stage5_60[1], stage5_60[2], stage5_60[3], stage5_60[4], stage5_60[5]},
      {stage6_62[0],stage6_61[0],stage6_60[0],stage6_59[1],stage6_58[1]}
   );
   gpc606_5 gpc4700 (
      {stage5_59[0], stage5_59[1], stage5_59[2], stage5_59[3], stage5_59[4], stage5_59[5]},
      {stage5_61[0], stage5_61[1], stage5_61[2], stage5_61[3], stage5_61[4], stage5_61[5]},
      {stage6_63[0],stage6_62[1],stage6_61[1],stage6_60[1],stage6_59[2]}
   );
   gpc606_5 gpc4701 (
      {stage5_61[6], stage5_61[7], stage5_61[8], stage5_61[9], stage5_61[10], 1'b0},
      {stage5_63[0], stage5_63[1], stage5_63[2], stage5_63[3], stage5_63[4], stage5_63[5]},
      {stage6_65[0],stage6_64[0],stage6_63[1],stage6_62[2],stage6_61[2]}
   );
   gpc606_5 gpc4702 (
      {stage5_62[0], stage5_62[1], stage5_62[2], stage5_62[3], stage5_62[4], stage5_62[5]},
      {stage5_64[0], stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage6_66[0],stage6_65[1],stage6_64[1],stage6_63[2],stage6_62[3]}
   );
   gpc606_5 gpc4703 (
      {stage5_63[6], stage5_63[7], stage5_63[8], stage5_63[9], stage5_63[10], stage5_63[11]},
      {stage5_65[0], stage5_65[1], stage5_65[2], stage5_65[3], 1'b0, 1'b0},
      {stage6_67[0],stage6_66[1],stage6_65[2],stage6_64[2],stage6_63[3]}
   );
   gpc606_5 gpc4704 (
      {stage5_64[6], stage5_64[7], stage5_64[8], stage5_64[9], stage5_64[10], 1'b0},
      {stage5_66[0], stage5_66[1], stage5_66[2], stage5_66[3], stage5_66[4], 1'b0},
      {stage6_68[0],stage6_67[1],stage6_66[2],stage6_65[3],stage6_64[3]}
   );
   gpc1_1 gpc4705 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc4706 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc4707 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc4708 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc4709 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc4710 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc4711 (
      {stage5_2[3]},
      {stage6_2[3]}
   );
   gpc1_1 gpc4712 (
      {stage5_2[4]},
      {stage6_2[4]}
   );
   gpc1_1 gpc4713 (
      {stage5_4[1]},
      {stage6_4[1]}
   );
   gpc1_1 gpc4714 (
      {stage5_4[2]},
      {stage6_4[2]}
   );
   gpc1_1 gpc4715 (
      {stage5_4[3]},
      {stage6_4[3]}
   );
   gpc1_1 gpc4716 (
      {stage5_4[4]},
      {stage6_4[4]}
   );
   gpc1_1 gpc4717 (
      {stage5_7[2]},
      {stage6_7[3]}
   );
   gpc1_1 gpc4718 (
      {stage5_7[3]},
      {stage6_7[4]}
   );
   gpc1_1 gpc4719 (
      {stage5_9[2]},
      {stage6_9[2]}
   );
   gpc1_1 gpc4720 (
      {stage5_10[0]},
      {stage6_10[2]}
   );
   gpc1_1 gpc4721 (
      {stage5_10[1]},
      {stage6_10[3]}
   );
   gpc1_1 gpc4722 (
      {stage5_10[2]},
      {stage6_10[4]}
   );
   gpc1_1 gpc4723 (
      {stage5_10[3]},
      {stage6_10[5]}
   );
   gpc1_1 gpc4724 (
      {stage5_10[4]},
      {stage6_10[6]}
   );
   gpc1_1 gpc4725 (
      {stage5_11[0]},
      {stage6_11[0]}
   );
   gpc1_1 gpc4726 (
      {stage5_11[1]},
      {stage6_11[1]}
   );
   gpc1_1 gpc4727 (
      {stage5_11[2]},
      {stage6_11[2]}
   );
   gpc1_1 gpc4728 (
      {stage5_12[6]},
      {stage6_12[1]}
   );
   gpc1_1 gpc4729 (
      {stage5_12[7]},
      {stage6_12[2]}
   );
   gpc1_1 gpc4730 (
      {stage5_12[8]},
      {stage6_12[3]}
   );
   gpc1_1 gpc4731 (
      {stage5_12[9]},
      {stage6_12[4]}
   );
   gpc1_1 gpc4732 (
      {stage5_12[10]},
      {stage6_12[5]}
   );
   gpc1_1 gpc4733 (
      {stage5_14[6]},
      {stage6_14[2]}
   );
   gpc1_1 gpc4734 (
      {stage5_14[7]},
      {stage6_14[3]}
   );
   gpc1_1 gpc4735 (
      {stage5_15[6]},
      {stage6_15[2]}
   );
   gpc1_1 gpc4736 (
      {stage5_15[7]},
      {stage6_15[3]}
   );
   gpc1_1 gpc4737 (
      {stage5_16[6]},
      {stage6_16[3]}
   );
   gpc1_1 gpc4738 (
      {stage5_16[7]},
      {stage6_16[4]}
   );
   gpc1_1 gpc4739 (
      {stage5_16[8]},
      {stage6_16[5]}
   );
   gpc1_1 gpc4740 (
      {stage5_17[0]},
      {stage6_17[2]}
   );
   gpc1_1 gpc4741 (
      {stage5_17[1]},
      {stage6_17[3]}
   );
   gpc1_1 gpc4742 (
      {stage5_17[2]},
      {stage6_17[4]}
   );
   gpc1_1 gpc4743 (
      {stage5_17[3]},
      {stage6_17[5]}
   );
   gpc1_1 gpc4744 (
      {stage5_17[4]},
      {stage6_17[6]}
   );
   gpc1_1 gpc4745 (
      {stage5_19[5]},
      {stage6_19[2]}
   );
   gpc1_1 gpc4746 (
      {stage5_19[6]},
      {stage6_19[3]}
   );
   gpc1_1 gpc4747 (
      {stage5_20[3]},
      {stage6_20[2]}
   );
   gpc1_1 gpc4748 (
      {stage5_21[1]},
      {stage6_21[1]}
   );
   gpc1_1 gpc4749 (
      {stage5_21[2]},
      {stage6_21[2]}
   );
   gpc1_1 gpc4750 (
      {stage5_21[3]},
      {stage6_21[3]}
   );
   gpc1_1 gpc4751 (
      {stage5_21[4]},
      {stage6_21[4]}
   );
   gpc1_1 gpc4752 (
      {stage5_21[5]},
      {stage6_21[5]}
   );
   gpc1_1 gpc4753 (
      {stage5_22[10]},
      {stage6_22[3]}
   );
   gpc1_1 gpc4754 (
      {stage5_32[6]},
      {stage6_32[3]}
   );
   gpc1_1 gpc4755 (
      {stage5_32[7]},
      {stage6_32[4]}
   );
   gpc1_1 gpc4756 (
      {stage5_32[8]},
      {stage6_32[5]}
   );
   gpc1_1 gpc4757 (
      {stage5_32[9]},
      {stage6_32[6]}
   );
   gpc1_1 gpc4758 (
      {stage5_32[10]},
      {stage6_32[7]}
   );
   gpc1_1 gpc4759 (
      {stage5_32[11]},
      {stage6_32[8]}
   );
   gpc1_1 gpc4760 (
      {stage5_34[7]},
      {stage6_34[2]}
   );
   gpc1_1 gpc4761 (
      {stage5_36[0]},
      {stage6_36[2]}
   );
   gpc1_1 gpc4762 (
      {stage5_36[1]},
      {stage6_36[3]}
   );
   gpc1_1 gpc4763 (
      {stage5_36[2]},
      {stage6_36[4]}
   );
   gpc1_1 gpc4764 (
      {stage5_36[3]},
      {stage6_36[5]}
   );
   gpc1_1 gpc4765 (
      {stage5_36[4]},
      {stage6_36[6]}
   );
   gpc1_1 gpc4766 (
      {stage5_37[0]},
      {stage6_37[1]}
   );
   gpc1_1 gpc4767 (
      {stage5_37[1]},
      {stage6_37[2]}
   );
   gpc1_1 gpc4768 (
      {stage5_37[2]},
      {stage6_37[3]}
   );
   gpc1_1 gpc4769 (
      {stage5_37[3]},
      {stage6_37[4]}
   );
   gpc1_1 gpc4770 (
      {stage5_41[12]},
      {stage6_41[3]}
   );
   gpc1_1 gpc4771 (
      {stage5_42[0]},
      {stage6_42[3]}
   );
   gpc1_1 gpc4772 (
      {stage5_42[1]},
      {stage6_42[4]}
   );
   gpc1_1 gpc4773 (
      {stage5_42[2]},
      {stage6_42[5]}
   );
   gpc1_1 gpc4774 (
      {stage5_42[3]},
      {stage6_42[6]}
   );
   gpc1_1 gpc4775 (
      {stage5_42[4]},
      {stage6_42[7]}
   );
   gpc1_1 gpc4776 (
      {stage5_47[11]},
      {stage6_47[3]}
   );
   gpc1_1 gpc4777 (
      {stage5_47[12]},
      {stage6_47[4]}
   );
   gpc1_1 gpc4778 (
      {stage5_48[1]},
      {stage6_48[3]}
   );
   gpc1_1 gpc4779 (
      {stage5_48[2]},
      {stage6_48[4]}
   );
   gpc1_1 gpc4780 (
      {stage5_48[3]},
      {stage6_48[5]}
   );
   gpc1_1 gpc4781 (
      {stage5_49[6]},
      {stage6_49[2]}
   );
   gpc1_1 gpc4782 (
      {stage5_50[3]},
      {stage6_50[2]}
   );
   gpc1_1 gpc4783 (
      {stage5_50[4]},
      {stage6_50[3]}
   );
   gpc1_1 gpc4784 (
      {stage5_52[3]},
      {stage6_52[1]}
   );
   gpc1_1 gpc4785 (
      {stage5_52[4]},
      {stage6_52[2]}
   );
   gpc1_1 gpc4786 (
      {stage5_52[5]},
      {stage6_52[3]}
   );
   gpc1_1 gpc4787 (
      {stage5_53[4]},
      {stage6_53[2]}
   );
   gpc1_1 gpc4788 (
      {stage5_53[5]},
      {stage6_53[3]}
   );
   gpc1_1 gpc4789 (
      {stage5_53[6]},
      {stage6_53[4]}
   );
   gpc1_1 gpc4790 (
      {stage5_56[3]},
      {stage6_56[3]}
   );
   gpc1_1 gpc4791 (
      {stage5_56[4]},
      {stage6_56[4]}
   );
   gpc1_1 gpc4792 (
      {stage5_60[6]},
      {stage6_60[2]}
   );
   gpc1_1 gpc4793 (
      {stage5_60[7]},
      {stage6_60[3]}
   );
   gpc1_1 gpc4794 (
      {stage5_60[8]},
      {stage6_60[4]}
   );
   gpc1_1 gpc4795 (
      {stage5_67[0]},
      {stage6_67[2]}
   );
   gpc1_1 gpc4796 (
      {stage5_67[1]},
      {stage6_67[3]}
   );
   gpc1_1 gpc4797 (
      {stage5_67[2]},
      {stage6_67[4]}
   );
   gpc1_1 gpc4798 (
      {stage5_67[3]},
      {stage6_67[5]}
   );
   gpc1_1 gpc4799 (
      {stage5_68[0]},
      {stage6_68[1]}
   );
   gpc1_1 gpc4800 (
      {stage5_68[1]},
      {stage6_68[2]}
   );
   gpc1_1 gpc4801 (
      {stage5_68[2]},
      {stage6_68[3]}
   );
   gpc1_1 gpc4802 (
      {stage5_68[3]},
      {stage6_68[4]}
   );
   gpc1_1 gpc4803 (
      {stage5_68[4]},
      {stage6_68[5]}
   );
   gpc1_1 gpc4804 (
      {stage5_69[0]},
      {stage6_69[0]}
   );
   gpc1415_5 gpc4805 (
      {stage6_2[0], stage6_2[1], stage6_2[2], stage6_2[3], stage6_2[4]},
      {stage6_3[0]},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3]},
      {stage6_5[0]},
      {stage7_6[0],stage7_5[0],stage7_4[0],stage7_3[0],stage7_2[0]}
   );
   gpc23_3 gpc4806 (
      {stage6_6[0], stage6_6[1], stage6_6[2]},
      {stage6_7[0], stage6_7[1]},
      {stage7_8[0],stage7_7[0],stage7_6[1]}
   );
   gpc223_4 gpc4807 (
      {stage6_7[2], stage6_7[3], stage6_7[4]},
      {stage6_8[0], stage6_8[1]},
      {stage6_9[0], stage6_9[1]},
      {stage7_10[0],stage7_9[0],stage7_8[1],stage7_7[1]}
   );
   gpc207_4 gpc4808 (
      {stage6_10[0], stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4], stage6_10[5], stage6_10[6]},
      {stage6_12[0], stage6_12[1]},
      {stage7_13[0],stage7_12[0],stage7_11[0],stage7_10[1]}
   );
   gpc1343_5 gpc4809 (
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage6_13[0], stage6_13[1], 1'b0},
      {stage6_14[0]},
      {stage7_15[0],stage7_14[0],stage7_13[1],stage7_12[1],stage7_11[1]}
   );
   gpc1343_5 gpc4810 (
      {stage6_14[1], stage6_14[2], stage6_14[3]},
      {stage6_15[0], stage6_15[1], stage6_15[2], stage6_15[3]},
      {stage6_16[0], stage6_16[1], stage6_16[2]},
      {stage6_17[0]},
      {stage7_18[0],stage7_17[0],stage7_16[0],stage7_15[1],stage7_14[1]}
   );
   gpc1163_5 gpc4811 (
      {stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4], stage6_17[5], stage6_17[6]},
      {stage6_18[0]},
      {stage6_19[0]},
      {stage7_20[0],stage7_19[0],stage7_18[1],stage7_17[1],stage7_16[1]}
   );
   gpc1343_5 gpc4812 (
      {stage6_19[1], stage6_19[2], stage6_19[3]},
      {stage6_20[0], stage6_20[1], stage6_20[2], 1'b0},
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0]},
      {stage7_23[0],stage7_22[0],stage7_21[0],stage7_20[1],stage7_19[1]}
   );
   gpc1343_5 gpc4813 (
      {stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage6_22[1], stage6_22[2], stage6_22[3], 1'b0},
      {stage6_23[0], stage6_23[1], stage6_23[2]},
      {stage6_24[0]},
      {stage7_25[0],stage7_24[0],stage7_23[1],stage7_22[1],stage7_21[1]}
   );
   gpc1343_5 gpc4814 (
      {stage6_24[1], stage6_24[2], 1'b0},
      {stage6_25[0], stage6_25[1], stage6_25[2], 1'b0},
      {stage6_26[0], stage6_26[1], stage6_26[2]},
      {stage6_27[0]},
      {stage7_28[0],stage7_27[0],stage7_26[0],stage7_25[1],stage7_24[1]}
   );
   gpc15_3 gpc4815 (
      {stage6_28[0], stage6_28[1], stage6_28[2], 1'b0, 1'b0},
      {stage6_29[0]},
      {stage7_30[0],stage7_29[0],stage7_28[1]}
   );
   gpc615_5 gpc4816 (
      {stage6_30[0], stage6_30[1], 1'b0, 1'b0, 1'b0},
      {stage6_31[0]},
      {stage6_32[0], stage6_32[1], stage6_32[2], stage6_32[3], stage6_32[4], stage6_32[5]},
      {stage7_34[0],stage7_33[0],stage7_32[0],stage7_31[0],stage7_30[1]}
   );
   gpc1343_5 gpc4817 (
      {stage6_32[6], stage6_32[7], stage6_32[8]},
      {stage6_33[0], stage6_33[1], stage6_33[2], 1'b0},
      {stage6_34[0], stage6_34[1], stage6_34[2]},
      {stage6_35[0]},
      {stage7_36[0],stage7_35[0],stage7_34[1],stage7_33[1],stage7_32[1]}
   );
   gpc7_3 gpc4818 (
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5], stage6_36[6]},
      {stage7_38[0],stage7_37[0],stage7_36[1]}
   );
   gpc2135_5 gpc4819 (
      {stage6_37[0], stage6_37[1], stage6_37[2], stage6_37[3], stage6_37[4]},
      {stage6_38[0], 1'b0, 1'b0},
      {stage6_39[0]},
      {stage6_40[0], stage6_40[1]},
      {stage7_41[0],stage7_40[0],stage7_39[0],stage7_38[1],stage7_37[1]}
   );
   gpc135_4 gpc4820 (
      {stage6_41[0], stage6_41[1], stage6_41[2], stage6_41[3], 1'b0},
      {stage6_42[0], stage6_42[1], stage6_42[2]},
      {stage6_43[0]},
      {stage7_44[0],stage7_43[0],stage7_42[0],stage7_41[1]}
   );
   gpc615_5 gpc4821 (
      {stage6_42[3], stage6_42[4], stage6_42[5], stage6_42[6], stage6_42[7]},
      {stage6_43[1]},
      {stage6_44[0], stage6_44[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_46[0],stage7_45[0],stage7_44[1],stage7_43[1],stage7_42[1]}
   );
   gpc2223_5 gpc4822 (
      {stage6_45[0], stage6_45[1], stage6_45[2]},
      {stage6_46[0], stage6_46[1]},
      {stage6_47[0], stage6_47[1]},
      {stage6_48[0], stage6_48[1]},
      {stage7_49[0],stage7_48[0],stage7_47[0],stage7_46[1],stage7_45[1]}
   );
   gpc1343_5 gpc4823 (
      {stage6_47[2], stage6_47[3], stage6_47[4]},
      {stage6_48[2], stage6_48[3], stage6_48[4], stage6_48[5]},
      {stage6_49[0], stage6_49[1], stage6_49[2]},
      {stage6_50[0]},
      {stage7_51[0],stage7_50[0],stage7_49[1],stage7_48[1],stage7_47[1]}
   );
   gpc1343_5 gpc4824 (
      {stage6_50[1], stage6_50[2], stage6_50[3]},
      {stage6_51[0], stage6_51[1], 1'b0, 1'b0},
      {stage6_52[0], stage6_52[1], stage6_52[2]},
      {stage6_53[0]},
      {stage7_54[0],stage7_53[0],stage7_52[0],stage7_51[1],stage7_50[1]}
   );
   gpc1343_5 gpc4825 (
      {stage6_52[3], 1'b0, 1'b0},
      {stage6_53[1], stage6_53[2], stage6_53[3], stage6_53[4]},
      {stage6_54[0], stage6_54[1], stage6_54[2]},
      {stage6_55[0]},
      {stage7_56[0],stage7_55[0],stage7_54[1],stage7_53[1],stage7_52[1]}
   );
   gpc1163_5 gpc4826 (
      {stage6_55[1], stage6_55[2], 1'b0},
      {stage6_56[0], stage6_56[1], stage6_56[2], stage6_56[3], stage6_56[4], 1'b0},
      {stage6_57[0]},
      {stage6_58[0]},
      {stage7_59[0],stage7_58[0],stage7_57[0],stage7_56[1],stage7_55[1]}
   );
   gpc1343_5 gpc4827 (
      {stage6_59[0], stage6_59[1], stage6_59[2]},
      {stage6_60[0], stage6_60[1], stage6_60[2], stage6_60[3]},
      {stage6_61[0], stage6_61[1], stage6_61[2]},
      {stage6_62[0]},
      {stage7_63[0],stage7_62[0],stage7_61[0],stage7_60[0],stage7_59[1]}
   );
   gpc1343_5 gpc4828 (
      {stage6_62[1], stage6_62[2], stage6_62[3]},
      {stage6_63[0], stage6_63[1], stage6_63[2], stage6_63[3]},
      {stage6_64[0], stage6_64[1], stage6_64[2]},
      {stage6_65[0]},
      {stage7_66[0],stage7_65[0],stage7_64[0],stage7_63[1],stage7_62[1]}
   );
   gpc1343_5 gpc4829 (
      {stage6_65[1], stage6_65[2], stage6_65[3]},
      {stage6_66[0], stage6_66[1], stage6_66[2], 1'b0},
      {stage6_67[0], stage6_67[1], stage6_67[2]},
      {stage6_68[0]},
      {stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[1],stage7_65[1]}
   );
   gpc1163_5 gpc4830 (
      {stage6_67[3], stage6_67[4], stage6_67[5]},
      {stage6_68[1], stage6_68[2], stage6_68[3], stage6_68[4], stage6_68[5], 1'b0},
      {stage6_69[0]},
      {1'b0},
      {stage7_71[0],stage7_70[0],stage7_69[1],stage7_68[1],stage7_67[1]}
   );
   gpc1_1 gpc4831 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc4832 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc4833 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc4834 (
      {stage6_4[4]},
      {stage7_4[1]}
   );
   gpc1_1 gpc4835 (
      {stage6_9[2]},
      {stage7_9[1]}
   );
   gpc1_1 gpc4836 (
      {stage6_27[1]},
      {stage7_27[1]}
   );
   gpc1_1 gpc4837 (
      {stage6_29[1]},
      {stage7_29[1]}
   );
   gpc1_1 gpc4838 (
      {stage6_31[1]},
      {stage7_31[1]}
   );
   gpc1_1 gpc4839 (
      {stage6_35[1]},
      {stage7_35[1]}
   );
   gpc1_1 gpc4840 (
      {stage6_39[1]},
      {stage7_39[1]}
   );
   gpc1_1 gpc4841 (
      {stage6_57[1]},
      {stage7_57[1]}
   );
   gpc1_1 gpc4842 (
      {stage6_58[1]},
      {stage7_58[1]}
   );
   gpc1_1 gpc4843 (
      {stage6_60[4]},
      {stage7_60[1]}
   );
   gpc1_1 gpc4844 (
      {stage6_64[3]},
      {stage7_64[1]}
   );
endmodule
module rowadder2_1_72(input [71:0] src0, input [71:0] src1, output [72:0] dst0);
    wire [71:0] gene;
    wire [71:0] prop;
    wire [71:0] out;
    wire [71:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_38_gene (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(gene[38])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_38_prop (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(prop[38])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_39_gene (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(gene[39])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_39_prop (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(prop[39])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_40_gene (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(gene[40])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_40_prop (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(prop[40])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_41_gene (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(gene[41])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_41_prop (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(prop[41])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_42_gene (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(gene[42])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_42_prop (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(prop[42])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_43_gene (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(gene[43])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_43_prop (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(prop[43])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_44_gene (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(gene[44])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_44_prop (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(prop[44])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_45_gene (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(gene[45])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_45_prop (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(prop[45])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_46_gene (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(gene[46])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_46_prop (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(prop[46])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_47_gene (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(gene[47])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_47_prop (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(prop[47])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_48_gene (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(gene[48])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_48_prop (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(prop[48])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_49_gene (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(gene[49])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_49_prop (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(prop[49])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_50_gene (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(gene[50])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_50_prop (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(prop[50])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_51_gene (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(gene[51])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_51_prop (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(prop[51])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_52_gene (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(gene[52])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_52_prop (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(prop[52])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_53_gene (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(gene[53])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_53_prop (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(prop[53])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_54_gene (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(gene[54])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_54_prop (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(prop[54])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_55_gene (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(gene[55])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_55_prop (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(prop[55])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_56_gene (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(gene[56])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_56_prop (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(prop[56])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_57_gene (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(gene[57])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_57_prop (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(prop[57])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_58_gene (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(gene[58])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_58_prop (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(prop[58])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_59_gene (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(gene[59])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_59_prop (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(prop[59])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_60_gene (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(gene[60])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_60_prop (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(prop[60])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_61_gene (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(gene[61])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_61_prop (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(prop[61])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_62_gene (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(gene[62])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_62_prop (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(prop[62])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_63_gene (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(gene[63])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_63_prop (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(prop[63])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_64_gene (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(gene[64])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_64_prop (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(prop[64])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_65_gene (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(gene[65])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_65_prop (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(prop[65])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_66_gene (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(gene[66])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_66_prop (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(prop[66])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_67_gene (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(gene[67])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_67_prop (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(prop[67])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_68_gene (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(gene[68])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_68_prop (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(prop[68])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_69_gene (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(gene[69])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_69_prop (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(prop[69])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_70_gene (
        .I0(src0[70]),
        .I1(src1[70]),
        .O(gene[70])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_70_prop (
        .I0(src0[70]),
        .I1(src1[70]),
        .O(prop[70])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_71_gene (
        .I0(src0[71]),
        .I1(src1[71]),
        .O(gene[71])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_71_prop (
        .I0(src0[71]),
        .I1(src1[71]),
        .O(prop[71])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI(gene[39:36]),
        .S(prop[39:36])
    );
    CARRY4 carry4_43_40 (
        .CO(carryout[43:40]),
        .O(out[43:40]),
        .CI(carryout[39]),
        .CYINIT(1'h0),
        .DI(gene[43:40]),
        .S(prop[43:40])
    );
    CARRY4 carry4_47_44 (
        .CO(carryout[47:44]),
        .O(out[47:44]),
        .CI(carryout[43]),
        .CYINIT(1'h0),
        .DI(gene[47:44]),
        .S(prop[47:44])
    );
    CARRY4 carry4_51_48 (
        .CO(carryout[51:48]),
        .O(out[51:48]),
        .CI(carryout[47]),
        .CYINIT(1'h0),
        .DI(gene[51:48]),
        .S(prop[51:48])
    );
    CARRY4 carry4_55_52 (
        .CO(carryout[55:52]),
        .O(out[55:52]),
        .CI(carryout[51]),
        .CYINIT(1'h0),
        .DI(gene[55:52]),
        .S(prop[55:52])
    );
    CARRY4 carry4_59_56 (
        .CO(carryout[59:56]),
        .O(out[59:56]),
        .CI(carryout[55]),
        .CYINIT(1'h0),
        .DI(gene[59:56]),
        .S(prop[59:56])
    );
    CARRY4 carry4_63_60 (
        .CO(carryout[63:60]),
        .O(out[63:60]),
        .CI(carryout[59]),
        .CYINIT(1'h0),
        .DI(gene[63:60]),
        .S(prop[63:60])
    );
    CARRY4 carry4_67_64 (
        .CO(carryout[67:64]),
        .O(out[67:64]),
        .CI(carryout[63]),
        .CYINIT(1'h0),
        .DI(gene[67:64]),
        .S(prop[67:64])
    );
    CARRY4 carry4_71_68 (
        .CO(carryout[71:68]),
        .O(out[71:68]),
        .CI(carryout[67]),
        .CYINIT(1'h0),
        .DI(gene[71:68]),
        .S(prop[71:68])
    );
    assign dst0 = {carryout[71], out[71:0]};
endmodule


module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    reg [161:0] src32;
    reg [161:0] src33;
    reg [161:0] src34;
    reg [161:0] src35;
    reg [161:0] src36;
    reg [161:0] src37;
    reg [161:0] src38;
    reg [161:0] src39;
    reg [161:0] src40;
    reg [161:0] src41;
    reg [161:0] src42;
    reg [161:0] src43;
    reg [161:0] src44;
    reg [161:0] src45;
    reg [161:0] src46;
    reg [161:0] src47;
    reg [161:0] src48;
    reg [161:0] src49;
    reg [161:0] src50;
    reg [161:0] src51;
    reg [161:0] src52;
    reg [161:0] src53;
    reg [161:0] src54;
    reg [161:0] src55;
    reg [161:0] src56;
    reg [161:0] src57;
    reg [161:0] src58;
    reg [161:0] src59;
    reg [161:0] src60;
    reg [161:0] src61;
    reg [161:0] src62;
    reg [161:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [71:0] srcsum;
    wire [71:0] dstsum;
    wire test;
    compressor2_1_162_64 compressor2_1_162_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc3f92e693f022592c92abb8a7d3a0cafb8110e1ba05c99c3b47bdf923831cd30caefa7c16840733463f7a4d4c9a5e37943f719b7b0d0590e2265953a2196b7fd280f55adb407f06287baacfb054aca61fc9d289371d5c1f7688de7714ab7a0d18fe0030f2dfdd8b0fb79c33a902f64f0d8df121e8cd71179f9e6d335f2e3b705d630f72fb4b48d8d056d5fc812e313b6242ab362a860c3ca6bc8270349cb8d0ff6c52f212fe97dcc21e45c9c6964300ee4cbddfaaf8f864a60742707f9cd8b68b3edfb17227f34155c9c9da152d587406ace60257a34af3344c86534ffe17df290f6f2d327afa8b790db59ba635755a43f1274f49943a937e14f300dc22eedb0c1edb232fd3a8633b6f8eb6a4c2c5c65e80650e8510b54dc4b4bdb2e6a3175a5ca75859e4b1e3842a5d8d14e7958735d6f57c7d772a491079aade018ca288b83e166c637e3f331fc5e32e81d04dc9ebc2cb78d8cc44c097d0a0e7129d830e9849500f4bc8924bad48f3509647eedc1c9066fcd781d6478079d70ad089fd8965fc5e4af5fa975482d9ba1b2337e810654300ac32dac2eb0e080e3e1e3566ca1c6f98bcbceb635c6c532f0e99fd9dabbd7fda3292127ed8034cf8cf005b8aa3b5d47208e0b0add6793cfe4a94d01def901875f18832edb693e221fa74de5156c9883d6c33a510b8e897046d344b6a44e034849aec2f8d8e98fc00ac277a294abf91bc658adde6abc53168568a4d176aec59496e3935b5d982441c2756efc78ff879e3741ff0488d0a58030467d14f246b867cfe4c929e9b393c7ede22fe5aa0b765e47ba045edc20bc76c3a42c20ab830ec8b1ebb158719f9829ad24ed42c4aad4547541841cf68037a373e7f27171eb8d04fb000998391d45d8b6e2741a17cdb42f39bff0ba75c25ff1094633be5c693b2e71edb73d26be05b3577f1582299df899e7af850af50ff4379f523123659ac8169e7e25c46e71945debf20f6c213138cfb38268d6f564f8a36850dad2f3e874c36db4b187f9cd707e92076894935ee2f3bd8a0c9999a2de322c06636072a73164d249549655f4fd072416e9881b64b7a19049d55916df2e0c0890251a1cf78f8c2203627b3d717e460f6101f06bfd79be1e5baf40321b386a82ce2301670bc4796579e36745a50429ea7f3e9c44522b51f9d6d63b9ce9e55c80a388c5ae88edcea39e1f8a34acccefbcf89b52b2ae1948a18968d788c762dece7083e8e6075f313f1401983d567f7373fd82d1b6d2d35b32218a45829fd77c44343c32cb069dce9f7f28227ab2044c94b0c8a1d9fefeeb209186a38e0ba4265d72b78ca1afeb7dc4aa555098c896774bae99ea70617a456f3a82a06b6d57a4c2a2b2c05421f186f3bb0449b4e88ec71b9cdfb7409c1eaed72db52d733ddf6ecf5ed7039252d74303c0c2fd89250e62db50032e6145c4aff811aaa5d3b9d2354562dffa61c754628f8980e5396251ac7eb5e5646c82b9f41dc833282e63403eeb5fa31d3ce90ef5ba032ff9125325915e6128027c307ef795737b5a02bdd87525d0e4cc21aa6f306db909637b642ca4a51d508dcd34a25a93d8538d4bb1a3f620bafebb6108c9a608ef0080573df47d55d8caa7c2f8b91e1942d0869ace37fe58a6608e908b98f40560b98c942fbef4a3b0fed131fe6b4a7c97cbd84291db2b1bd1bb890d26885c4868e48fb0b8e56799d624eb685582cfa0ecef8c2fc54eab1fc1e1286ca62f55935dbe3f05f0255e2189420dcf385f4373e5a7db83859a80a73071ec6d8e0e01bdf81b5ab88d3f69c0a3eb7dc51810044648a045c0cf4e93c83e26849d893d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h72e8bed8a58426ad0b882f71dd8faa8b758a28d376034bd4c0bb25ec6a36bcc8560f05a15fac0db4fbbf811d91c245279c60df5178e229a2322b497880adc277106661553ee8c945d636925fd981ca0026f61a495be67bacb98651b8826281e4dcaf7bf96f923d39e20d861775e36530da56dcb89fde5546f4be5c3cac43c2cf29f9adfb7a738993f4cef58a06ed3a6bb6fddd727844d68bca975bc123ca11ceb4a3c2c10f5f815b4370f6746c2469eea619e54d8c835f387451518ea8c8079c98c69166f39d7d122d2ecf4e0945d15492c417f040bdeb8370b398bc154d71cf223a5f171ab66418d4a27d23791c28bdaab5cef96558aa94074cdc41c80d8752ea65aa0d753f95491afeb698dbe8c41735ecf7524040f5ac8edfc6c184cd9b1b8a8226449c8ea108db3485f9f491857fe80a06901b59d394811df1752501e1acaaa728e83a82f01a4062cfbf3af0bcfa133c5909df50de9a27b4728e0b0922e4e26cf340b78642320548f88a4fce0e06597be00b3ab204adfa7c86f292fd007c15199ae01793aa1e5b13f5ba864f87907fdd3d759de14bab25affcfbdcedac7d64e3004509cb48c67fa50239837802d11af0ab4c27b14966638715f41dcf4a77663a1cd48b17c0889d829cdea5cb53d0f4e77426667919d0237f7ef57918f5f37ec3ae732b5f83f6f61437467373f70874fb47cfc9291336d9d4a3a5f4a97a962164f330279dee02f2217a5427d4b656dbdaf48812e033c7d95357fa20c5684317ec48e1e2df34c86bf5bc8ead8d4b334ef14ea48d445a396c148549feb0a67b9e902de418b22f8cafe7fa8347627fdbacd2a64a42c2570a763af79ddd252aea51ad41a9a5399ccfe0f98d3e294ad93300a7632213d41342ded42dfea6c63163e622ecad121cc3ce8ccff4bb3d92ee55c979a338b5d13409273f89a2a709116b1d7c84bdf8cc10dfa4607812db02f8541eeb11dac4a9f1cdba2771e960254746e9e4d0c5bed2eae3c0fbc464c56ce78c83505462ad198fe891038a55017aa0a3040e8be4965f822748d8ca4944cd4ac5fa56d3a3cc6180b9d75e0fae776a5a82388e9d7567c1873bba2f163352a561b7475cdb0e4ec9c89bf818f52e7cc8adcbfdab7926b7097ae1cfd99ea453055e48cd03289cbefd0b81d8af0318083fc1cac111d42437d293cdc665c5d000fed9ebf13aa30ecd6478a5f3d968cd4aa99d6da6b229469e013b595a05f0e3bc80518aa8598eaf013389edd7cf75499794797a66e4a3bf8c5d0f88a60bcc7d0724db9208e456faf24d10f2adfda0a78de23175a5e66f2382d8dabb93ab23ab6f457e03b2c0eb8d7d3fbe69d59837980918131c04bdb73d35ce72102172a82cb6e8187080b877d02ca5b08f02b9329c977e7644a84ecb124cec37648bb1957094915ed550858adb22ea106fdb497520d4a1dcdeaf54a30c497394e131ade7bce429daa785202d56f8580e4a4e931333375ab9bd30da5e81b5237f83a262b8590840b5c276434ff95c0faeac91d364d74f739bf192bfb531961255e7b237ec9a152eeb3f94a0cfecdbbdf8778fb1504cd9e52ca430e65e83e4eed8de0d023201bc9f36db67c97be612fc802db3f8b60fa61fcc4cd6c2c38afc2162168e7d4c355a2535c69d46b08bfaa926998484ea0ff1e4558c29e03748b0ccd7bafc8af7f10bcfac3a8b200a133b4d686e0eeebaab268e521b782cb1e7e04998532e609f8a2b9cae86d2155cb5f422f0427ffcad91ee7af3b39cfca915cd0fe433b3176ed8b68dcaed3fa94adf542ee8b410b84c87105a4a841f9ec9194d8ad91a21b68cd030c13b32;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb2026d156dac0a65d463d769b8ee531ba2d06a7141d9e23b3bf0ede89f57079a8f97aae9d5816aaa46822547db62a41197c38bbdf8a54501e7a38d43ba10b9d21055da4124918d880d3757eda1254b326700f592cdd3c8d5dafd36945b0de8043bccad34195b86b5a52abf92cf831bd5cf550b54aa0e40f7080e875e59ba0cc6d5c77014db3078bba9115a06c24d910c72ab3c2cd38b9a4901fc923fdec0377085fee07cfac90526661500ead12b248f816627de7d70a1a06599f855cb86f50f5a6612af789dd49cccb1d10f9b023c82f7ced99964cc26e9feaef6475fe35b8de511b466bffcfbafbca39fcc5775d79c17c54d7248fc774a08b181b972c4490be546c95b16459acac049f81140642b2b70011c81a8b4a5334b69f093bb3598f9d2b88d9b2db1b0b9de032a95116915a850affe29a5b41c564007f59eef5de030e3af6ec50fc5105aa57bba3202ba769305a549d145f34cf0f70cb39422bbe97e4fc9ed69509b5b5fd55cb0b4e7d70e05985fdd545970d98e85140aabfe497d7370efa59a0a3574b6041c25b620026e15b0e547442263c0279491902f767976c94f0b2d6482bd2b7d7ff62a8e581cf48bf50ffed2e740670741d5a1134d8222aa419f9c0e049f2fa4175bea2c21d887246cb6079eeff7a3a8efba71d97d7c2487b9774d7ded9ae97a246c7a4fc65e3fdff9a6bd401792b818d23fdb6e1026dddd4d4835d6107bd850454975bcf6b60feef5176e5f5fab7016e3a8a1899513766f53dd2976224c000c105433443c0c2a67e94aa9f70aa2d104ae33ed427c0a105f3495b10862d484946dc9573881d0ffbfb6d66c99b6b29eb95fb56174ebd863573bf373738a94c4da3115c75b7c72064fba1ece0039934e0052f718e7861841c687d07c69a9b5ba251b9695106979e3e66620143b05aea0e1c19f282eb27c3494cde3b3de53552e8e1940fc749ed420866be3a4e17b855c843a47daded9bca2b56ffdc79e253a06992ed5a349f0b21453e2beb3d18113f2f335b82d31666afd2b552f7956705693d67b6dfa26b465168ed3832cd0cee56b1da60864eec7051e5345716fd00eb105b5e6ae1b94f710f31bc7b23df391c5bd50e565cefdc169939ddfcd28b6afe5ced574fb9bf53c562c333084f8d901dc5c6c96d8689776785694baf225c3dbef59f4ab26495afdc5882a6b1bd6fcd9941c302351621e82009dc74194f3dc4a9fbfa5942dc54d9a11850cde0fd2a98c3e846a5fd78efd4dfb3b4a4d70529e3e533abc94ebdbb5cb6f3ee5f2c43e0457fd79a3bb7f880be281efbbb2b439c2bd7b9cb9f92c6e4b87573de6bedf8ff8d015b65a5966f11226c9f51aa72541c8d0615cb87e06bde6d6952d92ed7769544af45a56d1804db8403d0a1dc955d6d8ed7765424506bd3d96e0cc07e1ed55aa2b926fb8980092cda0ac664c6c3bf63a595b25ff5fd35bc4f25bc7d93d0a6e1d672cdea2ea821bae162a1de31e820a726fd8ccdd284593fc90739a52f3af0c4fb67ed0de871687efbbd882875b205a1422f4daf73748bec6af85b974ff7f4b81c6ba0b7af9bbb6c5d3aad6aecbddf76702cd657b03f4c59709d56f06c2f865eed85d27dcd717b04f590df487e50d342a5366abedc33c591a34b568a37f0ab862612391d586306043b137cc8a9604f1cbf802fcfa58f483e532f0dacc3f60e389188bb129acf714a4425c072fda1d95b7a78444bc112fb64c28f2c8c4df97174ff1f8305cf41b24b7814b54f0ff606691e56145bbe0d43ecf1935d1b79be4b680a8f9d47c97f8ff441eb4ec24cbf68cfc416e8eca510ad6be69cabc0d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1cea62bb210b0466b09918b9ef53c00fae06ef04d446c38ab2d19a70c1515e90c5c1fc7809b6e29294eae2e38118703e4a1bc4550b44847e5ba33a9145eb1c82618e7c104ec6eed8eaf3ebd48630e0aeeb8e0fa8c78274c62059159b75409cb92d0be029364acbc0fe688c42d31b2bf8450b2efd584289b80cdd231c279d2d77c9e077de496f2b558947b3d92fc06eeaf233fb9377d0c755b4ecc8cfc7a15378b3aaff7e6a6a577df64a58347bf1bcef987849e17106c1879a7981a68a39a248039c4470383d43059d60b114054ae8235a5d864d99e612604ad4e642909295b465cd0fb661d11a9d49b660c6a79de8cc4acf4e8584b5ca82ac8498ecb601cacda24246aeecb088a22a25bcf82e97a6c0a6a7d14ef83dd167e5229cfabb7199faacc01f2df77706981be91100686823d195f4cbaa70242cafa7ac73957d99b1580e6e10ada48ec8d041d5004604db42634e475666c5427c72fc4a66b79981e06299c94680543a63149c4166331a5cdd99bd7adc91d77b1d2de3e4d4a21c7ca08be17c22fb536357af384d0f55f79ef303ba1f7bdbd9f23a782d5d69130e6d6b75c37918316959ebce2a282909694f714bdd053084581924f91640b8e2a112827b519208980b641be8ec682f3948aab221e32d5bed123cd8b387b1fc0e41bc61b92067108fe0c7472bbf9045f9c04459c3559091ebbb18e02a7d4ad9ecce6efa98ca59fddd17175196a9b80ce8464a5ab3b2b527b7c895a6b335a096981c09ca084187ed40eb3870be683eb1a7d6828ac6cae7e98fee04bf7c49378f3257aab5a36cc97966d5b779330e31c6e1e4285a203935ae360b2051440d8ad59dede11661a5990806b579490d5af7a0255614ca289b879840d71374934f42446073d7c3c57cd683534cedf054d12bc4b2cd4f2190d75a26142a27ae16bf40a78cd20a5668bdc166592978f6785c64b11b44c86e68a58e8e738e8965e6e804d52edae215c5c4807895b8127e49d0d13bfbeda4f856dd31e6f73800c7dbdd7df75f6ab379b02cd9146624dd57e831ce986e2513e98619cf4785a70c7e1bd6acce088b3be76f6b5562e9ed24f6c1cf379062d8680788025e104c580e5111c31cb0ebc205afd9caee349a1c2d4492b912b2822a6e85a8e1d5ac25d51567189d3fb8b70087145ba72edc3160c3eb27ab84a3d999f75fffb12bfd967429c1d266b06a42dbee20695fcf120cb6d4bd6a62f16b035f2808466c94375f3e6b7ad97c0af61800407676fa00a57821bfcbf875fbf9a2dc8c6c4e88d08c611290a71a707189cb95db3a7f915cb51030f32760219c254d7e30ff0e804b9d911b4eac9668ae44c27f2fdcc95509013c748eb8f7a62982c399987de85687aafc3d3daa5b13362a4ecaa393779b5d833c2587bee55379de3ff49c5f7bd15a9cfb586e93a79d3ddcaad4d2c71c39a3f639e20b8ab23825fdea3e5bd236bc224f6177260b64c8ce5f22f58165246bbd99680e12eb12e9a43af6bc2343883e234748a52f85943ea17b8688db2f362a5543b3d030cdccbcefe27b736a4e14b3fb5ac427335318030156ef89eb426d432a70b0bc5c5688a0e49fb9a8922dabdb0b5f7d7ca0f7a49b248ac48719cb8a02dd1915560c2dc4982ba9dcb3f2e546e5554ad4e3868e7a78d7cff953c925f17f9e134a7b2896417d457edc2f0ac6b2f692ea40a3f78a70fa9946a85fd065fbaca90a963cac64a2c45fc2343c6a3969400f85a895b75cd5a4ad5733922529409ab6369c741d608a8a6bccb41449ecbbb02d6a295ceb421f7ce01074bd9d5c32cd6e1e236e36ec2fd1fba0d39128466d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3d7c67b94a93e0d42e10e7a2627716bc82ea3995166002495b1b126998c5aea05dab455c32d608a383550be8c04662ff424acf418c6f1e2df62ef5166e5a6bada9cfe1a21d95e37851ce58831de9fd57e83effad800dd4949d8157ceb30491a5cadcab97a691af14b064b7620d78ea9429d001af6dba5e0d6595fe61d2908408322347fde157ebcff1c5cd2708cb3dd2173a67ad6ecf89450f67cda8714bc82ca5b0aae0b981ead67295ec5c7924999940aabb701ad0a90af26a43ff76c376a65c6573f2b17197c5d3cc0d3accdae4e7efbab79bb30306fc61a116fdda66c964e61388089f3be7efbec358969ee1e3dc34d4ffcf317aaec6c9f92896b0aeb94cfe6904de49663ae44bedd4c41bd558b3cb7b88f6e424928731ba3375203fc4a7c5fda1e9e0c6689b89096d75405c29cffc77204970db24f85498ff4945fb1308f6f4f2232a97ad7b6cf26fbf88f711706db8a5ac9ba4df3fe58e8a3cb73d6e27794e2c5c867bd1b5a4ad5985fdb579f3b33e36ab4439f89f4673af326d7ff2c5d098c20c00a2864d4b25e342de6f2ca794ecb8cb5293588996ff8c5fb3d14d941b4f0e9ba1cb5c332b36b724435a52d1b84282c6f99ece0b64978c281e069852a1cf68f6683109864f9da8b2c3d2daf6c18fb9813db24f9edad68bb6355858d84b91550dfab311db74a4d8fbce88a30a00d8e4a5d0b0a4d3ffdc1055be151ce38873fe397429b72bebd3256149cf780fbc998a45211ca03ae3ca6fa84fdf7de551e4d251e738897719b1fc73e58d19f4a174e85f77e20b3169a76630aa548d2407018ced71ee96bc8f99c8a17ea52e4588460bad2b9dbcf611ad0e7587dfd1d11a6a83d05dd559123ccbe06ee53ce5632fa60031fca6581226ea266d723b575f04b9ba736c4128f4fce5a8a960b5947d7c6b7b849c71e70805c16d344733812c4e8657fc68788c86d4de28b7ffbe59a2a2bf187c138b1baf77650f33bd2492f1446eb13d0b6e19929e429337fbad56b5fe2634c5cd358db2917648c82d74485c03fc2dbe48c1491cd9088f39b1105622b1a42231bc36c1cd3f5b03df37d344d264769d42d04aeb5e3601dec662fe0ed717720caec2d283d1b57b0d845612cbb7df412de0d697aa8c80ec77342a07767e483dffa2b463370ff6ca4b4249bdc48b9b4d62839115f90c2138e882d6784c9247592c72caf03d3863dce6b9fdb37e645a28f40c0261ea1ed014569be15ac142fd74f87bd37699f733f849c8b8eb7a49d8ff62ff39ea84ab1f7a09f72148fd7f31682363b795a3bdbcc9d0e218195d23b63b0b2720a114f1b0bbb79280197078978ca2a71b7b4335bd58b989d54d0799a386b8fb8874634c4aac667698c9b697b46fec6aa7e60f1a8926917f0b37c738ff144aa2bc0c1ecb8a6db02cc4c4a169acf07124e53f7f2bc43b2f02261d4ec5723fb430c047579137e6b6269d1c582eeb46b58527f872f9bddf318e8d6e6f9f32d6e6bac578d723710000c562843a1e2e284dec51c5c3e2d61718dc94a1c356e04c7b8fdb8f893f84bac672d6110d7243b6ae6e66ee629664f1f1b5559fbc85a1763d743cc7473493e8b49ca4ced27c648aa7fc1cd2d5a8d719d52f4caba56e367f09fb7f11f3d537daecc8260413010181b76de8276a34730953f90c50bf2a601d5561a239cb1fdd2cadbd62055895af85e01bf6a01ea9365586eac685d8a9d3cfb76122c14630b68492659aaed04e91292f92b0904920a31eb827de552f5107d12bb93f06ad38fcd1afd24348d9d0e8ea8f6b06d331ce034121ff0691210c661f9a4aa8caa5cc73e541b8fdb64bd6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3a3eb72abd316dea18e5b26492f50e6ab6320d86448d8eff6aced6b4dff881f89956cc0d7e299adae5ef135ed4a730505e452649dcd2ba56d02926561a91fa2e76210784df8eea534aa860e33521ffbbe8e8f213a7a4958ba374fdbc2f1eb465faef7979fc7e8e129ec5471c1bab746dc34056240a961af1357742e585dbafcea952d7ee1126bc4d8d87ddf0911b3c7d86fc738feeecfeb31c4df8bc2d674581de66976fddfa9044c662f39b12ad56f0228baf43e52556819c0d78245725ca0114a5f463906b1560d1bcce8dcdb3a454efbbabdf6e1474cb68ddc2766c555ebeb8935a38e03c2f3a55e86f03c41730b5ab1d4162ca3bfe30ae3da845c2735b99817421a2ac85c42f6beded8172eb76dbc80619fd9c7c12961732ba0ab8477700dafe7a34886d3b70c2d535ec5284bab890dfd18193f4823851371e5b5d3ed5ec7587706d2598ff87121c9ca26aa16975330e51b595071d404271b0f9ba21c7da54f2d6deac57dd68a5ad609199fa8aea6fe00207ccff64c23f28c51a8f81f6ee8e154a0fa1ed03aeb061f31bc79e3fde8131e839b056f940a05c41d6ae7b2559bf462aa0d91536c354d958836b98c5043ad020aa5b30a75bc9067f5904ef98d1cda828d840865a9bd92d518f4eec76859b8df5387a91a80ffbd54f8b977dd9bcb07d6d8fd83e055e2fa7cc5ae1e28471e85f2a28bb392d1d2e7bfa816ada35a3404f4e04cd4f292eeff195e7b4e398e7672cc87b52a200d85d03e5f76909f18e392f45c1bbd04055e3fca1fb6b1c17cba74e5ed2b0f1fb193eeaf6d9ca5f8940868b3dd6942f75f0b21025a0019d987ce4b3ce73349957b4fc7c1a29c456149b2c28f62d503407b9bfeb98a375dbe58cd4617df25b00819d5a3672f4433aac554abee3d0cbff825b768ce9069e3195c0754c881f9ad7b2f64a8a7468546950d10dbdef8add32f94a275ec966b26c32bee4166325adcb664effdefbd0d3a0da542458f11b153cb4dfa610b77bbf747105260890a9fa41427ae60c112ab9f4c09e59fefa438eacc97e5bc49d0f29513ffdf6844a167ac7eed9a906ab57ddf1f7a6fcce3d2a17eb2336f7aa5b6e8bd49c56d97c64ac9b5cae3f3cefcc127d4dcacc6045db9f78a02b8779bed6453424697602acc3530419d85dc618597efabe49efe99169d11cd647e3a82d4ffbc040c1db946b8ee7125b974b65fbba4f3b5985436b01d8a63e61351d27ffd2c3bfd424133b39a5c3fcacaddb1a21120ede4b27dd2dab4d0ae10d63e6e622ea0c88ffeb61df26d065e26115b8bb22a0962af04780246af70b26f560f32525ed463407c9bb74e7fa5b954dfe9ab0fe5ac4eecdaf524354f59c39456d22519ea5d1c418daf95950efe54c614fb9db1b95c1d61104fa814bf12d6afa5f796b3b4a5a1380488bc851b5843e8a95aeec289ed511dbab86f5ec3f6c6cc582d510a99b456736c0e7ae30df8a137a780f9da3ee1058334d01c0eccbcc643787d26bf8e832bf36fdee8e07440fbcbfae84db0c10758c368a723c27ec162087bdab361a9e66ea038a291c5bdc4d5614b1f184f2bc8a4443dd8960882fb31e218c4d8d75bf9e4552dfe551b84e5c28cd44c8f4e9352b2f247711e92ea8e38d9682c87a2ccc0045fdb594cafb20fae7474f9f93f8fddf8c3ed3e813dc9065a4c641af1f54f83a86176ff71930810c69ac23f24dff91a337ec1714df3812a47397231fa94d1e47cda26421a16c95051307b6a2c04244b87f8c2c55caaceedec46fe085a2d2a954066529cd2480d73040a4fb01d4f2a6d7e6467e789d63e346bef0169bc6488202946865b6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8b109f96444a762d3464e1217e20350b8f52a915b8efb5b9c81c9486265aa65af0c97bb1b392a5a921cf9a7f528d2a9cbb70c936fc12d4fec7b3b7e6193077f33614e00441c999f66484fefd5e5e319faee34a0c5d218296f6bb90b4e02df3cfecd38f28b185c346f5b9e39bdba6b56f30c8d0c286a1e96e49f98a5dbc88aa9192c98de378012e57b897fcbfd215b0edce0967a1c67255bd83d5fe2fb998504f32e55d294c7733032fe62e2f3c95f0f6f228ef49198cd38dc29ecb1fa31eb0686e3bc3af0b87652d46a68c58359d19b951ec7b8cd0d1429b6f9c7f674b265cf9666970a149bcf8d31da39ef1af9ec35ef1a453e64e2663f757f874a13f8f136987467268e7b91f2555275357a90d91a0b60b854ba0907571c8c1e7e2054cf806a30bb6b5c7cfc08c577aa7043c0e12fc7129d65528b7afee36ba640b4fee974553647b8cd53a57f637e65a762b7f14831363e0f3f738f5ebae13665e85d36ccd17690468d7005c89f86a3b90b43667e244d6f55421bb82205238713f0af3c257dc8672b92d2116096fa36c195c9ab84bf86e8a93e53ed9c30fbd9e40c23175fae8c78e9825d7f3845bf9b5540c8b517438e6573a46b1fb1d2cafd2153f5ced54bdb4345af03439a17f080973bff8ca89467db3035789a38f2ac0911f8e2f5e9212e9b41afa63a2a4cf0131060f42c148eabaf5389069ee9859f0b0161261fb7d0abdc24154a9e22be835fa4e430b3ce2ddea438bcf9df82161984a958b8d51497233821507023197d33c5a596433ca7d7f9de1e8575cef660a98d0c63930ddf5f0a7aabe3e233b487b60a4d59a93ec6a8d3233d5e63a6d96a5700c7008b3cea29bc8ab0c855ecee4c2d0849bdf3132e222c68f98d451fe2ecc6df080ce988020398ce4d7a6d5e8d46e45a9e7fcd06e67c57d9239a65c9b3923adb69c37298d8b19f477d6d912e5395847904b69d6acc8b4e97cc0222b22f0612bd94304ff0b6df55a1d412e309ce90706481769d22bf98c22f097d073e56fa834c524f96277b5fe7915efc8bb9957bacec9b00c345d9e37b4a4e5069c02fb2b0b145c6b27dafb4db2e9ff8c7a51320b834e5326b4e05f0341b09f77dca84712f01be6b2e57545810ab7655db1a85e1eca301f5c549b49d66bd08292ef7d83a8ce70cb773f2db7424c4a7d96eb8f5abe1a75f4cdf5ca6e1d568407461654c6acc1091157d2653aa5441f4fa0dda7594c47bf9270f05882eb39c3db849b250cb937f80f8d4678bbbbabff07b19ba79efca022e635e9961f6500108fd4d4caadcf4f9495a13856e1a872a529c2c8dc06e86f76aa41f51dbd145c02f7061e98a4e061329fc2f1c50204364be57ec2cac049c2ee8009edd70a54fc1d9159654fc4ffa1f13d97cd803b6e2520aac160af843c9964f865eb90ae6a98fcd7146b07fdebec61c7033d3907b0454e0d10c7e60bb5b918c3494239e0006dbbdbb2fb3e2cac1d0bf47e38996f405859a0bf17e1e8236b4dda8c15a18e486086415507244a90e46a425c50c6d0d15a2e89fcd6c592085e45a021682ff072b13ffe45985e6ce6d129faec2f6eed4d0a81d9a1f59dd175a8027792e3c2bb024f58add765085f0f00338335c3efb22d2603558ab0714ada45f6a37df4b83fd23b1c745ee07350f45373785411a75f5bceaf9ab1d01b077b6033e9fcab4e4b27e66b3dc3cc72223edb6db5019f53f4e473d07bd0dcb7737784e22578fd3c3d485a27ed2d4a7e631d78758df2c1c5823a17e1fad1c557d0c9f53a398240546e075108a0b553cee4be01a9cd69c2e70fc228741bd189ef7031e4198617cf742c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6af3c26bdf46b13c96ebb0246b6754ff8ff5b14fbac9092581e20394932c14194c36c9221b1b3973d6c86e06e85b6fadddb9bd81c0b91bb09d95c37b25413394ed236219bd3e0ebf567ca675a0110c7ffd33f8bd543c46240c6d9717c8197a5f4313c631e97787cfa63ac32d124df24e0db25a539a10d4e12c6cbfd0da32a7231c80f2ae917fe18405b6d97aea38e35052704ee2c0e25af039655759101b9e38891bedeec6b0e6a1c551b93e49a9e7a9badc368d9cea9c0e65d8939733d670c0ae57ba778e8fdeef89287c95593f084410c94b4f228112993f1ff986da106c3e104347c10fa29ac594f7f3cc5bba89ae3752fd4005ca1b85ab8c27f96bd5dcf1b78a88382fb5feaff1c3dbc11d434e7c0d2f7ba1dbbee061d30cce094723242014603cc8b68bb350c3c6c7f0c6c8ac9b8bdd269f287d5a2c6d7b5aa8fb0db730604d5e15b4453fa17bc8061cafbd7cab6a9f18a7f3b47144ef07079f34da189fdb9fc64b63d4c9ccbf9b0356e15056cb565e3f98d9c7eda91f67d593afd9f356a7a8431637f1fad78d2a8399fac77f0bb197e1616156c43aa926d3c44d4d1f8afa700f76f291c6aa5f8e39f18e5d8815f113cd781db05c01af1d208323dd457f07aa3ba06e31834126ed915a9178b4abf4021ca227e6f78cd516f2f200bec4ced6eebb5676bf8703186219031bed3d9945600f07da6bef149491d2881f161679b877a9d4de9cd6b48e171c77de3e7920bbfb88ee8f4e4c21d4877673415566fbd208f7535412dce865df29db5bdd57b0ce4b1f99cdbddb17819c59f2fe1e5744a29e008a4236b854d970fdc52695aaa133ba29be83929b238138e4b4b02bff7ace6c8232f7f6ee829004eab955cba04c9804daaf3c8fc11eb08719c86623b867b02d5b6c5bdbfee751c9c32d5cc4f4bf17f57cf3acd89d57de110d821abf003af0906b24834408bc60e30e643392bbe895912303fc92ba0076993f74119cfa826f90fb88f40233ec99b63a7ff84d4bf81256e2898736907d07dff06839f58fe494318371c6dba73a52ad9addfc2d8674520ce05b046138e508e72e7e99a362c980abbf7a16c113f7b3554e21d17313662a56ceaee23e2eb3c9dc75e4fd302f99fbc748c0f83f30aa0910ecb3014772afd4ec7f103f53da74c4e5a61ff3c7f215ff7ab55c2fe720277714694313747a6fc6d6926745d219350562a419c7bef199ad8c85b1fd41474227556d981490bc54c74d917380a925b9a31ab0c15b3c3cbd63d317a3a8b65c1cf8d9849ed4ca4274ed04a81550b981d26d22b50fde5834e559f2dce26eaf607dbef4da84d1f7e0b0c6b24ad12d96c3a5d27237ff3fee7df416a79e2ef571533d8c0c351e11dac8056f7b3dd168d37064423ca92c919dc4b978a59b342945b8556d3c2f568b137647eefabe4ab036f4a80b4634d72fd40f50c65f2c9c67792dbe8ceba21041d95f16586c414a4cb444f02125b0bb0148cc84141106d7c13542f8db0d40119890f7bd61a95349c253663b8e2d8f07719d0685962142917914711df91fdb6f477813c4f61dd23b24756093dba0fb82564f6328cd4d4535fe3b714c6f9d4f2763189774da20b1306e1bf362cf4a6b868bfd5a20b10818f467d7b4325720239d1c5b55015ac055e50649a006b3a5083ea6a19b16fc67a856ba819ccea6e697e1c7d8cfc28ac67a10c3565830fee20ab4c8b3273046e90478280ecc6976f3a55e5c83e248769e063e410d37f12e61e3d2850b90d167d18068862f2444b7f0118efc4d0460300db916c9be1f54b710cb2d83f869bf36daa41a9907ac32fa6d8ec5fb21dbf9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h40aa4d0f5fe51c4151b4f90d3deed7770d3781b579b2722c390f46b9a1e4142114f43cd7ca5698b455e72c0b5f255cd21527c9f4198164d45f06bad56760eb35fef05e1a049a60b8c5d02e7251ae44b991b16d55d2dcfb71fe21ffc64fc7db9d947e5f308d7c1f8af6189e321d2d453ec11b204a0e7082ec901f124a5e76d60406f06e36ae3321c0b56c9762552979a5beb4d7da013503550bfd3236405ddb3d90321868ed980d4e5d8f4241b1c45f27d460382905c4198a10fc1bf4adb2b43ec618a01d02a2b459d873177aa6f0a1447860abca76c086a64f8907ef5b68db72e0601a30a5bcbe5571d878862741243898101ff271768557fbe32cd46c6488e1d6a4a5ac5d46b5575e071026d042fd66d9531ec2c31e3d33c2189087beaa79584665c1ad6761926030d955444d97e64b3fba08c8cda6d1f29f5dcf7b8692c727512015c5cd8e333a002dea2620aa752d6efbea3e3ef4dd335a378606cc93ff59e70cb029ba4a8a8ac86c1c7e39c0c86ddffe193423043c3d73ddd8cb452037d6213bd428ca49712a34ed094fc73c45d911e11499470e3208d2822064523af3d6e47198d19f55bfdc2d14beb56a39b2988d6eb0fa7bc6f404d381242146e0e0f3f32a9586dca6df809b7c951250fed996cdf6c473bfd469cb52443a9e31ff1524acccbed1cf39050fe72dc2c21b0728d65bb802ad872830af834c571aaebfa38eaee51b7d9438e6ff81cd2ac6130bc64485cb185d2e946b2e4ae8f46f84ccd2f36dbc6e3e8924cc21f37a57be7e3da8d935ed3b8e2601fb5b434d0792f3c1738a77b2a03246fd699d12ce4f9d4deb1e66a6b6b46c98595db700e40a08721304f69ef6c174db1ff281e860df7bb82abb99b81cb67f8c5fb9ff65caa2bf8114c9c3e209a1fb576de666e6bb986878bdf52888003d13f8ba65c93b0d36983d1b070f20b483ffd85772cd6be406b55b1546bcb4f0a5145fd423d30e57d31abb4872ed89fa4d84682b1d26e4d7b8f4ed69c7dc47b9321913ac2078a246e186106f6266e159ad15dc2f52e67a1d0321f515b42607d9b5b63f88708f0072767ab087aa830618a31b7a7024c7cc937cf1b9e47c0e20916940769f5ef9f566730a424e1881406ab56330ef556f24c1a973d0e1fbfd5e38de276739e32714cc78c07e7c68fd6dc8844f88ed706741a057947c8cfbdfa006191c67f79a49ccf9ec5c6f89245aba55bd8c07cc6fddf6895fd623273ea5ab59d09221454ce3b67c3bb9c8b20245c263f1ec6e28511b60b59b53c67f2796f13645ef4065d969cef6c683f35030e3f8669dd77603af1ba9136da994c02d6291af2cfee7919c533e486e99c6651981a5c0d7cdf666ec0a1e96266fb64e4e8cb47d78b10c7476981aaf2c248929004786b56fc2f3481403cfb2027945b273a572576bd151e8de238354bdc048fb5c6ddd74cc31ccfac5bb505d80ae04c216b2553d4c033a4d470565a243cf4bc6df60ffe421aeafe4a9ef2aadcaf44af527a40ba9f747fe6a1fa7384b9e8ded0846f8eb1cf19b5bcccf75026642112f4af06f2b8ef9560266b51df3abbe555ec93c33bf9c93822914eb42649553bcae7bdc556cadbd89ddd05d9d218c502a9ada67e2536e95559cc9ef2ae3b7fc8d7b159490bf75837f9cc137c378141bbb1b326e9cf3185659c29beec72fee6428de7d21956fa8818e4802dbac69202b36e4472998eee41ed361719a569c13abbc9eae41f84fffd4af0fbf1793434760c2852a88947e3490c6b8f913e023ad67d856c2b9e5f4f3dc4b02518034f2404a58fb4293bedf4aa5a1ab8ebea7f6300a7f08748591;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h5228a50dfbdf372ff4bd108411b8c5efae195cc7a0e5731f7ea1bac8785d6a3cb4db6732282cffa914ed35d4d85eee8440fa6f67dd9cfc57e110ff50996ef83487801e31bfc9d3000bf7c86363ee0300de881be57cfa63e3b5b7c173c91df1715b7f8ea1749e5cc0615311c354e10f6a421b86a033216ac5517335a97538489fddbe3d7f7f0caca3a73483e33058754f78f90230fcef642e876c97e0ceaa0e40d5f2ec196f937d87527faf2790c5b27ee9adde936d4e443f5ab835769ce3476ccec785f6795148e243bf0623c949f44d51e63157d2e6c882105728fcd71e11025ea9dc97f479764a59612164a6e94717f9d98f7361fd78dd28ddd395abaeae7058c6f066d40bfbcdff6f2704a03ae5e8d549ef18f8ef0d19db091ea3237cf300a5d85128b4aab843c6691d61d99d7ad1b79fef1eb323c3b53b3c3cf68c5ee7c8c00ccb321490e8449b0a93e0d84831cf15a063c3c857435b3fd07013c8fb6b851ef1d3f04a3f0e1e3882ebb23895100e3147a354e6ee6a4a3cf58d56df67362ff1ad2d37d9dd3b758a2f3065e5b8c1d82f66500ebb1db866ef09175a24f64b25c58a51f94ccfe1df4ddcae6a0af8e8958cc4f1dcb6b661fede90e44f70b13925dc8a3fcff3e3edfad22049a55bd0e8ac4b3979459ea36fb647e50421a59051894f9fc612be283fe9f36710b83e816b5d01cfbbbb718ad06ea9a7a32780e190c436a4cf8d5bc933a5d53badb3ad5af0c98fa5394d4cee3d54afdb2d1325d934d90df0a9cafff2daa45457595370d65da2327592a160ca6ed83a965d20c038aacc690517fc590d04b4c47b88aa32527b2f0eed1868f11fe9405c3c3714d709475741ee28cf3fecc8e3d5685ca029e762442165775704d8d5081b46d5a8b0c806b97341b113b282176b5f091f3754d7efdbcee397ca2ce37d936df7acb9dff0dd0c485e2ed5533c8933ab8cb534299a27d0093d00f7d0c26873e5a15334e382ab8dc8c3ad45fd403c5c2f06ae2e365e28e8a621e76cc6ba1a0793a462270048c6e1569804e7a029562fa9258a98a44641811f5cc58d8bc166b60206b9c763c3759905135d672b4599809c277591deba403a041e63e53dd0796a3d341d16e576a1ba49ac6adf3998c287ab3e575aad6dddfa875b3e9d14569eb516d9db90ff6ccc6d944b11e0c68dd07bd1e911ace515045a3b313d22862d599e008d03c06b2f761f6d7d15cdc29e512035612c8fbb721cc6c520095ae84c7d785ef0ddc8d10cbcb86fb03a73a48873d944b6841449ef358be25c93125cee496c4c7289653465bb0b2c04d1084f172b3f48e408954da820efefc4661497a490470c005c366d3389fbcf4876e50046d28c6481147b851a77303741ae998ec9236c2a78a3b762533b0a77ea5bfa6a947e2c4f548a1146afe5e491d624d11b13441382ca3ec917a50490fa7111bf5868b7ba0c211167475c3ab44159ddd1976262914fe58eaf67604a850e0971694732c8bb20600dbbd41ef261c087e32a78c4997d7edab2622e575fb8e6ae7d7e30c93081d56762d3a4c76894cee755fe848b89f85fdbb70b93d357b60c830830b176e5b54feab4d6d941bbaaeae1df29f4f8de5ea39aab98cc5dc82d54e426e9428c4039fc83a3ae9a3c5637f071757d18a268315e1e072f5d923fc76c3f795240957447b939076657868b244a6d46a13b1a7c55fa420746433af1d4b6928b6203e753b76419e8fabf3badcac9c4fa5130587a2027c07b3f465609127364117c41158c361ad404ad53c60abbb1586fd3cffa754e83c856bc311f4102a89ef6550928f21e0f9609b746d97945;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hfda3460137c3489928e074c0d337514a7310040f3c95f8c63368371935459143d9c3ba2bf62ccaf8e511210f950a89d96154a8fdd5a79959ad9d0a76da5b962734839b306b7da3fd69a02978951225ed9f591290a4c77354f689e992fb2b312e56c7381919f72d3bb06092e02f376cd713251f947bb64089c38c427fa6c18f672557a9e31572e4b45256c5d8f4c76a5b688d6ec8eb74eaaff48a89b07d1446885d5ea7f65d38b025df882851ad0c48fcf7cfe836f47cdf0b5eb6352b3e8b27fe8c697049062f4b7ff08b735307b6820dc59012d38895164df8c7e45652988f23c581bf235eb7f8d96b8811642d69e06649ba79f11e9a73b97d6e0aa014818b8e9be625f1b0f0c0dfa2b914f7b94759a583c46a14d0e3dd017139b1d33fb37d15f46f9c2278c6050e5feddad7e8ae51caa97cfb28119d6a67520814850ce94b9396459da71d043e3d4733e32ea4460a410dd36d5d3cb1060a88a587d6663d7d2f5625081aec704cd57a415444bd2fd52b5876aad0c981edc4447f03c9b40d8b64495d749e77b3a46ed88a4a7997e7cb247e52a88dec8a5a6f4080f4915c4223da976703eedffc4d85bfacaa13ba6b87dfea25b8455d41e64072273685b4a2e6a7ffb792564c2ab68b3bb55b28bd23479e99e1d20214d5e598058a02b3c0429e3c8461c6c401c4609d675a05ed8075bc5055daecf00e046eba6f145b67c74f3e450df5d74b21dffbf201edd21603cf6b9636050ae068f1af938f5fc578533d285590496561094b89d6b7f37ee7bf9945b9847b73b2b045cb1bac980686e8282f5074033fafb6a08a70ad4b1bef99589b5a46b7d8830135dc25b0a9b02ae579407e22093301999391f398d06b9791264277b10bcc7e0272d13071403952d11ac92710418d303f8b4a59f2f64fcb306e694c74d3b0c6b9be022c3a86522b5f26bc85133c6e4aee677d9d99b8102e1a78d13eb4cf38e7707694b5c8138afcbed1a908c421c4e474bc695bc39555348bd17d6a98a13b727acd0dd178c19ba272839f3f22fed73bccd00735c8cf36381284757c7f88983b909e687329e24619edcb6b4a632c21e572cd954e4bb72d2779361a1c0e2764f7890b241b34d5fa6f6db0075a8b0ad9dc70bac1fbeb6c2c7ba8057fede94e7e37031d805674e33afb5898926afe56c828df3c4d0497392524d7b30c545d332f42e2f5a6aebd4196ed4a6045236a8bc45ed403944a014456722b85f560619dac2606947cbbbe27c7fd7c1d9ebfc586f94a6217dfd3ef49ce2677aa6d5ebc1ce105f71530e98446791f1551a1bd24f4cad38267acf024f8b842f055e0f92b103db5c7c145ab3be441b09b526b92746fbca8320c620070af4e63157a430bdd5491d23daa89b1244b06e3e173f2f446cb9c3500a773e9298a68ace55dd01fade5a886b6c393c49a01e3a29dfdb29ded2b99e83666ef10ab227f3c454540d0fe7f8107b018e2e4f2efe437b127a126b520f17a923fc4a50d07e5a57456b6fb6fcbb36f4bd0ac8b6c1ee7adc491fa945164fe1bf70b1814afceea79c98f4c242c3cf19d8afed4e548d1da23505cca422a55dc1c59261db152456d79f7f4faaf910e057b3ef76d9611e29c4fbe1bd8a2da7cb4d2f4371178e5246f1a1707e62d82f8d3d9b4a691a83fdd556649a8206a1769c17807ba846d3e90fcc966fb02d509e560efeda23aa36258aea65afa890f0102ae5b0097da998d196f3f3fd974acf44d5b6f9f0568280d004f4d86e7609340d9d66aacbb1a7c84db4bf8e6ffede727d9522ff00fe63ef35f663492c89eb602681f1067d9d589fd223324ec9d47cb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'ha13aa13200eeb989f4fe5584f8f0b341444476c10c48c0456cdb1844a0e31495739364d9509043facf85c1c128f45631d5c6b335e2817aeb4de07c3b2dcf4b621fc73608aebe5a969b0d3649582da9d796f745e790da78c088a4fe349f173b2159dbc2cb70e04af3872a1d93dfffad60925f6082694849d8def4f5f82174703228572647258c2a901cff5e2ef38cae92ae87feebb9c66a059db8a3e1cb555505e8fa3d8e1e5f246a7febb7e52443a2ffd7795a8d39fd96bb3474de6a130042c434dd2fa07f96ccdc5c8b65b57cb7a735a9f0f5e4a3aa34a1d0648d61d95e8bbaff7c955abae10d5200bbe6ef2450e1ed16b84556b1b619aa949639b72357171a1ff0114b614347742caf30952ee71bb315f7588f1606a2c3b710e0bc323156d1b66f44e9ddd0a599f3c8858178f445cd2221f53c526f9bd99da34677e5ad0a9590bde40be0574bc3f2e413d80a38b1386221799f9ef56154db9a489224041aebf35ba3310576538e5adba60908e1f0e4bc8a6a806e25fa875f64a9cbeed5a322a8b078a19d9d688ff1be4b70b160810943c2d85f1981f567de65433a67bd67a323e44afa4473e2172475993c09259d20aa79db634900bb7ca63788c09c9856c4c9ea40134086dd31b28e482e10ba67c85712c394d6dd4dd3f9b3c8559b5adffdfba0a93a7e89cdb39d86ced6b3426ac122a87492d865c22a8e9da9c9e93df079bd1cb9eaae373149eb9d78f4f7b9592199657651de14016ee4a083d7a1a838bc5fa2113fad26fca00c9e4709d64fc916a807685b76d5746496161ead4b8e7b005e2e8786df86d34c8f810a77942f9366fd40e1acc1cc03bf3026769b527f6f32684605f3060bbd968d2c257da70e97b768dfd836fee18a6c28b2068cb6bc5a14b94838c78bddb438d849e60db134c77076aafb8e0df5478ae64dd31ab03a19ec707a414bbb465672ab39d4ecbb63eb7196fa177f780699acdde7e70d757c2f13f45314de5740a7fe78a7c037090bd51d96f23ea8d75a5df04388dd0c032d87793def4624e3b3d277339c6428ceea587ba5a46bcc9a91985ccfa3362d0f336576304008372f37476741e18a02958a9322575e063d248afdcb6718140ac0607c2f076aa000da6f44d20b5470f53a34d80199a170d732cd5f9669db912c39c1fece2a52d84d86c7d81f97e05a6e992ba7dbd5dd7d42771fab15a54752c6af4ca99e219bc64b09d058d894df1a689b082a7da0da84f653233180f9011199419332405df56d21ed48bfe34b12a7a85d3580714b9a120f4704421750fe3c0ad5cefadd9429ddd6612bdc36aadd998ddb0310189ad597abf9472a44d15eae4369868f394ddd3abd736b7317c3b351436f361a7e40cd6b9645073658d6a9203339c8886c7107a5c4519a44e33bbf6fa40ecc4ebd5a608ccda10dad5ba9713b4d5a39e63e4b5fb9d8f3a3299de501cd64dcaa598810235e364ff15040662d2472515ad38006ffcafb54bee863354b558145b897b28c9ff0958c4f2f61fa8ec3742aa88be8aa97f13e589d29e7409ab742b2bf2d3165f7cf01b94427bae7856dfd97534626ce60d81cc1cd4c6abcf47c160e1e2ef94148040caa5ee346ad005183f04b82a8a92978cd587c0cafc97762540e01a023438056b95659e4878f56f26ad4e034d3bf6aef13969cd507d653f59e445c537b9ba6e300c94b29d55d202f6757eead5cd9039da7295228598e0c8db51f4f3325cd15792eb20b4f87c81a5107d1f3536b0c8bdef639c21918ecf9fe26f75a634321f5977187e313cfff708e3ba5a3a5c433ef51fff9a94d559d83969f6ad486cb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h853a1fbc44d6ebee98d7461595cc07a72eb0d0ae7ab160db28c6c0b961f77ba8f86a95eaf43c9a8c3870309083568be700af1dfcec316940be29d70922e3d3307e0ee6f55b11becd75f203bcf079b451ad218da7140ba1faa03b3b8a51d36bcf65412e608302eee5593b17d85658f3042cd7c651e9b969d71a9bbbd54197e4736676d61cfbdb3827610764d7b707f1bd5fd1c151ddcade47550fe150878bb78d98a86c644e483314d4531463d29eaeee08d1ad433b8fc16807cbd69cea03ea0e76a3487a352d970322302c5ae403466a4ee1fb7b0fbf7663e8627e1786b9708560bbd97b01712c386fe4ea5e4f4bbae3a88d287f49f2f6ea672af21d3636e303585689b292fae3bff26df8f8e3db7fce728eb1ab5978da6f0216f4c511f8e74044a4a8a297480fa6d24527dffd5fff86dfd2459da04d435259bf99f6ffdff305279da57845d8c4fc1f4d0ef074bad3e852a380807f92296156cf472f822c433c1ab90dbab944936edd67663033d2c8ee966e22b398e0b9223fe5d946e7efbe4b164840708b8442f8d38dfb3360f79971c2aac7adf92114464bf8a1606a75c64af4212da535368a5f9fa67fb0e856897f15e9eb0afd2e6d9181ca2ea40463f0421992befc7da45213688a1726c7b17970c751643f0c47ce3d7e4340eedfed338ec904ac3ba27c75500d50da4918bcca2c5a5a38929332a5b31cc00c27cf769c6602a9b9d4f7c91eb2168fed2fb900d5fb0afa1dc1eb398508a65179ecdb1dae8838dd1684c817896f7ef5867f468e469b897698df51c9157096ceb9890ca50c417d53731162195f39996e54bbf57b4f717c9eed12171c4d4d4801f1fea64c97bed2e5205733d315f668768af848f9e19dde1cde69f68d854b2bbbf82396079b6e05806326938a893f12ab23571e6fefeb3328feb2030a7d8d644e82c755c31693026b2f4367baa99a2b098e0aba5266b59e38d9dc5caa0be25222a42e0450463053b65fcbbb713e890d72cb956e2a5a1d1d77320f6d6b82b4a6627b1ed5d35c135e2c8c2533747e5bc6e40b6d83ade1f2cb7b6350aa69b6e477b2ca94a395dc5b08310824f0183954a9a29dc87a67488d5fb5609ee19e9ae09d6463b2a4f00e369fa7356f13d5b0e0973d82f01aa080d3021c1514c967e9ed5b09fced3bf337210deb5312200200966c169b22e85945989eda66b29d14341b6193a4a31c89cbf0685ccafeeb9681ed3a9cae785f361ca36427650418e59e76687e706999413142e87d8cd23287208a35a3a856157c0e61507603b93f9c5573d08adaf5c873dcc9db851d058d1bb0b428cf59a08b9c06c5be662fe105b0a215de4d992a64b580736a0d9e8413eb6793f91d633213d98e4577039fc3162b95cc695d26c308477084d4417ebe9d57db532edd751a5c4da51c2d0796dba2acc6ba1a3d429b3d3cf25a5f029a377bed7f37163b2fe79f0c40ab2bf6d711ed18a9a6b6b0a1dc443b40db87006792291e60843144665eb21358cfa2107bd5db2cfa8426f1b75c590791887aa28876326465736658114d523c5c34aa14490d0e5256b244a23d0b637de99a0647ae873dafdcda25a44531a45a4704eecf790ec3d79e4a7d535b8f3287fbe4d2e4645cf918205f4be7855115a20d0e486dc2813301b3b662c8412d28b0694355b2f231a6ba7a7549f302af8b294a6fb4bcf1df0216ee8da6dd9269d0b16a5289142312fe7fa63f2c8d87d02a39e23541b8fbcbd7b7e11e807beccb15faa5fa9096470e9b6201a3928df98db594e4d9684e5ee227c56de1d57a6b98932cf3e9dc62a095085756d48b34d34dd2346a07;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8773ec5278790ed247cc090fd5e35e327b750da6584ec75806d2e9dee6081cb33bb4a0aaf676ee64a87654d47d1255bf1597610d9b022eeb2f79b0d2abf935dba525d8331ad1788f132d53d4d2610010c3052a1d14fb2bff8cfcb7a6b83d2b29a2af53a4a0f5d26ae1e644214a49ef7bb46938bc714c1eff087756c6b4fa2b221e45b201db2e6bd449637745ac432da875b14a392ddd60ed25da58db13fec0ed4d187372179c0e436df3d06e173ee98e693b7afbd895e28a0a2304910dca50110655c65d7470f2e44324100455a36399bd557f6167091e0350a8454072baee145b289e88357cf0e4e7d362e7673dfd25e9986e265c0a3c87cc85d29229e25f29d66f366d6ec07583d3f70476f0c0081fb4fdbc9f102c52e9adf41c3c57f189ee6a9aef146d7d632ffbc754d689e92fa69ad1f069e0e074bf13c8c403461c981fa1973e16b49afe6be89bb347d8a4e753c7ae7ea0c218eed28b2b26ba17fa82ddbe322761b6a2baeb1d4a5dbebf16b8383fca4feda68dc8e17c62bebf1524a409df9c759cd8ec2a137434e888414b8925c252a119b35a0c5745f8e037c7925eac56beff885cbba1071295039a4d5c952004bb677dae1f8ed97ee25470c5cd6bb8adbec111ab8af92ecc7e788fd225bb43086b60a389003aea91475657d6c1bea83b8cebe6fc8892dfbbf37f4f468841e013e8c5d9f21909a54b24010813d7aadc6939e8822f5b414d79171bacefd949572258673b8e233619051ba07abd08a57afc00dcde629c9100cd20e3bfa65d793b15bac592f2fda78e6d115d9615b024dff3609d87bf413ef42b519072ec4adf1336329bd96f020cdb4505ec95ab3bb0cfc820cd0a78863b965cd3d485ce92d4028c45c588f2ef40ab8cd31fea0d4b1df16319453c2308236c9ab8dcfdfcaa13441ff0f7bf490041694b87381289e4e05e3b8a0226f8f918a36f2d347ae86d3535004274c103bd811eba5c113c044ffa796469acd52fff7ba06e7e152639fe2acfa62b256eeed04687a0f4eb76ae97c5822d6bba09e73f1af4e954ac66fb02edddf886770a340ce43766e5dcb55707fae56c2e828bdafbfe5c4160d6137746f1d667aca33cf21ba7ae046eceb7a16e695dae9d5858ece30f77df5fdbd9b63fb86b8d936122f0c09417fdafe8b5b25eb29edad76145b59dd511cd2d4046b74080f7c90c707a73b19611f846b997354ea7240441f889a06ba3ffa156c7700251eace7f9db4c4c25fcc33529e5b383d9132bd622c83caafda78b11d5885d38ac504123d66dac9f86dacba744b807950666f0b4da8750664cef0ea3c79a42b93b4e6d82196ef4cf2e1f2049ca5d1a8854c5e71722083abbaa21faa6d94068657de9d4048faa24d0609d30061d7ca762bb007a91929eff80ccdd85b1a43ae4ede46dc23d967590fc18aa95f14237a53f54f2e2c4f865590282e31e29d207bb262ad0cd1552646ff864e351b4134b15304ed49842c979b15b57c9dc742c0a67ed6512731183c5261d8ecc2f1fad3502bb7dfe71e9a7b9c37a3d3b3ef67c2e4af2dfa1d9c35b717d63ad90213f807aaa9db60096095465b4bc851ca611ef80ceada88c2b828b17008b35aa0a42dddbc84c96e9ec53a361c6f9a15121e80e8a6a8a5a5bdfee84503cbb92ce6c14664d9c6a4ae63a2982cb47569ae27d73bb80775de70339b8baeb263b070011577cc7f1af201b5d9e6a7fce9ebaae442693a220b0e4eda2e20eccd93545567898ef0825b6c979dc81266c3c83991a6121932aee63ee920166e20c09feadcfb41aee9edbf4b04ffd05cd4cd325fe97188ba37e16051c3a35e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h16ccd66ed5cdb4f4eb7931f7f1adb956944de601a0a30b823177aa2d1c3b8ba710f1cd90dd129c0065b7dfd320dc29c5d6f53b9e113f4eb36b182161b474cc93c1e81995bd2c3a34bd02b712d7a9ba8a9fcf45de106329ab39adaf30163c3306b39fad0ea12a96fe9ee86fa9e8d46abb29989d743b1794fb1c2676994e6131a81c257d4a5278d5f8b5a39e62f09bbec09cf502c922dd8f86ab28b9fa9a0d214ff6b6078ab08cd078320b61322d388d015260d595e8db0157d8e21267bf46ed4d6d7ee60856114ee969852b80a40f3b90de73a22a08683e7c971d0a917f6732a649b7871ce1ae72ccf676c966cbec8cd381150241ebbfce97fd7aac4ea1208c34263594353a4a45985216647f008e19849fa4dfe7ba2763390222607e27f3be79a5fb582f62d92273f396fe225c978551d3a364c0714c79e419149269963cb1f1fa70628c5ecf785f3c635f8c73e46157624b4792ea919b4602a178ea4af5130ed9d29ffa0bb0b170feec7b779f290bcc7a8eda88370dc3aeb3122b6e8459c344fe32306c48f59d105e4ba9e211a18f4f1c343e3aa538a4277117827729de105fc9c10ec35e2d0e4eff6ea1b71237a364f90cf13e8155c1977f2f6d0238f49b5671c17a9689fde3f469c1e4ec5746b8ea0e455659a0d6eb34e291cc6683c81c65956f67f580df5624e562ccb3918487a62d567f26f148d56e2843913cb60d6712ccf6ff9728378b42f999b1ebcae717c9dc76650afa6b07a8adc5e4a0c8f1e3fd267f98436f3f7abbf50a64a677434b1d5dd182a8821ac691d5a066b8b23b41de1a702680b5916cb7ef271ba7a8b8c531b4f904c29cbe693aa50527aad092d98bc06da2a8727df19df61e8dbc4a2ef41297832e9c3f6a9e478b4be116caa81769c8de19bb9ca113a4c8ed32a13094c8b5aa301f30623b4e46236943c88c390cb4a0d5af865361b2bb967b7082e8d340c4a4b1b0bfabcfb7db1ddc902c1fc42c65e9c8866c7759e75a9a84919c5d929ff7b2c5d1e8de9f2317fcce93d6a9c38bf78dbdabe51c6f7bf8abff5299784e467fe2693b3c3f560fd0fab2e36b8dadfb4a2cc6da8309577bf399f1397d85955a0bdb45e4dec5931a76f3ce1f01406f0140e45984dd194276a4b613f31fa299786ac92ea0aed1c375677e300d1ffe60e5bb523aa88eb0fc221cc7e21de5795128588eb5e3b9c820992c129094540f8294b9fbb3784f3ef2d6a1f295d9a9837237ac0a02c6bb3b82dc7d410521794b1c52c8afdf0ae22f1ed97dae41923741e956e32eaca9ef40a9a60eab100c74c5040e2e379d9ea1ff9c2b37eb64f12421ffecb16fa2913285c9ed18d6d388080953d00df9f5aeb78d870f2e974cd8af17a350d2b4fc13dfbb75bec4dd82a57b0e92a3cb0bc73d8a2f3b331fc1037c397f80f5f6cab5cb479921c55b4ac642b11de832fd18a7435928bb7a32c005193733fff5f5513eefeffc164c3f0388633ccd8fe53dd6b6745a995020c0a9d486b89eda4601369677967af669e286514fa20f3b7358c031afef07dfafff979e32f099b734f11932824db3064cfecb804703fd1ae66374b854bd5e28e807a257f7c48ea6bc123910e1d8375c6442025dddefbf78d6b8ef037f1a089493bba29f3599e520379312ea1cd817c2da55d3da18e88d177cf0b467eeef10715886aaed1667054eb471e375b992d7e2de5e3bb1a902e73229f18f9b55036f48b7f2b2d5cc88e949e40802f18bfcca08da908db0d844db635583e11d2662b6db91176ac1c711fc52c59c809a6cf08a33c80af7b4452b6310ccbf9d9ed47cc2ff8380bc80b60e27c9bd7f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h77d206a39be1c5caa7784a4e28caf784b065dab6bed2b8e8a30010153ef37a7decbf50fd7ff68946ab19e4244570cb5ace72ed4340958bef1954ef14385045aa8fdd7c38c8a506f8258d3e0cbf75334f32b3f20bb44da2572c0999ef4d9e2a6eabe52a452940ec47fee1f760aef33c16a1580e659eac1401fac39d6a8fd5840d2bab0c354e875f22888720b3d1f1fe300dff7bdf330077e1059b3928507a4e884450bcf3ce75a2068094ea36297f7e6aa2f797f8254b9987cacf6aa26db668ff1d54e2a08d35ba8115a4724fb723c0c67a79f5a7cdd99461c42afd54b382b346e428a78e548d965c8dd7baa3f9451582d2e7eee1b6190dcb54cf7741018573ef09afbbd15690c2365130b605f24a86dcac295f7ddafffea1feccda079804dbe436e64bce1189d4f8a32df750ea09087296c0eec6dbc4ba5644095b04c80b58c4ba25c887c97e7a44852cc779e0ec074a5814ee677c6bc9538ffef96a4098ca232fbfb781ecedfca37b2f309acd57c49e50f83517875d19e6f8e7c947b9cb5ffad68c751ec6c39029285a1342b6d36f2399d98d67fc12f3a30619e4338a492a5f547c94ec7154398dc6e1d8d87892d7d0fcc43420b923b34ac0db0a28cd222ed12bbc9e2b3b6d716d3ee50d078201fd80f63c4bf57d305113fec14b238a4b0aeed993371ebc5bd5c5d825b740ae375d8d659c5760fddf547bce55c0b50728473bb1b498b449bd38bb35e9c5d4a5ccb4c66ad18fa3a3139134e52e62448ad3f725dcca232d63499fb3c92ab5c80f3b426330d8ac2905361383422066e0c9cd6147c810328e46a3befeb03050d70e699e7c9f59c8c031952fa6216fa54ca1f41c4a3ede07f9e1d54caa6171a730eaac6d23f525683f8dcf47ef965663c802a08a460ec75e2988081be0800021ed19909c48e98c92c3e84b560e9aab5ff201e8c5fd71fd08186588ec47d34f199b6c1c04ad66a0cfb4f2fb9f50ab2628a1dc77f98931d6225d94b13ab8aa579bc53f328a68f9c531fe5386119ed154a44f8838a1a9f540ff1a72f463a89895083a12526575d71b0d5d451374ab7e870174be95a9295c0584360be3bc5a39a949594a8baaed9185d956a286ad571949f1724f3a65c68fcd21795f925ad928149383f3c77b5a2a5c1914a2ae845eea4fcbb68bfb7c4e9d96d2bc44e695377861a62d2db4668f8a15f40db498e7c478fe92706f5f9483bc37371cea1470dd7ec036c5465a4b456f42e7837c5cef35a089dedb2a4e7e4dcd73f8adfb26afc7010778a15b0473b158393264aabbf859466f2537a473a08df4495a59a67cb378547d3ecebdf099f081244d5f174b5e90479d6e214a072c834ee84d1d2fc944e1acb7b6838fafdab4d2918878ec271f8d33a7c4b84b02e184603e14ff22b552449414a853ab59fa340932ea1478146dd727164c6154558a400ae2d52570e85ac50c3b518bef6c25610b1422f32b08a3c10c50afbbb6c7b5e4748149250973d6e64c29e3a84b0b93f0e5ea3467dcecceb34999c26e1f46fe00200f83d0eccfd9665503debc148367f5b7d82f7f2cfbb70b5bb727a410f3f2a7bcb4a216d7145f2f8fc75f045cb7a1fff6d5d52ebcb065bd9b73b3c7ccb7a23a7925e9ca075accf8f9c7465cd8b88b908953411927ac18620ed384e097dc3d520ff06aeb67f9ba2aa62c69741efda25f699bb8f90f008d2ad52b945ee2692d59e277a51c2864e727ab2b305ff789084cde7a0fb00b22646ef88d80babff4e582d4dbff7f06bfc486a84cca36c08e0d86a7f3527d0352706d499519d59049cbab1ad9734bdddef3de80adf173ef6dbdde;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h86b8b8e0018b6746ad845c9fd1f192b19e355bc50cc1921cb21e7a1fe14287c801c4511ac5b36a687d3cad725c0137ca0c8efaa2df8e05e6fa56ccbdd19a81d4648544b4950a07c5a759fa363e71832e4b13434b4f096947adb4f931736e7f4671cd21ca682ad7b0397d15b8319ec2b3ea884a5687128d1615f71f1598d36d9beb99b73be9edcac6b53d94802b56390d34f9c1245cb48b56c993fd0d3b47bd42541a80b8a42f22fe64fe346c5a326bba5874e5fc0f58601235b431848c9f29e7b9ccddcad2cea9a6100300dc06a233515e9ce4f7699a1ffcf25f4bbedfea74f323c09c8bca75280d65233caaff4e36ac38dc92720f69f117bea815ba8b70a0beab174684c684554016cadd7429026bf66c2bc5c8b2544f02223763b0f43b76c0013f3fb34bf57b90ec6483fea2629c3e0313cfced07ccd1c4ba0a3e0995c7107f2240a7410a740b19e553ae071ef7f1648ac33dd081f4c36399b649a4d73be7c4d8dfca306c60803ddf034c719279e22151c84d14b83133f9757d2de3dee5b97216dcff658ade9fdf43d69932f98243c973fca7d9cd8aa23d18b16f7c29307ec5a4c841436583b412fcc379e47d0ad474b4ac78f0fec54b7f07460dc942a514060db8c4f54cd2765b55c6bc87608c95de3d7e61d1a22097c4cf3af51e7752905eaac76305978914b57222594e9eba39d133fb7885070c08e0af388dc3ae14c49446d8c354b27a3e1e8c639faa101f65a652d1332b1e5b003f664ce8d74a97cf57071a4332f55f867e45aa684e4f422550ca5bc76bb0755f38e3573dc18494c237f0c4612a429453093d7da8bd36325c31a0fee6c4ad508c7c3f2dbe698b687c356b9e06e97083ef2c587dba4dfab2f094faaee12091d7a5bf887ff88ddef1bfd103cb664ed71fb7aed58ef05ab3240b091326bbfa364c76572ae07b3990a51b25db3715a24677c5d60f269aab92b3e9793910f565b53ad93faf3e785dd188756dad17ef8bf740fe782202cd8129b5c6dd26064ab29889487f59fb20921b2d3d2c9513006fbb4740a3c8bf16d59a6707ed4d97568a95579533521bf6097e7bf5fbecd96e0092992cb6eeea05b8d7ad897539ae64320ec706b8489de02619b8981e45c5a367adb2916cf3617bd5bd768a21fd9e7992172223fbf5cb1067bf0dc5b84b7682237ce5f58e903eace6ae981c92220ac87552d6df8c588722e6c7dbd1330fb59ef2256ca83c967f77319f4f8f75ef296efeb4276592c9a745fd21c974cfdcdc81319332dc46b575261dfd393052bedc72fc48c92528c2bfa32d805dfc3ef0aa58621a7d071dc07b38639610270bb9153fec8c2959aede6d4291159f3923384b352e40ecb06d8f2dc13b9822aa7b5718d00cb121ca49afb4b595befaeacbd3bee57ef7adb75b38ef0234fa792fcccad1cd3d0c7f6aafe7a18adddb813d0b82bba45f18b5c9d091e39a8faa79f685a6dfc571135a6df6fb270ab854c3ca2503593e0ba898db2f8f8f7355322190854579fba82851cb59ead17aad42064df62a0f68c8dd555654ff1816adc131ea414fbe90f073d1e1727e5a3b49396a5ef1d37d75754546bfb2d4a4752473b90639755b6c460887591e71ebd59830650febe50445c64a30e82e43f54978945e1c8733c7db61f6af8b3da8a63c7e30baced00f7b972814decc0f822740078571150b45963942142f4f988a548ad50100ff891961dd68a431e1194b8d525a15b191801f953846ea638ea841721d98617f9a91f67fa1c43472d3980f81d1cacee22c73040dd63884d6e96792324ff6ee3ff2b9efbf7d51b6c618a97d0d9d6dcd03a41;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h9ca5c789cdaf58d57489bcf318924415774589a1d9142bdce29d4dfa90365433a8a97ab877ac08d9c4f4db3b14094004a0bb2d36b11411ba3c7a48230a8afa64819ab205440ba7ae51cfada234c17b749bece6fb1f096ac00d73957b39c1b3b74ebdc7b6f31571b4a37b2bb66b9d2485fb5aa42fce97537fa75c70151b7f13e2e84ef2b70e1d5f04f274a8a05262e0442096d30f0c1f3acfbb64fbc9770b4b93cf78dd6c3ad0b88b0c7b2982dd3c6bb55372cadd61c6907d3f361035a3f46bc9b1d8a0966dd2a76f073ce3a2084b2f8e1ff57ab64d8f01081d8ea113af2379e07a760ba1bba09e3c7cfc7ed654be354afcbc027aa6f7df543b473fc6a144fc387f7d8485850a0491defc146c159874e921f89fed7b4669b5895dccee063631afce32482f218ab5797c7171b5d60d8b35bea86c62bd82e5b113d199b002082fdcd273fa2101967bf817a71bf3c43fc1e2cfbdd2e7b2d2f79bcefcfad7e907eebe531e19ffb91dbc8ac2378316f7f83faf3bf958915c5394c4f88992ad4cceb3f3279b47e3b8ddddb3143e6eba13357d121893685e19aedee2c19a3c1f6ad6b3a259bf0f64ae82e5f26222cd0044d0b8b766d27e0dc5e36e2b767152ac5d6194a5cdc31a3c40facd86d5ea24ad7fa12f9165234d6487700e06e5ff169c1e6505c8cc938469537f04349480c05d0151e0f08b0f78e15a3c81f1d98b3754485fda4456b2b51e31caf847a09630de56082c4f2ba3d5cbef1ca4af2537dcadae57036f0c7f973e01e52b65b8b22457d67790433fb825af053dd0a6d4d1bd1c64125d7d15632b5e151464456a66601e13c345d8ddf0da09bc177851d6177dd54d1f101ee323bb67ef671c092e60a0db42a34414d5cab0fa8f6e323a0a359d52ca746f1b9cb7bdc5c824fc2ce07d2f9f3b3445e35f5674e3c1d0a7caca0f05d7374d1b8b80c2a6a3803348f67e5b11b98412bde51645ea14c09b7b6451ebb94a76af56a3260a79abcb8b03b0f98b3f44940b743d00556786357ce884a34d97a809d0bb7ee3d9c5444cdda879528e87944a9c0490ea865d6be20ef95e67680913635f65582fe54ffcb8ba4727a9571bb23b0a42e706479396b1bdc511124b8c757ab5fdb6092788ab9d88091e1867839d3531248f10abd28d9dc0c222dcd51cf3126d95d00ffdf508167be8109086b84b9d82b1dadabeffb375157b5526d96aa795d667458983753a7e06403a9f685c4e6a90eca325961ba1bdecac8cf289620262d55f7c98f2466e66ea3d92fe6099b2cab92243b38864f74758e28f14a9310fbb3c2efd0b236fafea2fca861ebde991050adc5ca85f234bbd641022fc15ce2b0692649b993b2bee055ae9c97004d77a7eacdbd987543bce2383a54822d4d9f3020d8551483b5ccc49e654ab157bff71482fb0831efde47d5b828a731734968da049dabb610f2d51f061a3c8a1831a83741d1e44f42dbdebe122939cc0db05836336513310d9e20f1ea7be3a48e53ec7d06867cdeccf5ca51eabb02027a9ab37a60c79aaafc694c39a6546e109e1629695d53f37a0df441a8869bcb31d8487a305302acc566e02d5ab0f6fe625db648735cfbc53e51d2cfe5b02d8d51c86b1ebe59a77fbcbdfb49e9b8ce3d2838eb593dbf7f8777d9362595bb1e8bd14f37b801811c8d3696a2cf714677cfa9f696c532c8d78e3f8fcde2519d9e0df132d408e0729ffe4ca098a408a24dd836b85792acce24bce05e3dc037bb526a4a738b761b519a5782671be9190302c4dcdca1ea1b59c5470ae39c1b392039a154ef1a1b0ca6abef58b641524154fe57bf408cf70cb139d4e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hbdf0ad578d18d4627fc88e923bbd72dc455bddddb91f11759c4c05c3aeee201359980a1ce4150a14012744554cdcf349762193ff69fe9d355d57cb85e82fa7ca4f08a7029699d43c577b400f87f7e875447a988e54d1a99f11a70f360c00f16d5c7c26c8c46a2c89010293cef077514f335971ca481598d047f7e062bc18c3441cbd6a338ea14b75a7ae36efd058255a89ce3a4bd3fa346ea64da68ce155be268aea231fd84d2ef0cb4776b55a2ccdf7f371bb4e87f7b804a9ab4b445e69cd0eacb981d4bb39e977313fa6c68c4796d2a14ab24dd1270784182894812b72da92f7a7ce2f336f84e0b0e76c27fd930c166f421199e869d6b6c948524f69f9d045987d29a2fe3655b88ad55b3df1b04ec05236908de7acc1b44831e50fca4a08d503dbaa6bee83742ad2187fd6608a32e647aa9a93b6e479c7d19fecc26aa4b80e8b33019d6c2763b9a3dbfe02f22d13a884ffa11ea255408cad8b26c9bc3fa10b89f63c319927864474193401426ab6465c0492eb355321da3094d5597e04cb3dec98e10879cf30dfd9b16e9c0ece546904b1ad5077710c143ac8ecdd7558977d20693348af7d77cab81bb61efd9dff6c1ac3551387679d083c0d0a8cf3347d6716db5ab108ad23b67417e2729238295562ab26a60319f5718cbc783522e05ea5f2615a229c7d8a0647a14518475e7e578d6405d28fa7d8adb626bc3f9de8add666fc9fce1c3358943440f88337be116a5476d5d591484688fa26abb9fdc038b353475aadb60323a038cb0464320cee5c58fd37c584086b85e5a603fa07d3445b318921edb3f046419e2b9b7e98f18947e31bd3a26a9e059c6866c731b87205489d0aa544ed19314ae1afcac233dd0edb2db53769e0335c75d5685d103b40e1a636619b65dae38531e3cfc40513d3dd3fea863f4627a426e5039c8f92456145bc86bbb95a14b5ca0929eb048acf1399fffdf33f94b4b5db0c172d2cd63c1e63b91d505ca675aea350073e936d04af153c54c703a75aebd0e50c73e6d2b0f7fd80e474e064105a7697aa6f42e8df5a436b265feff6f9b831cf7ccd961fb1d981930ac86d8d694c5dd48c0094217a3e10324ca4af13ede6c9a769f3206b19d2b7740fa5c42285abd427aa0ca61ba8dc8790b2851afb8097fa3ab5cb84671a6a476fecb805a442efe3425071c47ce2dd0f1f0f8c8337b6eaede4d249c3c1aaf652818717209e1a4e56fe9b039acf4a79b75e283c99a4e2f81e6aa16cae0a39eb82dccddeb695ef201df85f31f889b156509398dbfa4135476fda00c75e86a684cdd11e3b7d5d36911aa85f5ad54cb93775ce5fdc91eee837f9b2ac45eafb4f07483a46bd0709c8586def7a7083cf96bcab896c349dd52d69cd060a0349ad15bac8f70fef22f12518e1575637dbd9c5ca4f8a11c7b661303ab5114fba73a53e69aad906550fe821ad21e52609e6b13b8efc3af3754ea7b56007c33cf747f1d75c6bf67df36b6f9a104a98d08c74dc1b98913565fd4f424fc91a752a867565b4728d910d9e12360b4d1c962e38645362f8910c29712f360e94260f47aabf2ca4c669d6038d3fd39133e43f5e5196e6689fb8456634189e8dc584b163a0b381d2a1452947669a2bf1f4130e32d736d26fc8f8ab3c279efdd14b07fb33ddf0cbd023c6d757b988b6afc1ce0edec697ff629bf73d4aa62edf1860f49b0be38305d32210351fc4ceb0c79acfc4f88387abd9bb7183254c3edbe5d24e94430cad3773ad24e95684c0457cdaeea6a07ecdf1b08204117d594210ac935057c6b20e5d6a65d95a45d6ad9b932184b3322b02760a356f58;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2a450f8ef84df3057d61c227fc6eb3a1b4819c23f3c3fc468b6603906346393093e1b57110189067b7bd91f42c4526fe6a4ff3f139e5a7ed4418650cff90643dd0e7d4e782373cc3eed13d47d696799d01e3e24c5084d5666db70d8d0a6b46d71581641dc010818b4295ccd10060fa9742e9f2d71fac1b0ae0f9a06f09b24a0dee2aec6c8972b09a541b28eb666dd0e7daf30a20bac5cf5ea922319ed04a9089556734dfeeb0d9bfe91e924c756141addeb31de8f1d8398d204093cfbb77d701a4caba9ff5fbbbe73cf878c7a25495d6c2f75c005ea4c5dddccb4e717a8f4b5a73276a53dd092d467b9aaead26d205331b0145231e192de103966d339c4884087abcb92a125e606080810a39143dfa39d6ce754a2708065d2845b4b0f860241b14f211c0a9d5886c1a146b288cd3510b8c334e84fd441767838f2d58c1d56bd83ee53a99ed9a0ffae4ca4a432f8cf74ab7e0bf75b2e7882190beb3e9dd7413ed38306bd646236271ece1eefe9c9390b118c147576f02a9b1dc22926ca6bca33dbc971a8525e6f4dce098a2dc57e68436675defa2430a198c4638c59d164280c284527b82fdb2e721232ff8d5cfaaad71d4f6bf21735a0cdeaa78575bf2fab45828ad064e79e858b209b024d69ef2c613ccbef65a8da94772d91e20eec650098625560d9100a40ef462bbd1e6f5545a2daf33cb3cc82401b11b2b3a3f1b8d0901907636c3a01a7f55a2f2270a88aef4d529b0d8fc9ef47708c20ae03ca5c615a027217a4d7aebd2f7fbb72cee7a080c5ade1f67bf7799896a5f0c8cbe9626fb19a0f03a1ae20e652db3b908946c91e8509b116ac5c2df1f03d33acb4f8cfbe1fb862aed3a249215e9989ae8e12515a69eda060e8d8f5cd1256f1c816af6d8767c6720626484303667b0b3b90216dc9a7431d6fd8572107caa3969cff2ba01e7a900a2edb5de9d61fed979f59bb11311cfe41f7f5bab1039464f6f688d1c6fb8f6a9404e2ce8737087ba959f5d8244203d6905cf39e3f4d8380a769cd4ba13c36383f58a5ba6eeb77ef6fac1783c8e367b431e9adcacd05adb497ee4532d198944a8a1f553a1b6614b18d08716468d1772b224a838546a68d04300dd0884ad9854e6c6559ac8392ea72ae0e13dd02cf320d64e166267d91535c373292c02ef3c86a43c2dc37a316617bbda1c9166a10362f62011437e9cc925954d342760888f3ccf066a873cf648ac0c0e9b69f2b064395afe7d0d19cfaaa996d8153bbfff2b94ff58cc63468837a4bedf18672b589b27db419d82e462329510992454a262d16c8bf7ed75d639d56e65ee9a42aff5f338d1745a8a0d23c4972a04649effd6f56d72e6fce57cccad823b7149cd7019f7af53e030eebd26d699731991876f8b6f272679acb17410b95a3c1872ff5223cf8b9daaa006c62a6b26bac41d072de7271c7acab0425748baa443d02886e20449a4eddc0ae85f1106324c4500529579a98833f15e68fff5f06193977e62556cd0830d7e574942eb8b2c44e02ce04d057182b8be5041c852645fa887f84424a84072db76582478cdebe17ccf9c38203160d0481b2f16d27e63575224b6d19774e822e08aa5f19683de197a440bd7be4f71595d3dd375715d8fa37f69455109016387152b01dae004598db862edf7f061131d15ba1d4f9c9b61b5476212c1a794174c18fba13240fbce55f8e6adc88ee2c613b420233b46381ff398e53660d61a4c605492c7e4fdb81f1d19506139fb8fc1f94b4a5665073f078fe796b90e00d92d76f401b1b0d675c30a143922bad2812cca681b3a835b172499db4faccc01723977;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3f28aa82301ff38ab26e5f6bef77ea7557abb8d2cc518fe4495ae795a33c688327d2cc7354a7d8d597f0f1245b1af776e73f94e29306dac5e18873621fd7ccfa8a9a9e95d375c718ecb32a25fe435d851d7965cdbe96bb54fdc63fcf4181c1a85e11e3bb1ed65f344070deb041f79d1b6d10b1c80797d0413b8613bdc90325a018936c2bc4828903fcea822d1fb5866371c039c25c782b038538733a7506a9df06ef8d0374a36f74f9cb1381807d7ed44a5ee0661ee9ab46d847b6d899fc881a6e18ac48e115a3c30704a3154ddf0c46f9cbe50faad6c359d1f98a8062384a243b76b59c79f562c3f5167dcc7e394e689c9e4a440cc8912e5a66640fb768676e7675da542b63c7fb2029f9d7aa8ce60558da0115db1a8f4d764a3433af5b3274a63ea017a13fd189af29fa8708b904b30733400744aae6290a171b1ddf8bc5b763284c2463bc8ace250cfc1b7f3e1d40947ecd37cfd62d187c2910568370130ba4ff352ee0130715f89d5da7b7b931b345026303544916edc8ebcc78f79f889a71d683fac5dedf864c4ffbfde0e5e1402c827d061adcd5040a48b2adb117a13a4498050f8ec4e3eca03fc3b6f721a1452f24b7a1f368c60492e71a87df80aacb31471ebc98015f5e3b436f3dc8ec3dd6fd487ccda3aa6f9fa9fa98d370d00840f7fb208f7349a1c0373de8f7ace6de4118792b8e53ffef95392cd46b119f9ee2a4e015b25cdf74479684e619a8268f6f2d9c549f231cf865bb3f73e914ab4b7fd614665cd748301d82cea63f0bc7be89729df6df1708148067844cf519237b92fe1c52cb6163f72be44c45e3c639936c85ec5863090b14bff029d327949beba4b57e36a2970145fe484e4b85b36b2c72a2c93477beb71e3acab8c25265c9cbc320df67f603aa3e6cc39302eafa57f79ddd59c200b74d5190590e0b33fbebc71790905746386b324af2a4bae5f1c3d9915a6555b4f1ae8ceac45a2a87cdb3bf195d62c5061a9e6de7d63de3a93f42ccb32a92e535c9832faad03b24cd03a1d7f9ca19b624baa5e0d91233eea71654b4e6fba260a365a95d7f42a3679e95ac872fb1e135ffcd6e0e1454dd18795aa56652be6af840c37dfc7d44acf2f1deb9611e902716ddf75cada9a2f46e42e0efc8942cc527d6578deffa73145285e18cee11d675230726ddd24ed2d75f320c01f3c25f80fd84da57a9ad83ea6f23334dfed62c8b7c802bc065b5794a7ba4dee488d3627f771134d2e8ce2614e3e7d1d4d62b88832ae3ecaba91ce85b80a4fbcf6aae52042574a7770b324ff46a3f379cef05f63b6c212a4d5deb96715eda5b3257692120d794cd0bf4f8ea940c7ddf19130d3b9c61d56ada78c4ea6174dff1168351b49bc2663289636db0e3498ae74e7c90cf30664d21afc808a7a7902899793fe9e2601a484113472762e2ecca619d7f008144750b0c2b9409b877bb00d3e1996895c7b11e654c14c0f64b62ee40f3e70c719948f60d00691a52ad7e10ef4848457481d229af6ada25964ec48774eb7f1d32509e9417410f482d2f6b37fe8b34ee8601f4d867c6d26e0eac5d87a1510ec1ef8d4f4dc3b0e222990a2301d18576eccaaec6987f3517c59e1dc105d2d781ff1bd0f4287a6c2f62c6a7b42c352cf6d74c4d972ca9f206a8f08f4a92ae18b7099a90830e34e81c0c0c99bb5c376549a9d2d0a4e07261f2c9732f8677d7cfa91712d216cf446eacd40962f542fb17c72fbaf0c92c60be31da395ea7996763459a0274cec464f35fd1d7da34d68c1091b03d1cf2feb3279476c892cb23008e97d89e3f96b25a401bb34361ae3e2a785f00;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2570132c9949fe6b40c97ff3384a3624306278268258c8713e1546aeb4a7bf033816f1eb841cdb03aad80cb53c3628c923ab27d4cd1571586e8bdb919fd0641c9b6d102ade1032b473345acdf619886bfbef899476136b50ebf36141d3329f9eeb6d7349fa23eba1551ba4840958a48ae72efefa72c0582ea20868ad338501f14825fe09dea8fc5633f68aa630860ed784da83e772d217f5aac204b3e5b6b051ec661ea9ba4189d4592886f58844094d61ac8d8f03e3c4b61f5880c85d00476d9a97b0720546c287b5404b2a12e5e043f3ed7b691e22ad0970f7494bf9410bb797431072a7802c4830029ebeb8f19713810e386d5578a59d242854e838937d3699b6a24df5896f3e36ee52515a34269fb0f0fc9c311f20af8b3f4f48497069367a33178abfedb6a716cbc03d4d6b5528f773d8991d27593ae0caefdb12192a1634fcf93fa61dfd8394502c6d459166fcd63c812e17c9d8133f8387b1d8cd652061b1e396ed1defee8494ddc5a769b0a21d30330aa632f30c9491cf1b2b59371cfebfd3f2507c3bb0dfa9b3c2f2b340aa740c4f72bdc52469f563b5dc8d5d4a9ad9bc70645124da9bdc3f6ea5ed54875d090e542459e8f6fc555de097495221037318496271c01136b15756d0757e38a627c0ea0325224891e39dd46573c75dc02eb617213e9304050667c49d0d20eef29b3b5e25eb8dc79ca9a1de791e0dac36eb28382fa4e0e38a70aebe9023db5494130b86b2e0e2b08f1832f3d94a1a479c1d58b3f0d031fa593d1396fda754d9b30e039823bc9c1056fa200974a09cf0b07c2ba0e3eb8ce01354f18e0977f769b454e8b7fcc81c0c8fdf509384d2c13f57940c927383300f71533ca9ff91b4dca0a6c359312997001eefa6d5aba63eac60230a063c7d7ee4b8110c0b115bbb8d37b117dfc00fc18d9c745402a30ee423e8acfaea42e6eab726f68d904a9a8e39b8aef701664dbe85d7b886f3f4cec23bb875781c6e50eef6520a409ba210a136b2f4375648b7ae87dd84e37acdfcfdbc7694062dac271a71f456109e39ec188a567bd14b8014b2713f111c4f7d2dce1299b3243fae159166d03a108c14e4197885d9fc60f19dc87475c85fff89ea990d10137e2070759818154b44d38121a5212f81203d44aa7b3e10b4990dcb00dc8cb44c1ccc64fd22b8da7618af25351e34c568a63e9e7b11302922285d3db452372bf75c4951711129397082a1caf4fd8ddaefaa90fccedc71eaed88d38b2e1f0fa58d4f8c83c14dffed7b7805679dcd28f73178bf168f13c466f8cb10259c62b3781db3cdb028a876fc735381d9efc42e5bdc5d49668dac12a080599b21a248f7827576e1e19e086194c8871eb63a97a58df8929a077e33be598ed2928fe045923d4a90734df6c6069b37d71dbfb519576e1c7a9d78678b092f81e44cf00296d3a83195e72637e228797b40323cd586187f57580b12c1f42f88295b7319d9da22534e969aa0d0e3e0ac5fea3aa9f838f38a35311de30bffe6bbf53cf41b389f61b78ab90c2ae9976dcf232a7b25bcee19facc64c1cd57f43ef03de11bbc9f59151f05e071f111d446962a8704f4e6e6d0de56317d33666e83e55c5c0652f70652beff0d0176da788aeb87975379673ad1fdaddfb7ef37fdc9339a99be67c56861086066d88570db0db191f82be0791383d945f0cd550c57e0588cbcf57fd0982b249875f128dbeb4af7b369044c10c1db0bf21e3a4411341febdfd88b8080b63c31cbab3da191f23cb17b0d0591282d82bf91f3615b17e34f9f33eaa0acafc9c3e2c347d03045340cfce4762b09c0d7e69f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hf95118e44fe0e4afd803fb114c1a5a465882eaba6df7a0ac347eabf2c463d356244579c628612f52aa88497ae815dfcb80850b43c6bf6054ec5d3b4aa1323677b5d80f9d1a82028e459943157c92e2c682630cb5d2d33d6ed2e6d4ca0016ebeee9ace834a9117ff260cf4029f061761edcc02c80e072e37373191ade3112d0ba4337146726f02d2ecc6a5b5661fb45ead0666af2108caf41f8830b775c3f9f3c0000fca1e866fde7c1a458bdc65850e4f482043a713f5901a8847fe161083f72dfb6afff12cad8968b675ebdcf4b8404cd38cbcdab3dc9296e89c833cc71c74b71004f7e682e27c83299841c858a0c3a42e925965013e3c04b0cacf6edb30198b18b5afc749bc6df01b19aa93809949345450c2cfb5ede5a89df6716aa510365b54ead178182a0d45c1f613a1ab03c0c51cb8c0c1c82670bfca859b4bd1c4af937ab053a9b98571e8d90ebed71147b31b21affacef735e846f6719d518548444a7dfb76faca918a45324e563b643086312c405993149c98f9e9859dc3d7f2dbe1033a3b2e530282a97a1feafaf75bd66db4b284aa10f8c236b205134e99d272ebffe04b33daf059037f2f12c2c93e19e8039e567ce49d25cad870ff90c30bb92acbb6b2ffe514bfbc98fd5dce6840e49097dd1aa5b7b28855d23ca1fb4980ef50d2fd699ee86b990aca6951c18fb7f92ca60906ea2169b29232c9eee7b34959d4bf32dcc3fff12c46ae2c4c9a253a2ee440a9fa77df697ae36a88a00d523a2656e2d91147c1906e0c7b1616e471811453c4ba3bf9e5f093c923bfba88695ddfa1e88e781695cf643f91890beafdf24986cbbcb49bdb13c718d55d4be50c396118c0f71c09d65a1255fae6d574a6fa2d4f7d682f11c28b22f6ae75cb960c241cf967511da501da752f2f6cda5ae743b4949f0252c4eedf50e3884f9216905a7ae1c859a1894d2e68a6e1876029d7f3d0f177f9569dd3dc3e7fcaf2f6e72ece239a5f70ffdc330b8e6be3d8e2d7ffb507c4235f25f699a9e278eca335766f5685aca129bee316ff3795b98ca0bad184d5f4f8fd8242d5e6bf44db73351aaf182994e17d66c9933f0d7b9ec81e101ff1d5d16cbe486ecb5fcd78c4865c683ab9c7c40cdd92e14c917c8f947ea524b2836eb14fefe0d6b55086fb5ba5a9792fa81d8b8cf8af2f1a3b705920ece89d1d9cf686d39d9fe1ee359b9f6274ceb0351e33ff9e0d780fb9e179ddf6415c96a2242951240e2c0b6d7b9e6f5de6641c15102ebcce86bc6d5334b0f0c101fb4185fc7880b9611c164fc9e80a483f02b9a166299226081fae34dc4e9c6967c39726dbf8a1a3391a13395d16795e4c813481e95fc13de9ad6a79c78e48e916a404e6229eea765612272f087683980d8028818a3b4c4d0f4896381b05badc4783261fcdeda6a5f24d75ed1d24176a7c4f820a823d72e2a5110e1b49d4d2e76d30d5fc91175ff8a89a99d2b6063101556947dc8c42142a251352c4d0e46a44bd0d50454b49d91d643d13f4de8b36404173cc6d7ccaf852d5ce2cffe116fff79fe278100f63f9e7895db31a20ccf646ebcc5769a0932d2e18f58585fbcf8f21b593960391f223d7b64c7d88f607aa62dffd9cd7846c13b18debeae3f77a062bfbd4c331147af192a35a14c90081464944b05457d3b53fcb9c4a13a136fac82f601adaa5ae0b94897ca528005712e839d5aa681edeba0a4ed8a0b140a1ac8128038442ea9368e6c583eb3496c37b92f30f9b47ce2b96c18f84494e73d41558db5d0a9b5fcf924202a4ebb6ee5c24197e8cba1aad76480dcd3cd54ed053a365d8409e7dc51a294;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h5c338b397464d29ae47ee467691b4f18313c9c97a7e9a70057c5993fca834672b777f95a26b761fe9a1f87355c1804fd0a089d72543f64aba233acef5b4f97e1e181d410cc760b6630cb3157098b2557baf437915e8f1d9df5d200c08b35fbdc61c75c0ce81e39a84cde58d3e260a99316ee013b887bf73ef478261ffd811b1aa53d642cab3831bef7e7af88dfd07934076efdce5eae576a9f3d7dbfb9a007d74244ac7bfcb20406ae421ab2c0ee90033ca92ab2ddbdb15349aae56f943cb479cb4609175e9b29773ed23ef424f3a3bec54774e32321d6c15387d05a12d2fe174be274c4c02063256a8f8c672ab27025bbe03974f7b42c45a795f81e765e04670b5d791fa36fe278948461dcf5edf48734b11eaaeae151dca0ec5fbb298ad9dd858a2af3b4b08ec31df11d7031fb0222328573b5603d27d13dc7e515322ba1e576669034abd7e3a51e2f424ae378e54fb7bfc1efbafc6c84d5cbd14fafc98f76b3866abce04686169b3d32ef23ca465f729ffcc2542af577e6b53feca2eaf08d2737d40f2acf668ac1593e5c7dd94bef0635d428d82a898e8bab8fe97b730ec1cdf5bef567da117d0017a41c61c6fe0a20c3bc0563fe679430bb6d91dbe35d2e98f37ed8c754a13c73f6a56998bc92bd3720e4888857f075975fc7688d10fc734232b77d38f03b79b8a9094f2696f5b3260d4b423817a6cde16557a90cb0ba6d801237d8924ed15a136ec152f5baf215a466faf252fd245782b0e4470aa2016a5a7ad3764f315d157ed88c6626ad1861647455859275ad63c019831478ebc8855b36f53d78d56d3b77d70b85081e9951b97bbbcb159e5786e3b4f42a1f6d49b184a365b15d21a10df5098d78ad31017c936782161eebb4579903b658796a226f9e80340dc8fb2de7c982e0a191bce44bf666478850497bb599b59496a242d7b41361102f1f4d2dc181e3605cba5309c724a9be15cc338e5b5999de846ea8cdbf262836a85b74ea65d978781b8f174195e5eb113e81e0ab409b1aa334ee8f39eced24a60f1885ec21106e0c752637865064210bae2f409192d8559765eabe3922aee3d940d6a755785e0ddd36da08ce9e2f1cbad3bf161d60550ccbcae4fe9b1a7dcdb0470e429154ab5bb1240726de8f14a8daf14e8b3e4751cd5e9cdc16c27527536e908572913976edef7d4784c122726619933529f3c95be7eb8382fb7fc0617244451c7740dd35d307b2cfa7088b9221b89d09eb2e4301f67d6b4024ada0b3feefc07af3ec93551eafee3a342139d9c270f8dc07b3de9967291e6979461b383fc91306cfe19adcf611f24a5d0b48cab154236afb74346e5c2fcc3b24fcd6dbf5546a31c5fb2a5a886b50e7bd32fd2f218ef32ed6500cb72584d592320a2bf972f0f8dfd7d0764df06318b544501d6986e207733a44487e34b5f46ad24a9644e2185c8bcc9fe59053f3ab4d00af08b2398c3026b3949c83e5db12775036756386fcff91927448e0e7cbb0c13a5ce4bd5996f5ca755e89b66db46c3f843c71b2ddefa59ec4974fa1e0465d625fea4446a8352e7bc17e602fb42e853006c01734fda9c9e3796d1183f8f224d53c57d8082939d3645a12d4c26860b75c13ba182178aa533aa8734927b247fa4c4b3a4a870b014932c2d7481349650aa1eb3c6cf241b8f1e6ad22f0d2a8921798a166758e5131b3820d1a1a4e7a7cad2eba12a0322515698eae4e6d9a71148e0dd5aa4f6fe9fdcd072a4139f6b413ac998a7230ada9a52a27f39f5a0d20939c7354078fd52153f79f7f600f3bbcbfe13d84714b819b9573615852eb5eca85d76857cbf5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hde151987d4091809f342ad0126d8c56f20bae104711f0af46474a5a0a8844bec584be5026e7ca94aa6042895ffb3b7475d34118d9fce5551a2624ca0dbed6cb898565bbf85f4a82e74045549d675a3ebb06ca56d7b80289ef541c16acb1eceeb17978fc714cdf25916d03227a7be099e040be69ddb1742c54b425114d565c255c252107acc9b35f00e6e2daac7074e6f70c88fb8512ae4a5ae6743fd7c3aabe6f48093fae62d42eff934685edad4e51351563423698732a42536ec9131b8e5d671c204565054894fb97b939dca95e27bda85ed91613c6580a978f6f483b8025df559f37bb0ea2ce08350c6663292679f11272c7470075e067da3cd5d6306edc6aaca5e3851a12903c15e8d3e8bf391ffefe68a6b241dc6691efc76e4d1710e2a1376cf08d095c5e6aef3643522298cc3aded69eb3ad125650257d8b64935adc91a36b6a7b80bdb0c8afff93dffae42b70a4cfe9676aa41a647b1c115dfdc60cae7e5252acf5bb69121f530cc5959af36adbb478f2194955f6341d5dcf6c119390d52fc075e472d80dd84da3e33005a1b1ff30cb7d00970897c327da94a1b77da8833dd3cd0afa8589c7c4f6defcb3f6036da80b102248be7928b4172fc6a48390c48402ee5748354c0baf8da8a4395f76952ec40a9e51a91860acb6644fa25e94eb45d12ff2cf1cff83c5dd8feb0f164659c45d087b9c3cba4fd56a196ea015ea4188512567d59c134d89461c431927cbf3267f692b09fccb952108811afb0a67981e7aa8bc24aa4eb55a3b57cade63a66797ba46f72e09f8efbfb258e5862caddc0f5495ccf28ae4ba67b948ec62f86b0995f85e3720fc8fa7c0282ffd55f5ad2de9789be7d412fc3f94c2b2a9b0d2e07669be4241aca101944a09e720ca5f46f7194a659fd348ef1b22ae314409ce825b382568b99ae19394650835da7da7a8d5742c11cc4a2db7c433374681fcb3b6ad3c011f6f1cd12e14a4cccf7b0890d1a1f93a585ab43be8e112003cc32623424dda3c08ab9f69fa039f1904c7fc3d595efdc853a5c3fdd3ba6acdeed03fdebd11a5cd1ab9e65e69e1a22cfa0c41b5dab65aea09b8b61ce8d640dfb5ab6f9c4d7642c97b902a0349fa190068f05035a490d10ba5dd48e1d1659ce3c2ae2bd0c6daa095927e1d04ae2ea196aedad20b50eefc6eda6657baed76a896caa9b212d9985d9bb9f12aaaf6876b05b5fa7590b211c5670d7f331720870071716ed442897b66e8cd1a9578cafc2a8d402d714918fabf359dbfc702f9049e152284c7a0ff9c3535ce433080e066f810756de728d7c1e91fac1547818cd3815e077a0a63815f82fb65f9dc828f2d288a62a7c3b1f8dd76f7ec50b571388cd9aa3f844eb984110c03a53e9e22d2466488785dbb1074287c403a1a6bed02d85df53a24bd2c2dd6650c32250007ffd3bc72a37000c137fb1fcb40a05c80a462ef880bf461de9ea61e9d1d87eb5fc4f110dc8cb588c1850416e5fc23af531250e5773ddbf673791e3f183a87596c464d3c804c4caeaba118f179461b6e6ec324bc8e973f126ea9ed37e3382917e370f150fa67d1854373263073b2c2e41cdce01fabef6e8195174768fd571564aa38268a1b0fc77b9ca374149e40a70902774ab3f1c65dde850fd407cc468dcb315ba919fb4ee4aef70712778f1926902e5135ec6923af1a844295b0fceede8fce5a778692604123efd48c7c54b651a1a9723c6d96c9dbcac5090863aeb0f53ae5e464bea508f97a663dd1b94d426f5b67be9977a64f0b37d9ceb627e580f73dec2484ee878e61eb764b3ea7b3c2c478a6a1db61379930b0ee4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd0b2b28ae504370837c42c7dc5fb616800bd49579f1b9514103a6e00ee17b15f5984b11954fcc57205230f5fdf0f4e54b46e193c2b2f8e926c939845bfdc64db89bb97ff1e57a499c2525f492a59c242720750630fdada0676e55c7e5b86ca7f8e394e6b09b0e7b4b578ad5d0fed00469733c29ff20b7f5eb7a3489a10446865526abe51e25bd4e31f7f1269d90f5a9c262db71ae00a4d4c6fb5ad2e4e2dc8612ff5cb4ee1bbb4df84e1eb2d58bde7bb71f8627090fe0386695dc1e29e0b3cec8611859d8d74e00125f824f5a102726f50f038e0fc1c62e1741b8cf5960e0be5fbb425cc759e1cd217e43eb965fb34f5114de735b0358beddc31637ccc6064f294522597f92b558f70e213ca25f4bd5ae0e8a203e5fab8c2f83806fb0c938ad933a22bde7d8d7ebd6cf572a98801b1f926676841d2581ce7f94b4fb069c3a7bdf8f44cb54c276f4c20982bd1a8950a2378311a1d9d7f021adcee90c2e5ec4b4d6d0bda1771571e1b417a03be0b0e91a3c8a92cd870c5649ec139ac31a5b29e17aa8f7ab1a1174fa8ef0531dcddf58eb75a5b8f70be2b6f55a0c053342ed532c567154f17b0dca1c821ad540c72cca1f0d95987ea1b147cce5f9e3bafa03c79e47d5076b13aad8bb601a38e807c2d557f6443fad298e3325ef1329b2c6df9313b726678940fc399f53d9211d4e99c536c32ae742d5550b2a01744990b3d1cd8d5decc4ab53b4a4f9f6a76973df1ec49203f61256c372f516004c7dd46dff6304886c5dbe90f924a13d4098efa49602907ec01e86ef527026c78c395c639b2d740123ac52b1a5dc6f9402d0a7681c9b2909312f2e54c4ffc762fa67e1bb90ae2ad64e921f4b9b3126ed03bd6c3f7c1968dc47828417722813e511427056073be67d2e546f8690695f32df4dbdf811c07d81267df955e8b9949fe5fa3293f9e178cc4062c6c9f1980b94049e811661530f7825f42507cd9d90e3d9280967a7e6f8dc728d8d94e2b0ee418d209abfde66c7b5cc9f39b8c4e8ad2af4d9b87c1477bb351da917056f18e8df858c4d6f132f99d6f2ef8d6b300ec80705419e6acbe7a1432163f9aac57ca2175c0d4b1270571224a6c6e4d8fff097fb40ec12155bf32f2bbd4e73b2b95b34897dd41c452660ab25457fa7272ebdb0322cd209c235a069ae65d55dbf1a4a07a4f493540031a70a56a55f2289fb78d3dbb519f27b51b68340ac8b5f7e36b55fcc94a3c6bfbd9358ed0d3f3cb6d3ee8d4ac30dbfcff12c06b22d76739c3e9ae538bdef6b152bcc26bf968df6f46d5d6f53ccdac638c25760d1123206fe43a3174243ed67d026d5f24b95dd645569224568eeb392158167a0ae3a2cabb0455e274b4621d1ed66fd5037c3da592634b754f4d17709e6b55c68b1e8054a853f90f5af5595db5056f63b47761b1da65019e95a643c977195bc604ed824a003cf39561e851ff45b557a92abe7de14444455f076bfa48eb23b036942c4e174d3cddecc9363fe59dd4d4f11d80c5833860358b4847dcdf127a82951ac1972567799aee40b67273649006ddcea2bd4d60d44c90505d64d208141661ce5847c24cb65b94205ec91b9463a67411c42f8837ac689ee7cb27c1331740624794727784546c83427befc712b4bd1d8c903c2bbb2ac28914bb13295f88e4385c308408c5fc7c8ebf556cbf235f51fefc1f66a98c8f865f4eb1ce06a0641326bd412ea5d3d87767777a8c6d37fb46831da538bb96342b5b6c3a66c5c817bf94610f3e09a13d9a40d25b2d0e3b587e62d7ccc98541e8748c4c411d9b8a89c4d11276b25a3dbe57ff5db704a7b0f8e48299;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3c709a51bc240a8957868f85b022d2b8a3b0857ea8dea5852aa3827031102b0f7373beca24d9ccba628a2d4ab1fd5dee95a155819c21ee856da14f190e691714eb3c480252baa77086b936f0368985ab5c0ce479780e77ba7b386872cf37853c690ebba0aa1e7c3b4feabd71790bad92610e8d66227f2a3fe8ab0b33bbf11fb55f7a908247ff526cb41d84a0a4afb30e627eff3af6528fcef700b7b7313d8fcb72a0f98aaae56bce89d16eaf39a4107f053f57e8e52b6c37506023b7fb283a9aaeb227e5ee53818af8f329f8bdec3a22ce90bb54e99c1cc6f82abca25be671d9680e9e9e5f9f8d0913dbbaad324e062c2937304b6c0a3c98bdc2f353744abce6d3efedd6a6a8624608913bab1639a699f9df46787273e01263d64eea505ddda6c0400ded59820abdf275e4971dca750d5b35265aa113f08ab91a965d823461e82005e36d2bdcab1a314a1dfe2ac626effa95d9fc41fbe8af9a5fe7e404ad0cd2511456ba674a962c3bbc570685d16d1d69394b6a0db61c313577d73b91152571d8ab88e8bc8d19f72b4d0cce56282b697cd696986638ae1ca0064654d8c901a8ee7c903955498e10430d097951079499e0df8d275425349602b98a6e5cbd197db9c2575e5310abd44658e2d925c330d59b06fa7f748d45ef2981c232e6229b017fde89648e1d589f46ee3b1390601fe07c52f3161648054087c7f90f7bb77d1d18dfc1c060e44c5f02f24dd92363827c3bdee9b8d567713fd13c2c1736038ac4fb5b416b1953ce1f3b009d22fa150be313f666e53767a5370428dd779675a9673d9f74a61885513dd81648fed1ce08f932c292703869301e67aa6252703ab73ad171a8b445803000f0700c4f902aa3fcb185a48e7a77df3417796b0041e54a4dcadcb63eaae982774c0cd8a6a7a1ce48b294027dac7c0b88a0982ad7a305c1a952fcf4625d30763ca704ae1052413812ed358857585dcc108b44bd9be46ce07b0ae0f89931755f9767f007aa613aad5d9b174b231e5e8cbb64532b88b3e4bcabbe16ac775790f03c3072ec327a8987d1943f6e9ea43eb0e81208ffc5786d3ae0a02dba821f607e03b6bafff5d8198421033720a5745f2bef1ee93bc21ad9a27bc2f99a6d859d07d848c506d35a3319629d422a1405a57c290cdcd617cb3d807fb4791247566fcd3fc7a780e9bf0afee952520710569cf641111a0c114706e165567ff53f73fb9116689aebd4424d74ea01cef4559bcba561ec574c6705a1fbbb38f51d947902beec4322f94301e8dc0b7db68679b41d0040448d0d4d7fb1b3d71ee68ede8a3741d00b6400ee9b8f0d76807e1f3c919db9aa7539de6c5ca3a36099b893ed196a9bd5b70373945e94d5102e2db23170a9ec8d938fc3823d1ebdd25d8c7faba6dd3883ca9c5c32bebaf735e0e9cd9faf4ae746e4d4c82de5585a36c9c5d930a7d96ac3edc9e36776191d437ec20f3d446ed91a98a9d4cea8da54f0c655c645608c8b8878007bad62afec58c8df981592f220cff6f2a0b6c324834e38acba3b5aa822f719711b37543f1ff91e854f223c50ba8f0e520e159811d888740fb1e216f67e24b03efd209e1d191a8697eba9edc7eae5d49e166f2d1052e00b34cb46b7a2279c2d7e83eef8ab86b03308ea1cdb8bb850be27ef73064d4867613a3e403bfd58b397a434aa1eb76a3b5703dbba84a7e1ff34e07ad4ca791824986c70f46a82aa1da3df1d43cf7762df13bd369eeefa378baed61cf42f1cd8735817b10dbfd8b7d841a1a4cf824937e7b1a9b287cb49a531095c54fbe1bb8f3fa434c5ec0a7661bacf3a0eb34d49c6ee;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h27dea5d2ac3da9ab1be073c2f20a1509a766c1b88d1872d18ed40d41a12c59c432a0111a7ded691216874aa4bb6746c5a2de51ebcacbbecd68ccba947a219f8e2acbd13a8d985cebe9ec20dc7c1dc692238072e93e6e52c37839d0cc07802f74dc1ae3df4050c01dfb162209b3b37f86a626a3e5d22f26f8041f5a28c21857edc560803461e0bb4d335434e24a04837de93c197a6497215e2eb3c7c5d7cfff2e5f74d990ac88aa368ecad259164db55b7a9c95dd0b95ec3f5d2be3609e71bd0b8c5e58f3981eb45184b5d815fa9dd1361e857e155a5f4dffb348e9417f9be70ca9f787dd646e51462c8cf95af24b1ce76ca8fb9d5302cab883106277b147c8bad706156ffc4fccca71345372ca809323414327d11e361f0465e80ac57c74f18d5d2b4716ad1854d9b056920a5f6f828061e873ea18583ee81faf31451a492eccdb55208db8cb9ab59f163458eab5b53a2a016eb4ebe96382572fc5bbfb5d8abd22c27201ea8f63cf49d5a58951affe428abbe2a6ef9a458b6b38ac087838e2c4e5ece95ad4f345e5baf7bf45f71fa08824d0fdda34e1f4cc874978878460b28a763bc84dc8c2767811b0106024feb4a368e8345b5f453fb4bd0d16fc6480a70320ceae15328250b6d2a6953199be6dc206cf2f654820b2f173b000f5919af9e0e1ed36e0c406e257795292dfbda0b010cabd04c52ee915aa959f1c8889875606b950b643bc8c6fb7f6e83c0043eb1e7f08c46f2d5acb35941473a54177a847214d068ae9f89c0f8ef9a1a27d9452329b28e24827a29ad91f318c4b7edb8c7b5625caac7ab4f597a22748a72969808b07dbf2991dbb2cec35b55e17ea17c1b786d097b5b3a581dde45d1e8b396a0b52c02f04c99aadfb500e06fe4cdd2339b43ec70f016e67e49e2164f482cc3f1168dfd7e736c7368c4f7e4d8a483cbd6d8bceba178447a1f2c60be6297055eaaac7a8463537a62bcc2a287b108ac805780a334fd62d787129a64d0fa99e80533676dbb4b6e0df138b5423a68628385c5a88e853ed1fb32b3163f21f1659c2f16d93b0cc07759f082c4aafc714a7fefec3ed4cc58bbfad8eb678128da139dcc2548ddae6a58caba5b6455ee977d397dc16503b8e66023df3896899320a4ddbcd90544787c3d525e834fc6e32e45d3378b4ecf4b626c075a72e2f09ea8e04d060453e5a585b56ac0b5a5d758c7ec1d6a8b2e714e0681aaaf943e873daecae64a3caa4f8197a3da412a37639a53a48e94a8d8909acaa605f456cd1fd0eb99177e0b8b44ce2bde1d42a94b16794d669da59104c309baa018e682aea5723ddbf54715272184fed96f72f05bf841cd7ec75ac7fa2bfef31dd226290fd532ad2fffad7a6e259de3a2151b5f75515b51c8df48112b09f56aa995fd7403cc20f8e93516148c40bf2d4ce372f7e0f7ed6ba5d22fb931301cfd0a0fc17880d95ac967e070d464c2d2e2758d0301b821d53cf84cdcc5993e55cfd98f9f3e6d951d8275ce04be8ac78bacbec97488f480f67e281161a8374fca7841914c45d2179c40b8ea8a170fe6d963874cf70aa222a7bd2f954b5b087cff3683037c7ce8cc1563a1bffb57039ac05306094c6642b041ac4e523843cf1f80bd094d697f4831c03760bed075cb99dcab8b98c642c23bf89a0b9fa7974f4a780a88a0ec7eafd87f91a724568a448c256d6ed7485c6894684ac8214ce2e8094ca98f0baff457793e017682332b301e4afd9236ce7e284bc0a3fca16de15a7468a65454589effa945f92ea4497a4fd5c0b13c83011659e5f216cb2edb1c4b08fab265ceab6cefa77b38b98a67c81c58f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1ea43eb519cb28ccdbfcb9e08b68461100fd63a4509ba9d61eeee9d26270d73d3af114ff5932fba56c800420fd304795ef069c1b736ab2a08f7a8d47560c7959df5f8e687449cf064a1dccd05d6bcdfed26dce0a05a81b84d2c9f221dd930a61ca3319d8f94a7fe6656bca26b5bfa4e91fdab0aab9a69c381456c47deaca96e4a9b6ebb663dd8d7956b1c8f19c0e2b507afc12c6fbacf1ed02a2aabdc55b832d80a0e256687e2e4b2f9811ef1a298da84883204f9a61ceeb88ce432beb5c90f19be8a9ed795422c3b11a83f0ce4967567b952d02e9f23c8f23872c52ea287370a63989d330a3dece772d799a4fc9b475cb41fb13f9f4dcb983904d8f1a777d61b442e243669485b0f9d01b5b46f109252d335d63d2f19bf41bb35bdfe695eb26ce34aa68d49b8be7fd6e8b40ac3e240b543ad9d8170af526fe1519a8148d9d040aeff110ad4f4c0bf9b3ec7ebcada68243f694021bbde8727263ef7b263c88e60986d32fc4f62b1156932ece6b48a83279eb9432fa2d68d667af6aa9a4cdcce728dca0d02625bfd1b89fe98f40949974c90fa80558a852b3144f7aecb2f322eb3977210b31867920535f2848aa9f78d21d5d554e0227affd30b7c36527f1781615dd7b196fe3f1bd9a58931be355485f01dd2f03d2b9c0e7c3bdbad0711e50871579821d2cbb76b59117075662805c04855ba6478fedf0cc165723bd188b94b95492ca9bd99291d16b935ba7f457fc94da1964e5a3be43cb44f7ec6c354048ee94b44a58606efaf369b2a867b90f305e2faa21fcd8a77fe7a52cf3867093f7a6f8e03fe7783b90352a69d917def9f9f4899d6d11e4baaa94b0e085d665ba4d5859e56aec2cad25851e837a845d9ab0e0dca4663c5a7ab95029b98280541763788bf61325bc9644c8a84ee87f2ef3df3cc4e81b781b1e880f545b25b560b45fc3eb78541966971fdff1ecd66077beaf9a3be04f172054fb7f9a3ecdb3fe3fd49ff5e565de8243be9d5c9c910799f5851a88dbf4e9efab1e7385c56ef32689ea44ee750fb70a44e14758e29cc4cbc7b4eb420ff0155446368ed9d9971e9c834ef3b4c102433dd0ac2307442ea53202e836149a131636a0ebbf00994ae68da9c8ad3980967574d93797618daa421ed50f64564488bef4f0c4e92bb7eda47db5033ab11a6fc5f0aea3b618b417b04a05629a9326c6745eb4ca0189bdff3fe9f80fdf08a0612488af94f83c39f9b14cfd0ca4591fe99dbd08d8e1426bcee16abed2ea2437d397df089c8be9c38a1271eb23a761e90771e605dabe2febc3a356499f1f67ee4d0d6a9790c291885f625f2bac1a1276ea9941857ae5fd6a4821551887d9872057133c6d676c09209b251914a92ac71b5781861b27abc3b226cbf0136307e8828678a405290abb7d0938d35fd4a1bdce5f197dde76803156416372df0d9aaa0fd09fa181cab9c60b8ec8f26b5e0d82e6382518599100be44b710ee386d0679b658ed43f052f0cf16cdff69ccda8748645583aed5e84bfa258e9400ec18149ae7037322fd7d6c723c81724077d14969ee3b536307288ce12ba8469536aaa6c3cf35ada4c1442cd1e7b8817ebc5f4a30be974bffd392136466dc2555186a8ab1434e8325fa2c2171352e44dfe765e679532dd2cfbeb1ad806e9df1262b4ae94dd89a98c28c31b6fda070257e9a99f68298ce991a6855b7b881831beb506f587202b1bfc94c19cf57c84ad19637a99d965de5b0e0da9ebd310c03043dedd61cb7c1d97dce74e85bf4913a3103c5de7ddbd7e37bdd51a42064230ec8546f14d1a2d70e684d587f6fea85ff4a7f25f60f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h37cb857342654546f16a26a1d63ba923be6bc480939b1cc9cfa4054d9bfc8121ecc3403e2c6048fa02d1f4834ae21d8715b3b61c5d79eab864cd6893c17e077fa4f1a9dc3e5e04c4a3ea3458248041204050193371caf8f1b68f53e1d9cc20a61a65caf8b6ad9c3f6de093856ece6b45abda285e169a037d38ffc6b92d7046ce753b511a08aba752162dee5452fc7a828ca8785901bfc8255849455211ba7a9ee9dc0d052341412aa6c0e4a8d658fe65c4cc7739f7ca76699d7bec14a7623096f8af54f9772c0c03ad8e0bdeed5f1c816e812fbccf759c60a77e2e4a78a7b987fe47603a29bd7d3f46876b96843d6fd80d8314803840a8277e9e86150b2a9dda32ff6c3f4dccf8a7914448b4dead083c5d0d3c8c43f0de1f432ab3d78debdb3536b2e1da121800cc487d65104ecb587eba990671670c5116111b65002f7a115f438c65fc10daf4f29381ab76c7548e8940b89800135d41bcf06eb1897fe274d42a188cf80fa846b5892c4bb4843e7eeeb5857a7fe5979d1bc230c18147ca59150ac6f9ee5708bac1400faf1e6ccb88a21998263fb023e745d1b6e99be3de0186282a10d5c9c19a4f679a820ad20b930e02b31166461625d2d68cc53bfe7f2eff16985b83602f80e94e06bdc27a96fda97e5ee13f1f9c7bbd63183f031345fe3bb38fec0682c9a21d76657828889423c12039a21786501cee0da60b52ba8fdf0507be94347cfebfca8bd2ce66b01003ab85d71b4597d722a07983fc9ee4550c2a8184f24f9c2d91267f9aaa491f6fbc55d999d2adb37946799b70ad6c276e960afdda1252d69ab5cc32e68ced88c49d2aaaecb926b62a3fcb75f4e86f8eeca6fd23fda744299b53e2c9a4c48e47e37f9c52d1a0e693c9ef28e9177584d281a5eae8a35a1947fb8f6cf97319e3b18d94a2ffbe4a543b16fd163e64c6f8c14d9bd4636a717570c15d34bf5a08e0034179dc2e5b6702b9d46acc321c246b9d79d80a5759ba4d078589d8a9f5c8240846154b1be5dae0e55a3609d3b6d1fa2cc46508c100221b8d99dc3e090c31753dd0844e0b7d0e593734ae95e7b0b1a0db8c79e874dc5a5b4648592081f088d82ffc5846931e7cdde168956dbb375fc38f7509d87b5ab0cd485257457d4799b81dc66c36a2b0e8f03dbe1e66af1b4d5470b2a92175ca6a1a421e25e129b09334fd1700a409009b9bfe1d41ce9829864b88c885fd0388878fea77c4c9f1956f582a2a74ff8b24b48cb76fc925e99d475893df6dc11c4a3be3236dcb6c824c81333118d221b1842e966a415ab4fc0ee3780a5d53d0111a77afda5a3b6de8f238655afaffa85b4a42710c9e3ec3cfd0ba076766dcca5773a8001eab58452698f7ac023bb3ed562005d4bcc0b8d54a9a1b55f26e1b15f50529a75bde3bd28bf1fb3c057f770ba9741eaac5ca4bd89b05fc2cd24a0b21cea99625818f69a986fef51491c2052f35695711aacab86a38d20250705ec4103e770115ce65d1d7a7423e8e28d113f060f1dd1cbfb963f54920813614ace8ee455f5e5fbff5987468a01e224806027fc47af73731791ea9c8c66bcb4d896f3aad45bb8ac77fc77f1a8028716413261f5c71a41be85cde1cad33b16485460a6b852a63ef9f165ec06e3e2d0cc76af1a7843714ad273c950482ab9c12eb6c149ec9d209ebc814797ca1541c6e30362396677def000602be0480d8fa41bd735b20a0f7053dbed428320a1fc9dc053981e583b52369ee8e70c043a2c42dc1977c6ceba8efb45bde361f87eb374d23b828e58e5c4b5139c05873cfd3808bc3a11f13a84ac4335b30f7c0b75c6bf9a8e80828;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6fffe49d65feeeb92a053ad178018adac08540d895579c76934891c0f39dc2685eb151ed5d01b5bd2d6cc8d0d1c5c44f593f7bd464681338a9b0e573b0ceaeba965c86a9416eba2a345f9439f1546f046d77260e6a09c2f57ab01747dca8fc75db2e595cf6b52e6e60ed49cd5041e62b9175ba1d7ef9ee6fdb1e5544471195b73032279d76815cd178ee21a3df00833b8e025dacb950e9be5e0d061ca563fe5cdd76124916872d29818a6e7583c2f30c34892772757e9047854f3886afbab23c115a27fd869f84b2cb54c5377729ecc28dfa94077a31f357bcbc8f4e8c290b609e4e4dad40dc2bd0202a9af7aa2d73e2dcd0c32cf41175e4447520ff24807f74f09e51d6916809fbde4f2703e5d840a92a133a9d03cec0c6522c4ed1cde71842d3108e40f3be20a30e8df28051b543d0c51c431101cc2095fe83d8c9b2af518c2729f43ad9e8c235f99f76ced3d1a43adc718d14500e6850d3e32eaa91d559df334ec2052537736ae23c3f40af4af778164a72658613764dadf3197af4cf5a644e17bfa8c697e2dfc3d951f6a7ebbcde30320c9ef678dffef46045c9744976d6b8378c929478eddf64fe87e2e9581de8ca7df44da2c7ca07c478dbb38ad855a61a93504376085edaa140450d0464336dd01a2cb2919c7c1bf3ec54ac979d1440af0b1ea7dfcbc8067d0654ca2688f4853ede4866e896144ea1a61a2984692e2b959fcbed96a08a05890209b6e2d75fe6c3f1448a74b4e89ffaf524fd491d5741876a2d698acc3eae0f4cf4d42afce5f2aa05f6b2c8e237042b06d40e812ba16b5f90c383c5c3c0e18e8a5f1083e882536bb21515b09f2bf16777f3dafd6c372e85eda2b51393ed1761c68a571bb486eb96c3411d77a3561778af7c02759bffe929453a38b768ed6b593239937791bcca71f339ed9b13b5df821da106237d03fe069a77dcacf17a1ce33941f93f928bc8729680779479131d9f97f897a3024f676c0d8a512bcee84ca5847be5241742cb98ac176a4f118e432a3b65aa3695d04d411f6efbb365ba026c01ce492ee7220a4e4bc392623fea11707c814190a185f7502592605d981a59ea6a4efbb5c7a4d1ff801f40a7cc3ee7596d8731283d6d3c1f7b2e54afe9ff5c911c5a596348157e8a9f82443965e2c5b93097f56331077d18f52029b6602ef09b0a25ddf5cae24c3c61a530e4e7770237cee19f49c16ea8dd4191d3f4169a12e0a7cdacd36088479af067663b314592cb62125388991844720c973ab5e949bc18aee29ae109f1fdb89c5fa5717917e8009baa3ef319c98df2e4f7edbbb94d7cf30155052650deb84ed579dde310cec49a408bdf76770b245129982c2319f8f699998c9b6bd3ea18217547a0df8d7e676ff4436dbd63b6748528e74999a0a59ac809c8dbba46bed84012c3071d757cc1c88b4cdea9f0dbaa1ce701ee334598bec18494566de1921146c3cafc7acc0ebbe7bde5bc3e9e8a76d68d68809e3ccb759aa303887625732099b45de9efea770001a2428b720f0f90ca17657642ee18751c9267fecdfd24234138879b4e061ba14b20f623c3f2ca5f9ba6aac5d0b8310c4efee032b9befc705ad0c0ae44a0c07e5422784c09675d06276edad542a413a2f87fa77ec5a4afd25b864b0a691eef2a7cf51a5d7336f6b79410c87544cd133152e84a3fe5d99e42a1d295fd2748a46213a1a4574b568e01e69e231a058e7d68fa0c8397a5ab1e6a55c77fa722ed186f7b6fbe327676a22fc4031e72a4d1742c492fdbc09ebda91b12b530ffa2373af5201a128ce53725f0c5a21df60eadb9a18900128957453e58;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h432b333e7adcc71c5a652c28f44f2e1ffb432c8bf743019057ada3541068e0bdc7007c7a42c218e6296f9929b51b44d07064f1ab12be27d17149fe3c41901e72ce3df47804eaf7ede7233b8e403737b1797c62f012a048e6ea324fa45a11cdbf46c2d51b879302075866622d1e0ed66a821a7904b57ee32345c3e769e00e041bfc9001743a915f4aa9fd7c6ce5bebf16fa2935488721f793f79ecd8fee15a85d67c8c9338526763274f4d7d94394b15348e78368e6bee528c0cd49fbc57980a89db6f67996177f53e9e67921309d566a1e1ef0d37802d2c61433351caef3a7817f857aa136c2d9b5713eae5b53fdc0cc30886ec91eb61afb4444ac91966acf4241ac63a1d1c98baea69722934029ad5fcc14c5f5dd0f0728362884a6c3b0df09bd929c63adaf1a5a8cab912b1fbcf6d5357a93a583f1b662b0e003bafff7201b734f44fa128d6b7938fb11f1df78857ff921a6d0292972f623c744184472d8842a0ada74c958140b49640dc1dcb6881388cc8ae337a98019b72e98b2640210a35e47a605f7cf0a5e50991f1943625a579cc39af593d26b2124abb2b798550350b103d7628366829d2704bab1454dfc1f03933c0947121b39efa2172a1e6a6d25b6098d13406b6036e56455279db0dc0cb1fe853bfbc0f4687fa4094df4e1fde5a0723b5decd114e7d41a10821782c4464cb6abdebc28fc9d0e17287c3128f205d0e82a6e59ef6654a8d32f4ddc5b716064f1df31543ba7bdad5068b9859ec726ce444344849fa8ba2fc7dc8d74f62517a983f7f53fbc89d244aa4f540243cadbd1b5cb84d101bbed1aa7f477b4ee997719d398c33b78ff8994aa158f8a1876e15d80c1f942da1d67f6641179760adbe11152c6e41994bd127b08ed25e361df7e6424abe30a14d03f4fe3ae25494e75ac04a1fe916bbe9ad7d088827464c5eac31cd9d7d473cf9ab0bb7d0169b7002e8c5bc02d3f924302fc51a29250acfc409f8e5c7c5ba932edb9c2924c85471fe22cffa624d873fa3f549fd77fa6da4376bdbc2a091bfc8aaa18c77330855e843fcb520cd40d50de0fb5c6da11c5897aa5caec16847dfa42d7ec9c7e5cfea58452165f81c5f59d14bf2a342964e9d1e3000c35b8c7f96c4190a12916212794aba6af390becd55769e02a4e604d16bc83c0fca1e61506e8d18313fa16bd1bbf90c833ec5fee5becb8804d4bccd1e27528cf24be00b9ac03c72da6778b5e9964b330c12da332131b1bca5362f50793809e85cb5bf0beb761ff5df7ee69c6ef1addb0b34a614f6b6faa78bb51eebdea06d149089b23396ca567064a3e6df2771756189779f9b26e980fb9dff555a5ac2029610378595a5475107d772d11b2507460c0a01c44d704c903d5e5d41184b779ac90df15463bf5f4d5e46e7043aeb47bb3c28e9ec28a77fe046453cf0b451a452442a821704a085a08cb3f8670b9b8f456625db3c6b65fa3f755206c71db4c01a4c7955d503543ab9efa5915e3b1e444b6cc7de7916cd050844a88c8405af040793d7ecb726b4c91630078798390b6f5d53d9aafb2f8463fd55cc28b62dfd7da2c18feb51134f9737ff91238635d05487a0ebf30b5a929e055a1b14ad542470d53680ef7e88e297c88e41f376f045ce64c512c8caa51f9a8005efd2b883574dae5740d0c0d31a38c44bec3666da21ff2838d2b85afc9f0e0a0b24040666d7fe517c53d971bb029724c8b9588be1a35929e0beaf374ee3e8432673f5f809dde3b2cd26020b124ae8ddbbb6b19b964b31b284a4c8a12e4a84b39237c3cd00ffb695aec161b3a277533b5d0bb820840249805dacf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2ff2c1cf29d91f36de0026823faed7a1daf875a8c9622241ba67de0c132a58fd7c64c61034e60e0fe27672ac4989a399398925f5a185b618c947171b57603bdf246effb8ccf5be748a0dd28a093d85aadd868b8f5b5e3c31a8e3a708b689fb285376f027a72da1c4678dd4a6f8529f2309c0de6b970af454fdc28ecc0425539e8f720759f537d96e2180fb854ef98530303447c888a81cc4e900e64dea52eea4ed9d35b12edb030e5521aeb9d825b800fd5c34a315938e4debb96f027a969b7085fd5ee73403cd857508801cfcdadc674b4640015ed828133994cceb8f770c4e8eecb9f47ffb5d137808b3432723727f91115cba8f1e7ceab245de53bc56d0d48d870790a2c984ed03da276ab85955bfff1820365048bb3fafca12cfd7262a2371f004f37fbf99c836725dc99b5843abc33a58580b067eafd8c9518e0ef84894bb876fed2bb18e1e4b53c8b19967357aa65d1a2190e367818fb46b8dae75e29f40ce4dd42b33174391d55a69fc0643c9160501243f18992e03df8c5020102c6d0115471c893139ea8fc7e5e3125462b4f2aaab8e63f97f5a83df5b7f11bd79914b3f7fc2b0d7434b4f6a39f753f86dfaafb62f53335fd980ab4931aa76b7fce70c5354a498a69e226e000cbbda36be7fefe4daaba932cc015dc819e7292d619aa1d24a18e2aef064c314742a47af89d264c75c917804ad3c88a116997c2b575292a7a1ba558bc05a8d50b31201f1a58d64b63d06746860bb82dc60d84e66776da23f6f7f33089b1cac188570cf9ffcca227a68cd7b56f33d897a5d125e309a9cb4c0d01af6dd227a798164ecff6e0dc5bd4129842f25acb7805057f7f02549af11adbac64e47c9b11115c7ad23a4fbfaeb1d6bf4141d511a8ec75fba0166217aa27f59b3c0f2986c7bd993ab8b972012b7f2527bde3ea2f2ee0cc4f78faff11780a6a42d6a240255357dbdb9032d4ec03e163684aad669561ad72074ca56f01a24d9e739a56517abc6a792d1478fa89951524d0b9f184a1037e675bf60f6e472cfbeb22869ed4f40c5cbf16e9f33f5d3f2edb9d9818e2793ec9834fc8c23505ad659b590b0ca4b7890ec24f3380fa14520de6f00a75fa2770941e65d3ad1321aa10092c160c7248d534cd3f166116b7044d375985f13a7b6cbe2aae9c3fb8841439ca5595847b936ab89cfbbd88ba400afb26f67d77ec7bc235b0217346ca18129477823a12b051c67c5a867d758f9a5dc0c1729b805f139d0c59f092b227e5a410873573e43c1c2378964e08b265892bc1a7d9d9085edb66bed7b126baa2daf19f1d32bf849c68860b90d93c10dace0f12f0b0e252a2e08d617a25b4c5f992337798767d153a9515858355b5f0736fd49d493cc81bd44f8fee12a97fb901898a3969acfa3544b1c455a6729542e20d089dd803b1f8a0625a4e3c291894dbe5a08accec909809f17c083e0bef46ab2ca5ee6d0c5b5e9be7191fe39721389d383ff1945194c490b8f3956c713c519b6d78e8865dcea1d0b58f1c4aa6e76edb1ba48d8ab7300600c214a5e6778509484391502f5f09a24014cd65973b67155a14bc58d9be1e85ceb08ce28ecb6ce7554a4787165822152ea43d1eea1b9f1eb2d16a88c930dbad8069c1cd9cda608b127fa68b9dd52d2f807ac64a8254b171b70b8e6b0b2290077b2b09770899670bf33d2eb14123445ccc1d8d073a28ab3d68aa9e05033351a578d5596c0784a45c126d37512ae4d4a69752e39aa86ff202347486c94794a3f0c6931a2cb235e5e5db4d6d4ada406ef351dbcb4519bfd16e4138dd6138179371d55097e7b2d7d8f84ea1f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h68d8aa897e609b3da2e23c8b98a6a790077a9789762ff38daf9dd7799e4d4575175050a23ade42f32412f26dd37b4ce150afd90af11e2aeac9ffcb422bd21a1a0d2a82dc7e4272170f362d95bbcbf8ed9c6f301d3b2dd8d38d3f001ed48f9ab911fcfc47af2cf0222c793e576b011c2adcfea9973ca3c846b2e368ebcea887a30506583277285d8e3ba12e67d6b7628bcab4b1cee252a86632dedeaeabd01c999415e321d1c7abd081de263bf8b51ed3e2097654892c85553739e11605d674edbf5a08a79fb89fc54130422c77113bb65f605e27105de325e14dcf0070b7b451d89c21efd78b4aa3459b3f6f032f7252f9da0f6d29533188e00690f734a11455d0d1deb949ba62bc5d311e3b12218a428198de7e89139fc8329f6d1ba0b932cb237315be7edd51ef8ba683720cdfe958966ea7783c3431d3c33f23c92e9762b2ede94275965bdad12835181d4c4da38f2fa3d2b1a85c27b5500ca99fb537290847dbb6d0e785df8b78f1145a2c53e41fab4f4dfe000ab5497dd4c15b67298d5442fa67d0cb6a657598277f00bcef43e1a919680f447570af12da898b8927d44e9f259f15bc8371222a322b11480263892567b0435722eb8f6cb964c806db7e07baca03e8e3804d79e6355c15897e5cd528861bbcc16a3eede7fda75eba4d411d619b41d641b8587c48e1c3f13930fdfc776a4be1feffa81a9e143d9e2b897ed5faa0a6a8e4fc4a1bf99813abd231196adf506f1d8a948669f68d45a65fef3bb6bb4c5fbfe3ea8d75277fd47b967a536e2813f4676a6f37751dd248a4910898a2c02ec8aee8eedb74ec317fd96fe2485cfef8341c11e633540801dae7de02dbcca330d4d78ff90d88b67a8ee8ec3554ab1346ba49f8fd484ebd855ed5ac6980dcc57880b37c900266e387ec6719902d634c88b334f045bd3e37e41707c607074eb739ad6ad7ca9cff838890ac85dfadffe0cc9f70562fdeefd9316d2543c64c4c7783e541c0c9499472fefcbbc014900e6820b18d602769d1372348d40061089206c1137b270e8f89a46c6c70b91c8e464d62333e71e6e92b123137815695fe4ce09f080e344bc6414571a1ae2175751955e8dd24696b9ffded5aab47481fc95257df806b2738bc758ca1d9b540b725d3e2f7d6952242fd7fe49f464accd51d995c18ea8c7a2afdfa93ad629a64c9c7811e4f507cfb112ad44f6282643f981c3f9ed76d3f6ae61b12cea7fc81fc387b89c403e3f5325f5a65d676c2ada9f95d801df5ea5b53254d03dfb9df219672e988fac6d7c1693866dc236dbecd6b0d5ea3fe22bf259a2acc094d806eef66d65826bbbac9a36ca7fd23516798e3a0e7244982b068c50941a86bdc8b4bd63ee5d2994c03a81b7772d474881e539d483876180d27f3ff0352608f04b92bf1588fa3d127fb2ac38c817062f447f85343a0e688b5cb0a9b2a50df3a5f72db3241a9c96205fbb97deb157153cf4351f6d349ebe63ddc6be166d3eeeac1b38edcba25629f3dd1005372474980252a0be4fd09c2a44369b81e2b12ffdd42bee7a6c9b7de93a5c1aba82fc9676fd1ade161e9c4f475881fb7c22a00101c0b09478d0937adbf3072494ce94a4e4e44f82a33c6beca530ecf4a62b31bbf4b85e4578bdf087be524d4cca6f3abeeb2d8a3ceea0f55cfcbfab688df2449fd77df67d9bcce87aea50f601301cfdf95d5a572e78a49aceed77352b4e78831472c5c9293ffa98daf0f5b35a9ed420f5822e1605976d0c36265e3eb1c1640fb0ce877964e50d554d51e5250155ac92534b9568d877775087f9728c6d594b86a03e00c6ce3334378629;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h11b19b95c1205270e60d4d4b8baf0e03f055179ac45f645cb6aabca56b56a24e9c21acb0de7c76e3a4a8a4a2bca457d279f58a35ebbe82b1515565012c7288ce748216f0076b821887b70a5c0c8f1f02494f10fef764119655dbce5d29549759df8855ae760029bdd8f740b1057bb27c726e1f7a6a220891777a63e842b429c2e8521d862346a8283a4974c551b9c1b2fed4257a5813284224ff9f97c93b2a488b30ede05ef48b0ce16e46218f85bb6a6a68dcb31994b567326560d14f371e5c89189c906e3850a84c3b379431c43c9995f9475179a393bdbd374fd0fa9afc916319f5414b46ad541ad991a5552ce3dc62d3952fd8570c388d079300e7efccb616b35a2f7ceba9495b17d2f34828cd69bc05875a75d3beb9ba88956351088062509267e1bb0c7b43a9d7b33f3283f2eac471839da3c29b1cef48aaa0e151dfeca70b4605742348a369e815d86c521a75dfb876e33f0a7bafbf564ca75b380cb876d12534b0a39b18eeefefc3a59e531d9708e6625c891bf84344d9568cc3550749c0264e6b9b116b69bea7e8fb6245cb6926a1348bcd320bb0bf9ee53830bd3e152b54c40581dbfa42547e64f23189a14858b909a30d5f11a80e09c9da11654b50c4b51249892cc4eb6d2b30e860120d3da3d466c7a771deada6bdaf5d1d185ddb7b93287d77aeac69946f09452ae7a6d0163fae4adff267965d1b0cd9dd9c114f47c59e6b3074fc1aea88d0934bc1fc15dafb939e644d5ffeacd5ee3f9f3584ba06b0a5aa76ea6cb45c810b291c8766461505da77b4b411bfaf8d0d190dc31583bb605b797fc2f530d7f2e63cc4df115dd74226e470c44fa91b282a18415ad40f59cb2b8e3d19871d6f35576ee7b8d965eab10b4e0f9984d33a6d952f2396139f7a7ec0a2dcbf15cb906d32ba0374da5172360582642ccfeead7d30f7099ebc74bdd919a5e8a58bdf674b23718d301fcb0855accb63b648f8eaa83551948508b6929849424aaa6796c12094aab57307d8eff3a1532634a451f3ddaf5a2182a2dffcf554ae87538814dd5ae3f8f8e3292014a6dba2b6dd9d2ec66aeccb91d27631cc9b79aca18e6ed4a1943aa9909f863d9b8dbff2ac1e1dbc6f7629c992dc6a9255c443a9e0c7288a898e9c6bd171d4bdb28c8c1fc21404eb1205aad3f629e7328fdcb4d73f27175e0c1214955ee86e5b5db5086b7d762ee5bd350cc947261bf803ccfe7776a39db33c69bba32eede4c5dac4cff29454def640e48c8655c6391a358245d4bd27959cf738812c565948eb9d85764f3e29249296589c978c18b3d1923db29d164de69a7b7443a063cbbe5141dca7f4a55f02564be60a37de2febbc1e176090bd9f000ded6d73ea20f39e09edcf30f2e2057b167d407b569ed63749dd8ebb36723219466a9d2cb02a4a1f2a233870085cfea4a1473e36ec5f3e53547aa82fc4ec9c89ceab727e44feb694f8283b57005ddf9ec05618a26d09c6ef6d4ed94effac2842047851f1985580452b6f396365ec674f4850eed345a6e82cb05e3927fb817e58f0f7da5d936396fe07614deddb1cba28290e5ae31f4560a1d46f2064f2b396cf54b54f6f72a629dc3c4a97f5889363deb67baa0264c1d3a9599fec0750644c61636f520db96f4dd6ccc2c2dab29df9eb41d26ba613edeedda4e463c6b98e0b65a8843e7eaf7509605e3e9629c068b7f5c40439b0dc542ed5ad0a59bddaa90f2b124de8a43872696b230645901d01612819abb8b5b084809f58a3507c71ed72dda0c0838eefb6cdf3094744afb6adbad89e2af0a44063a637ce127f9c30fb338620c7e5b6fc232b93;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hcad56696f57f90968d085b7c8074f0c01bf334a95ef239d206c718ed1cb5f614f3ceee3a0cc658d7e8e12eb7abe400fab9c74df618d475af3d61351ada104039b2131105593c159b2b1460e2c889e66e3661955631c3c1ceded54db58d677da3cb4a1a67e9fb162681626444761e78066376cd039333ecbd863983cdaf5f7dd28b9898df3c635d4e8e38b6ed2796e3221f88f0a1e7edab317f7f1767dd98a830eacc7d3b44f2901c85f9bcb50fc0e3b9e65f6e8645a090840838cc58fac3efd27e224d7bc632b132cb5691a174972b3f87502cddd4198e13797c1b9d02f2517e9301b1e569c0e4d98af8a2d642fca71176deaa4f3a3ed65d7edd9eb0cc04c956611302f98b45e90b10328a8e0beb4b3533fdc6def2f4fb869867ac4cd4249f26b02cd26bfb440e3584e88356002825db97169f9d13118ab2ee9220b890a7a6c3298d9c29d96d47b750553582bb02bb0d2e7cfa634dc1ba461c59987aa1eabebf3ea498543886da45fe7197fbcf18a8c0dcad449705fae5d10a62c06e72db934c91a9aa6ad28dd37eae24fbb361cf5f453bda930621d5792fa6fa310398f5d552fec6a52f46b37c5d5ecccb1bd6a0e6bee337b16da68061c66ce05c4f0ed6957c8bd3c1ef3f47d6c2eef0663a05ece218c0357d307c0baf14b410d42a5f44ae95ff6d5199e868f3ba03d6bed1b1ce169c832ed2991e770337f6b67a1f6f14d55adb1654a0497309110be50fae47d977c21ca18da02c32df6bbfc364a118eab2821d5e8eb878ce97b4158ff917c73324f97c9cacca6fc4b9e1539c98070236a51aeb34c2a1dbf77282bcedc9e5c9f049aba458e3527c48b5c6e3858e343bb5260ad352a49ebc1c2ca6cff1536ba2facfa8a6a5dda263280a6ae46272fcb56f10701c4c2eefb057bf007775c09f700f93007a7924a06d341838405c5ea05728483c5f0008fda3409edeb21229dd5dd9529d049270ab0e0cb007e48a58bebf233c207b90d7d167def7ff82f3c2a8f408f269410ad3b3469c3d944a0544b6545819980dafb8da8d597f63768c30cb3624420b5282c92b4a23f0b6c4b516ff6591c3e7ee1b3a0a4ed867b307acea5391a9dba563f625de29b45dce484f3ca75ba02f8e00c8fad6fbb50861951e89de8eeb24447835ec692aecf26d743d832cfa3320b0bd454c8fafaa4b1729150366e2a5bb7713c79ad24a33f135955df75e640517310395dbcfd1e65014a96bf118645e1b51b82407b5abb48a6d80be15f8f5640df0ddfd26afae34a520fd625cb36c5da5925477f183ad59af72339613469340cbd4e47dbed811b7398e365cf5678e18ffddb03a399307ec479c327c8da89d425b311dc90f37cba5be8104123c23b0bbfcb9361a70ddb352d80c4434a7710e85b978cc0b0c6bd1d5b930473369a363f2874a820682545684397902878101609591c7fd936cf2b978a16ab100bb404333cce74c009e67c11e0b413c7097cacc1bddda8d5df3cba892a279731502f04845a0560782850a19ce16101a7cf0bb97446716005dba65f16ba5b7ea4a96afd3329a03703a951ef46ada4ab73fd4110cdef6dca1afa17c69fd0e1c3ba2b799d5db1da0319a2b6ad9923f499f2b1b096ba095202f176814dcca3b70e5f6cc8e4fe67971131054bc955424f4961256362f8f0d2a92f65932c644d8c59739400cd53bf8872f67e67441acc105fbe8883cccc65f7652a439528caee0fdae8fb091bfa856f36478b8db702efad003b766d6f13ec363b9291b65a3266e981445870e9db93a39685036412faffc3d79327f74751df87702b527b8dd2850cc66cdc8db26ce85d8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h49ea7b0b803261b5cbd2b4f45af4656e87c7092a06dc4525ac01c20f0a7a3794d0a09dfa63bc6cb52c49528a928d12593a28273d5b3756b6e0bb44bee9c8090eefe9fdbd534f6065966aeda119b984305c5e20972c6fa6a3fedfa313d3adf55a3d37f125461abba290a924eee35d2df383380ac412288c7ed12624eb044b76efeaae4562ca03688e6223e6d6281172d4ff6115193cd5af7494c3354a2276c79f0e70659150027c91e780462e474a9685ee39e54151b4e5416f8928c1c358f5ea105d70896d34169edf083dbe2c690ad9505602d360afc8b4ce54231ee90796ea7396eba3ffc0e3dde8a89b0978127ff76138ba9ae5647412f654ed0e9398aa5f06c704e6affec9ca1e80a6c0c8ab5c24c3ec87cd8a5c08a8f696c8aecfd976342271b81447d41e83b20ace7eb2cd4675bd254b8895d92ada5358f5af7f51bff812c8ec962950f7c2c9a737002bc9f9d03b6c373fca4b925e91b7e3fccfe492a677eaade589b6fedb514109fc03d0a5e4514c92e2019e67760c7df2aad209fe08bf1aa18d775f6674ac39757ff4d791da042b92050d47fa20e2bab4d6809225772053c8cbb474b0a1a839c9f924d6f55ce5c67756b793cf93a0e40b78a9840b2ee0292e084439661eb68c1638a6c2667766d5fd85246cd74e85e2d567fcd2afb7233057a377b96ee127448309019be4d1e02e540dc68aa4914314e689b98ab352204dc3f9922566d0e058772d66e59876744db952e0ad7fdbadf96a4d682b3042ac4aa7910664f17361a67119c58b60c286a48b3c3fe04dfab1a5a9f18790cf45c7ba4b358a5d68fd3bb4cc80c4cbcfcee720c6ac3271cdf975ee0071c74eb2d40571482ed5ebb4a493720bc04d20533ccc73b2a11016272af6fa4c27c37146213e34ee3968373fb1f3d63f86e386cea0cdb51f2e524576ea49988530a7a415361caeb1ea81bcbcf8c1af5014f3b25fb29bee59fe261249937d23f9704af1d9103aef95a425fe365dc6c5ef34e35f84d5e63a703f5337966d5300de3557cd28722b51b4165e834d5d4369e30839f6774b64bc924b6ca7689b869ed359d21684ce1099bdb72b0914ae8e6dbb804424cd3e46492a4121baf729259fcc1e51b43e8c729a3646e07a7bf3cda95cacc3b895be93b3756b1c65c651b947ccd2b303b273b52f43ce4bbbe5d59ea7fd406271dad59f42d6e9578039c7303a7e4e7120e391c13690259a23fc03cbe5dba5e352a11e16585661fdd6ba5ce2910a59382d8187f83719aad5c236f7cb71fe4d3df08e4285a0e89974507e567368ce68cb0615edef66724d843d87c39d4d35b22f19090e0a8b28a41ea53f077c5b33fe184bf854d1eb3aa221d093d0e4a52a9dca9ac90126d86448c25be99522545d8522275445ee953ab9f5183432c5e6bd83b0860dcb7c0b88eff9c5bbbc6e325ea6cb2c6f0128a4e12ebf1135b144e6ea9a96d84cbffa9f1470e1a0f75605daee4c348ec4ecb7320eeef20cfc5388b0c95f43d920f19ef80d932e87d3b6624dd38e3d2ca8c715b3c9ae7692807256a00f1a9b6f2b54f0f1181a04d2a8031a4d5ba886322755ab2a89004378a6541f7b668b48bcff7ab7d3519874c65cd6e107617fc4ef922556589fe96f2ad780a0af23ce2d6585b9908d7838af2a52a873e491bad7fbca37ea7d12e32be2f9e815c7e55e509ab851a576818edc4fba13719bb8eddd88502f6cf3c3265289d0b18975f939510d1b13d51849cb7e004af8d3c9fb092c83073c7825be6e55654507a5e51dd0025127717fe39f18caef65ed253a84873b9fa4a3bebb3582a6d6e24788052178deb897e5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb7655a7c3349847999265cd45d1940cf033e40b60dbf356530663aec8f3491f8f6f7d7bb88d6c666e2b37056470e815e6ea7fafab941a92192289d3e83da71c64845366ba2b249944ba6d579e363bf0bf22a613aa618ac0863f455bcbb198c37e7b7738c2d14ccc1da389ddf16e818c8c56b81f74b1670c8550084d115deb860fa124b3e1c746d1acbc72be9ec4a8b1b9dde23ebf260b56e99de5a0e6eb5c3e80a670c5510c2689cbfc401a5a58e81f2c36fb92e80c0aa2ead994e42ea558be731681e6ccb17e169f0c8605aaec82d5318d75a5caaf50d5ccba35585def21cddfb0f3e28b4206b93e79ff921fd18804a6b11b78d1b63672bff766a16f6f15841dd094119023b469f198cb47868b0aef2056cb91d5b81b8d51fda25bb314a75aaf7a655986d20383b91c898c341520527cb12582a202b7032183d0fdd251f6ab275ad1fa02f606b2724d8687421323b8694d1bf9f0364ae2bd06252b9697adc7cc272dc0c6aa57f48f1a445bdda1dd15a1ffb9d80e04785f9e07d70fb34cb79d49b1fd441d8456f8ba1ee56ae58d3853562a5683f3cf99ea4f48ef3168a2f8168240367cf95bbdb3c398fe80fbd22668a8683b1fe0222436d0d99bd9d2bea2bc5fe1c8c1d74a7db06bd961294bac5447e694779f5acabb7b86800bb7ee1d53f74f9e7a148224ff5c48bf630219b0bdbce761774354de37b5728ff0e83a7c687e65a5f50f9f373c4c57e091fa6b58d02d358f097021d5c503a019dd4c38554f813d888e2e9dec03722e3a6c30e7f36cd402639d247e6ca1521c19fc69285fa5ca1d8d6231d511646ffc286e742a94cb611cc92fa99f0f759e2a3b5dc4a55e9fe542552fcdc8b4ed61587b2627dc45876ae70011cef27cc3a0184722ed6935a619d0e1613e6160a0323a656b3ff5c26020af568a39192751d81b7aa31db8a173cf23ec87d968d80ef45936398b4f18b698c7641632a6a068a610b6429a45e1381a2492b25fbc92122ba650443dc8565451d5f70f2e8fc3f921266b3a2d326f46941c74fe1f27f694ac8c4f002edbeef0cc71f61a426dbb517bbbf7dcf09f412b08d9e1a705c9001d89e4b6ff055cdce61b0cb295c458b3091127c80bb3a5daca0865e105b0c4c8d49b1d536c8206d5669a4f2ae3b84ad5680a470b921358445cfb4c34b8bc0c5409fb45179f96d2e470fb89e2f3345d5e5ab1f5f8b25c9436ab4c99169575a6c32d52e173d7619a3f218b4794c750a99defa6764e6c366d9e120cb3a975bdb6bdd0f99cf9374742949b99d0995d2613d4e6502dd60694e0741d53528e71a3587f30cffe943a9270a4646fd4ee479b2eaca80b8240b28f231acc5939ad1aa43808523c8de9acbc663b251334064dd1cbbc0c1242b7486c3b3f454e308389d1c8eced81624bfadae2228b24750458da263e21b559e5b1ba53d482ac40840af6205c623cd77c22554a1bd6cd0316f7fed320ad10d026484b203b67e9410603b691f60cc9c537c7ce9cda7cfd2f378c8ed19da3219dc55e5a05a72018104ba5100916c73716e14c159f111beb3fc592f5d0919243bdc8ed20329d25c4cde81d5d25a79df4d6874514b106911d480f53371253fc0fa2eac21d1c956964f2f68afc0dd9e9607687f8285b414bf0b4f6e6e7bf1476609b82508c6ec119c076c42ea0fa4b81e70a5ba64f51727615d30e29284941f65e3cbd9245e04ad77ea953eda2c28adca128f8d9120c35dec2870416433b9c91cdb457c68e2d6b3be9c7debb0f54026297d0c807554088d74686bb0f54074ba84ff5a792498683b28113623190f5a48a3d8eb7218a0656b5c12;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'ha9764833b9c94d6f781da660cdbced32ddf0fa19c33c4eee75b242ef7e88167fef97aad5d7cafd99306c8bd456c56aec7a91529c476813092841e87fdb4008bf15abd543c62b65677eb69ca6faf76cae6d8122bd0f6a74578fb4f2574f88b3952da4d55444f13bb11b5f9c0d355f22403e3bfeffac2ac84c97f42bf75faf692d2179069cad15137e935103327b65222768e4828a6a48766a7c239e945741064ca16c9b9379786dd35578e7f97a37ad8a020d783935d68a915f299cb0dff63f158a41fed9a466930465e741a68c55ef9498cf06acaf59d2e11af104359259a621b555d607214ed53d682c3ce8e028c0d91fe9598d666304ab669350122076cb0346352fc2506e6b3b025fcff699cea37feb5117a8a1a8db2c7fce4fd2340c5684019df1b4c829fcb03bd4a3688fa0123305848f488f17023c50dfc06f535387efde686398bf117ee2208893befd45c1b5b3a9f5192cb859f052ba20db265fa83069407451c9d0137224b4e4759daeffdc2fd485c4d8a0e1b8e15d4f680ca0f2547147ed19a0763eec7319bdae59ac969a57b6a78e38d3faaed96f059dd9176086baedec3ef3ec4713c11380b2c8995ce6ec03c424d2d660d7386c3ddc5c927d3e0495d1abf974a260da92b59a0dbb8f7d47445a793c6e59d5f2dba4557f7f940c4bb1b2abde1fe9103f37015649201c3c05309e8762d7defcf0f0cb3fd40c4d3ff9785e4adfba881a6c139e68aed6c698f220f49a2464284d294ca139ef6ba6e50ab9c4191f6c30a7ddfc6d7db83e3da1f05649ea42617d9d113be8fa1f80880d0a78e057f0eb94c3453fa22dd6d24f98a9470cda002a27d535dcbd0ec059458560133ac0048aed0392e70de573079757be6d07cd2ae54b87e1930ccbf69fcc5e400eb6cc8a3fcbb5b1e5ce65de7c4cd6c37746a771eeaa36116452b46c1fd9b2a353d91ffac5a50cdb8360b4ae3dbe5c186c60dfb746ba456600bca567596c5f3da5a06fc92e242f097de62ba980771fdba644c38730ae278b8a454515a75394ad68a4169b410210b34057111b31b7c43f86a045f58536c791cf3882e46ff83a09503747ff90db8a4503484290bbe12ff10ece601a493b491c81330608d819edb62619867f8374d8989c22731fa55306c84f3efbe830e8331fa9bb9042bad15e626de69b774a36026e30658e68158e8397f2556413811c2cce1df93dc8e91d899fd61ef22932e9c681e2f392a57ea821e56ec6ffdc75deb484ac28be12ce665fab02336fb6d60ff55d86ab3f61c2cd5a436831c41c64086974858f47bf2c41fa0052d5150dcf5b81c6652151391956d76f3b201abf99e9b1fb9e05e7e51004e2b30872c0f8774a75234ba24e05f6f76ea8ba206fa565b484c5bbae9ce26b4c8dca352c86c24c6aaae95b454d33070b8ba34325b0c76eb28e5bd1d94e053ca6dce6224910a0dc17148a5bba08e39cd436779c12b9fc0f378218277b8ee3ec8ed092931acf868da6278c0626671826a73849df7e0f232c5cf4035ebacc503ae2dc7b46d8405652da9585aa60a9499a2a3af3705da99baa0a44b15450000a939348e430dcd658144a0f60575e459ba976fb3a189bb5ec58a8251a94400bbfaf3a2a31ba8227e6a966bad9ee18d0b40e75201e48ba6b146727fb58f83b1fac540702c06596f3183c8aec688858f0e6e2b430ec19e20381f7d9d6d5b2b04318fbb7fd25502858ce9dc92b9047ed48cb36dc49f7fc8f340071e0ae45f755a6405531af3f96e04482bec594b76fde5878f54ebc183e7702632fdc0ac11e8e0e194c39f392fda75fdb469a9b4e8e53bce8645f87;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hf9c02f8bcbc51b893aba4086c5de8af2f787636f661074b1149a6a0a1be410daee2e7420bdbd418e6481e23b6ea2e6fdb732a10cd4f286b7549f4b515f2173063a3e1e76694982aad19cdca264a67b6f084c61838ff3cde1ac45b2552fc42a4d1bb7b235e0b21f376ec4dc509f71a72e8ec7d6e7b3274e40da28877a9faf4b7e3f8fb00a1b569d898e228825533fcd5216f7a545c936d138ed35e6ecb4f01dc59fb3a1eac325903a82b528990becb112cce4a82438fb17a392b26209dd787f93edaec57328420c717c34c4e912b71a6366ce1130c0584b65f10448041d8664b5c9a23abb08adeb6b45762e1657b7a77fe479b5eeaba56b75e3d028bcc416baba4ee3c2b46ebe80ae8309ef2962d34c0d94aac94168f05da39381af742865d1c8b3170cc1d15fcd35f9a4c4b289bce219e3cc07932ddcd8e406ef68a364f808532b480a3ac15a0aa2c5529562d9d1aceb10e99c32cb46e126b959dabea4985a43999f03624a4f402f6f8d1a885593598409b61af8e1205e2eb3b2a057807ea705a0a64ca2a509e0c8a9d4d03a259803c7f3882c1d19a98d2a64eab8a65bcaa4b9abec4f0ba61d172ddf6e816d2280e1aa47e4a2a766a99a058cacda8ba7efcf4f763bf4f9f36c671f63e70a1f1e1ebcba0540d21f61ffd64f7e277de6feda157b761b5de8e58c0fd166724a3a0123615cc878c292b46df63bb5ef44c0a2a606a6893ccfdc2c928c40e3fdfc81fceaeb454164edcc1c39cb3a33ad91e5fe18edeca916bb931dee6596249369db191bcdd6585129187b5b8233c447f0121ad9c181a3da4f9d7cfd495425c0a382df727f4209474f6a98ab3849b58e5bb3bac543f6d586bd896d172ce9d213facbe725c0d31cdfcea200102cbc7f22d5dbed5a7c5678e9c4de2dd3446041e296f788ed06da71f6d7d7de957b6116161d7cdd20bbcc78aac2518564f69549ce13afddddd585868ac3e56bcc1632044c352f606c0912fc92580114b79075002bc1276c30bcff25d9355523248fbe35d3f5a0f4a22dec024c70fc84da7afb114e91ed86552d6c4e8c7748861cd31a9d521a002bd1d2025d69bd793389048ffb2283f3838940bcf7edee3f438db39cb16180a6caf8f382a28c68663b1fd66d4128185ce28c5cf3daa0607102784c2e4bf96ece9b545896831e924c4d5787e19e33a73f8047e4b0deb0528b35a9e9eb0a91f3f99ce13a3fefe6d534450e762fa8f40d6a7300a736ec3ba0f3b6b1c5359ec9f9e4ae2c8a41d8807c92af86a8b7eb098c7e590db457dc04dfa38b67807e739328401b47b68ff7b002a7331d49eec0fb32d488b567146ac35df8af824ee59a0445d2141551f3b6e2c00b6d656a6598f86ceede8fbceeec3f6a59a1fd4396f24b32c7348bc7301cbd73bceda9ae8eb4200e3b80c8e9791731c43ce80cddcf006fad28b5d26fb6c54784140594be673bc092069d7fdea2eb7fc854bf87bbb43d2f573e146b829ff9707cc993b12474efeedfac18a222ca447fd938d13303bb7e59110a4cd3ae902bad71bf3d923ca2b28cdaa89dcfdd1fd1ed43b84eab8a1f83b9bfece209357769cff4940d79c6aa2a59861fd3d8bfc864b2d597bf89a1603530c1ef1000b803a3af7627c24de251756e53b951df1cb8e6cf79377bab28caa4b4aaa2a0b197da604e3db85ee3504efa12ec1d00a584a7ac2a24922346f92b3a6d8c3124f66e3a91f2670ce9d5c537966db1c3b0ea70533e20049f297a110daedfb953b6eff5f804dabc40eb0b667d99dfe7e9f9a375fddc80b50df0b2dd973df885a84f0a535d43124f1736f8bb20b9a59cbd1271e363;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h53c29618f5c0aee42e29d54840a3d2f28056cb7318e03ca73b947d86ce9e8ae5fd4c20792acd3ca62254e0ea8f02e5f7bc4ac40419cda75275c16cf85b99a4468b52125f54cb902891bd1450a2591bbc7e6f69439c0609d4199341c111c050643369eab4f582eafcf0273ece0f86b84461cd2c2991b9efc809b79155c8dc3457336a50d8e86ed8cd542c006fcf49a2960f5c8e4345ca1034fb1cb598004c76f73ff0c67f21dbc635430d778725d7eb7a3e6f3171a3c95a9739b1176533ff283b89f99d300d32a5d37c22d618fc2af0d96487e90f6894f1f4705d54cb5dc9730350fbecccbefa44532420284224b2e5da3a98c13c8f756d62944307719af6c558d8e28c8dee886c8f0660cd6cefba746eaadd765df07758407e51092e7b717884a51acd0d365a5efcab6f881b3866467876ccd5dc197d678ffd4bad0b407660c68af6da4a9c5b51801e0e069f655a93697a5e93fd095b04da0d0762a76b5d0d89ba596b8d472025916b26cd4d92cbc7cf316a7a35d68dba6a71fdf17e9809c67dd842ae7abbca27d76a24db84c5b53f8cf2d33c67e87c5ace8ea33d16e34d604d134b31ac19f69b0c258b7632cf0cd294d32c44f2dd19ac4eaf723e14793fba5389ec447071874822273d0c3688e4bca14b3493d35e29ef6f9431cb8e541e7d9aaa2c0e3f91ca68c45b6fea42fd4ce362b9d2c0a83e5054d1c666884ec3c97b727b6c5b39a380b1556f84c50038b3b5d7e52d5d426517c2a77c1610da4c166298d2c4588e599c9e280ca6813077ba3be45e2621b88deed080f344df2c5063e260fdffc4e9356193e4fdede9f4f1778bfc0d39140da9f32f1eae5f033ef8dfcf9d764f7427b2986ccac28ad2bea61e659c77c9d256c7025791f826634360c89870e916ac8cbe7aca5da28c8000790014b2dd6941e49412408bcd072ef2198cbdbbd1c3f82b12b3164c344e22fb52a393b502b7f6863bec0b38b7fe0ffeaf7b36ea8c2a1620e5e875cfc6242aacadf529896223482d42b44813a7a7181a34cf98ff0002ceff4cfd80b3998d2b0308a6bea578502565b5c09331be9a329a0054036df2548c766f456fc6fa79dc2d050a9573d88baa96752637578574345169d491ac3d22eb669efad0d3b30efa2cdbcbfad3b538fa80bf1aacc5af477b58e7e18ae97ba972e3197786f5221c54e99c8fd24d3dcafb9842832b924d0b68a9660360c95a342df4eb59b6a3d2e16642a0ccb8216556f017d8036275aef40f8f2ff7cf0af9c4e28f3d379dbbb989905b3952f4a282e65fa3ad2224c6cda7f1ed3ed929b87fca1416fe8378c73df20e36d34f32a67ca36c21412dcd2e8fe9a9e54b745019955cee9738356e8a706cb99bfc697b46817fe1f8189a12b80a30169eb07928d15444859cb1c8d44445d9947e14a989d67efc2f608b6226b0b01d80a8664943f13a2ad52bb47a89ea00817b36240c3118b0add491942c52776bc3963fe8028f25cef45d3ea59531a26fee1d9402e701c5751e237b16f97290f2cb98661476dbaabda552a2cb399877562de58ac213f2a3735d16de87ce625fbf5f3a4d34543aa7f2ce0027a6edffc0176ced2d3d04a4b46536932843356b4562e2a5c61a4c0d136ed5bee66c0f8e848fd405502902358742a86a5fd4043a8fe8e113a0af89290bf5ab3db6ed22dd88a5b77b27ae8356b866beec06cd26898e8a6a8e34b291b8be93235a6c5240742f662a7408bf124e36cfa24e155905a7b83aeaf970c83a0dbae4a7c05cf16279263a06cb0d964c46c8bbb173ed83dea008c12e532497d3ef575fd067d701642e11c4ae5c141a31f864;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6841df512138d9c038c0b2d6e451e0f684e2ddfa18e3b2cfc60e37e05338bbbf72368041d666baef1d8f20d6c0c6eccea2d840b61f835338a34c6d66b3f51f4e5b040217ecb9dd897531062f84141415293645e81914b0047f73f02793ef9a355dc2b477224cfd78fa90379d140c0b19f78b54c9e75926daaefed1164fbd7e036f33a68d3ca3df30d95f6c2cd2289500ce9d4f8716bd3d0b4b1ddaf91b9a0a0f6e7b5c5ab4f3a74fbc1289251fe751f465f47d0945bd3a1a8d4dd5ba1a2763170d6ccd56d1b7c531d0e92f7adf5210e0a57e9d29a0a81a503659b41d508d3a6d3550590a0f4794e8150492b3efa0e5e531c90aec5cfdb50d8da86b3beefb201dc4edba8bb9a8dfc0d91af9bd5ed350be83d47e9c424c52e8fb934651d902720ec2f361b36f311300da676611365282a1341b283215ca4b767513ce9113ccead873a3773d0fa30d61549a9886cc9c15489dd9bc866c7b30000fb1b3b8a5274cbf42ef1ed26995d34276bcebb78f74792f257f2d069d9575736c973592133c3e7ff4b2fc8cf374610694087c54b017441320b8a57da762b56850cc4a8b41edb9b61bb837ddf85df07e36a0f935df8b06b969450b1f911576afca0da64245ed70a0930977012e2486e2cbfb1e2109dd54d95bd056ca5c199f4aa7c80af70aab9360730f60be9b242d54d023a3b94f2b83a0efd732a87a4dd205df2e5308d6399f00ddbaaffaaa66f48dfe8348649ac2478102e0db2f6a7722a6e40c6cb3dd0ebaaaf6395a3ad573d8859415c487ea2eb781e8c0ed289485a84dd7f9256a23741c429eb1638c34f4c06277bb2b44ca1df0515cbe50a7c82dde8b13506d2462e3649c610cb2fa550356189377b1490166626624b7de32301aff740a9887f04285732e2f2058fb1b6a5583372b689111fccb8b2d852f318939711b91efbb9ede74604b26d56af2c4a42a60f992288cea47304aebdc0150192ea06b66de16136957172a802c8f7f3dfed9213cde899bb5e725cb55d3ccd4b42ba45b24e4da83316c2cb6fc8ddf973ddf70b8e98adcbb426ee4cc76cf04775aba1b749eb4dec1bdd7ec096ff9cf9a7ce1a07df9d25b4bbabbcfadee7ae23fcdd196c2c0286487639b9fa581123311ffa0256df79e01799f84860a32d0cb12f03302c2702c7a152a3d898db20bfa7a635e67ea59cb8a2f5c5e657ae01143d122c71e12577be025dc3a2dfc9704801017fffcaf4b76e2fd3c7f9827dd529759ea01bd0b717496f2067af1e092f4ad5b6302a18a6a6886fccd99278737da7709b83268d76d26ed25303bc2fc4e57fc23c32a6438a279845daabdba605a93fa0cb8d08e645d6921be7e49f2680145caba5e8616ccc4405899b199b96ce4b2cb158a89629651f7958a56f1d8252a68b54911bb0fd65a8a5cce4b83a841c04868a3392cd3df19a46e2f788696db6d1999569ec87487b9a6c6a104ab4fe07e06103c25e366086f8ac9503580b2a469bf18ed2f1daad06afb44fed9510e74e9a21bac1bd96d99c8b00d4537ba3f6d1da06eed326ce57c822de74ccfa599e7329bb161fc72109a28e9c9f6b5175d27f24ff982444da762054d7e4d927a129d4d670fd3caca6724901329b2c16044bb9cc46c888b20a883834f1b9dd2bacbf4323a8bad2405e318ba3278fe6fa2202fed797a86f3bcc8f5e7c59a69f89b1485bf8b9a889d3e9e8ebb9f3fb58c9cdaafc707d5dfb2749f4f59c9d6c447e87fb9028d2a34966dc529dc2c763536fe44ec78bffcb8a419f6e394d4f7da5f1806aab2b9efc4ecffd193fb6130f5cac6270fa9b0ebf547488132ae82ccf075214dbd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hfff172ec192f1ce00e52aac1b5a7bad5a0f5b09e2fca067330c31965b4f719ddf938c6ab0ede26527b2ef48583b5d594514795e0e6101c5be069f1af24b9d464a3ab69827c606cbfe5515898fb00189abfb8345c226bacd36c66f38deaa9b3cad8b51948a6367b212fb3fc11903435e472143708530ca4c56d7d99391a1fcbad9bc2f5863b288c1b20520a0196b1ed06e7c981e8f0e510a793acfb2a2865d76958122807aafcf537b91b1e4c4f50245bd71d48b9ae3fdba5432829e73e118c4ec7b23edb3ae18049b5f80c644c967a91ff44f4c6c543df242599663fd090a21555c6fb2a7e0228adda09c8828fa4bf3ae80f18b28ecddbcafc5a6820ee559f8c4d78fd56349481059c6cd2505bfc9eebe866c5dadcc23e89891a2d81b0863b63c59b51342a5263e0bffd22b34f34853edd685a7fed85dda53fec5800f0323ba195aa0fcf38e96860c10462f75ae1cf7dbd98976934cae0322aaa2c85afe93cfece5bdabb15516b02c1df95e213386e38abe3bed8b8501471f9cbe159f11711519f965b4ab15d01f1c69e3f95adf69c69b1371d5f8d4618a8919488bf096e47975db6e5f0785ac42453569de92374bc37939064d0850b56325beeb97c16b7b146905dc26836acdeebc768588d0b1f8be497c5f8236f5332871a0120a6b71939e9c35604b9c35471fcf7c2c08d1b07b355cd1ff0eba6c189c7344e252e7b838a5311f4f61680b5d477b48dcdb1466d9cde157242728f58b4f4e805476c4a51c03fe386441fa1b1afe4eb5097fb9aa04fb262236b5fafd184f1789ce30cde1c1fe9a5b73f26866b036b33efc1ebed3b6ddb247e08745fd3d51b28ba58430cc8840812b1d379e67d8826bb2d9273326b7f12e343491d38cb509356798280f4230d926a5afab4d593bd343952cc7effc02d5ce0a9434037492c5a86cfdf62d2de2cb3c31e3fd481c1e6cd181c06c6e3bdec0634f3210e3d04e8437406a6ed040869392b68e8aed528d200151e58b0ec784a720d72506ff20a1a743b1ba374dc1797cd705ab4ddabb377ea05381809f0d1b7f81f05b694712975d6fb42d71f84f5b003252a179ecdebd0330f49e86bdf9b12406e5166cfe235adbf148e407ef6f343bb8db8585f2554a2b6cb4962b617d2c8bd7da0194a1a0fb7043cdb0c6cd2cf08f201d3eef7d6e0349c652bcd0a7332d122b106f2c3b1c669eb1fb655c3edd830174ee255886ea58fc3685013822847b5e67b20c65506de1c6e22be43d4d30c2d2e685f0f60a43f1a6ec5cdacde88906b93e25dc6c9b1ec9734404505ab4c171b5f5ec47a8fe9d251dc55dca36f5d4f2524b100e4e4c1847f212dcfe2f703ed5e420cb735106cf4951e88048053b90b419b38acc57fd64c407215744cc3b7626bc0c51cb073ca8463aac39d5de70cd1d8250f34611ba54d37d3483c91067956e9d6b0a82e96dc80f47eb13b7accefe9fa7e6f6077b12ef02251b4399ac2b4158f24418fe2676c18b778f213d5f420e07d1ef6f058e7b11a1c1c0530dc61e910bda9b9f52b26ec265cac72ae24bab6979cbbf18619ad03431a645a8e4f5462a524c21c1d81af5446ac8cd3977e81d669154736e74f8058fc27c95f8f25d063e2d645d1338881948997186996dd255c154c5fbcf29fcaf39402d316605f6e9576f62e72e4bb19c060b59979f6f34c015a88fe40734f15669416eff43638f1c50ef1c8fcf30458d657e9bd89f7b722c4ba1e368b8fd8bc5096157db78b1ec14c8f0cf07f8b10d28f594bbff6788c5541def18a0a837c9ed54855d6adc73d1666e848860094d43489e5cb1e4368fff370f47d6f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h4a9209f0b543e5967cafc69eb8d4f1a82598b06ac82be0185c4e03e48d0b6c7548f4c77b6eaa50d5c8b4a7248b42ea1663381f9f362b659fe56b89838dbff4a43c9432a13bcff4ad290f88327da4841cff0a7cb9bde9acda8295154869668125b4ccf5050ed3c80a368beebc6af34f6cd2893181feea70c6874e836756a437e72ca4a703cad76c9967d01764f37d80fc8533b1a87c373aba483955b9028bc5ccf752a79cafc153cbb8293de705dc0a92f3cb2646cd046c271676d8de989b79a780aee520cd063e6c25fec32786f3302cca050bedb1940084d339192b6e7ca1e0944a6c4a74dfc57b4444b5a7893f85a1cadb00b0cd6f3d688f8da5094c1bee8afc58c47417e35e0794b058a835a60f00a1fc9e79fb49594e21f5d8886ad6e553534b33864a20f83322b3c6f4806c7be1262332fdb3ebb1bc309916e029bd64e61693ae109bcb96dd2b2d1fed7896c352c9c48a20854eb8b3338238e1c8efc667556458d6caf90c8145cedcae4023557cee05f08407945fbca36987af7b8f1e23620c50fa84851edafe1d8935b2f1fd6be0a0f3c7fd585e0f5fff734a3ce49833515c959b447c3e66dfb7f3a28df36125352e39091957ad9eb36af3ddc2f439de9c456e9a262224794eaaa96cfee83eb2ac1f69c2f545e463cd1a4a29fc7f012787cf6e5421708f40c649c79411d4dc2c19dcb4aa303388f7ecb4be23c69643a12366980278655a822c8b3abf65e14812f729f542d13821de142c526b99b6728e9064a189b8573103596918c26746ad6ac767b1ad700f5e2527c952b34314d5d318196f1b7bf43e553af70c4f6f70a3124a140f05306d724bacb9f14664dcc4581877478bba715b937dd27f7a914ce33145634a4839f477f6646ce7caab6b294896f03c82792e2bd9f986c1fb6caad6393d0d30447e0065832f0fa812dee6def85f9206d040532ac1259b7cf7159872b4be2d4b89d7b8751a30c0c5dbfe4fa36021db9b958523839fbece95df6ab01a82595f6b04fff8371dbe678e55fe1c01d4c0ac83cb3132648bd4747274fd8998de0b2455f7f78fb5a08f1e4ab6e2e99d8c962e1c8fe8cc77081c728960bed009d77d77d468cd57a0545fd4efa8c697cc8a18965d81c3d4552572699680fec5707175a9b25eb0dcc3929f1e3ee319a5b58f568eb3772fc03580e5b1c993efd918608cf8544aba8f518e40cf68be6033e9a01cc9895b34868271c8ba44e7a4d7390dccdf7b8bbc4c3f03b6d1d7f11b20859a57466002f6f8d967ef68e23c7289ed4905ad4b101f161f8f9e40c3f5f3a858332e659328a9065c176bf97cfa9abbcee35a078a25679b9591f43cf885e6b550f15e3f452e67ac96f4bf6b8a62d9d6e0804d83aca1abfe4d3541891e85ee0e2722aa9dbbdffc4eb3e382e52ce194b418711780eaf1114b086b3215bbddf76b6825b4eb96e5959ff444029ce678dcebdd906a23bb4e7813b2e4b26520c15962184768c48e6881583454353391f3333fd1a828e2db99a89852a76999e9378f159c2b4a8d8c2368bac0c036393356422337e71f2d8ee5031f8366ccb2cc4ee720d5bb81d0aa2be30b459390ca1f82b4a53df26197cdd30626de63d0b472b10b4365fecbdb188f069f4b98e5911c6531c2919488b0933a6abcd593127539357b17724e6a04e59857ab4a510e98ca361ea4d06845af8e067e74b5e9826a113b7655fdd86ecc07b13a7d4d83caef8930b5856cef7d016c833fcea8c4ef0c701065cb06bc0befb152d2818f412344619569bb42d4ae96a6c828d831a7eca50959c8f26260adc27f4cdab8d8d1796e31baacc32bd5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h21b62a40735a5df4d7c7e0f1be8c75f259a8e0d4945e7f51a0b26865fae98f80c184b1a802c06f5403cc37ac30d7b3d7ac4974204d3d48e03e1ff2a6a3b2321749d5fdfc937d62dc4b38a9667fd93875c70afc9c8016b2b1a47e756bfb41f6a6119c740b0c4bf4209df2e6c35254612c613300998f46beb0847af87c3a00d464aaf0c3b1c01310a6750d0c7a272521a7600d18b8eab6537f51555451d6f4b0491f552e56e98911d850919da6334e21688578f611119898eacc0cf36248b0ef3d2b859ca7e8bf83d39d0bda6cf0214fc86b038cbd2ed3a1a19eb6ff45a37adf50d2e85a06b8dc598cf0e2595258348843ddbe9503c1c62c5eba21c8bd2d7ea7713341cf76e073ebb2d7ef70f08a7f1d42e11d55486a01be0481e61fa0590af89c98e695f587c9f5dcac7fa38405bcf06181955725a3fd797c8740c8d3c088ff8b1e0c48ddab2082be273cf6ac629a1ece11689eeafe24d89a903a3263f8908a5f215456ef5e67d5dc913a8ed84b5abd60d760ba0cdc1e6de9db5419be9330e137899809bacf21a042b7e51a831059b157d507d1360fb361254cd7add6cf068385e33ff80fcf28c400f5290e2bb7e421f581f708564c024d533dba9a89ddd642bbde6808018822651d1ec92df2ca2fe3898c4dd3c53d6dd0a50d830db807ba31798ac226934547212d68a6fcf325cecda04f30797e5d514d5c91210c6f1152cab4aa25b5c165e167c7b8a6a1bcae0cab26886ca7b709541d8b7ecd77b7cd8432ef4441fe22351ad17404ee58af658b93de852f08b6f66182cf4772255e850c4ba8d791d12f66c48a9c6db7b244f58b119496f40380cf995438765718e34ee061aa98985ec48e730162a90b999a57827b0f4e5f48f9cf2748a536b0cc701cc470a20d911d3b6c3c7f74f9f306487ca0ee593f2a748c63ba882cc7ff7bffe7341a3073d5da1dbc0bc865f189f05d1d7fc591addcb30fe55288841de9f6689807d17b82f5d1becdb1614b17eec2bc6541adc14923352baeab0c4293513d3bf12671b62e7712d41ec4e4685f9db67e20cf1e0a8f85d20f1bc13874297d035f3db5dd010d63b4548e8421bd11947899c48bfd90788aee551f7e4bafa2ceef509dd9e89350245c41a6c6796f1529458e9da38320f5b467744b4974ce8dd394e154a92846f041576f8a6ed76cf658dfb1c967a753e720786f904e5ec616a3707c2e4cea16b4e9d0666857c9575fd8a7252eb60cfad00e51a1a063a5a731232eb23406e5f3fe9a3a95b223c2a70b84bc105dc54cff43864679aa596d94d1a91a83269acd57403b9a1a782f7c03f40fac580c6982640c5aa57b5945c8f5687477abb2437f99ba7927127898ed1ecb870e7a27941a4a5ec6a9e9d61b05007b360469694cb231a84f2ab1731c76e2b6cec6c491fff94cebb26e6eb6a730a0600de0599cc63f4e6b11f376ad0fd8af7e700db75c1113809d46c501c047eb7396b9e3aaa99f72a39643b3cf33a0cc4675e33a2dd9c78eb8a22f1a547e9e2d00573f47b65f68283a7034a8b058e1e6a3b66658bc15693acc19d47c3f961fc8176e3009d7663ad2e5cc6b2d00536b12da10f9cca8870235c230ee07dadbf953337b930b76b94e2a294b87f8cf6372dd71cde1bb6db0b73090e21a0533af53d5e8ef7c5926c22c1810cd3c477d2b2369a35bcf8d3e38a81e9cdc8f28253f17bd97c99c1465448d09b578b43e82a48d2ce87a1ec1d16e7b8fb9890090cdfbea742f842157cc22b46f3bd553ad9cdae35febbba3d759abaa0ac0bf6ec3225bb423bd16048f06266e7670b9652b75b588ee342038423f0d11fe56;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h88f0b2780232a8b9beb298b230c9506188b0efed78274fa26319b98060eb92347ddbfa78f02c8b856c004cc85b1ebc7b7866331105e29873087d9e0e3d84e3e9fd7c6e5d9fd148cedd139f5472e83c4accac7c21c717daf6a24470a80f7eafb31fa165f05222dbb64a5d725276ce76b9ae2bf07f175ba2f1668713e618980ed5af4cf69b60d8f24b481baa543d4fdbd747ed8abe3a3a8d1791eb2c6a8a59fb07fe93d19d7cdb316e2abea91487fbb69ea4ca4dccfa7d78bf6b93741316612f4e9f746d40c4fe3a936ab8c3c9e707d57a8ad94aea1f80e64299df482876474063a2b7ae6c34074207dcc2eccad05415f6ee0c75d7c20801059a3e1bd82c7e117e10b54d7c1aee32b8fe2efef9f9aed33526f69b2f6f53622175cc3af51b120b80479222c511c66fc4179cea8348c4d71977088d9d21661068567b1b4e892207b6d47f3c1da2a0086c61c45fe847d720157cdc519b45d635d8b9a74eb605ec6d9acef60736652f20367a12cc72ae59462393b62a3c821198ff6446cc6560595950923e66d5c15d61c371d3ed77aa56532d08e24bf15922150f28c78792dc3fa497d2fbd4aa4f56f273e5e34055a0e63921b2f802c546cdd943cabe458e456474fd3df1c8efdd4f1b47fcad889adb3b66a5df063b33e0195e3b3cd7558652702685870a9728834df9ca6cd910c9130a055348bf5f04edd947a1f8bb16ce08406150c2b9db376055be0c5df4d0c5ae467f4d65bdf44e4a188c78af83b2ce08b1347fcb6827b1c37a7f4de4b31ee7a64e174ecb3ec754c119b41b905e8b8847a3e7cc0d8eb106ad7d9fd07a677ccbe50efdbf31ca539207baa2f5fdfed7cbf20c72d3af5f84861d67ef27d65f37660c3109e41be86c77d0076b3ecffe5314e37f22d02a3ce1ab9684f24ca5c7877e95c9e9e5cd738f705587d81f55b8d4657ef42a87ec671d7412b18416fd13a617d20908e7fb349b56d843224b0407c65939e026433c77f42dd2a3cf306326fad98bdd356794f088ff54f66c2fcd72fefcdd6f45bf5145227d5a25f2146e803cd52fe927350b3aba5f739b1ca43ec876329fe2716e49888742c5b4fe0d6154d0d8c25a930ce17f57892539450e7fae016196b3aa297012256aff84d500c57a8127113868f3975d5eea73f9068fa1f207c0abfbcabae68ec8d5857485d434c64a3578bf144ae72274de483af030636f6475b8e0eb88989b84d65df530451746bf3b102e9a37ca7da424a2db201b8537070a28829f24d2f622bbe5dd90a39e6200fc0c940fc7348455868aa98efe2aa69b53233ed68fcc1ecb67c5228999ccc56b1ac4b43b4195e87127b781222efb54a443c6c8439141420a5952d9a18a89a4dbc135ac39b8c7cc465c153ac7627a3670d5297ad49e63da94f036604b7ee9c7a2361cb36c6c174ba5ac0eea338a8880fe431a00a6a466ce92052a4f8b82f0e8e92b697e178194a1ed2d589263a28e6043c32d322aab31dfcb59b0afba9b39d064e2269dcf603d48469bc167c2ec3f776c27118c1adf59321e85f634641b8f16a922871b517801267582dee618f9887b06d5fce130f3d8265848d433431f7114059c74a5eda78ac6e965ebfa073b88fdff708036137153e409fbc744dc3ebb07c75d35947d2af13d1887aed0f013560b298ad1291dc4ab79892d4436b2517e3466e77fce84bf4b0cef9ff121ac818158d5249fda4f9bb051325898c189eaa5d27c63bb162f3d9e7fe1b4f45be37a99fa73ba2d0156a953630ca06d1c90695b3c75376201f5693bbec5b40b678b0a351e64f03ee126f57d438ecd9b4411066cd1cb98989b903b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hbc3d35510cb079497236163b3f7ae180eab08d90af743d456bc3dcd86d5900b4abb2c6fd7c633ec0de478ce9ba80e1105e1b80c6e6fee2d1204d5426583db70712f450b411e4b200165c1b0cbff19c2d9d7bc7aa192f1a5ea104acb5e8c83813a97e599c25d9cfcb0f4405240cb3d8d32c1774a5e45b363c5e82a365691bc1b78bcadcfd62f4f9a06e9901a77387c5728cc8a28f82a022aed58695bfa9813591b46b1b9ebcb09927814eebd3380c7250d11b11f9deae61585d53eb26b27e090c4838e3582c2e252f6b15596c72907227dbff981a829f20cf00bdf341d60c58429755ced2587c98ff1c5d47bd7d948ea55e88b37840165c8fd992f8da32f654f92f24955dffae8316299ded8d5e509052ca88774db6b688cd7a77c662628b9448ca35776139d07fe4744398afc5977d4a5bc0c631670d6e2a47939f1445a52efe43296a21adff5fbccb18bdaa7d1b87bc59cd247de193185c5b52f381338b9e873219ed1dfed83d3600f4e71c6dd618c29c71681f0fe49c215541441efddab520d7110136e06f1bdd05807583e5f85b16c81ea48d4c3e1fd5434e8bcc063a8b7e22db1e1175150ad4585db1cf6d9ba36be52a60baef2dd5ef26f75fe11f31789bb72a9f2ee87a104136dfa413a1a2926381008dcfd5f5d824de364c46f51ea822e33bb61004c39f09f9e2882abd01edcc760419a64a2a1457bc0792f6cc126eca9e81db901a4a9e096d419dd82f59f1b35948ebe6329ae8c790af815dd18076ab0defc75a45fc9b56b5c0f7c94bf55aa297330193c63df41fe4b2a0266197bc9aae456aa731c3fc0e5a59c980f6c94676e402579c44aa12f0f43fbd4de1952d02c89a7558c028028359c23de43a032cbe7b9cb0c3d2ae35620ff3c129d8e055cc159a9bf33e33db0dfa4635d7cc9a610b181a1f85ee6f8f4dfcf10ca00d5997033e58b81c0c3680b2be240f223091ad9b5a943dcc52d2eac83b1412d8d54a68c1db39c283b73d6ee85849fa746a3b29163823e317b5b3ed9dbe488f3cb1c4ed4ac968855bc389ec2c4c0696f703e9a6073779cac0a178436f0aadef09eb0cfbc938a4c78038f7dfb4f638079cc753eb560229ebb5bfaf17512aaf2c19a0e6a2ea07e24bd3f74a3075c7314056c03bca9002cd86acd2c55151a4b20dde95d88e9a060e4fb61d73f1df8b8afc818aab6e425bd8034ecf4831cfae1ed452c32eedb14f4c236aa5f6ac6498b464282df51fbd5d1aa19a0360ca0e6cf332b89f284996652e0b37fc8fad73e4abc182d86c69270c292f1913518ffc08648a30036ae5709369dca8195d43c583f7076facffc4a652bc36bc38eccca5127188d6a5448d538fc59391ffddf6a25a8931bb6e50ba1f6e2d4648e7a1a829d3262a8eb4ea41f1aab36c06ccabbcfb478dd93a31a93381276d7180778787f16c7d4c8ba0b12ed696e7349c3337f7a83ece37ab17211bd235196d780c0fdd851c0cb8de32106237e51fb5ec239ed067a8306379bef7e035d42fbc01128e9967d975f746b2adf209c51e62f5e21be88c9de5b0a6575d7dd8049dfa16390102dfe65ce2183c865e920a1f76845408936992192cb4e4096856a3ec12f8f1e0b1224300bfa4165c3c7a5962473216b4005197a4140603bd9bf726dd3542dfa7788bf9bf62f5a063eedbd92d8e3639bd9069a703aad50c8c3896f77133bec693c1b9d91a5a67e69350fa693a78d40351a1f040d68e8c183eb1fc9e4804f7f04ab44eb5c066aa09820324cfa3d7e4ea87428c66056c876f7ca347d5105caf32c60ba95f8ac4bd0cd676f70f07a02026feae97ef75dc42530fc18b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7d64d6248ea9699d533eef869be6b6797d087ee89282c8cdce54ba8e88e7b4ee84c37c82038001e942e588ef6bbe744b1208e6d54844f443c7c50f16c9c88a9af8fe14d76683c1f65d7d43895dce95c19ae762b459b191b182cf5654781d0d9fccbe8ac5b5ebb6d61632d92ccdc5cda2ef60c88b67a468c64680c20fe192d6003833ce1b062b19169edbc7895e425976042f790e018d8355aaefc875a08b1f90de0578802712ec716cdf83a72892351e79b4d5e6188e3e8152c8a9756ca02dcc8f3da436bdf4abf1f87d18b6fb79b3a32b40eb2b69b49830545692280a33bf21efd9889c16a8d4e867204e377c65ce96fe7e5f78e8772215a7d4c9ad1d80cfd411e95b04cdbf3c61914aeb1c54c66668ecf629a6c6e59d38a4039911f78ab32051afa36f5b3cf4710b27c7ad86aeceb470d92ccb63078c2efde59cc73326b29dd2c6fed00d475998bc39fd17d18b1c4684339549bcc3665c6c0e72b7ca4285ac2cdd53a4caebb4091c4750df125bff77e2252df374ad029baee80fa6d2d82f242c292e73431fb5686d4625d78691eb94d1b3159873fa7cfa977ef0ad72d8c9bbc1e3040c589562ea7ce0d9b337ccdda12b06aa2c068764411f5674d5a3aa5ca0d47a2bbc8136ee6abbb0a6fc3da45b2cfdaecfe366ff6df386ff68d4103e374e6f02913a728298aebb228b405eed896c6c9d98a8993e9c2588a0dc684080faa3b549e278c946f70a8bd9f475e48c42f0fa8695ea31735baf3f09be0b25e622628c7084640659887970c6f8b895fc983c4f7dc50d3baaae62588d06cbcaa311abc3d91d100de927ac4215439b839519265091c8a517b23974351ed50314afce2e35951f34dc0152425b18330220667ec1a4a00bea5e5801aa2f9b8d96e3f08f80fe19ac66d80610a43cc1c5e67498f467146efa69c87d32f638d251780be43385fcb97ef18b5d80cb1ee78239a6889c924292b5469973d13186fa1c818eb401850fd317cbb7834fe004e7ee66fd2ddee5546d176ee6281b0cbcf94705e721014b42e906ffeb477a97699c4294c55246ac6b8b52b265fd91a7aa58b3d1d4edb932e713506dbbaba8dab4acbe9100ce26a7ac9b500ea293fa62831fb6c5e80468cb8cb379cd9698db842015611c34db3c9570d498627e31a7e0a2e39b5b1741128ed84360e7c67215abc8e41959f4f277f3893819006fd37e5ad81b6b895b502fac89e97b6f698238b53a4be484d4997738ac0dfef2cefa4f401bcdffa4f6c440302f0856c6bfa4a279ba3487c072c7a44fca57fd7137c46909db9dae6048076dfbe98be269cdb27af30df9d972a32e36657e5b19a639d8fed20b3c3d458c1945752404bef1bda5e288210025fe74adccc020bc7d7caf18c66c08be1258b458a03d683ad7b2f2c4c3e66d55c610bfcef55f24dc283f466471f29a73234baee7a7d276371faaab0aeabd8228994633c71d04715e98907ce8fe944c6e2a8a950362432fa98af19d6ff3a5365b9d3bf24364fc68134d2cc17c467e749d519e231ea86f088020fac1fa764502151740dac90c809d0fe957e3e9c5ffb0dde4565389e6c98873c8becad05fc7e4e0d56de1ff4720c555881a16adf991287fd09f2a11dbb96c3b68b5be2e002cf20166ad6688a523e11ac28957a6f0ff9917ed694151ef49ce4ae4b0debbfbf20c6a1b4a6b39e349cdd4a9d292e645a7cd7feca49cfd7837ed8e8709a43deb4ae5f6008501233e79844f4db981502171b39d637420bf569ef00bd493c1aaaedd7d2a0a6b6173a2147efd77b95f4517b0c3500a466309dcddd0706320736c8ab713013a42d71184d8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hcdc717bbd1f914506555a3117ca999e708a4eae4cc798ab1f8eff716be2f8494f93e219fdb4321370e7c7c06ca71500b89b3e398d28c56a981932f97ee5c3581532280527151a7e11f0d293b25b201c2bf7387630e09af2283ae8059b3eebc87c1ebf0d1e09a791495aeae1d05eae6097ef9ee15039d72a3ca329c9d3a303f8c0dffc743a02b07937b063c7b916d62cf5149e9cbc72cef0f35a6b259d5af1de99be63126187f93ee2342185eb9f893e44559e380ca1c9a6fc5873aabc5e84aba0396f360fa517a17c46c67c3667b67e9384a77e73f1e69b8984e0def9a3b394b5ae8796186669d5185dcae1a7d7cb2e04fe8939c2ec30f5d7111098e044841afae0131c36174d556c57e99fab1226c27396600f29566b7e37a5dea66ac3fc11295531f6233ae5268786a59632110ddf064d772d1f7f1b14273b68dccdb434400d0c3901288d381255577344641830ccdc487cf59b59297706e7778d0cb395b594172c4555ade86775191a4bb5f2cb6f8a562d1ef10199e2da9053c473099d5f86086b86a82abb14f0f4671dff6b156f4af029412b74f45a3c5b92120cdf9f7b43f2c9f2b3d1fe8f4dba89f890c69f23a339010ee879418946b8ca2acba7552417a521a83b60a29185e758650805930698c52608f892b26bc7cc3d1bf905ebd4ace28880b3d67af57846453a4e7c9672555b6494ec088d6126ea0877e9f0e3c4f58de9eb2c4c54d6adb0fd455c12e50fa57e5806ea44f81696168b53f2f66d8d07c8cec9b94edd445ff899615ca5f573fcc097ae00d7efcf41d0a72100ba221f721e6323ccf46c50d02bd2bd07df4650df1be927301024bac9210ba5acd1c0c4945c912b1260618c9c4c7ff7843ba28d8e87027748678824c11dc989ec67bee3f682b16d4b880f92a74da245d2eebbe13d3cfd05bf41d09adfa55e8bbc283962090485d71c826151bfad1433713bf5df0e03e66612d900e992d65f0ded0ec03c348fef1e2b02378bf9119530f8a696f50e9d47ca2bd5d1e1202c428c2f8740dc2d897ea58fc0a4f3d0fdf516ca43647ca8b6006c1085fe4cbc4125c571483ab0adc05bf53a3b956932796ff4c69d3ac6373e72a3651eef2334892a33d979b1008651875cd5ed8f0a416b07617628cd2d323b0eb1c01fa26ad93358f6dedad224a27a9fecaa8d1cc3c28e5e10a3fa90a8ad3f85fc750fc9d94f5240f236058e415b609d5f89e9c5a581167af16e0d72e1e74cd3b6ae215208d882e28825935eaf2030c0247298b0e40bd94028bb8295d118a1139338434be871f672d36b567b3b8bbf5bbc1559092d2f3a7fe1a49b12d4b5f36ad7c42f90d80d0286d9b7fb9d121ef9756fce8b3fa8eba25845783bab2e5c2f855d6446c97f3ad2c9f78d2e1959dc7531396ba6e0e7e69bef5fc0060510c4affdc7a8460f2ed68e831fe6ae263c85ba8694a8451e745974b99ce52159fcf8ae0f82508272b515a7d471b0b064ad5be3928e10cd2a2567659a4b6822f85b4fbfe2dbdbb238f7bbeaa6a0d1178da6affc708f268bc7c3c881ada801043613b565026ed74c1736df7fe67fdfeb337c6b58d0d4c2afacaeb09ef10d7abe4c13cc47fadc09c3913188d179e789a420fb8aa4bf3a0ff44e1a15adccb480daa9532a2c2255c13588e63ae22ac27027a31af9f088879be4d5d360b28189b47ee1f1cbf897e42a49499671c824d283a3c062dfd78fdbd0aa2fd3ec528baeed0bb312b564d985cd67a565a7f90573533abcab32d7fc774188b1921df68a2b7a2c370bd359f2cc2da56cf103b8f5defdae1dd41b647819d67e242127c991e3c4ff665b6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd074b84275fa87ce975be583b0fceb7d86227e436263fc9ddcb55d402585951ec6262716c964cb569bd198ee26479b02a5c6774323419a82dd1a19183e92c2b333a7ee9a469427c6c7bda97f1bb150b1c82074005caf648383a143a4f57dbf12f91ace7630483c44387668d8bf750e294a89c3e66e79dbf58117a022f9b478fdfa270b95944951f2ca6a13ed15921b5074651121c1e3dace1b18e62dfdd596008246e3623b98b607a322acd7b460df644b5e8825314d6107551e67a9d84edcb83e0d9091f095c24fd00bdd6d9a10a2af95c874a2acd2260493f4f3027b3a248b838afb69d6aeae0fa2197c382f53a337743571587312fb645742da536eaaae48c9b59cb10886ff10e9d44b40511718355b0cd7d69279afad605f3f70c12fbc378206671cce4c5f861209c316a44cc89d850e55f301e8fbc08579e2d27af081a614b2bb7ca5a3dc309a93510b83a0dd0c7a548955e56c7e0c4e454588326db51b79c8303b95293da3b899a83243b8263000fd6e92dbd15d63c9770fc867afcb2b0d3620b45390b0b37c8680fa4aa664bf97bcb8711e83081aa3c85e9716238f7eef08f3d827103270c2db3ea7fc886c08966fa32a69f2c4024b0cac6d28147cb5992ebbb4abd7fc125596ea70e57dc7aacb50a1e9f057880db5baef3f06da9ecd5d3e6398c9bd8749b4ed16568e6de21bc98531168f51822f20dfbba582af31a253bfa2d5b7370c6a121ec2e32a187763ffaf8a47fe9635af03a1dc37e1d5a010d969304b42e68f1d081f745a6f24f62885dce1cc9157295808c4c8e8e7f5e83fd57ffd640ef905ed95eeb5a89b80954badc6894343bfb8cfa3c30c598dddd309d19ff29a3d6ee33d51aa083e6ff8e1b954c28a9c4762a7acee1b1e65a60557c5667a1364f74d5105f26e33b5e24daa0aa887499038778632d265d28509e5d31a34c81bebae2892dfec48398057482b727b5f75bd5c48ccf1cde44d4bbee643f6fe453c728305102c5ae1628707ab018aa9e53d1cbfe1116f3dc72f190de8499ce8a7470452b34185e3b2e423e7459a9898cf62b61601126427f572b2614682fd506317d32880c93ccb0c78ec876f8039e6bec2bb02fe32952c8075b00aa50f51717ff61cb9f7962f7988efe2001b273f079df2c20a65679faf491d522d7d3098a0e2ba5985df48824fd31b1a0d79c46adfa800eced36618acb78a23aa53afd206e400c37050a97922fde569962a1532a7fe61cc890f0e5fcdbccfb9bc7aa72b329141a8e7b1543cd3b94462108769aaf62040a369505435243513441f27237c1681d058df553c01fd3469c15059e3ba00e97d7b032f498e12f92dedb8ee214d77b59b7b13620aed7abe96bc07ace9ea1e688b6b24221accd3c0acd3d6df9c685ed31bfb390a09cbb0ed0f82fd94ec7c3cc41f94b4f88b535d96eb54a41ab8df0caf03ef5a4427b51c26ac6653658ad9d770231bf388a9f1a13bb61328fba28acf9ebaf40dec2b6996f16fa037550ef22f820889900438684f2b27554d8f13c5429f5cc5511345b744b3821fa24136846140152faabce43eb91a29d9f5759281f3675cddff7ede57d41814f799755567c7c01f7ec1509097c118e96d7a6114314ecfa340a0ad94b7fbc10206a2628f934c6640a795df1d2888e9ea4b18028a2ee0421a3fc286ac27975c65de67212376d557d8c2ffb4861ef0e1eda8b16c106c8b9facaa80d1c9779536aea7ae3675d3f34a445c650ba686a9aa2b861046a2df72426a5e15fb45aebb36719a3db9756d3ec4e0cd6931f5a84dfeabcc56bbaa74ff5e50bfc74b8ec0578f6c368c5597772;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h33254a9df9bc663d0772a57d51468db3f259b572e089a83aacc7a8881ff2e6567162364815e940c7c476e6cc77fe9d7120c6d51f6c1a94bb47931680b578a7e6efc8a66a875477fe5c4658abee103cc7232c58fc0bac066939c512d8861c70a279e554ffde1ae8746fc6d6c81140f3d61059c2837a9040d5341008fce1dc96e11920dcadd0f331e4fe61c4764cb0a52dce2a8b1906658598888b0e7cdd7600c2d059bb35167fb3f2605a43400f83d221467366b9dc49f6f19b4065abf008017c2c7702fd2f7fb67d692d08e85346519449f2f60b0c1bc62d4047f733be302fe78b8933e00b9f439e11ee0eb9f1cf116385c0a9f3ddb144c6f42a54dd794977f4d0338633f4cfbcd7edd75a0551aa5bcde878f4e81a9b48716fc809815db28617e2fbfde812567c6d4b0bbfc068aff006439a35593c6b9b27aac0d35b7f9aa2660a1619b3987306e76714d6907433fc30bba07eb363ccf361c8d35ac41ab1d1d20e0e1fe55c7248d90e3ff7058c81e5d6fe166c30b5d8e759fe88c548a83c789c3a3f1ccf3689e85e663a84f7eaebba2a8e5df465d0919da0c8e106e2c0d389c577ecb52c5e057b6d70d0d5334cd33d778a6f2fbc26d364175cc3dd5acd14436269aa302fe4da1f468cf48f9ecca49396aa1f2f4c2c350565212de02f89ce12832727aa019eedc81173c6abdebfe53c4aee10808fa49e8ac197f074e18857f79a61b1a769fd6dc94bc2dd4a46f50f11c29ca4506b33c1f021e1b18982d42d3a43dbdee988af3b9633fe59a5c7e9d0b48521e6ad3be10bb61dee93303d1b388765d189618202a0631958ec6f9d1893670fd9bd6cd0d030ce54d8bbf5802fa892dec1ce5650e8fefa1e3011b9c84fb4feb38abd8c0ea64ca475da4993b0fcae97019779dc6d63c0f800a29f8adb1b03033ba338c6678a81e087b46fbe1faa1c12ef3d3ab866e4ad2ae677e9421df7849dbd3023aece2fb10395dc9c66c3fc07690992fe5401af757cdd3f300c6bc6eb97835da59ce83436c2da755bb8093045648f9b5d73d9f4bbffc424ea65fb889fe51689f5989e916465fa8490d21d68a161286e434691d6b1a115e4bede04066de5c8db04fd627563c447aedf3b79c93437be7d1ed4d2724d1b130ba0a64e7cceaa86fe420c8db7ce2202e9e2d451a5d6abe8b32644e0060e843d6b3b1ebb0b86a2fca96c550e9fb1b7766bdd4cf4071626792ad6f1890af634982a2bf65c4ac098d040a0184b09cfa65285474e4d3c8a89fa143c5cf7624accfa58b02a2ec2439e4ee2652a422b71976dc0074eee91b3ca2c3f3108d455bf87ed09a8301cef4dc17d7fe9e9da5a906bfc61e2182d286c7896f1bcddfe6fd23401192cf45897017a4604f87c226db9fc21802a3a201c7e510146c9f3c98915b8eba7004e8a3fb2dad22cbd0bf274eaacb1df5efc6b6feeb436c6a824aeaec5b191981ddf554a54be62724aaee63fd3ad3447895cb5b4ea31d8a705bbdac6ec0266dbfcdaf7fe2a0b32e4803aeacd4aaf4ce5d2c90a582826caaa26eb483b5eef4c133896bf81d22105ec288927a98e8f5012ce67d85f6dd468ff76798076eb266eab56f519fb176431d55e6b777451e67cb659487e03bf64803f508b40bd1975d6ddcd7fc58a2db810701ce1c53f1f5146f24b860eeb2cfd9fa51c02ca073747e369477799ce92676c652b9d699050beb62d819276b4e6f005a9ed9be5c742fb4b617415a74c7cc94611b56fce85f4869242fe47977963e7743f4a3a5ea57947515caee2c0e110174151b317e5f8863f98952e579061e7cb3d9fd5a950b06012c41584ee5843edc26b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'habff5bb00565558e293748f35376669d670d5a885e2125c7fc038680395724285ad0b24a3460bb7edc193a7e87ee2914dc94e70b55c5959bbfe085705d2d031ad34be8cf83b3a45744461ee516b2b0102ae595f552e0a2a499fa0106a5c7c74642ebe02928890d2a4705af4f707aa2612e4633e7ab3244eae1c596806ca7e5b35f3d678849c582d2f682e0566ec46de425e0548ceff3f0633aed89663b9ef6181fc7b3834cfa388136c7b7a884f8251ef259d7b7d091258a9dbb42fd87553a898c0f33d17bed90b14ae433248150a785f2807341d8ae09632f7a6750342da9a4c565be1f55c86c96dcfbd5eaea46a0f116484bfcaecd53309d9a2d1eea06a604faa6de810a437baf7b501c58b48cd7cc98b5b92b5e41531cdbeb287b62a996343a07a962d07acf311c5392dcd3eef37e78e2ddf50dba263ef97a2db78804a1c84871a0d96193c7e32bef16140f5735aed34241812ed8bc913b03293c850719d455818485091ef53720ffbafc322fa0f5d60a7594430c3497a334e3c72ee3f7f5bb8d3f0f2f6f22b321c00ea3d93d864cb51bab3292cfe2ffd748ebbc26fbb379ac26d8ee316679682019189fe1c6ab4b189d37b00aa768b3818dd1f32dd5b35fc074e0a7f55dbed482a4ef3e729b48890d402fd4155cefb8ce4cc184fa8958c1d6918d654a03d4bdcd898a80eb588fec5e34d57bb6eaf9806a68a89fe52efd68c55a0a8aac6428734de8ed567bb35e7f721f2b6ee3e79cbc083dd319f7d4f8d342a600a3158bf25336f204c945edf7ab6bd9ee4d5df8d0f70c0e8cdcc8bc943d1e4ea7c777cb8dc7158f27131581f832426a0672a368a8990b3549abbaf3e8b95bdf1a5ce060aa4d73f98f7db2fa82f57f08f0c75c2e8907e0f2dc4d3724f293548473f8cadfa33999e39ed9b88343449ea7fba27728e93ae69ae37cd3a45925b8939dbe7068b81adee8ee696655269d5b4ea4ece82566ceee1753ad09e131e21fdbc32590c74034174add0093f324e7efe3a16c2ce04a81382a64682f5c2199fe83460d752ab1da084a606ffdd8bbc1c3846c7f2a07568ab6924309bd6b4caf58c9b3cca8c52d287b13d1a805392c427d8333f60ee4539c995364af459118717c34cdc09d579ccd71ef35cc82d37713adc163663291c0c751d193163e39850499f90b8b60ddcd93397f7c70544ef9fdd11dffeb09b81a96a266bcdea4a5287c52a4cb337a3b6d204cf421c860568e055fda72d52ccf1beffb302208c26a164480ce2a5e78904c955daf48db93fcad8ec1de52aad9a53f13ccbb6392a6b48a1363ee0ccc71aaa714b5c5557df6774c84887e8e1121f66f9d7289a78ef16cb8e0081d067a8a13db496e27c4e84ea892825292bec5e7ef75fb6954e0bffbef809ea6e05d38a93cdddc1d217b0e205302cb4eff84ed136c399db2fd24eaf659e800d894d75adf2b7803c207a6a02c5db75c45b5d91b82bbe50d8dfb4423e6b65e8e4acb33cc87cbc7e8ca06ed6921da63d341b2e161d0f232302b95f140f1bbd49a35c382ca7c74dca63919c5886036ff57a22d20d5807c9519d75ee38c74434188f074dcc05d9361a9d283a34ce323a4f60c63d1495ed552e3d5520e4f518dace15f293e77cb6596a86c420a55acac2943745632cc4391992e934da424813b5d3e05bb3dc9b2b28a8d2d19570ad2ecfe207496bb77fe8f3c1d91f8ca423f10af112e4caf52b9586e5d2c18c7348103cd9990df95e80530f01faad3d4ce169e79435642421f7b6aebae86a55dbdacaebed2ac63680a5fa7ad30af54a63d81fcd99b6eec061e948d5573ff074c3e01a07666;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hea0251255edc56ebdfe582934c742b0c34d5aa5b7a9d675078c8147cda7bde2cff6e60f64ff5dda34b2316bdc94553f6520eff41a7d6392655ef1627a6a46252000ecccbaf9029b96ddd6a473084e74a0179be0a937ffb18136e798253640b2f17ff0a82a1eccc3a54f5443d72f3c5aba8a689cae25befb6c876537012ab6c0de5b465f4af609419551b448206039ec0d62b89d7cead23b45a6cbdafa934a6db21e236e86860d26dfd2d7e319ae93cffa10a6b8f5a2e21fc98ba2d646406e907bc2602f0a1bb74f15d4f619f55ea9a8312bdf7ff414ed09be800ec55aad2f8cc4456bd2ed8664989340cf5661164ab3a8d11a7d35ece7736c4f28a04761e00583c9e750641a94fb81c4dd7115a43ed867e2812231f801fc896278cc20d123bc3b029ecca7596f35a471739d32129a6759610679d9a8a38e53bf786566578e1a153d44066dea809145e29b4d8ea40c42a862013609c8da17550f0617c0b3b73435fe634a73a02c92817998a129771ddca627896ec2d28a181c9b6dc36b98216de429d31ea802d93c8a49c2b77a299278cf089806c8ef0ab32f2daa60b5100781c4637d0be5f5fd426cf4f067d829a94dca776562c53fe818f8df224a193e9410bda223baf56f8051bb52a9eb34d87e88bd21b59c8daf674459334b3a832dd3343b94d7bbb76c0b30c84b9e6caf43e0be3db7660bb16416e919880a25bb230973d31297fd54b6a1b8d5564ececaac2e17acda834df4798efb0ba63756eeee13dee500eaed705c7bfac5d23b1c87aa4bce0398edc0db0a061e6f9226ad13875a68412ca0fe860bc59effe89f4e6ea951a53f920c59d92869b3b2c29d431c9c63f73838694b193edccb17b838811d50eb17801ee8efa1c136a329a89dbb6d5c7ae1249874e2f24192ce66c264eb4be9718990b390607997c4f7db6b97ed631dd85693e7111399873a775a12bcc0bf58a9f4016f8eec60e534f31325d4a63e37da6a4112ac84731021be05dfe350566e1345d27bbb1ff7ae3e104a21d0b44b759787dadb77cb7ad9820747905069d1d96b09534acaae6b2700c7a18dfc1b33c8b0e8afbf7cc12543efa341f2382e1f94a02a56776b08a239a9e36729159916c69c75cc308dd83d997896338ae7497fb9cfdbe52acab677fa68d38364473384016ffb9add63d9d087175de852bdf02a0a4cda3e3598a24703c0e78477c3837443c3d5ed1c151d73a913489192eaf398f006d072cf7185c919b5eec08cddc57b561745360a9a14f4f37f727f53a574c6c40f23dd0e930bdc3bde0cd267cf9a6c6e17a58a1cf0e96f21b43da3a84d51c950aed7e6f860f65d5ba76939d92db59d746c2a709e97fc86063760c79c9c5ebb2b6369608f58ae7122713e71de7faa26870f44207b1bbb34ab5639ed6fbe7f13141f4aa172eee9e1f63f9160d92a227d20e0979b8608397e9218d65f34afc90423005577975821d3f9fb70e1e9ab7f07fb01de74be6399995f56f68b4b9e9ba32cd3decccbdee72bcaa9c0de254c563a71b7bbe18fd1be28781c7bdc2d88815f6f5312f92f8c5a1d79711c2f1691d306f4102eccbad990d0ff6bc340f572c5ef3507a30cda8f79dd320831bd2ab8a1c96f1ae2f9b28fcf7bfd1dce7bff167c695d37737f44f72c89705d4685f7191e5490cc1ca1ceaf68bd36419fde24d75baab7956a36eccbae75b3a5f03c50cb0dd3f4981b68d777a7193ccb7ff80b841cf1ebbbbe6833a296a23e4f0f87335e00dd118ca289b8c365e9d75732770cd4fed7358ab586eb1caa6a5b66eb7f69db9b66ca852ebc19356e98b1fd9361e55aa32fcc563bb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb07c3e674c0b31f1b38f27328a9a8bb3ccbf5bbb58cfb110a3a5bf3279cc5e1d8b4414c77391acd75f1184ea76002491a49b0cdc5f1f81109abd49b3c704002b21476c795c6d197cbccc2667b8370372935c7d3ada4ece542d62d82fd522a7d6da917f6f0998e610f7e63203a347040545cbca59bf8eba76adc26cc4f636c21aeccaec246a369163f68395a4903106642d3b4cfaaec1902c9bb9e24b8bbe9908416c97615280c3a97131e4bee8d96c953ecb0ae11c79bc0a09cf88eccde9ec78fe4a71587c4dbb7fc43427b32852736a5474fa8f315f565c3b3293dc723b84cd16a930632337f43a8e955543a5804b59e21dc2f32707d54c1783de61299841fe56e57d01648f1623a182296b99082caad85438a75099287cc2cd152b8c27ccbf0c7ee3177b57d2181f4db6dabfae19539edb5db8d30046332bbbf2ae07da70869b629cb2d00300a598990da065c58d7e62690c7bb1e31a4d1f7e28a737694de70b04d3c709368889af5e6ced98975d18dd757612fa5e42bf96e00edaf3ee306da4c2a32a7caf8f4e237b62b83cdd9c422cffadf90434f5e8c65b4872ffe5846bfdc3a3288a9fc94b213dbd1bfb726634b0aa5fa961754f867a5ea14f63610bdc1d4b310cb5bdd5042af9f673b82e14c739664004806c5dd2cfd30eba039062446fc9774659d76d2f1175b621a99717f36e8c281cccd2de02aa7b4f9c7cc189b9037081bb21305bda30e4e20b052905bb121bad47156ad8d7e3e66ad640146f38ff51cac126284f8cf573490e1c6fcfd468d5c841f93c12d66b4916424cbddb2f88de90acb7c7764ad302b18a82f3fc32fe61aa27324750edfac13ef91632f1845c27f7789bbce5a3e2529ef494ae236df4b7ba7717ba8d0d7882f1d15adace3d2b2f4055d2d4cd03a37bc749f41165764c2aaf2816a30abd83d228d964e4661c8405dcac46f808dc8588a7d21ef5cbb9050b8ab5d35b2c04a97c4234942aed7818af80a313324fac3f505239031907d0b372e852847282fed12a54989fda505aeb13cfd00358ac1046d1b963ac4cc12e6080bf2c83d42c917ce2d552dce3c668426ca8e2db16336afe95e3c622ede2fc032d6f7e66be24e3e3b7cfaeb6c5698067d1e258bb9f3b82fe5188791d770f0c610b0d28cf88b44f5387da912b7cb20516a6a1961ec05b793271dbd69850b30f26d0a8a8bec6e3f11e39622701036c1c94f1da71320f539a8c04081077133a84f1fa7a89369a0091f8a2799128d3a718cfe59aa70ba65dfec5631e814b0138844e1f93f441e2448ee71e3d0f7ba44a194b230e8b10647c1b93fd333b4455d248b48418ba0a19c8f4be4da05d9c64dd81819bffd68006c73cc3dd04c1169673a163e6e4f4b1d4d395f4a501c202aa2a4644c8824836e57c88dcac1744450019ebd8fd5d3a42a020fb18fd7e4ecf1d2ff0970bb764177a14510faab8fa8130edea378b945673f1fad545cb8d0f698c0db6f186da97dcb17b234d50a6cbf251d10d10a5bf84dc3c33a32d6c7badb5bf5728e0c4a52ceaa7f85dc806c844f6b6c2853efd727d815a0dee2e1e86236a0863820fe4c311b71107cbeb010ad1163738d658144dcce17593b38a4f141ed8ee152f4b8ab1f16267ff8550dbcd31c2c233c96cb4020dfcde1b9ef3376e23009195b47d95ebff7a83d84150afb409938b5ea4a21aa123d2b92e06ae336ca664c0304a06a6d747ce5b52807867bac7c60664b732e271086fb58cffb94349b7964884b8d47c19c6fdf6903a6c7b60148b2ef1ee404e936a79457d45cc05bc9c243509276581c1c4f2b423bde0ee3f57ae3fc823;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc87a230d197bd22e40bd095c01d55e2fb606b60782e34cc4847dfd4ac4a39e947e7fba4ceb53edc717541eaa6644406137abdd1abf51daf25baea0b6b3dbce395dbbb5050fc3a3a1b62016482f206a17a3f6980cdd5d598d8515c127c813e61be5848443b11d9fa43afbe7ebe3d155c5df43c68372881fd06cccc5398beb2bddf2e1825525aa16c928d7acd9fc91a4e8a5ffac2e1c392bc757afe6dbdcfc07d31c5337fb680c7c33b93dd7332b975c843944356385d30a9048d76350d1256508974406a20d836c56a8cd6626f73461d78d1dfdbb4256d51a6beff0be43cfde3112a2303a012a472ffbde171508a2cf1885b24f9327da18120bd5f79de4d4ac6843c974679f7840f169a156175a51a847c5df03fd10e7c51934e048e8a54f3d56fc2b6accbc505d972e38ca69fa71a479490351e18515bdd7451f3cb1f9e4e8377606aa70954d596e7674b431b9e37e4076dbd20ce3a49adc1c2519c749b8f1a80a3fc53c4946cf98b17c8ae5307efeadea7e6a88bcfc05623497ced963cbbbfac814c050d97a700303747210eed330a36ee4b2db43a48066d69d62627e9ed4d95daf72783625d8e6c16a2e5161535f25a32c05681239c76aaff4469f11e8cd70b0051a53c81ae48303946d15716915f79cb770741b8ce9dc4949bb97a9d5869d5fd094072d59a17fb3453c916685eabbebd0fbc219b7f37fea9910c97ef692e51c9e0e458097a1f9acaf64454b821def300bac340161d541ca14d4e4644571f35f97c09346ed068e7651fd85510efd4fb181daecd09d79c4a3aa63c31a639c42fa00c6199a59cf54f263550cd8b8a9ce61eb84c191cf946decbb0574f4c1d4d7579b7d547069c8c9957dbee5acada65042e9fcb7c50352bc3ddb4c7fe3a7a8326c231ca143deeac7cfb429ca5dccef70f2bb8ffd3b142565ab32a6ac15c20bc193e4a796fe91532d8f351eb50e7a68b430c6ef86f87090b6e40e338e02f22c4cb1a48597f0abd9a241085779cabb79c006f63df1bcce1356ddbc2bd15ddbc21c2298990bf775679d7170a335c72aa9ba23077de3cf5f80c98be4875cd43526efcb5e8567f63448966a3d75cf20ebd4feb9ad10af8638a5bd60edf2272d151b24495b0e392027d9ae349f80239d65af4fb8fd517da4e9defcd312d6a9120896f3e2cd4315f81c8ed83065db2d940555c70cfb28adc463fe3820bf471a138945cc87865c4c228d4d9b2cdcfc05fdb88ea4c8dae2d15d473f770594458ef7bfd10bb2df72ce05b369fde715638a2dc5c2f37bfab3645aa4d701fab3c5a256cf6520c0c51470717047b7b1cca38dc0917218bf859fe90f1c9f2934f2dbc5676cf651b78a1598b0be985e834c3136c35c6fb9476a641028b30c100608419e4c6cf42dc907d40e76de38872fd84128d3ed0626b014d27957cca4cd849048af3fbb1992f94e1463f1592b2d1aa6a42f3d2dfad25d833fc3b0afbd5eabeb05c28a50daf99b2f4581ad00952b468390699ad05197b4652afcf48047812d6574411080f0b055ea56893b3793de77d115722b3295331da6bb2723aa00127bffb02ffb52f29f2334d74f2d2f786194aad9bc669bf39259dcbc9e3f7f632f483407b6867056f240895d26f83aad8e4897028c8ef228a5a1d0a08e467ee329ea0e0eff7a6f8c95ec654301ac2748ab188c7e67ab054ce21de4ae7ffc1be548bea56b0fedf3359a71057ef79032a30c26531288491eca08c0adbe30c0d06f704f5ddea6d8ddfc3336411c52f11c30ba323c92fbbb617f77d9c12c36bcf0dac7bccec2e028fe58acc9377965b856f49703f89db50a6d4b03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h13293ce290330341d9ad7b9882d8cc4f788047965f4c909e64df16361f596e84187273311e6f844938f96a9343aeb688b558efc3da26ef82cd1fab680bbf4266233b3dd0ceb4a5ab4307624aad598739e3e1413da93d878ec0ba8e88892f4de7a3ed962beaeefecf321a999566506487a78eee161c39571d5cf55101caba677cfc02c080e042819bb323c2d718ccea4c94117139c53611cac936271ae5610d06ef900a1ec7dae0de6523858c80b896c6f445720e14108c9aea99aed512d7f48be8c8726dcd22b4d01bf008aaf326f835969d77f2eab5718746b7e7d5fbd15c9ef8f45e6dc3f75d00b89595d62edb8a85ebc51442b14952e89fe89b1b8e1ad10f74459e3f9deb24ef9812e1fc92de72ab690101219f8bf318b64d4ed1a0f64ed82efebc1577fe59476c4b7067dfd368c7a5fadbefc96e8c35476acd46bea73bc60614b1a2611ea475a7e1ccdedc423c4ad41f643831756dec51cbd206b345e5cc7bac819c5b09fafe7a43b69c98ecc6355fdabcc0c6420f2aace4bf17aadff1df59372abc1d9e50d462a693e16f636ae52485e774f64bdb0c8ff25a6f0555d1ae6b81e30c7a5b8843a7993dc4f208ae24e3fcb092d57b98ed17383ef93adabce9d9ca36754beabb8905022e753930871eaa28652824c4d2bad43a55211ba6b95437a0db9e74298424661b5226719aee08f58af00c77b7dc6f38104bade326d9586fc7a6c9a1fa31e2dbdae41b07e5c4768813081ecf2227ae3a734af0ec946eed65fec02bbcdae17fe57d147b0bf33f2af08101a9eef082fb34e81a6ea878c6ddb9db31b7800fbe65a23bc7e41fd726d065f8bc46933c69a265213cff0d7592cda079f94046b5f82711552e8a7aeb60acf5b48d8d98a690805902e687e7c279fdf1f3e69255ee80f15ccc217848fdeadae8e454c59aabe399d03bf3231127e41a6fc799646b4279d436d0693b8c64d95e022d20717e189746a0267126e3f7f63917a39b20599c704de2aff55e906541150593986ee4fdf77ef74de0cab31b19def4adaa1deaf827897780b6d6993e7b4958ce749b581c56be35bf38886f9cb2625c5136220a26599e6cf26af24cfc37bddb42102c809c9121e5a57709c479ece34a5128f191fd36bd72d3d457d675d6ff0dfeb58dc2c8007542e5fb115e4997b14b1556d60706196bc0415494812649467ff4c0a75546dd57ff21e58646edec02d2a8825d5d5ec60a6b82e0f267c606eda82f715c41a535824252c0080889d8e342d2a034465ac2e642f8978475ebdd39246e60ce2b3c523f5ab1d3bb5a2c11a758d1fac32baf4c7833e86628bfd492566303c6f599d9a1164cddcbf602478db5707321157c4f7f5dd689bb5c4895a0481ceaa562f4a4d301fee260a3cd5868ba9429700bad24ad32b951d97024f45cc1e461e8e9e8ba74f9d8f58b5b17674f95c3cf6401f40f4af5e042fc88a9956eb489d404d3fd033da17ab439109d3252e18fdf83671f206a573e4700fb9fd2c8a5cd0cc5ac48463be96014c1b07cbf3b8ab271f4a857556ad9644a9c9a513c31b3b17ebfbcda2b815ac88bd7b2842c1ce5c62fd495ef34bb96c141022690be4bf565bb3a4955c641c000d47a4465050b85f93c40be90f811eb84bdc835f5add3c2102eec8cd19922e4be93a3ec89fee793a4553d16aece3e29034f905f9bed09db36d68982efc5ff85808bbdbd756af1b4079e4c1f3194b1c6d44ce77c21eee0d023b66b1e93063d06a236e9737dcc78be49c92479a498274728e3f656d52b9072cdcda7860aa1eb68d0279912b188959dc9c4b9c7b85a874cb81c0bff49aa717f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h202d9a6f9fe48b970b08fa5d148ec4c17f13bac548a746980442931b0046ba2cad0fb4e7c6132d9afa4c1daf8e82cae90622a1f0c3233fe3f31ca11b1a10cf22c06aeb14c050af7e8f26e2cf74b9c1da50f24fe607556d87bfed79cc33ee12fa786e0a11c062fe05ac39e480bf62a2790d8c71bf64c7c412174b973cd62faae6a572b588ae8866ff5b1dbbca3ddd9ef5de04a5ff8684344dddc6f0e6706a5db28390f04e40517c8d6cdf5065dd6a5d2bbd1009899dd89da7850bafa70c97e7ce523633ad89218cdd2a02b0acb0e02f0d3a99f6a1181c4feb81c7bbb4a9b8a70f9fd17ee201643397fd92fff2513f0e5d8c00b8392830b52e44b4dfd2c88e35c213c0edafac6b88b9fa72abcc0f35229ea40aa8e77f76c51309016208526ef4e664a69a20ce5c90cfbb74b09c62c1044df0e6b942e378bd0989e46bbf4b4007119fbbc64b61c59ccb450e212f06a318213e2105016b2d268c1feb438fb6e7d3c60dc2911482d551d39d7287ba641994970179d256d03f2bb71565130fbf8c3b6828221cade5c0e4bad417a66fb85007736762b8e3bd9dfaad08bb8faad9755880b20bc94acb29b0e3d066eeda92e0a0d2c5cf13c9ad1065b8d4a286e8ed12bc5b4b6f23e71edef9d91b39e6fa28773302183e4a203fb3dc5e221a249a5fc7b7fbb54466d001762646533feed2e15e6500d722b6b5cb44b2ad99afd49c9d217b6a6f6614624ccdbc43c22d227d4dc6a9faaac78290d63c237cc83cb9ca5255bf4a56b44d4190c97e5d851634ba1a9c582685b7d7abe55cc5472cda89bfd850b52f18308820957850c2c1a7430bf41172eceff11db7cb1bbb5319abe93245bfa21737984597cecefd2e3c297df69be5c27c78d4c5613fc0a5bdaadf6243e3a99bcb7e7c2db206a76d19ae9af1308dd596db0e7122be23da8aa2c4aaca8436ddd6428ce66b03c1a91b5bd58eae6d387fe7e26cba2173e3da634672bcd9cefd5d43a4efffefa570ab56a18b2f3fdf453d35a4bf1ee1014d3d6c012d3fe00d24bd6a91e870e5df4e281b5356b356765ab83106531acdd2ff6dfb0683c9024c63745e474b5cfb298e73738d527823772a1d6543af4bc3d7f5685b924b6a819a296a0596c307e3ce9e6e262f51d112a997d69a5f0edb5019df573f67c0ed9128818382f52153c158417381dc26406eeb69afb28ef4aaaf3f0f2d78243a8cc470cc971abfb3e705900fca72949a55d4dbb81280f29fd2e7508c01e38782ebe7ff7b5a713683efdec21e671606cacaeab3e11b4364ee1848780596962110ceefa2370ef6841c46c91eec23f3ff1a517ff10d40cc030f366346ca637c9d877d40fc056b6914716ba49e0aa824b3c146c68714e83983856920ac5e5ad4e3d0e36c2c531ffd505141ac74c1cf9b56db2528e528c3a58f66a55637162ae77b6d83fa88f3126d6968cf3769daff1ffc7fffacd1a4941ecf5806557f81db37a559b1d48e4b490fe548e6a2e3ea5d78b1dda477f08ed6954591acf3d5587c68a38cd075f9ec45f9b435f2da4df5eed6b1e07f4d851769745ed8db70122179a8f4d0dff45a11577d635a590bd927be9dbba2fd29b748d1161bf67061d7f72bc546e84ce63753a81d8bfac26be480ef5222e7cd88fa3569b768fa0028bb163db1a9fa624b350b18bc3b6840b4293fdd29867082ad44bb6b9468cfbe5145567186749c3f568bb56f87724d86c0b519b7b06f04c1c68f34de1adc6c068e9004b433e96d91e96d38aa8b18ccafb654909b9f828e56221cb496ceb31d9001ffd325abc1675ff605e784b1bebca0ab6f3d0bd2bd5193b92a39766521;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h9e81f859295785d2bad5a4131e3a62230c3e7e8e2a3475bfc7631b39aad34108953a57f7597fa1096512da0f97137b6e64afd21b7833f71f7119dca575869503b17d8ab54abcbd21bf1dcb621dba3166d83d31d1f3ac68691da55ff5cc94354bd782d153b00bd6b1e951dcddf1c8769a0e57ffdd4b58652a9571be432c4c32f3aa079f6cc0db7fa0152a846d9c6143fd231ffda07523c64056118ce98b40543b636c142272931693ca038186480ec26e22a789ff0630d7352435d1448f249b8e2c2b0de110d8c545620785677e3eb8967bdbaa3a6b6ced7b9c554c98520a41dd14ecc29be33613720833e8c8996f56a72a1de88c60967164579d93554feedb84fb728b063ed13439539efef0c7b0be7c6f7dea7d9d62f6cf6833572e830b7fd9783edfee16cfde58bf629260ac5b06a839253006374cc4cafc545436feead8e266060752d0de15d461fa9d951cea2723bff292b72ddf668551f5458f9947f98a77a8dc6902652e047330ae7aa0559fb2a49558ab1bda758ee74bae18660b09bda783910a7db89d4a59787b41264396aba653df57ffbbe3bf4da3a0797a59e266f71ee97bcbeb16c04412e81e32ffb43b38baaac2c994b57696cdd4e6637e07e22c05bf0c06dfe36200708f9511f1a96dc20adfd3953b2cbc286af50ed35f409ee8ad8a88cf6abb0546bbb01004c0985c830a885559045b0d91b8836c64aa066335a34949ec20dc6c4313ade4fb4bf679962a83e4285119074fc6341550d6a9e6dcbd6aa116a934590908be077e6552c380439672367c1d347071ffb1e9a6cfe9e43b9aeec1dc1802daf5d64a088cda0d4ceaf948e247f67415ad9ddb24b5aabf2143c69d5688f257c5de5ce9cd21921a754761405dd4a818853ccc381860fdfe2becd7b724b160b2313d6abdf423a701142212754180eea13e9bb061438bc1e1f395a487c88059bea3c0cd58fb13423c8f0fbe7879b178ed449c6d8ed03f7a0d7d79096e01b5cab7bc1d626a241be5da8b1686eccd66aa7f488ba220fe70b6e24f3004ad9cb7b0f1bfa2bcca187876c6d35dbe74de2f91ffb7141aff4ff5d37250435956dca77c3d4dca1477eb39f647f3b00a4d84d6ee9c5dac2ffa90688864e8adc3cff8ad15a125e4ef9a1a6a7bd760f0f96a77bff7761b7302a9f3ac2b5b926995734f0dcb59b96ec1eb41ed680e218d5e45c447c55c5ae5e0dc8f7ce93908200208b2f14f8546169acf698c342ae2e38aeee4ce2d033e2cbe37e75097d63088e7d6cb7e0484714da056c661efd383a38bff6f755de7d812e25dd117454f17a652c636b2eeeea9e89a4718900fcbd76f04f1669dd464bcef8cbab7d8eacb468af6a80324aa1c06583d266861293f85ad4fe722b1eb84a99d46a2a1c3798ecf1116a9f513c372c051500ce1378e90892fb046336a320b8cc928875940ddb7376f5557c203c1a3f76b45617f9098ef7ab963b1fbd85ff879d9294541f450738ef996e908a125fdff6ef87339950ed953effb1b8964315b765612f78294eb706d4b746e9875c4ea89e7779c3020590aaf5e9c778b3b61fe9749bceaff8e215c2a0a06223caceba62e586073f623a3a873c64c193d156ea188ec4d07b0f6d23367e0a276e2032084e87ca077c00094594d0882edcef4834cfd9b01c291bf2010746033ed01e0fb6760f15021c469d1b4d568cd01826bbdf4eeefd2a396bfe965a5fbf2cc37d5ece1143eab741a9920292131ce9321d5f1629d1bf63eabb67c18bd4416d3306cf1b0e0cb7c704df5946a4e937b093da5c4db9689cf5b705a7c5bc0c889ff562e79063b91eb2bdf1d8c99;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hcd3ddd2214ec0c16b05c3a7ff552ee11389398e55a919a35507049960cb9ea696b52e55c590c904153c4e0791c92e53f473a0cdab465c9f0086efa73dee252009500536090d1d6f2ee2db614ffa8363a08e2b9faa85852438f0e1f158de0954398d764f266e93104076326ec9bb0aa9729bb6b8299127d57b1892b34e9268cef3209508a61b53ba887940e40a7675e56d3baa46c1d0a6259da963b13f5464ca88c729ffcd38608a26036274d0993a1c44d329f83777e5c8fce8207d268bee479f5ca8013c06d923601e745f3e1d8d98c455add38315d572a2d95d136ad7c848f71081aabdae46444635d9ba7aa49b82e65b290c9a137a2d1a84c4e651b48293979ec9f3de083b1bd0a4aa2c34958d613ecc495820c930d8b20029720f8a8f8b3c912573e37d73041502a5dbf91f6477984d4b3b461aa65953f0faddff432a03d85c88e30cf7c1fe7e5ea6a323c0b1bf8ed696cdc6f68a07bedafca5fa8d8771a1e770c1f5d77aeadffbdf2d27429aae32467a3e5c5599898071638383510687587183026682fa952311b9ec145236a4297487f91e32df74ff379d2616abb5be1e00dd080a8d5c1a3242df45bbe332148d5ac18fdb7157259ebcbe80f0d9eba3980dc4f3770fe0b27177eb483ea63106d21b1d8b351d24b8fa5a0797748bf7ae0400cab4361f455f19c2cc93d34b3f58d9f640a7c3723d6155bb3529e011d4be6dd68e3699b82b8c2958232a3c0c928094f11aefe6e8002e48b98587d9d30419908b6813ead1ea1050c8ffcdc11360ead8297f5145baf3b9cb5dc80279fecfe95a3bfa0b62c39750ee5b73a4a7a48ba613860a43388065d565b2c2c2553df0ae05f4df4295f08a62671b9a816756b7df8d87b57625f9306aac7348e43d1d0742c25ef98706f64124df11709b01ca029d36b2eb1623fd6d75a989e2dcca2e7e684d0a30302e871f14a6162f4e4a66b692ecef3d1ca3950c2dbe907dbfa15e46f85d2c10b507c168eb8e47da270501c2d9c1302e3253d4c7e7d958ebe63fd8a6a3aa4b1c9f1ac18b8ee54d3b82e2342161bbccd07dd34dff25b8a2ee0521835782d9094328c2e9d0fcfc4f2396cfe1d953e52ba806993f062898df37c01cf71c7e3b77f0a5fc4b8026719c670748c7f2cc1002289deaf708d9b8a440cc8d8d0e7c43f9fc5dc3d8460342aa9b7b189b5ff9905dd4b9befdb96c36cf95af2f59ec8567556c02699ceeee5cb7385b267144d2c41063db7b4432281342f637e3b9d43a07824ba6f8320f3687532fac285dd9b1def99eb1c66119248ce8c77d1265a2fdbda0c6cf709dc0bed86f1a83822bb9cdb8b21364d4c0111271e88a9bbf00b95aaaa03f853c22161e83d865ccc152a1482815674d8b948cb92c53cb1c63f27887e93fc5dcc0f6132a817d351802446e8f1d09741fd53792c8504875d68b52a03112c56fcc0a899e048c488e00d51eeee6bb46c671b629792174773c0810aebccfee4bed5e3a975230fb3fb113b0b315179111f03ea4e75218e09558df2d178afa4c11c5014b9d9c97e06b673dff03623c55ade32413615b20637b033da195b5d3f010add78d5a6e1aad30842359d1672b45e90b5ae23f13d7acff00f638ef9f9f5638a25b893fae8c93e2774dd7c0038f9c3224a1783d7c870774f4c0a56d2090bd622ca0e77ae5efab301e87fc0f81c6c1646335e10b9a72e536d2c4f65dc8cb54697ed059762eb1ef41d7df520edfa8fa51c99dd5c047ab916bcf85e4baa2d0badf3005ff96193accce64fc95d9adebcc8e5243fe252ae19a1314b83200deea7be534dbb594f1e8e1f9c7b64ddf7af33;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h9102d00f2794e9ca48a16b05fe4c8986db04b3e498f8428123dd07081626b7a172408a9f213ceb277fd572001fdddca989e75a6c3db6fba260032b04e1ed472ba26b81ab93c0ea6607923ab1438302e022e48e2b25c8efd61aab60fd508f31765960448eb7ca6bc065b872709477283801d52773ebebc63a7c46affa678edb243b323616baa5b74dc63067bee0b32ee7b1f3aaed0ee3af1726e40498521451a0f33354d6fcbcbe41585038499a7cdf4feaa0562691f88743fad33d271331cd75c0394084706929e9adb4690450014352e8b952df5cb2a14986987459b3d31e3e0c128e1df3f5a9f98a823d4f7960430cd8d90517b2ffb6327e1be8841251b0c9ad28f884b5b456619f6d704a5a42e07c4c84a7368b7e79e98ea90c9b980371485c86b9ea73068f52ca4b7654e59f4105314f85bdf09548970e66b070d75cc35cf78d6f36cdff09e403fd3b9ffa8f6dc6f87b0e092a57938086ed2b6ad72792b1ba3b4bf6056bd4ef1e878acac4c0818e10c5d6319bee89348a25fa548c477d9038c42fe9de6626497e7e3abfc56300c584e98267bee21b683ed6b76241503222106f8c14a64648ce0f040eac0c7e4bfd20d461c5bb3003ab90d30d6ca7f1363992f0c3e4cd74829ca075e5104955c0926430069d22f2a0fecf1ecf5feeec4fe019e88a59179508bb9498177765fad535b996414325dc030a36f31a44a6744c6655f2c8429dd4f952a0b46314a02899d8c73255bd8307ba0af8c186b92e51d0b0e3bfc7599905da5276cd16c4712a0e06085b0c35ada18f4c046bea54e3dd7a4f7fe1d3f3d33cf0131ced303eab735860ea9d2e8283cfa91fff11e61c5780ca5f829b581a0bc0be212fc772fc282207ec2374a11f9cf5f6580cc56601afcbebd9cc30ba335f1a52df3149873defbe7d35f17a583608efa91cbca873b4a6cd31e407c34b0c811e8b012cd6a1c64bcd53fe584ca39557464e27ed7e19008429354c54b74903aaf257d55651dad60346dacf68b367de1d949599e995e9caa3d2dc5448e910b19821705f599bccdee1b2be3a43820c925144f90898cc618b9a422ce95a5b9502e109061968aa56c22310ba65bb3cec076bcb7b2c6c6fc324abf3b22c03915d5b3958ac44205f925cfcfa86f92fb127519d3ef67d472eff33c6b9c12ff99be988e1335993838356dfc1e981db1b2fdc30d1521fb03ea1d31bf836ac678d1abd633d79308c8930adc2e00682ae3a77d568e4cfa350567d0b7752d3dc792e4a6074cf7ab53e873bbe4209df19a7d6a6d72fbbf4883ed8301199061ae8a0074e5f0d8814fbaafecb0e30bdb5f0d2e84f0d218990e6159cf1a6be1c3888ea115e626173bf07f346d510566c21650815cbdb898e364712cbb4bfa293054274c650d82bce43cd107187a81ae043810e82d2bb21ab6160714bb6793df1b59d684e45d6cb1aeacdc7f7bc54e1aee1b5329ebe337bd5696eff239a2b31d036e9fe3b1d6644a98fa0976c6a22ee34c4f56288605bc712e6a31c469a038374a547e0076759f6f98e26f4b9cdc4ec4210bf86ff9c835ac5bf69b1f314150ec3f57cdc0b9d92cf58c18bf2334ad03cdc93fcc3f3a5d4eb4409bf545ce2c9dab7c409d2220c6e14dc8dbe5a8aa0c0cf9b9c8de4b687e35b3122ad2560daf4e6f41221c8409ed3120e90a8aa22b5cace188acff57a3e51788fa20acdaa62c94f534f8144b94ded92675248b8ab283727fd337e493aeec0a6aba29bae05f959cb8e909ee52bcd5784daffb910a2de8b437afa3f26c766defc080003dd18a598fa618e16e56ec6e4b59ee3dcad44b1dffcf837e797;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h59763702c26a236c8a3d266d7a2f200ee1ba62accbf5b2d55fdb5e1ed5747aec80049730ea8f67b5ec47041791b6b0975f385bcfd2d49f882dbe9e03cea9b227cb1c1dd1aa9bfdedf233d2d52e0a783d3938e23960aa24b982c84bf53957ec09dded1371ed151e9c0ec6fc1f014da2529d104f0a3b6f197087d1c7848a4d52ea544da238ce8b96c5827d93ad23b1843a70b87f8ad58c4e23ce8dd83c3dd1679faa7e430d765323e3a76a569d876e0ae0a5e244227f1c693e765d393d63d532e898610242080af75a2529c6fa221d186f6878ffd16943bf88fbbd2ed699491b8b3c4febee5fb23281d9d5c3a7564a0ba5cc9b3bddba2f0b31838b983b9307ecff9d0bdd7b1feaf06029cec68525a59c023cfc8a967e0fe09ccddc492db921152d1ab1d4ffcc99c919b4420e8cdfd097140fab0575e8ea5ccfeb1901e84f75bb3920e99b06a824ff7e642778b29bbc9198baa2b5beb135434c03986d5d475e5f8513e944029451cefa9cdbef4f885b7235036f3399de9cb825c7d283beb9e81d9aa595ea18bcc3f2e4684a895132c982a0c3626f664b71181a00f920d0230df0350960bbd1c50457672be7be2e94bac167476566307a2f6938708907837f6b2156bcb509b9ae8fe169d41cfba0429eee39352843ae8b7abb00eff83ed88cf3f8af60c30e495a3ca72d057bd819b0e9cfb10d8410dad833f3aa6301178ad79a018eefd30dddc06d08430f313f383e6eb7b7928a3792be0c46a9b7591d255c4ac8f6d841f1ff00fb646c2c8cbf5f56c8e35ce8348e959df906495a3ef23b08755c8faccc5b9d2e331ab3190a06268adacfac16f2d55abaf7d63d85e568d1bd2bc6bdcb090ada02de8cc49231914c5925c594fc36b23a49411425527c522a4186cdb8dccf48da677c4146a18ddd87ec8cb02ffd97e81c0345814b9aadafcc69a9e7c4c5a1f52276cb4852780b85fe2b6f6924fbda10794e0256f8b0b83e300840de3efea2c62aadb1f910322221df101db3e1e4f7f6e6437785841a2eae4d9f60863a42e5c34f4fe68ac623588ccbe3644529b19d158f4be665fd346c01ef2d646c4b401dad4d837df622968f1b6c9bffe43ae539ac4593c29b7a05712f5ba7f924dc322dd3dbdd07a92a31255971108357c6078a09113fa42635cd23d7fc942822dfdebbbaa8b70beaced7a1ac1c183952e177fe344f5dda57bcbf732fe80370d02076c2479ee76738ae377fe3a5cff73db7cbde9a92980dfa60a3094bb1144054ceb30e2541b09d4e6bf92f34aa69db37915d67e0cd634ab342d26577ceb8c185907f00c5aa82f20dbdf5dbd638952410871a004f1d0a08aa8362868578c8f3df27b6a6a8746a8889fc821d2f1d39e60d95fe5a9c1141bc35ad9527035813bbe67986963bf5df1062012516a69a70bbeb4c70c8b1a645e5db9332f860c9d8eae6eb07ded021d7d9cb648c848878d09c944daa4614fa33423a81560d53d89b5606f0e26e199fe1b75376c754c7fddccb61ddf1d6663671bf3df415fe1d543bcbab4b43d2304bf0bf686d3ae9dc8ff1d5c40c597ac8edfca587448d185644afeca2a2ece09533fa13544016aa24ccc5089cf66f33e88ace0861cae5c35c0a0d68cb03f9599037505e83805095619310dd7d0a46568d545f4e6ad09c99017493ed8fb3920941748d123587fde486f2f60d4e31291cf6c1ac75b7632810595db7acd3229cf1838ca8b11d7fe523ee1b6fdf8d7ca688253c28189d1c7a10b2c7377277bd852006b817a18c0db89bb8af50e5b48f79bd0f73b515aa09f15ba81ffb365948cf0dd829e95fdb7f03c468888ba8ba49;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8cfd31349d9b9b4211e9cb39c461fcb458f7b9e5ac61859f7a37744d79961baad9825f2c7258530975608befef37c5811f5d64f54b1f9ff1e6dfea44d27b5d7ea2c094d9bf70ec4320ca0ee1b30eef5d7c4ead4d87cd3a61a1742ee2187ba6fd24fcc14311155b2d9adc682389071d79a27027fd6c0a1e89b7a0d8f1ec8252086c3d66e644c2ceb5fcaa1d73d4d4ffddd4979f5b330be52e2710ec040445b7aad32ce15e464c4f2a8b1aa7e97c53364338092f455f085ab9e3a05aa16c333b5db8239f3993115038e3f08e0d1ce44d06c437560eedb89bfa9e22fd19aead9b9ce2c7d9c37e69c3cce560944513472f5884d209e1d8aff9d4a3f590615cad5f50e7ac514943206de41276ec709c724a73f1baf3fc19b41096bd150add00e1a0c25221e6a30480989a8623ff3462949f92413dacb45256a5f3760374108a2189e66092a807443594eebbd95142a844481736a93263e1b2acc49ffb0e10600c892ce7e0c202f1fad1f9ba4c520d29205a4255d6bb24e4ab9c27f39cb86ec21cace1bc80f4e444d921412ee7d142477c90c58672287705ebac1cfb3815f44016f813566a1fe24c5088580d651aa4da7cd7a34156b6de264258da67615062f03c2af976b5f44245f901db4423b1a2441228f3fa84a22bcebbfe649405bca991672483ecf4565d8fcdedc8897ca955d34b75e74c4990543d6d22832c936badc826814c181cce1f51e12daa5e3f79562bd89f1f379bfbbbcf28c0ea10faae224b57f424344e89ff8736898a56ada29ba280e4321847a4bf0ce87a8ee086789142b5f89536ce6db88fd453a4ed5b11e12f1b45063f3bc618d4daddffeaf85cdd75c413f3c8d3cf3a2d84c144a59e76eed7b4339f2dcb6d3a371e5a2c5044e5cab3add2602355b8e0a1653c63eb18646d06f2647dbd2239779a0b9edb49e08ff7d56fb0dc95258401d9efa939fd7b60510994ebd6ab4e8b68acb7710f81b7b2aca42239e6b9fa7defd8fb063657e1719221ce4c5a64c132a3994399a85508f1a6be42b1b9a0c3d47956bf702c41ec9856163ec73efc4564ed921b1d9b06cbf054192676b641c9cb22e1d3005b5233bb53dd12a7a7b0b16e05e464feb2c485af594a0623042f22ae14456fcd42033522e7c01324fc64833e4ad6e066d0c7312eaa6d90aeae5ec1ad26eff0a56735dc79b3370c93c57ede9ab2eedd04758b1c3a889fe279d69eebf53972b988e18bebd8b697843089b3a95e408c16defac40c73a8b5326cc7e301f2e55ed5374b09231940dd4d395db16e906f492482c9cd3c2d5ccb6c15a64c3207e6fc5bab8e3305332e696839367be04fabb25b99ee5c57e65467271c0aebbb67e1eee452fb5c373616ef0d4cae1e5739d1be11e4d9c5ad6053595b5e6c97e74ce963b893247af3d3825a8f03ea391cc0f72a2b7791ecf89aa8514497aef059ec4b53bb9fbd9caeb09881abb755ba4b2b28fb114d897e85bf8eb439aec4fcd63d6307815c0ff6aec7134b26acfb1cc4810a1dfa69f9e8477ed75c39a1cbfd5e1ac6c4e9da733e15481db2c6c7d274163a5b94bda17dac397ddae399a5359da422bb9c1dc70d2999bd1bbc27d5523e1d462d5d76cae35a2815eee19ba541ede3d31e8c440028b847742baa1e9db2dcdff18276e26bce01a208c36385ce449d1cc69bf8bac617bdda984be5e0f78da59aa09c953a8627b17fe6e423f2a777a013555fa657bf2c43dcc6e830ed0b23ae04d95da1c8fe2388f362f602e561bb26871e77ce5461d172787c617f1c283b32075a0762598b666862873c0a80053e22b697618b34e43253b422095de8aca5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3347bca4bf7242255eaad4f2bc321422ac491cc24c630e8eff4c9ab0dc0cedd39899ee9f76718609cd095449121b1c1530aa77ca91d0f664c529e298599c0dfbf4b1fdbcae1e82e3ea244428d1bd620f19a0d6bf24d97820774dfddefe61b087b58bb4eb96b7c772f90694d3bd9325177809c7b09452a7f6ff0ac4f3dde73ee2a3f70049c895f21038925c2f35afbb7692f6308ad9eb7b3818190877dfae11516405a2fd1feeaf0154dfa5e70cad4903e942db316f97c71d90f1f133b7437c323f0c71b8828102423ac470f038d688a2fc544b1f7a2390a134ed8156498be639d67cc088c86a5ce9e1f09c8b2ec01fc98f53e5ba8f6cb1cf1a0845995a8a4fbcc50e5c423e24b6cdbb59bf8c344bac43efe046ddd44acd126c4e07335b7abd50635925f3b2b7c5c29568c1f349ac46014c4e855ccacfa7dab8e35aeaeb3f84f134977d137f3392963014dbfe0b4de6f2ceac5aecd6740e37c45b951ef608ad9833e460d533c1920b5ed3bb83d7d162cb570996953d2337a12ed71a83d8ff5de1abf03d29c47044cc6e2296985846f19b1d536c01f988f3e6c85d1e488a6be9991946f4a43de81fa14b78ff626e52b97fc2854edfdfbe7e0d1d43a65ad2d75b4538e1226cab46caf1c8506a3a2938ba019001e9f424e42c345d4b68b7f6fc880a21284691dd9fabbd157fdefa1239efecb526bfe7aa0e172a44a57d3739c228a79defc9e33eca46ab752e10127507f0e2586ba0c2876abae40b30d8c799ca977289cb66c864f2e4248907a488b9b2068433fbd3dde90449d23e8f4a956d29930a2cdd9ba208114a317ec298f4de80d7f2208bb49e5791df8f3d295d4734ca671ec06fb665170010021660968795352cd445714b5d140bd37bd12d462d3fcc8a0a83d8d0d6adc314e73b1930baff1e5f6587e5de116a8e2dec2cb53155cead1a23aa86c23f588343156ab5040b4443238bcbc68b3cb971d77c041d883a7b98fe451a1ac85486508338a85f426400b13e98f6fb6c75dc8a0947bbf4181a474cc8bc4352f129ca33d1bad2d79b1b1dddce4634b67555f3156978d8d83d4dae929f2334bc445d5b8789ba3c22f9c15a40bf3021636180d2d19b3e7dc9edbe34097d34cd1984366502e868971f50ca88109e5409de1e4dffa95e5eb4e773e82cded86fd9c9d0d79d2ce9047743abfeeb0ae75bcd164e8422f2ef406abd285af2c0f7ac1d31cc0dbc89a9abf60639c09937a3eac89dfb35e42c78b271e44cffb0157641908716959638b166ff5ef2e6f7140fbda6728a8be1a262fc005b7be92ffc10c04b028b6eaa5af6fdc8f4dfc8291481a56d0bee55b2731a44f2edf7bba44f985cbb0a6f62006a6ef4f97f96a7b423afcb053e37d93da220cea8e32b65a1066ec806cff48abf60e3c4150ce1cd2b5374dd659557dccc9c44e8abbd895907f8da17c953f29e15aea4c5689d6519b884d016f524781cb8b02f00d762332a5fa561d11f81d970c6a604b7c7c73b13d9fad3d0ebcaf278b6df84def368c5cf3b381ee9cd892d7a972421c06116d041200b4a7968c9e30648ae7192e59fc6ceb75b7b2159fd4f55a57fa3e7dd3e69add79182f61401a076d3b439c7417337d85ea1ff44ca3a50bf95ffee59cfb177047c08fff5f73b5323cda8a0e4fec8b169ddf869474ea915b4db271ecb1fb8984a329b6bfee8f0077edb72a354419e259c3874ca6507a406f1cd419a140a73baaa24c1d905cf2302d3d4a8c243a54db4027ee78d552464d434e05a499ab7cebcc30afb01e4d1bb86922bcb3e38686d51f534152c8de78b6c3d7cba9426c1e458ee7d461f39;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1afc6f7a6ca2001781d3e9cb243b74c7f5fbb3fcbd4975c732c16aeab02ddf21dc9686bc74e3161b81478ecfdb76a59bc96e1577a90f05c2b3e669d5ac3fd777f0f81d657029243ef9d231903a9b67f703df18ee2a66212c94047050e0a4497a4c775c919b20da0e5b2d3ae15d9cefc3ebf8841b3903766b413e01f6580b0c8537e7fb5c8896a8f97a63f007926c5dd36d1ff1d42696bb824ccd21f34809f38c63050b070d53272ce07f17fd8ffd06299c8ff220b193dc3736298d4426f049a1c0fdc70ce94f7a52bdc716666528f209805ca100661e9d730dd26fed7917d40aa362e37512eee850e8331b9b0975300571ccdbe87beed694d5880ede272aaddc754694fa1c0d7c2b7f389bee81565c6b5d02ebe881569a61e4927a9f7975749331c1642f0c19227f539735b6f166e010aedab43b30afee79dcd20879b87ee439c019749b9b375c88fc7adc0e7152b28719f11d99c38b9fb0dc6dd4d7ad761caa01bf0e1bf5464953d992411e310530d52da5ea667801e4c389d255a9ddd9bb4b4f7f5de6deafa43e64632713735a69732e7e02803067f3ce50b42d5509042dd4197db2bdc4ebc55479fb71ef01671c04c5c8853dd18e4914f088394a9cb906fe9a69844fbd351e5e97064de65dc7e48d266d93431d171abbfb16e213f5b63fa1b6b4203e570f6211e5f461e02415a0560bf135c0b9b559008383db2a1bfb0d204a40311712a9c16cf7f0af6b00e7ad77a8ae82e909a796e104a7a160018c9772eebae069568b9d80865c8313f8f9b50cac1a6bb49da3fc783b690a922febf6f8dfc377cce27d77b2de5dc23648c2f52112ca33edc935f008b86233e25541fe39c7a0acbb473aaf0e6711a9193a4f9c0ae213d3c713d3fd1f637f156e8fec383a23cebaf58bd0ac898a3fe8ea7f4c638b4f745bbdf703f0ae8cb4c892fbb137968a1c8aec08ca79897a607d1ac82c653ae8dc632879fdb39d72ef16ddba0d7475abde03a94d529f81e36646cf0e1e070043a2e12d8b8d3099851f8c14e613f5e23b012f8b13b0c9878c150c7101c147cb0cf2f3605bdc758eea9715431b3e0057caeb81943ec00d6e175c7757a888e5414f82a88acce520c6fbc20a1a9e7837e63a4cbf12af9d8bdbfa092c05e50dbda00a1ece71a5965b37584468541242c01ebef20c013c50d86c6d02a3ae0449e40b821cd08bd92a334a8afd42deb06b57230f705558154c370e028cd2f15c95800133fdcfcd85267fba4ad3dfbed60f0af748590ab1113cf46cd8e920932796efea25fdfd97fec2e812c71eaced06ace9d57b8ada5f2217e587ed3e1edf8d3cc9e11d992aeac9dac9546490022f4f6de8966657fd2445b402f0b2b3fdd76953bfee300aff039490040348a1d632b7c27be7f91be614d749d8ae6a2ddef8123faff612ace60fcd2e67581a32168868acb6f2ec6b27866101221407a0e1d385365fcf8c5b9089f0ac8e81c9dd2dc6a1de3908ae19533021d639cd7f43e545233f4a8afe4df7e3cb6c841f832f281eb40a1c42399cc6eae4a9ae50bec7889d1cc23b1c7e5b92d0a4c03bef7267addbabd9a6ee9cdeeebc9cfc9d185738403af5075b60b288ed57e5e3d1b82149ea4df83d92f56e75023b73c768ce33969ce1dc15d9fb3a7dd7a93235a832a3250e361dc1cd27e405f18b9aa05b2539ce7ee00e904e23a493c45619a52dd36e57934b22390aa7a90f26c44bfa7e319bb11cda20be9cfbe9c20d39ac262ed0077b911cb7d8ceffd12b9b357ed0c2d7f4d8f959a209d324ff0dff8f235112e3fbe65444a49d930573501b57144ecb676b5df20b92d90288;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hdcbd4065030bf6cdb06407745d32beeab2e568bd927d6f2fe5f82598851d16aabeda80bebf2c8451435906b0e13ece0cd7969281cc26532097b183534133838191b10ebbfab73a3804a3e517669916009a6c465a42ef61bf3fbab431647033ca432c2090313eca7c60d60b67370d15fc4096ad5c8b91556007b36d09909369a7526ee5bc15eb691a94377cd73fca4df976e1f7816af99e224fae59a2464cb82c1aadfd3eb4c7239a44534244d0284f10ee589b72b549e2a814e41ea4a5e995fbdca3d858b48f26a7953e9438143b6d0e73760adf0139515907562c3105d2587f2a7f458e605a81b0d42f00d6879f74e8e8b65f1c72f6f7eb07f3c04c42022fd945a946cd3884d8afdb3989346b6a504af7295299d0c7813de52e2e4f9521c1c0082846f41cde5495cbeac80474e1edfcb04b19879cfe356122f865e36f98f9b4b482948b6913942f4b8282cf4cff83cd48a2019567876e4dfb171c483260d19fbab8a3c7d4ae818df6b54567875d562577542b9c459aa92faea37f565154900dbd0581fd513bf35f83fb17b89fe51d119fe5437922e167cb5a8f1f84cbf44fe38306295e47b85af50b52c9d418509a9f6f3df6a91a8e13160e99cca6d77967a848ee0f2993ef42dcb204fc7c96345570e9fa6c22a95d0c1751289a3ec7c70204ce4a28161775120bd3f8e79494d49a6abbc12997d571c9eb2f1923f5b4e10d4cf12b0ac1437ecf12a1dc8566d20a53c9d028641ca9e90a6d626e4b357e78da75e2f2b3f318265dd2d1f40fc2e7addf48f19c4de839e85122ffa584dd683fc26ecce07c67810297fbea9c47c156b32777fe6da74778c8aa7b97a2f972f169c87e81a0d58cc0220478ae6430027917f41de64d37f64e3ee590432a08a5bc9fc5dd05000676cc5651d39f1e88d727c619b2f8e7367ad3b9c6effa4a086436b8b07a8871a66590bbf736987e2807123eae8e9a009aa07dbd65a8ea69e6232fdab49681319c4f9cb4d833b7c09fd8a13aff3c615be643d7dfe86df8200ae8e226c986c9e8aaf6b2504d086798395dc3af4e79c06a4f24aaed33e24622b1a2a8a68b5963a275545e03d1ab487e017cd06812612d3724278a29a654cfbcc2bf5324c19d90453ea0a747e3831abc6b4bdb4d3e446ef4f196d40855e6079914d1d5b0631722874c7d17659a9de91272da5c5c203798eea2c217e4d56ad7c232c8198060f727915c264a3985539045c6dab0e19228cec33ce297ecb556b75ae1bca8948e131d54bf77ca553787f98867adeff7021577459afe6f40c4b65ab574cb8e9f91865cc635ea1ddd0b111e800301376ed2f861e5b7f16442b4d0d4ebb29dd21762506e28b24110a4604a53fb34d8aff68535eb8187fa9cad57730af30e5842341a8c71406b897f6d6f2132e79acde697112005d620dd21586c9f48486f8f1010d922fba7e072cf8b64ea572b6ac19bf57fd0f54823d6f651d55bed0565c641ddc2561b1aa5dc67639efb60e53e598e1fdadb313abc3ab9654a7cdd002837a1dcccc0dc8c53623c2fd47e4907d3c5253fbea5b91eae626ebf33f8793c65c0f9a567889f723d17a7935152f32d23f2ee3ce04bf461e022135668c23b6a7c8ef76a288551100d9dabd787e106cc1a2a2184fa5c5fda6818eae3c14c9b06417b5e9323827a95919147a5e1861019bf863e9a52f8e6044e8d9b97d955bdfb48e30364b50c005d3e4b230660fddec3f0a9668f0a3b314cb0346eea5f72abdd9693d00749096d7bb9f9553e6fa7004d2f50f03339db065dc5efe9c515301a3c7d68bcd739a17a2eecd221d76f143757dfd9e301c666;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hcb9002bb29fd0b2c24ef0a3caf8c8a7beee1760cd83658dca3b075eee76191ae1c300c793f98037c1741e05a41ac5c8255894fff80d3f56a8a8967ae128a37930d9cbaa64293d5974ba73e62bbe873b82754c06d5c40e1d8516c09a4d7d8f7b23169194ebc09edfbe6bc02f0d2e6be3a612aaeeea6cfeb39c4c1cd3ee3253846ef142ee0717cce3d5d1dc3fc972d19182fb411b5981e113f08ff14803ea824c971412ddfeef552aa2b2788e433c387841d2925dc747907586f1a6cec9241c0638a274fc264e51fc15bae31dc7db05fd604eb99bcddc3c0da659aea58c2e84c0bbc64e9807807b8e48d31d620b8db6b2669e7cfcccaad391cdacf665d671769df2aaf62bec3b2058329206d4bb0ebef9a4dd21fae444485aa0e5c7c50c2d992507a9dc296cc96f24bd771e62b0a846240e1797b01b2feb6810822e3848d39088baa8d5b9e99f3867913f65f99e6567512200be2c250c8184bc381574d8795c4ba93f79ef83e6444d004a918484485e8d2b69b956b54b1b9769e57ec4e591201809c03dfc64bafb54654d9bd3f9b89bd04c409e97a4aaf6e7bdb50e81c29c2d78a4a5aae5085f2b015baac1d96f9b393517c6616b09cedded1a777797b544eff0a32ffc2b86ef732a9fc877121dac6a7d7886ae6167a158c0772ea6fe4ba6f01b7ccaa992ebc6ed8dc99758cb6de86377fa37451af787f35f6673f5da01470c8dda610890518a1e80661218979d97cc48750fc9275eb640302b7afa68d5cbe2f2113e32def37b5748e7163fd34aa9be5d6b8b663c2ab7faf41adb207d4c1db59e89479fd4f72b3a9b331bacc6829397c13de35ef2feec5e46866d72583ea80f19976b188b32aa6adf44bbe22d0facd508dafa1ff13e2ed3d0204ae31fe96bf1ca5637d2fb9546dc6d9f539d53aeb185a07ae78924dfdc772fd2efca1a4e14270c97c197215102b4db8a93c5ece8a2d764a26f8500ff92004d304d4759bc378defa2ccebab79cf47c62d9a91e3a463481c55fb4fa2434475012edd02d9f796354e68636d988c70c4a04176e383c06dda92476c7998d964dcb6e274332dc167833257da1e31125fb743514574daac62e4ec10593690ba4871b5e71d8d94216009ad259b91e2fccec187ce5bada8fc28949096e901ff759f832f867c064f28b4b22c8896d9543f880a308b56c33ae8a9886c39add9a09456e4941a9ce201153b7a83125061bc4a0da467b5046924a0a71a1f72b97ea8277f15a95c007c02d9940c39220378424fdb58fdebc113fbed42615aadc45aae6fd081080f2aa04098d5ddaff4bac5b50cf018eb08262b3426128db7440c9915ee5d80e510b65b11a067cf19de91ddd5fa1f6733aceba51262b662e3ae07cdc1c562ff36dcbfc8004a8e77a4f7a7fdc0f32e41b9af5e013605d09c82c254693a7baa3c5ae5c5af11b82be1cb9635170794f8b12b04868ef364b0e77108fd66c92942ed38dd1450f81c5c768f3062afca14a5d9fa3c2bee58fff15485a0b92bae9caed1947d915c6fa31f689733523693d3e5dc6da90305b0436ed415b75a79c44acba6f644a30cf82c14f5f643cca676e0364a2acf9be7183f5a6093f429257828a5690cb23195112820d730c9dfec8a908bd6fb010781d08db8eed590e80d36ac6c6d6d6d8d449214509788631d00b083f09682ca418153e8e49f4bfd86e3ae84d48f363d480e355caf7cbc9a74196f44dd722379002957d6994e17f8d253baf9eef48f426eda8648bca70141d2ad71113e006b3e15cd53376e0a9c9e90da89d1bfd50917e404403873dffbd1b2a5ab123174cb5748b8b5c612a3064;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1cf342daac1ef5ca6e4a5ebbb856ac3fd6537c986ba0dbdb2ebbf83bd0014aa22deb75fa15dbd63be104a86cec024cae998f97df0ffae07af6bf603886b015423ca31a5d581f5894007e156ad55b737e6e6eb75ec7bb7f48d03a69fef935313664895e4c2ad0db5a7f5ff02f6abfe077624bfbb7b78450aa83922120f7b07366099a48e32d723bd85c9ccfc6a40859934449aa812ee7523b62cecfe5a4d453f65af627a3dd84eca2e0d6df0d4e0663fbc6e4d03c1117c1859e646e931123e152acece2661a0a70b5f05c656c3439f977f4df6855ea3258208cc3755c692fd1400883bdb1b48eafe477efbe8dba31f5f1e2125eed8642030ec72aedb31bd0936b5aa2349ee52ec3e9ff72bc06b3be474e900d29ba2f0fab24526b0cf046bdcfa2a986a1ed72433c989b7a08c877c29f0632de4a4b1c64684ac57971df0d1e085e94a5317827de4764a957224ef380c75b01c90cdc065c42514b08d277fc1ff69a00906e56e3796f27a51dfc2fac49bc1bca4d7301aefbe794a359ab35e76be230cc995aecdc5ce08f837d3d0c116033b5675266981beb51592ed3d124aa9221fe16109924ba7128eb4ccb5a21b62ca066294639a29b8b4deed24fcf916c4ad5ce4d64464936a634ef97cc0098bd7126c3da14f746ae9855ab6b464a277d6ef38c4fb428303119bd5711ccc2e94c173f54d7c2db373edbde345611b4001c896e2e67936aa4552e545629742f66b687ffb5cc06525da9ad6b2f55f479512a845530c748966012f337a00082707081928b2f9e9145dbdc0daa3937617fe5b3686a2be3d17bc206f56149fb28ebd1660f379ce5dd24af5a92a611096550886a2953d656e0b5b18b10f8767cf0a703d85b27613cf2bf0b9a0ca310840a7c67f12157319e9b6db060f2272847e5ebfe651d8ec08c19b80c478f228e9e57cb15779e967b4a5f82662a4ae9b574ce932487656b178da8f8229b1ff1c27622adb0cb579f4dc667efe5d5a7674e8f26192ab19d5cc5560432e269c17e1f5b73c8b84b4ff45b5fc87370be4b55a903aa629e1e151f7ed7df7672e682c88d80ca475725301a058e0f3f75bfc1554f13bef182f22e8a369b9b1396c926f73f14bb6314b4ddde33d2ad2a42f88262cd57111830f86ba13912481b5827f7fd95960c786980ef8e3664e15c64156d8c2dd57f810c78fb39f27c44c4d05c39105f97f1fdaacad8be59642cd132968cae269190d4d8c3b159cffdd2625147497895ac8005dff684e23b40bb2126b93adce16b3ccd77786e9ca84c1b4f1d08935db4d0deea4518a9cc15ec6c5b928030450bbbb54d27f8c8b005e6f806b77fed3a257a217a08502bf5d090f6d74a9d59f3655218118d2c3e31c8315b24bd143239dfac6b0acce430fcc066c471e705614e553122bd0bd721a419a819333619b7efcde724d950493d6c042bc569ee1c4cadfb10fee75632639ccd34fa5820434df5fa49c6d4f2fcb5e3916d2278d59d97d1b215b414ce7ba46111b045c0d5e0ea90a80aa34f822526e1d6b9f54d1d8b0a2e8336bd84300d399a6da15808b13a86060438c2b8a8d08c6075aa7f64f7f29f8448005fd25bb0b96b3149d92e7fec739fc0163f6fb88eb80de36078b6a9a8b39fbf49f34099c56c4ec03afa3699919b950b4f5f23b8c0a2bdb4b2886bc2219e4fbeb4a77cf5c96c177102ac5d41cea61a5576c087f6c643270f4bac17c0a61731e85392e02a72af93aa72ca7fdfdbf57faed68b1e4f40fcdbe2c367f11c1ffbaf005a19804c2a3727644c20b96b067b9db27c79fcd519de35784763bb938c554400c91f93ddcc4543af;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hec20d1f2ac775964fd54cc8b3dd4e97c948499a666190992a018b9445eace44b36cbf2911b20f8f1966e1a57361954c9bc8fd00c600006546c34ed552d390ee8feda16acc11f266a9bcf5eddc3a551d0aa94ba3915609a5542eac38e2f3aaab2be4c26246ca8b99cc2794232103fb7f1585569d12016f9d3834dd73910f3f64e4a66ed3e8462eb685c6f02584b3c0483990d6eba0b4357357957ebe13f6c17915b2a9a66c747eb687b51aa13b60bc5f9441add63429fff5b9b6deb283903a0f242ee07fd27f52741fa44ac4ff5e39348a30ea01c8abe6db26f4bd9dc91b5d39dde88a7153a3fe24d6eab22ec584946041eb69bf88c3753c612d97e83b1bd35367beb76dfc564a6ac59c12b8ec0c7fc8d971e1e93680ea6f24be2adf96e0899f4d789f10db45ceec83a9f3877ba5abd9cca44f5eca224260bf5c148bc01defb6842344dacf191bf02c6eb8f07f7a98f8fc1c51099e889be4488550f034322e39ea4659665560af182b52d2add46c6526c4803d1908c1a4a8ea05322de38ab64c63d2513a566c54a4279bdc8f40432a853c8879f3ffc5d91abc25c91cff17f09d11fa900c9a12c04e4e5965c574a0357031592c9428dd43f641b8e045b0ccab8bcf195df53fd8289bca43745cd8b006ba0563377dc259fac21bf2349f376286efbe076f333ada9de5e4ee18112a9886f2e3bf444373268211285dea133fcc5aea763a07653f772794fa77bc381865668e8a5e80071199eae6b73cc71e2a9295305034b5b9bb55c451ef73f6755571d1307ffada84c9ee39ad194036bcc786215354138821bc356ebef09efdbec841d08bec7d5499e44b03c6450bb24e3e546ae32fd270ff8573d72fa0d9a292de2eb3a8d926f81ba6d8a849bc3b3014c0fe65de50511b3cd78a0b13cc133b8e677dc5f0495d6a1d521d32809079e222d3cfe67965a1a13855c175b2a300717db6f47a40edb620d5106922b0bddf7836e7bcd0a4a8ecaef85b260ffa30602aac88777b27fb90b38bfe09e513921d405d443b586a672b01ca5c96d040a2ef14e49aa1c95981da03c0a64ee6a67a3eedf2ebb0885e7f008b77692d2fc70627ced062a55e27e4a3d677bb3a0b426512e574a7f1657f1e44fb755c76271a23e04326c2398aa79c4f3db466801baeadefa2ff398229a3659ceb4a2f6a15a707fa3565d54ed597fd52f3d04576688ff6c59ad61e99da8659a10dc1ed975df2f8d7b52a543b23980c53042a558a37e57897933f590c371158d0d09cb3874540316c15ad809c015437f1fb7cdd5cb4d0cceb9e9d7ff562a600d458cfe799fe2aacea17ade785713ef836e152122a4f210c358b5ecc564e835da99a72b664d9dd9cbb01c0311954aa89162b790853fffa82e78642c548eda22bc9302ca75c58e068e2f1cb67dae1222568a7ae385fe97950b3d3b5c61119b66a1efdb05ea88f17e878e1d7200fc0085736638ef546861d98e61bbafd0c69ae729fa33d1fa4cfe950c797ebd34c5311267d59459ca8f20da2cd9d4e0880330c1e8013a74d19c0c8985100e4ec0c787461c1e0101c8ace76df1b5402c85b0294f41736ae6765e7799445bd28f1bd91febe406b951718cbee017b6c7ab6b23204270b77c47dd79f35c571202bbde117c6abf99735ebcf6fa353a954c3fdc5472dc5e6428c146df345aaca1a67dc490126c6c378834cb69d1470b26df06b80d6d782b29f66a81989a0c47fe39990333c60d17c98ff31a081f1bb32225d99df757f888b09cf62d63d75c22478d70d48311e5b8ab2767639a3f7dc94864fdfac083f004cec1151af9d6e574ba255b81a92b4f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb488fdb7a31cd388b1c94c872e83afae04fe62cdc5af14a45ce314b884dea136affe31c9928d457ac850887d2ba37f9df8e2cd73381b3d16380f9d9d4eefb377e0d5ee76615e839dbb2d121c4c6ba54122a354a29cf993398fb0716d4d785434e91df2f479f515c1079ad8eaa6d75e9b25521490546fa569b8f70fd22ae49c22bdf796e965edf1aa34dabd2b1bebd5571d9c0fc69d9d25bd438e2874e5aab71c4ffe59080dda78aec401d97e16f45636c4550e7d9514e760ca936848835d57dc7d3eeae5281ab2fe749d9c2668370eee81e113f522fcc200ce89388d9076b584af0271f0e21301c4e1645ef477c3faae5e553df0e7853f8d895719e466958d3d813c556df7e15496850d01fe8c28ce6bc2df6e242d5d4b518695c53d16afa2e8045130fcfdc0fb28e6c311acf906a3390cf85c5c547f1905eda33ef5d065a6c3877715cc906958cbcaecd27ca6068e5b92411b7dc103935c8f8744117eb9a42f36c0273afc81cbb1358c87bb6a74f0f19748d490a5bdd9fdd84a5e2ab39cf3afef0a0451f1ac6e3cbdcc4363565be0331a9f35ae31b13e48681285125f31704f6713cbe83d584dde24250a582adc383630266b80781624653997e3958b26e56b16eddfde13ae173adc1e1cb35acbec64cbb4e3aedf24b17248a604bcfccf4d4fb3a99e2fd0774f1b445fd658b0f866c0c3ae05636bccedfbf77edb1adabb44770057e82c9c1a9376cfc348135d9dae6f66ea0b0a2ca578e751c4a5ff6f282f14cbd3e2f6a000fbe85e3e731a7349339bad983affe952c31f9fc929496dc9661332605da52e0d8c77a9ac4b1f5d279798a5582987d01465f3ab792d3080fa05f6cf0a177da1130051352f063b62621d9e6c4191c5c0d163315af442da9375b8e5c286cbc6be1583ca65f1a659a90584332dee527f2386cc39104ba01dfdbc7debef18489ffa7e2ddfd2f55f6cf064a2b98a4bca01e79dfc769e50ca9e919fb821f90ac14a66e8127f3e85ac5bcbc352eb0e713ca25c7724c5c5620f79bba670ec60d1c4a6ae376de6e7cc5673aa76492f84c2361283e9260bf845c6e685b7d14f73dfe446f6839a79fd8639414b52b0e38ebd0ca7d11c0eb43896ef36282977b1b1ca4ec35c29e325660fecc8d56dd32cb49f6a3cabaa4cb2bab5bb3af8f79edb6cf15136cd6eccd7e8f3b5aafabec5fb599fb59c1a24615cbb467e47d508636287c888d07febe21639554206c0ec82d917388f4ff0c690ace16b7056a2dcf534744fc0356b6afb828849c951ed3d2689eb24c138069aa13674fb22dfe6d05c91a670b26f9e2b278e027d1d8d1b3c0c278745179890c305be3feb8de5bce7eeabe599efcc64f673885167442547cb43d78f8e6ec98e0333b15e46e014506bf1b8fe0b30654c920a24b3ef153a08a962c845ce3e32e03540c594891bf1f5e5a5c1da888abf2e357926c47a2d4f88f616a31d81f7900213642015fb94cb0e2258754986ab1464c9fcc2000e1822cc66b68debfc2e0b5c73c178115707d398d46e4217287278edd2680d3c9dc02bfb2a30ef134d4df8c0a5bc96517649a5d77fafc05ce94dd308d4782c34e8870860539a06d1f58e48917672002e2bdac7d5da662bf46ac11764c838a5dfbace0306bb527770cfe28743f92ce6f52ebf7cf6ea82356c2b45e6cf761fb8a901d2710699bab08a285cebe394eb201b2f14d968a22a5d210878b78ef4fd38a6b23f90f7a74b369ea26eb7dbad849d9d07c500099cfb6bed0280369f6138ea3d5dcfbcb223aea70675b01f424c62a7649dbb5020603aa915bdc3cb973153e3a40b6ba97114b4a7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hf49cc1c9a3a24b89074eb3f00f7d3403bb4b5c594deb55dd2b1db46fff6912a51b65be2cb8d61e0eddbdc8f33b37e20d9b483bf248f9a42e2a06f40a3d06071ea4ecd8603fdab65f1bd2d5647ad73def4737821e0aa9539bbe61ce2e9a513129b970ccd7219cd8a6d5f313ab4298add9d447029b38810889fa1040e83c8b153d8b6453f13db593113457f2d0d4f3656a0e155f13db4452d6e7572d3892701f1bf9da23f44afb60a43efcdb4844dd9f6c1923de09d66ba4e9f2130ecc65d5efb75f77b2b2092c15bdad2eec8f4d5cc5e200890fe8929cf55fb1eb3a9d44c2ad8dd72582a7dc5ee114ba209d74606fc9c243356b37fb056d3ded68e48d89191d59ff6d675d90216ff3912bdbfd16262128f852ade29ba23968895ae4499b999bb666900e41f7b9b8bcb1fc46520f5bcde050eb75735b5d9d710a6e283859162d8aaea9682d09c7e2e3655f26c23289367cd58f67ab3c66f3acb09e0f9dc5a15a668b78982946bc4c3bc7e017e36dcc342f6a67d7b50a0af55cb696d4d88e23564b93703f9534995c42dec3a431a928e6099861f34ee398be37f2b33223877633aa929467a764e951866d9ae202b250f10321cf43d8560699d0bec33b5c3a8164b9529a95c92d7d704204fa41a1b07ca1b403ea95c79f9f1f08d1d40f07b4f156ddf3c23e1e67d7595d1f374f8309e6cb9f49a14c7364de009f787f6213b89d6bc7d14a595be66ff1096794cfb1553635569d1ba8473f18e9337befa7faa8dc45f87fe0c7ee5461b9944c898dd6fa18ed936ffb3abecd480dee9023206394db066727c3c5a4bf9cd08a9a89a609ff8abed7dea709ce760929afda41df5e4429ec9533b53c0829946c2b9b75b31df8e1ee5e49d44916c639f824eb7dd4a224f4ba48d4e5c05a867774fe1ac0b500e78671e4556414e8c941bfbb6b370eba6a91182f7d47e156b25dfec40835c12857569eee1bc303e31528a4c255f0bd9e46db66dcba403dc75af00c2e29f5656a216bfef83769b15ee5c2e538c2e7d1c34206f0f3592af386a3a4b06f9c8a5641ba035d65f83b3a82da33ca7ce62d77e828ba0e05146d292a0c99a76aedea988223761a64fd30bd6afede88be3320506c55b044acd39c635020402b3c88ce31248c26e6f725631e7de3b8bccffe634bfd565cf4a22d4033a9c7129530b4de57c1d7033e7fa11d7dc15b2399859e45e38d38505e270c11bc2453fd68804897e18c3ea143fd67ec825ec410a1b2dc0820c3937441d82e1446fe94b92cc2bed5c19874351af9ff71bc256f462fea5f8a4c36fadc9af4991f5fd0de1091b600777e15bbc86327df23ab3e1a7bc3108bcf514b331485b36d5a2d8762eca330cc35bdddb228deb2211658de06b713bc728672d0b5e8000581bb6208dad7871062b3161a6ed3b8576ec20b84bf30dc65dac9e6c7f4a206c54cc76deba0b085c7cd1064221b5ab4d9f77c4063e180a7e553c3443de76f81e115c1d14a3e9409fb4de921980b53c2de9eb62cb19b121355ffd76a4f7ac12edda30de75283d2fd511cc98a3c49724cf088cc1cc59c5d4eafc51bda2363db2aab9f750eea70ce2d8a074717c7d66993041c53cd6911812d58ec94867f21dd93a5bedd0105a99b806e696afc1c13483cf0959ea25ed68645e4eb2626d3f28633f2d34a17a48ec759e248b168c841a49a971a5b17b2d81a876ea593204e9078252bf8bcc000279db1f548502414a88001384ad01e713377ea8d8801ec8f7d935445a87239f656154559020712b436bb2d6fecb9b7225e210a96d20a69cf37cc2de892a94e6a01a0f7e539b2d026bc104087;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1ef485f66018de1341a9e78fff880d8d9b4e16c6e255481af4ee681fbda0f9e4c56ab7dc519c484058ddd729515b80d32bd50c298ade50958198c0c933beba653bd433261efe63d30621d01c688914b386ed570922a2062f8f7f9246008a5dc7209840ab6cc3d84ba4d8288d12bf23e00faa69284df6a2b898f4f4d05746663668be9b95dfd45a58266cf61fb1d8fe01378e0bd693aab4b37d10f352551a1c5c6333af38a9268a1c8d81ad97fd5b04f23673821248e003f34072b65661ec7b750c8218931d94d67683a19005569838a8839cd6978f1d60275f98ba9e3d5c2b1f020638f5d3714d7a82424f0ec189bcd840d14a7b36bfaf3a17d5306b979e16e2a67fe474eb46b57fa7e0991ad0dfb5004a89b2978caf8cb96a2b0620a93437a9d1ba701f880285bd4f76e31b99dfb5602f4f39ff3939fdc15b693348ed7a3268f26fc4f58a05cb3fe7260d315cb759e5ac6e1b30fbb8e1b7f8b3819b1b585a327d25db80abad02f3cae67e66e44ddbd3a54e274c021e4bd0305fc6f913b7e0ef77613236d804dc22ca0fc643c60d1facc8647e08cdeb4ebf05cc9961f4e920312007cd6c6a1fd2434b6e431c7e3fa0c4c99f54251c60c9f6c4699d6f8c29e282b49e5f802868d5426f9c524602b74832bc71f78e4c1e392871e1ed9725eda18a88b8bf0c143355725e39cb49942dd2734f6cf50245e06fe9803e349553463d2f2905d4c932c503f1b7e2eb4d4da45eabe5c6bded2b183a93e82abdd62be736aaff0afa3a823294c1d2301338c00e800a21e72e189dbf6829beb355460691ad3584c4488c3ad6f69f38a094a582fe7ad5a86657f21cd67fc4a5645789a9688aaf4b07128bb4391db659ea7c62fa60f06705ce0c1d0a44bd72f6e9160b1758f57d0c79b62ab4483190cdf893247d1816c910689b85eaf19ca86a6ef12bae8847cf4f9eb254346724b4b169709f3aff2d0dec0d0e7a2b3a99a38c2ef193c2bbdcc8fcf58685e22a06b8a0263c5693e559f01f7b537adb20fdf79668339b82a85b5d16ea51c7a3a82d808c9ecd74d52416cebd171545366ca451d23eb265d40338422b2efad0e316a2f8c42e5f4ad0e5e381eca6e663754b5c5b2bc2d99c99dee71b02b372b2b1ebc14d0a391472f23ddf156561ea1ed876009cdc6f6a3cdedbf5c99add1a68dfdbfb86453a8684f8ace13e15f55f0a33c644aee603beb8b91f52a21a46b51b502f82b79a2a4dc990d95c4f0a933206edb7a62b2fba0ff682a050e878d803276f22fd6ede3146c4bf8729d89d9d998d409af318742d2fd091d20d3d18741b48d3d33707de9feceb81d568bad54dedb1f09eea1b75cbbb9691111156079dbe153c599eccae06d52c03d54c351303e08c88c1e1eb1d411787d76b1c8ee118020c050135b96b437db3dc2cd56a612e79784b78021591c56ce3494ab642403463586fb142673e2f111827503e04c7a0280b4a5bb342cf9d36dd8fdf14a4a907df50f53a148cdccc2804aaaa1780fc51cdf1c5f9b316701a6340cd5bb6c20eb44abcfca77d6241885c870fdb5b410c380e2aa3ab5c1481e581af646770733743c9ac7c3dcfa77a9d2244c87012d78f5ec03c27e2ccc7c6a6daf9716cd21bf24f686473a0df5cef9562444f01b58732f56badb4fb93e624dc1176f70a2829204da1f5b611ded4a206bc8834f4d779de08019b88a2d39d82a8be534c3c35218230fe784a7121e2308f5e60d948b6fc054d8ff9170e65a0f74e566d98e651227dc7ef0c16df7dc47354aaa02a15f9537831263bc09343e94e5a45143f7b6a67d249090a2220075656df03114d0d6f27;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd35ae28076152acda099e3aadf434ce02af55e4f4d0e3111da48dbc957ebdcaee9a4c2b0f246c8c10d725c7ba4c6cfbe6c10c75e9b26b588495749fd6b96223185fcfdf6e45eac0ef96a647f6fc11dd7feee4819f530d8dbc6c9e56244db30d1f2ebf4ac6587fcf47f0340b6857b4074bba9454547c17d4d76b95b0198a59d3064345617e408319505cd89cebb0e03cc1c0866305143e6690ad27d65fa4a15c3be36d6004d13f84897afc4de5c375b058a2289fc4913b5159e46d0eb34969782f1e1ab68f926f396e3d1fcf10f32afdcdd8d542f366379ef66da9444e2540652e5dae9ac839fe6b7936fdda07e7ef885e100116ac7dac27544ff18f0c6129ac934feb715d4b40bbc923a0ec4f1e86ff4b33e90c5e25b1780115625c0fdf930766d2534c600cab8786b90b59872ae9785a5844b605079830704d1fceac29b57724974338a47e5401cb8b3f9e578673096e01036ade8c0416ae090f240589d08f01690fc3ff7396cebf6d108684d3f6ff6e5aa72cd7632a2ed18d1b3a0b9b1746ff0be2c3be64b52b58a89ff08ab79be791619644ad0e2cf48df1ced4929a8ba0143843cdfb47de602249d16cf60b1a408c7f2242bc95b7c5920eea60892261a86453c82fa2b9a14781bc01a6d5a053256c758ab8810253d55c104045d3022ad1917206f77ec6e6700857183f025f662ab4085e028a1c953f4c4540d369724fe6ef13cb98a806b0033f0d8897767ce155f78a0bdbb4a3130009ff10ac232b771e1d8ada85507cabb9ea47d0fa7d30d78a88ea7a0d9544cde71cb0fb3583ca0393d26c1ff043f482de523c0f6f3eb84d305e2e200013a4f4373073b3f843b8bc6cf74d201d1ccf0a87249f725b06fc9e1d95f246dd76f7ee94f5a09ad491b8003b5ce4468356c44419d85628a94d5c1d3557f548d38eb8c49aefb37477b3345b6aafa2fc536146a77422b4bab4bd0546082e793cfd441db4bf40ca0c99756b940d215eb46f74a8e4bbb00bb960686f64931a3b53eb27a1deaafa6f03d6d0d875c007be52d1b13564706d862d62b20bfa246641d87a94339c7d642061bdcb31ffe41feb56b76976ea36bd7419bbb92dbc51f58453f388ba1515c68aeaa2e72de873b8ad75f2a67dcbd445a25e5980f6ab7751dffaa38fe1d87cec3ea85697058f8f3bc3afd5f7731a530c0612e0619e30f8f68153e6700a5dd8e41c12850192d5a6bdb76054a0ab935ae27a26b563a8431ce1b5c1936414ccad7a2ec1e37b911184603e12fa68bfd0c53d36267f9be7e46c4e65c72fd3e1e2e0ef18772cbc930e0cb235130111457ba34bb09f6e096b491dc1bb39b6b301969bd00163b3256cf44ffbb91e2e8311992909ea84ace6b6ba0296a86d69a4e25f8772839e48f0d2b7f29efaef5a97b44e584efbc6867da7d5c5aab8dbd0d90bee1cfb87e08c2266ffe8d5f960a89d7329d8d626fcf4e28a73ae9aa94d56676b9ab25f4bbd11bdab7634254927dd3d3cb8d43c0ec5dfabef1dc7069555b95c2fbe06468255a6cff4d8033347ea7862b7eedc12ac10d3ebe26a9089e537710b343fb02b44525cdc05b2b7a64e83eafe7e19775a28fed216ab24162d013012bcffd624b6d4b59954a623dc52f6a56fbd8c4571c457731dbd0159dec15297da4f0694a535260fc1e6308cc0c9aefab5f50d113056acac9da3eec944d3e433efe8e3a47136fe43ba022f0c98f53f8444ccdf57df07ca58f9816a1e5ca6f660dc6505590c2f79c915f8fdf669f385284f990ac87aade69e830bfa8d7c6bed244ba9c0ae8919875022e7b53790729e7d24a88628d9cab4d44ab0ad57d61;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h62fa1d02500b707000899815ed00fa2bed12ae2c28f8488d087502178b86a9b2aa9a31d7142f01f0626bf9821247debd603a7e29b6d2913868a7d297ae2c575f63f285b5595bc48784f817b0f89d567831adf9c4df68a743cee816b3d150cb33cb1b73dffab662dc1e9b3066afa63bf44cfbf9e6b858851f0cbae9ae45261edf04c5c15070976c124c01665613af9eda1cdf1e010f8b7fe2bfc97c01724d9d67099a567de7b1fb541e3b55cbd8964271e2544ee528dd04e7f59844d049cc1a35fde7136ffb2884a5ffd47e428683d2d51052cb2360f684e0201bd2508c95ac6ccfc7cd5fe8fda88fa6eee862d5b730545443d6e7342fc4798fef3a8878e127c17ab3a190834dc4819e2882b59d7f474a47d18b5e10c60cda68f5ed8e26ad99d038bf05ec592011be1f80daf59a09e67bb6b3140a0f3941bfc96d1c60ff60ada470300d7b025f1f66923b74c511c74253af989dee94b67f9e852cd7f0ce9bc86dd47045606183fd46b17a6ce41347ca4bd17f135fd28f18fe118e5c4471c9e5f7467297742a100ca5345bb2c9c58d2c4c8580162032bd07c1a3a28a3c42bc3b88664cddd087549b745feaf182e4469d42f5ed95086eef2b47fb665cd2aae99a27e899b6b460d0240073e41a75c32cb0c4d5ebf9631f0e73e1ddb1c698b9efd1615ff3ebbdd4da5db2a03f2a3dbe308572748be8438ee8d401013690f1d5c604b87a3f427170578791da091bdf4b9bc9575b62539aabd59888d89e415ad4c2d0bc837b3d1231223102d11a3f78043d61f60cf170b7f487c91f56f5d4cd694ab0a522945f9df94434a176c0ae0fbbc39af7cf98ed64835da2a84ed766d2bfd162902b9d3e22b9ab78b0526de35a9e3c482daeb9d229a3c10a427b0ecd2ad4004535a0a205471ffc9c41287f54e45ae07d8693e7a3303cd469af427a7887220a26b0e842065c98d90b608fd5a1e14402e60bb9cbe93320c01a34b165da394243269fb375e4a444e9128a02ed53df425fd353667288d9b6041793641038593ede52086cf604695a9f43d24f643082cee9e64310bc7e1d30626bc9019bd96f5a04fba6e938d5918516a566cbdde39cb1a611e288c57bf03c65b2a5dedd18678644e45a3e7fef2e022fda50bdcc8d91d5f03fae40981c214f7fc12c01780629d86648052cd7b21fb602457530e49b8dca15ac722124b69bb20117640ec0f1a43418de59cd682a14464b736d5dd08e45cc86a5d5aae37f77819ec470c3015fba76c44a2f809ef4ccd81321b383947067b4b125b3d2b0cb6ada9c380e48a2c9299b4cd59c38d12c0717f29f24329c46b34ff08ebf4c3a5e706cda4a264cb3108e86165ee52887a7c9c1181e8795899d967d6978c18c45a7b98424f6180a0c154e3466dc53299d579c6219e4d20bd42f8efd973809e54b3ea15d265f8d7661a66715f924020e1f2c480c8518394f388aa1e38efd2b874286c38e43e76cd8f411695ad7b4e25266fb83cbe4c6c422a426b9d12e8cf98c27f12cbf4754fe4b7a088ea6c7710de974e5965021c76d89537943e92a2157c640559743cf4d3e7e010d7e8d045bfcda3f8d2075e1ea7243adb6fc701859b656d02d93838258f5ae6498e44dbf045af5c63d1db9b3405848b957ce9dbe4d0f7392931e2c041a9f9768ad00a774d2b81e2347f0e9ebbe84788453a9c41548674e68e618eb97762aac4ab12adf60e818fef0be8fffc5968b63bf6a356dcc8dff2073f8dd617a46b6f8ee24f473eb5dda06780e19ec782fe12ec6792675da81422c173b0432c868ee96d2bebbd994df2423c7f440dc1327645f2b65834e904747;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h20e7437e10d1f0a88c12e757ba8e94db4baa578e4c8d886a17c5385b743ec595ad9e1ec2b2c3f90ef1fe42d0225af27c7e64bc889818747a7578f79992aa1b893fb139d3130b36f5e71e93d7065559eb9639e5f8d74f741706f04cd1e122dacfa323c1ae6834b86395944587510ba60230661671d9856504b5f4dfdc8c5f9945f7c446a3caa438b027dfbf31bf5697428bb6717a983719e53f37e36d029d7196905733ccdbed6fa6b10f387aaa52880d68982a37a82ca82116ee9d9715930ad9c8ac1557343ce21f7969df114f004f90bd6ffe077cd19634d66241f7f4e2593599ff613263a37a375df52491e804f99360e1a33c9c2e03cc5ca66ff4a8a9dbfa380913c9a85b806364fc2d53d02278b4fef9df31caa9097c9a597b076ef12e7ee0b9599e7eacfe9ea0498d611f0cce0d93691726315ed3703172b782dbeef5fd48a7d206eb08de880ad06c4519660abd31cbc315c268251ea2f5e4977e34b7764e1778240442e14c2c2b6220a280afbcc5d044267a771aba8e2669c22ecd2eaa1f9b08e5d40201734bc31ddcbce2eb8b3be90b13d1736f7e1e18a847a1016b06a0dae7365593a8a63b212067bafc41db4e279f0237a3584b5539885bb5e0f4caefd5f3bf36dfe7674a95f22ab72e638f35b60e5be93f35784640a19cf05205c8992301b990bb75fde731690aed830e485214539b4f70da03d97fcda397a3ff57929307e8a19c6a54a165fdd8f3d926c0aa5a137229b98497861a8ca4c6356283d34c866e4f4e167434e86295ccd6a53a7776910c8c7abf5ed375f7b8be2a0065831d9a30ac0af8e4611a7482c84fc1df4ec8a1786849cb193d481aae82789c005759cb8f305f5f5cc471045dcfc341421f8230fe5cb15c5e40c919d6e6aebcc4e202c531e94f91121ee1b9fe9fcb63d3d2ff85a65b9b415408653fdbde91427e6b3e25cfc0eeaecd46e97a12b8647007ef7ac29185eba007d711bc1f9499746454a8de2ecc80fa87730ac766f7cef3727c0c11e0873d1741147a4ed4d0c1fd1af322be8d11eb23823a415c3028624ae31f27282b597118b5a951d5bd0139e73200f3b576b785199713bda6f1c992b9cddde2d1821517a13f32dcbe646b9e5121a8025a2cb0f941bd7f8047ad0e3e1409d2c6eeff9a6b114a13d977bebf91521b713bac5e7afcd23425de13e3783c49367c0d377c65a1476142f32a3f06b164b4d5a271d0c27259ac7890d11b6eb3e3dc2ecd56c74e2ef8a0286ddaf062964dcaa611b2fed06d07ba68a79a6c6c7fcdc40fdae8fcc2f2d6d4b296479da10fbdd0c48b59d71d49ba95a52626e9be63d2662c4617b3849174641e4d8c671041ed3d0908ce1e4610b4ee48fc586bfa830020465fe93f72a99dc9255fcbbf4893d7b4c2589ab63778f2add1f4eaec9857381c2a92d786271f267047c3cc6e4ebfa77e1cb6b593068b3e3fd7769d3b4b5b9154644146c54ce294978385e98edf45fafb3e2951a7b7af255d10deba9c3f32b21aae71bb1e2436165edf8e7ed7243e117fe3298027bbef37386714a56fde8389992c5896c28a3d30fee59e74b25abad58a79bba9c7fbbbb286f88e4e0b417eb79fee740c02899973c1e54622b3fdf8c4e8ca73f97055cf8cf69201144b1cc971b0b55ca75232cf852539bc9957f6b2c536a7aa5f1723877a5aa650ee27867e260eed078b2f5ae4a669ff38658bec8e6c28855646207a09f4ef8cbf3f3bf15ba7571a6dcf33e1a0e17dd9d1390e44a93b15171cf1a6122df334d657f41c546113c9c5fcf413727db5094be9d2317f9559576081f6118914fd4477e0087d9c1234b2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd87cfbe7831556df027a74b5f2e8cb5fa257a38b8559801c4ccf832700d0efd2faa1a9add78b7a2b3651e8f4798736b8d030f48d07f0431d2bcb7938dff8f7bf671bc2603f906d962a7aef72f31f4591061545bb3e50fa967567fc4446fa7435b6005ad6fc8f0c35aa9faf634d1b363a44c14bb74dfef2b2f98fe6b274de0508c1d0a3683a7992b4f9b613127402a94bc437c21c53e04fce9b6bca17ff0cd21975b5c937510efc2ae5423bb5903c5921090133799f9df8f8600309b1f4ca9e786cc4e8e6401fe3e646a21b31eec232054a853137c14dc0c5e1d779208296bfbc3d56ec90a3f743f604905e3def1beeefc6dca49d618a5127438589cb6c826eeb93c2a7edf1f9e5521fd6bfd25816e5e242a58e9c8d93ef20307bc1ca11b6fb7a1d9f8620433460de9047961fb2e368cb779f8bb26b7d1d44331f1f496fee555f1e703884a08bba845211ad89e257435753b495b5cd49b38c8b52ae79366d56bebaefcc37a5a3b615bd35c5d957a6088263f76febb6780067fbefaa67365f9531240bf9bb854709911d8e032e5a57c209da758e8f2decb375df4efa623b9d28a202bb67cc48fcd8d1313c0980b7e5ba85ac1abfb86cdd2777f0e582db757741ac95eb92449a46637c1c55fe4571313eabdcc63eae0ede8bb347d10f6108a97d953a0d022fb08ecb6e5b8caeb55b34e60d114927377dd0bed5d379986aad3886cdfcee28092ac14ad8bbcfd195f35467099d30c55a1773164977b83ae5464cb72e0ba9bc4d0758afc6117f249083b805b6c90964723dd25cc2223cfc2c7bea38a266fe643e58f083a4e83847c1f46af675e9d9393678065f6ed177586733c761e2f9ca4f3ad83f20fdabaa2f275a8e2fa852896d42c31c3c6bc9498adafb7fb9d4998e13965682b47b18f01769e9703637d8f36e65d91a4b9bdbee8b3979163759b799555c469b99b3d151aef97dc5e37d97912dcdb66df17a4bf927fb60ada321f87f8dbe3bf5a463084996370bac1b4e0500a1a66e54a3e4192c48ba26738cb49cf99acd87682590d5b672a2e316089924d11eba34c3da9d44f4b1503279fd1303b32e09d2679b76d4b55cb021ac2eb10de5180de8a91265d3ae331f4701a35af327e31aa75442a5afbbbc1cbf5ecb76bacc3dfad35c92e1ce9798ccb03d4adde13894f1e9ed226cfc7f11f71f58cca94fddd5e611a45e49422d15d5769b4d7695dab39cd9c9a167356c6350f3408f13684629d03a24a1cc0d76e321240dbe25e6b5a19829e2e6bf0ea884a6459f26cf9f19c31d7418a89a5e868c2cc0c0a74c3d493014abe9f4146df738ed84e6e87fa0031f4070f2a0c1fc781e0d44960a99abfbd0c089fac68d7ab368f2c63f9fe4651b3955de2a3c995ce90a6e422e7159be61800adc010d45f45a575dd146ddcc7eec9dbf141dd65b6901d9395166ed3a896ed572fcf222d0b7ef417a7027a4164ca320dac02af417100113a709441622d6f12dd3b95fba140f5f4eababf547358e98a44bd27f899c8f2b5f1cb7316f2c0ce5a9747dc477b5829825e141394c1a27b4e8cab4658d80df1a19d1681cdef633774108282dc3efaa05b30df51673cf3e222853799429bd64e23931b577dc953e4798e7368b2fcee23ef86113309d0e9e56a5980f8829748e264ed3672e8c1d854ea77bbd5be94836c01192b1855c9a957608fdc552b7b07672e24b41d6be5b6f85b55a893c3b08c82fa2ee3d922c2f6c7063b5c650797ec61ab7120113d5b3ca33c511df14ca26f368b4250e1ed1c85e2e55d14b4bd9bdca38992505aeb5f31cf282bfee5826313ead22726a6fa369;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6d7b6cb14677bc470809ef21bd790830bb0d6bda27319fb8803cb48be044cda3ceff90957addecd14775fd92fc59320f4d8c5a2928bac6f219f5032aeff54388fae9298881eea8828f8ed77e44706e13e4b643a42d56d13f57188a619a9896c30f2146abb9555a71c131e2ef06d2539aff6ed93c776d988e834b9f79e781f9aec69351e8af1096ae70803756a2f475401bf80fe4c4b240d95fc0c3e36b0b1f2f75a607253cd6fb0e732ba7bd1b70d2234f90af8aa1f4f401a6f7fa7c554c08c817f523919fe8ef50cf0031eefcd39da5c20b331c7de6836263ef0af5ed9b5d890225a0eeafb6c7bc20284945b810f1e2dd983b2d69e58fa9dbbc039eab45c62a66d9d7fb8c8c3d3564dc69e9b9b3149685a7ed400fef0c7380f4ae3157e6e65a2e2a3910467a1f5bd57fb8fc5d60b9f3084fac47efde60ca10db2b66b649c158a5f2267f9d6f01394e7ffbb2ae8c1cb48248555b6a531e2fbb840e0921adcf01611ac54fae733472e5ef5bbce4bb9a42f5231e3594b9672f7041a7f40f90e7d26da939f86b85c2f8897405c467fa6675f89e829f14b05cb0c29aaedfedd87ec20c14400b8229324aca3050c35fa644be54a592ec29d10995eca7119308690bc1aace32bb89f00ca877d05ba68cbe6984d57160d7a34f78d9b0786eae067b4ffc5f8d5d2d182b7664dd72b6c61090d0733cdd79431a71ed76b0f3cd6b87b5cfdd74e420f9f64ff7456901797f49a6a9c3a4adaa350d66fccc795a83f51fae4f11244a07ceb2af6abbe29c39edef962729543c03cbb927a2e0f29aeef4a083bb24f643c67a72543390cac57dc178222251a003deb069ac5f7411ccf5715a12801dfc384f742531c3e24acfc4a00b37a960bd8da8eab22e866bea772f2c6d8be29c73c08baf3cf2b1afc2895bb86ecd43c8e70f1fbe7e199276f63fc97d3cae91476bec890f5325732c8cfe3906ec6a5efb121c73b341c553606331067f8d414d2e6253835f5c7f2e452f8c9a7d7f968366a6f649d5767f8cbd2eb11f2deb45e40026cba96f41a563f75fd61b4781a358c4c5bfab528fb5f025ec9ac660e1b3a9598859a49a2a88a92cd0b0dfb1e2cd9aba4fb9b0113f96d3e4c318a25b00256029e20e48cc10cc671270a7836a2f0c30e64eb8ee3b29e399d64167e3e7702eeab3d19de50b3b3fd2129ff13cd7d1f9d4b8731c0a6bfc399cb9af9ccb8cb3bf4b9aa143a9f1e81be20d4dacb1793d88b74387031e2d1a8722ee7d95e4dd02e5eee5dd1e554ecd85060227ca4aa3275178aa58c91f55929f621d5141494cb5e3424adc39ffed54278f5948819af1f1614e403f53499e297fd204bb8cea468083da6982ee5b5c5179af875eba9ca38d1a6dcbe49f3c70fc45fe2177a92bdb837792088f82528f833e68204edfe4c19bc674775223159c99fb3b5e80f57339ae0b122bd11f32b225352293facd854f89e7ffd1731782b3cd5150ef0b920c8b3154821067be5e8de2b87c01af051be4a4bf075dd531a5d4d1acf84d716aab337057c1e96442412dae8249de4025f02987f3d6728c046114b7485f7fe026e2e2707857378ed362178bc2f9de2c2278d36d71be8052cb5cbab0e1a4de27a4bf263fd422f23fdb70c508d06ece0b6382285b703f651d9dc721620169cf27ab39f53dc1cffee96346c564ce177a97213f6a3e5c74989ea66c7a9586b7151f3be7db50f05ca9fc02f45890dae4077cdc9b1aaab8a12df3971970f98fc5080cfae6cf746ccc7da090cc69165df57faaf67155f8ece0917f08fc4b2928312cbe4a879208261c470e5997e89cf79787912ae4b23b82c419;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h43411990d365445dce1dedb1833d972eb1d0e9ec66c229274e6e9b2a6e55c552047937aebbbc1a24606f9e31b0044a93498c932f4564e0e603bd7372fdb0b2cca50bd0eb16f00d174667af962d0b76e3b2963e6b9e84c5706683a3c0253b9d6bf003d52ec54f42e9bd824ff3fbd4d28cd8cd8017bce17530727e6f7aaf008848d418ceaf12a7d44dc1b2933ded0227b9b92ec8b5a375963df7518ca209ae711bb194f7dbbc551d014406b7f765036bff7aa3b683293372af61effda00965b7b6ecd5111526c388fb930cbc63ffb2bc2d231f9dbfb9f00db1ada6c63c8c05505b1e298321b8b893be6ad53e65cc6810d6897b48f0f6566deace215c53c3312e40b0086336e9ef63a34bdb20385b728eff3e85afb6313f726c92e80e69eb2dab36f994ad9923aba224aa2eed1d4a94051ddcaa88e89e486729d26d33a53cb945d1c1ff0cd3fb7b3f117b7c3a1351d12d25dff42b6b225fd12059f76445bb53ddc62f0748fc34464b062bfe46db3fc8de8148764df144947b9dacd9b057d1bb3df4681191abde47fc4b33c5ef033396b6b5b7f1d7c32a8faf8f27e218999554a67e2a1606db93b269cec15be6b4581f2e31c71ba4c2094de79788c20b4d82e28978cd56b235ff12dc3a55c4619799e9b9f4fdedf0a0795823d53907002a47bd4ebde217fc34f7e03cd89066980c4ccfeed12f198bbed9ed17dadc24dc731a038c71167d2d64d65be448f93c7558bb772acd9ee6e013e5f92ee9bda46b575bdfbad275ea719bd536366af966f80e0a401dbdae80c861328f108ec600ab8d196d7c1fa2ccedd39db9ce50f336eecca09dc08479c2d0aa41442ec2bb9570d083f66a7c6bc83da5a7bec4e22d16171c7296b8cce755a57aefe85dd8dbcd765fd11ffd8d5779e45e55a01a32e75fa133310fce91df577b1fffa672d6135c7264e627df1b3a7ba4f62cbfed48b614d3ea3a0a9e37d2a25f24f025a7ac9ec111d4c43fb41016806cf6d8b197eea74c3bd89973f7325763e7d1da15743876d5dc1544ac7f83dba06c924c605e27f01572cde21ac85bc74b34b953b573b72b32abdb84e7d0438712e1e58e14aca45422fc099518118bcb7bdbf89091f7df26513e67627993cca4acebee5a1688e18e756d0be62be231d7054e5fa276c69d7b90a829dcd774ea57cce5b00d504a474a9d9edb049564f8a620000311a5d7ad8880a22c1ef4c20017f09b36d600641990f192bfb37a2990b02a6e16e825f46f88794b13fed0a47967800dabe89369c4c960a6b8a97c89e03e65726d0b2d1243e3927841fa06f45eed0efad7dea476782d5a138229f2fac787c5918adc62f053eb8819d9080b8466efd8f1446c95f577021e4dd229b5947f22bb518703b85a32ba57c1c274039d5f10b60aa5844bea8d974cb8d4cfd065a1f97f33e3e84cd97461b20d660dfde1965b8a0e97a6d30e66823b5cbfc6642d4d3667d001681b6d0c4cd3ef4c31a15c5640fc8aa2c7042e34abcb858a29a5dbe640fb4a287bf60c948a3b8f5727a551d1bc6811581da7d7e3d1a13afc9e50d77a3aef1dfcf5c1838a9348337af3b1a37f0121441d6f75c9984402bef3cb664d0ad3fc47435ff085f602f6449fdae3a8ec27fd62848d2aefbb9923d293ed9be84164c09a0187b712369c1f372c1d1fef4fd9d69908f245bc8bb17ba77e8f315e7f2f91dd38e524242ce2cb26cae4178b17c94baad1341211d582ce4bb42d8224c796b9a9454f9bd5504d6a3c5040e0415110fd4c1579489c305d2e0faff51af1e4765e0d45b432a052586aab7592f941b645e8a2af0f0ea21d45064d7a99020e18;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1f2edce9dbbb888c555e08955dd453419b67c4601a4234b502b9eab44762993c2b959bf2034cfdc91860342925dd5e3119098bdb29e6838be138c402d2b6a682d278a821e69a771f2754112f656074989b6fc8b158c52fdb0437a28d2a192ec9e94ba8c503036d6461fb52ce6ec1a5bb6176d5aa49d4573d4b404d5d3f236344bc149ac7413d1e0923b10361e04741a173b3a3c9d2ff560c04e8d7820d8054d7d5248bc1dc514e6f849f106e3816eb9887fb645f22ac5aea578431cbf2f34e0355f651c7e6bee3073ca5eecdf1be63d14b0ea0227973e65ba8f05d77d28fccec751ca37ef6e995047cae44e9830a042a72a9be0c542e34bd74ddcd66c0d37bd828376a3293d4c479837d492c34dae739904a1262fa4c528c256c0279da107aba819efa68fc154624e812006c871c5fcd490b05e32ca2968f860a12b63200dd2da37d257e5356a6fe3d14c9417b3c88383650a2fe7f94add1edde77937f59c20acdb29f208a0a97802afa230528923058b4c5a872f726689c097534baaaca52fc3a5af52c3068435837f2c318191beafcaf33ebe3962afd1502233ef1881245244f0a8efca7dbdf714e34f2cb110a1e6815e8740da6c1a007accb93ac64c1c255c64297c92aebe03ad22e94efd441e57661c47834d8806331fc27672f8f12b6bca6e53b6037dd7ee96838fe279be51fbb8e217817cc31352345dffeb74ce2919157f021c37366a1b0a9e81635135aeae77a02543671e8a5393a639bc178fb1b7df5554b6526118f68c3611d30a4e057f91c3f4c2944f721d7538a8b537e6fc5124e57dc688974351d123e94a215ecdcdd158fd3375b893326db49547c428c933a295a7a519368250f1eeee8d4ec3baf444c55b625f5309ff13caf44f50bae97c5fced3364a23674074b01972d3e1e1234f4e13d59870a3b71a8911c7c34701d960af2b390c03c3f9238cd427222a9adc2909003e668a7df6d603637b1c225763d8636b2476748b96fc8f2bfee8b6192e9385c0a38f73b581510cfc6006360ee506259ffa9182f7060f3783e52080af81e5ab8418b2997361f2792254f46fa3b44e65fa13b6d3353f957162858f41f0828ba0133336d2c011eb8a5558f5c10d268c8e22e0a0e7f3cbe31debe2b9277b84b9d04ae98b7658aa5a60a55d014db729b6ea7d647b587037ee47656c54b7a0c8610b3061a02657ce9bb9d59c4fb4353ec3938016ba2c4d95aee268b1ca960a7f88f67a876769fc994638b87690d92cd5117c6d22ec3d23960a31ea83df8b658b4466be7a01288d4fa0a3a880472f3d85daed2558ebe78391005db9e2a54fe32ee198911125618cc44d28b87f2c3362c82844982e33f7179ceee6806fbffa22742a7d5b1c5b0a5bbe2908c68aa64f704df1a63f7f88ecc124fee172544f901a0dde27e3a924b171327b663473313ed504e443a63943dd6d34894cf4f73bd075241208c4e7dcac0c79e2e47c5793a0dbb034cb76f4269110e7c836766c8b75c7309b7b2a8190d551ccc3a9e8ae70ae14b8ce0fb41f1d42432fa8fdebce69da006fa6acad063161ed2780ddb3496d54552ede946f6df6ea3f3d61b5ff9c3697e0962c6f82cfb28a9b5653d83cb554ce4b5a46cd4ca22e26d2fbfa016f85f830072c6648ea9dd363e01c48b57c885edf2444ff305eb6c5c18a8bbedb38b87ee6a906d02a90aef367e6189eb74d9c7239aaf22b336d53ac55b13c2cb2375d9e03ba040b3229d090b4a29fb61684438d112a1e649c2062c6cdb37349d90b326385cb7a471f39f1a9951a1a9fd1ebae8c10bb8a4173af87ccfa9b495006258d47c0f7368;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hf1cb8782886eb4d6a2730bb2f1726ed5604229d7aa8f8175c6e38cba7a4ce3b327e1847f965f960c33b9027b4233e71dd817cc6a89422d5315fa43678410af4b20a6fa8c5a7f411429e2a4d3ce85391ae561678cfbb9713d59e4829194e60234e9399cf1a745e6c6474a2fdd437a350ff8810ab1c1e9b7ff5e6dd29dcc43e0e9ac8cf125d80be92a7613bf930aba96b594c59523f5f8398ee8f255c91412f7f9295d3bc76d47d19360f3233b9faa2d3ab3815f02133922cf27726a7007099610be189ef67191ef034963d596f905ea12d497f334ab13802599e96a1cd96c6a77d1cf1cd774c2efb6c83e46d43c4d9eabee69cd1eb30bfe9d73b22a68ecea0bad82381871f4cfac3e91928a56a4ebc606fa0b9fa158e78f7f983a66d15bdd7f1f3ecb5f3cbdf0be39c069e54dacfd7f5d4a366532e210d0c07b21e7bd24384eefc33cda647a416baf6ea5836b402d3f708706396ddea239909971c2a1aeabbea5c9eec45e60b63e9ebd71bb776d763a7ba5d9dae680f016441cd6f81a4e3740a2770917aea72c22436af2a55bdca2551a9f80acbefd8044b53ea5bf771826b261ed16b0c364f41f5bbeb0a5f1aa093c06346de7f4f106a7de51761a68e7f6beba5574b53c01931e897fc1e87a52d28431280926bec741bef92f6151de26574279da1cfba4ec2db356a43a9287d187c7637f2d8476c3dc953b6cee6fdf0fa3ba8bd5dc7e47dddff8fb45c6608422166364a91cee6508d19f6e5bc24b0236ab381ad696537ea2683d378d5a509397350b42afc4ad6bd47300601d914ab2627d39094e606f55dc9ec5ede828475503d29b2a05b338ac2ba9e26531bd0287e16b5a67dce6ba29cafcb40ed57dfbea325080f2c2d13c9fd95ae1d74580ca5ec11d2c557187de6f4c83a5da1a3bdc7027871c8282ec5bb1bb08ad5011d75931bc565b008ff0a30bd74af14dce1cd3fa94342534651377f662d5fe0bf6f7e608ba3a3f960f4d37ee2e29cecabeb5fd73763739bb05a6902f7b923c447b380ca5669eeded94d6328504b500368e7d8c766ca0b3c4d2d1c4a2afd6e9384682db55f3314308ff4da18e0eac15c738234a6d3ac8e0f278c8cec3e217c49f72c56106801ac7945e22eddf6424bb88986f32d2178377ec3d14032f3786f2ed7f51c0545fe32b6e207329228c43f20793e36ac8799910122b48766f98d406c4254848e5318e1585fb28fbbe49290f8f1a18074ffe44488aa38247587d6d63891805c32c2814668a05eb106e253d3053930d857d0314fe359ea9cdec0eea2ca7423d65e5f269aa025c6a0533c0c237cb6e32692d62796efe24cb7483508daf7b9ddd137d992055e6cf8bba0515dae59b0b7339f387b8fbfddb8913d091c9f69e700240f36a678d1a5828a36d562692653900a9fb798b0edb9c9ce0d4f6cf74f3e478f00702170d72b7b537538ee90858297d2837716dc6891924ab0027931cfa417c260f3aec1a11168197c589f4014e103c024043df34c8c04ee4af5ff8eab1597265ef4e629ec540465abf8f3291885f0260ffc91589700e9cc72719680630c73a63a033eab9513c592e6ac2ff0325408a812064ab79ec19af72e2480b281dfa0082f62cc695037e16297284554ea3a79876937f57bcb0b1351161afc214fcbe458157269e4d051c166e2d13befd44089f49f9473a20cd52da60d440234c18411ccb0c54e033ff5df5f8c5d18e6afb7b6305c0b9c5aef01074f5a8ea593e5b21ccfb25d21c6f162dddc57421513dbce6adefdb62968a0820ffd81840c8fd8bc7d1c6879ab8888f3d663c7ac56b0ef429b2afca2fffd0e7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hea662b0df1d019adf6896b7bb5a5acba3a3b9a888d2340f9dec8fb919a2f34ce821f2b55b5c390c7d8b02b3e73ddd12a0de179e56fedb18050dfe4ad268e30e36f5ba05b438e1cbeaf4bd1f4c268d49f497d5edf6f75f517be41cb443e628ff40a95cd05aa052d5a23b8bdcd3891c8e0d3f4bfac4d4f16a752d65b265e59d6cdfe5780a39e1d6a65a54ed1b0dcf6bc0f8fb65d682e9f600bdc9dabd4f03c2205e013b0e22f7af032587fcd98628cc9bc6d11d7ef445ceb82d4f0f52c0dd1a7fcf260fee8999f185d6db744de95549a7de6988f3d49bd998dda4c7bbc3f21f84dc67a2d1139343d045e6b9e1c9c4ddbacf3a6880fc2a60281b5e0bb742cad7c7961ba40ae206ad60390f330de78bc210f8970bab15b9901577dc9c9a6672c7cbf4b8c2fb8f4e1a86529b2c2faaa5ef363fd30f244b6d9e0e14bf50743f8a8047dbc34211be512c332d86e9c7b2ce82878daf2808e42384b1a3552a3260ced9f3af06dadb016b942ef90a53cdb81aa4fba0357dfe00c848488bb50f9b076051e46033a6e4408200cb84553a4083974ff069517d71bd64250d86a52cb6b958a15a8f25e19f1277cbad848e688c19bc42acc7416faaf734fc2a3d7e92afa5626afa5068e37be62893153728fb4fd1255f12ec3d6942de74bac3ef8bffd2ee49fa02a7b771424e1ceebc6eba3aa60ae2aaeba7d2cc18a8e487529fe61d085042a90952951a181b14c1f1401e48a2a6bda4a12eda0f5f27b9e08b5a0247feba2028206f4f1af8e8b3256573e7e94332272a7e42de0eaa37e0c97eaba695330d83104ab267432970343e09446bb1ea2d909ea1a1ca2503fcb95ead145fe1697cc6e41b7d2647b17dd345e61a6bc37ef3ac14093ad619df96a6e7f25e5da8ca63031dd9e95b4b28a02f902a5c9dc9a26addcb61604ab89e5404407832ec1a5a4333a45a229a84e91040c64203994321e4035e9efbee8ff479ba08eb437906318c4bb4efcbce4d36f1591502cc676fe3f9ae3580b5607e511ed576624fc2baab4d80bcc9f72067dbe7cd9aa0e910ba6421fd2b60e2791022b8930c106d3b7caed6bfe5383de510ded5095ee13db1425f061f422a3c5dd167ab66aa75dbda628bd133f821ef7924b6d85a66cfb1d185e2f9675069358bc259695db3437d350ce75a79c0af37882e389bfc1fd030845f84c9a7607acbf1c2310dc3e41c72a977bff29e59e70d719dab214054fda0df5f8c3c0df638c6efc39ac5c511c9a5c75e411ceaee7cabbabb91a6dd4e4a9c195c2f787cee008400a98d3a3a389c93ab5f03f23d781961da5b332f7a3bf5eb14e355a8b20e09656b6bd53d100c9813347876344e592c65e4a01287eccfda19716fe7141395cfba64465dafcdd04c25c12c99d0cf9c8c72b1b9b5c192293cd48b3b15e5a0a37389a4488c64d3471d534b30117769036babec524492ed92b737eff046ace2d79f2ca9c0072d1ce9fb0fb59912463b50ba2c79cfc4219c96e13818ce7d6ec29b0dce8e5838bf33e95734ea5bec269ae45a5f951aba14f602f54ce91d97b0dce0d9e3aa259980b985a3527c321da105f499307e24f26ebfdd5388a97f33295afdc0ad0f47637d4506c475e7d26bfe4d3b4afe33afe6ddd7d7d1737fe38c13747529547ca3eb34ff05e53d674dcb9205967277d73dfe780a22925e234f2357a45287b3b1032286eaaf53f2dbea0c0aaefda24fe8a0c3a4841366fcb055dae00b855d9ff76d5a235fe0ebc4872be65f2cc86698438868895dbc5c4e6bdb5868d66229c6ab1b41eaffe7101ad88ad84104fdb7d12378da021d25fadd89feab28de0c9e4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h341c0e69391faf43331c9cbe2ff96da5820ce27bdc449d5b305bc5ba069680c22b6fdd6cc5ba4f192596151f1eca3b0a384613d742f69c5ffdc9331ed5d5f8011b40eb570e7b1285f7544eb7b8131524748f023f8ac13985847e24a083b83f722cedf400cece5faa2a3875f12ab2541b11cb5eba8b0efc6937da1aafc59c9ffdda2900d4fdc6e62ae066150bbf6d2820fb9546caa392976e493cad8db48d1878f24591e7e9e18e6561bc3b273bb0b80360a27a71ec8e2f247cafd39bda8ce96639e5e0f2f43963ae0775f865cba5241c5ae5bf6e0ba3cc747fc4920f513b2512e71483ddd875cf142913e145e67b18bf11776929498b8bff9e58aa13faf4dfbc57d3cf9c6f7a34d7991a5452212d424949d2cfb7bb6ab04c50b19cce540c7f980c6da9b2090030e4e8b7f9d6a515b75a22172c52985f8596a4de6565621ca698a1780c195066749c5a494f3277bd0fc226c93bdcec150f8101194b2e0b605001684054eb3726e3b9836fb136aeb34bd010c1e397f27858993d6547d8610d833d8f25bf01ff2cedb23b2d5381553c07845f2490d8eeb3abb8967df5dc7bc379d6a6cd371b9e9a9336719b8637d251828a753f316b57a9721ae32ca8e1001d9aa842963590db26efd09a552c3690f7f06dcce042b42d6f764ee78b56582df6b29116308ffded4edb0d05f79ef20cad836e3196b3c1e49ae2a98229f7dc2abef90906c779b673a8185d7f66615150243657efa6994b6ad9c736d28167f947067a6f639752f551d8dee4f75e23d96443755f3546bebb75a7e0a9329127f91939813d5954615574e0a48c1ca22ffcb994e5307628ff3108699504b2ae1779602438f0e7c777dc3a91b866f9ce715008e54ee12b26efd8274713d46ffcbdfe1e4654d1e8ee0d0b6f238c9cd169a1ec1f58e6d958d591f6c346a554f7a9fb67e2a83d3edfb25c718a75a597019362f2d8402288c46ecf48d268a08e1511f953a548176ac9c31e20f91f6d476c7dd93424a722845a68b0634e37e9821c4cc9840289e1c35cf5ee452cd8537186df3d71234301443c3363428345cbe7cbca71dc2cae289fd6d407a9f0b6cb572bd36929874f390f8deca44aa4c0a7d35218ffcc4302ae0fe8e25da11922199805d7b6548e9ddbb3c9e3b8be8cfeec4c9c5a5ec206cd398e6c138d55cc8ace199d9224ecbeeda49adeb7b1fb22f597b2eec1fa729894219bcf70d2234a634bd349c25d6f20dc3f702b72f5b0d71dcaf0cc0e1e4234dc3f06b18fce08c9865150e3a51db15fb0d515d6d98afda8cb1767fb060c96d9eb98ba4669e8f41148f659518d015c1ccb05f6d132ae396d6a95e14e2df7ab1b528a6cec46b5dc6bf0b71afd3f6f867f1e683f1b94a9cec7d14489bc92b1ad6f7659f141672ecd872f92315fdbfe068521b70e192b6113e2dd6ae6ba3c1df23090c509bb7e4f59164c86e3d86053017004d7c769575896de7f77a6829cd6354ebbf89a901b04cc8dcd2f1f2e4a86c7e852abd65f4a7f02ece68198a496034c4cfa420934d0eda0d7b2aa1e968fa96fe182c4473d1c968d79726b9bece5a21c7583639a8a900b20951aaf933868dbe72e064e6307e09bf8af5b54baa3b79bd73613be818df6de5144c595ad0d0b0908ad372df363e53000ded19f6c4ef7a44c167309e0a38e1a76a90d7aa75a4147d7f054eeb6dbd3b5112747386eaa8e1ccd9989446172ed896a17565e130e14e217fdfca6492694f33eebc8d9d0506b09b0a2d4a6769e6463175668ad6d9df5c31e41934f8bc06041276665675d17cc79efb8cd5791f6f1eb4a11a6ce31a9b6e425d2c56fe1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h25791b1aa78f6ad222c17e29ac803fb8f93ce154d943b2c5bf12ca9a0c1a5755c231739bf8447f05f67a7f492cf38e93c0853399475524a7b2e7255a1128a5e6e095b49e7e3ac6d2c067e8deb5971b75d9b3f6a3f049839d912ed6f95831a26876fefd3c0a13f104a86925a176a85c5cc3f0f30aebe452c38d14d364064f52c5c5c203c762d9d80260ad731b60419061b281bb31ac889bbda84c75b317815ca716bd75f7719998bcc4d10ac93b6f92a220e246991a170677c65955bccb1425c8758c38b88e7ec2dfcacd552cbc02f3518d72fa1085de26c4b0d02e04eb927deb9f28aca27dbb4cce6e82c481d510e4b6eebe3fd907eba8d54f9c465b917d2361e6cc95a8d40be91b1d71b572e8ad315784eaa836df4bab625da440664d4d7aeced171b56aa2906c1735bab93bdf92e886481272035c27c47877af36c77f935e7aaa2969d9bd934ce79f5da5845e539438652407719e9ea82561b3e5d1c5dcac6452eb8410d42708d492ad1eda518d51694831683d69d2779cd974f307f44d5ee40c9724f27833945faaf7a4e6b43e39653a830549237abca6bd44f20cdaaac19c789b31a05942cc3ef63105cc4629b11ede4f392d4ba07058466e8250bf365d9162e367b2d28e9a42a6d558bdd8ba0531e5330e597536fbcc1c925a57e48d12c85ede1e9f1fe78091e02e34a37114ccc75dbc9796bbee80cf106350610f75483f58ddc2f760b622e3936db4418e6f1465b633fd555acb2215f96c8f6734ca276c0c48f24d55665b7250bdfabc25ed76438a09472a0cf6994ac1292d38d3edd1e78d430a4f21762e4c57f26d5274c44636508c88a36918ec7e9401dd5657ca67047006185e09be21efdef41aad01ea8360ce04987d17f2b7f636b893eaf6acd8bb230dcee8e1c768830d6f11073fb8b24206e3b8a93bd67a607b3f0e1f8bdd0c56666759fd3934e0f8d39ac8b7df1f1de00f4e7038efd0987d3beb0cd5c0c23e56fdae05f0a3f5fdd6a06fc9cc09222cc9a704dce795538ce261d02c1e0fb41fe1953af53d477440bf9d65092bdd83a1fb4095c5e6844e6cc16b3a6982b718285dfbaaecaa36cb6f43cab36dc70b58485c90a448e7c69edd931b03fc981ba96e7903b39c043c2ee411ff5444e447fb67e984d96133bf7e1c7e48c01b101ef069ac13a10c8fbc8c594ab5c9fe6bb3d060253e30a799c04aca41be3005e1ae82a45255b85f25c2fa6e8ea6be4bd7ec8355ed771b868fd5422b941fffc7aacab42a1fb5e8437b7a7ab2a04d857706218d3a17462eaf11f3e3cadaf593f18eab2e7003550cd4917ffab4043c5cd88d4e8b72d32dd4cb8d2f9daad4ff07a0b70d52c915e7d754c69bc104b7f53ffc369075c0b489fe8050b128f5cae1146bf594aed936cd2a5a3301b284f31cb1c73c10872ac8b6728f10f467beaa05499d2c649e7b703bbe96b3f9f42e92c566e3b906e91507b0487f98456b20242ca385755f6924b8fa77f546fec613b668ad2447de1dedfac2b91a68ef9f913e04701745c405837bf94288c3de021eddf2e226fb24a16ff8d550eeee35fc0931ce395bf0e0ff10f3008a986dd78adda2b9019ffedc10a95821239186760f19077c811db07b7d289685d6608636569b63feb8fe3d8b1a46e0c751ed99926d26e58b473f007cd9b5bb168432787849eb44a68aa287cd52a69b4d85e866fb0b777d525e7ffc1d64a48b3b7592703d3238fd6bed7932c2f567636c088fd7bcf867d31730c70300d175967e36f39dbbe4b2646ee2e5ac9f8473bed12d8959d5f600f23ffac1c0e4c07dbc431fbbcb9e631e880f9e0d9a41f584b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h669211373c9c3da6dc1eb51bf86f09508f5f2de7a33946a2ed8206116327b41ca4edac5733b2a70b82f961cf52e24b32a23732f9b2492fd2ec8be984654b097c42c9ffae45a6ba466605f6d70041ce1f46be4efb57c3a189b463efab07421adf04542d674ad2524333cfcc4df176addfa07cdd8c65e8e39e364948c76f4f197d7298443042e01d445bcc32be8d877006fc460bee4b4d2e137c9895861e4757b9dcbeddeeccbb7c67295ab1802f6bf47ddb00da630f93f261fd83769ff2836953b399a91a145a42a2f16a1e0f413882b560706ba3e7311183af1350e5950ca9ba9ce6c1feacbc999bae265db9b84298aaeeab782e774f3fad9a6f522e3de7f93db47b2eff7eef85f5f27768ef9a1ee458cc795c286f9c35bdc8c03459de654c05ff68bc6fcc1fdf35ed469dcb9df7526bc7e87dd2ec133454b19dc39b218d2d3152946dd0ba1e2194d4f858667ea25414bfd4af3927b369eac83430a62ae4087c848c745b3e1f3566b2235ea3a61a945481e7b07105ff3a13f1dd8b1522996bcbe19e30137da1d02e4c7d92f9bb29fb4c52b3a33e229020cc21d8627f5fb6899081d14805476e627df9e35da08ad646a5039630281003151f4a624156f2154f403da500056df221722988596d030c94cb466b57639cd79668121601c96bb9b94c8d5b5a67ce6bb66574cb6ada5fc8846a745883512c8ddfa595827ccd1915e2a19afb08c3241de99abb30a828e164ec13ef630d7d9ad2f79e079d9022bdfa2eafe4cd2e407a054e26567d483807de5b8fe0494890e69b90a6684a91a38e8b33fee47f2a59f72e2e9887b0b9b8aa25e23f9838e96ba750499d043512b2c6282e1cb9517040c9b8abf1aaf2c8e3dbc54eadd4dad3881abd32b2fc8c6c4d5a404b7e9c172c8d026b6af3deb8b57a554073725176418387ab1748bd540d89733eb73a43f3f5ec12905076da9f28be056fa8c18ee80f26f688c6b13e0ac41c736b121acc61bf601036a19637b7a219a5fd2b3075f72ebc39e5b8ad99e8cb0a51f94931704f9ab1197cbd388cabbef0eb53648e959ac1a8828ce12ee811b234050a6ca967d956e9f53c6e3f642cf3b56902c34f2f3a8db26bb3c7225bca8fe8a69f6b5472b1b0647392554b21ca5f5f1bdc5599791e08ff6f90fa143a094c23e604cc9e4f8427827a357f6b5a0b68c31cecee603ff743613874c24f1429114809279d087e4a194d9b1b6a891342c0846058d8a92dda1d1d3d39e3d1dc0c5cd9b348996725fdefc4b92ce46263bd7ec034ff79efd6125b71880ba8fb58647dd838a37278085e255dcc33f101aceb2052208cf57b21f04dc9ef42234128c6696f1e7c99779d249b528c4ed0f40fed62ed7f96e9ae65ac4c3e8411aaa683c00eb62d02278557844a3971452f3b5ae9cc88d5517c495d328a9fba26da498154fcbc3ea0e2aa972bb56b0faabdbaa0b721ce6623535d2a9c2074bd9ac08b204d4a769de6a345521ac9a433b7d813b0ae449632c7f500bf22bcb062404fd934f0ed4fa03d284b317b0078eec4ed46938380b4e3f623066f96dcc1dd53d633df0800f1b166136f5563f60a40bde33c88b1b2ae244ad748498925cffc4b60406ed16cdc89c2acae83982e4949ee4bff50ab6de6397250326674114ac2f4b9ac47547f26d376784fefd3d510f25e1dcbd9a662e55100fe455cfc94d1d0422d05135537ee1df8bebfcf9f1ff1b63a981a0d871b958908c1670cedd4796e67e1cf278b8aa3993eb21aa5504e827667de02167618e385151c23076ba9ac724f75ee329516f3fd4c651728b9349c90139e911647637ab1321329;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hcf91f59936e4b4da5c5bacc6139d729c36e63af81e2a208f9a74dafac573dfc274dc9738f6a96e8ea86a37e1a01702166da5f91e7501d7480ccdf6e72156b5014ca8d79ac82d8dc433aafd895187ca3f0248fa51ea327b90b56eb7b4e91d37651d659db09bfffc9d654655b1699482f8070b31380dcb680d8c036b20ec078ddca5cbe04ea3b6662f6fb3a5c84d489d945e01cb5f78eb8f53d99828bd28182b694abcda1b0f218f386f3edfa8a23aa5658c1cace3ba146ebeb5c6757f03b8c3f601f6697b66489159c11016f3a1034bc5b8bc53555adcf45bc50d00957bd9c90285c7559a8cc2d8a9978c92c51fc0c488cfdcec7062b1b5116e7fd30eafbf7d985d8e7606a2e5393cbae1c0f68814877c5998f09cc321fc2b3597a233b18e390936e9920ead484586000970b0a34c0e744787013729cad9de375f424b1a1ffabb1643f00e74392aa378077a5b9967bc7cf4d0a97f348a420ddb22948cc70407d99feb5dbc1442bbfd85bf7c2468fc889b4c4ae44b9ceedf6e2a5f4fa8706bb343e63e7858abc776259caa70c435610c659c553f8f0759db2b83c22bcb6fc79d0757ae5ad1e7c377df52248c78a6ad3a2dceddf3617ea811655f54608441bc831c34404bdc19676d2f604da0945dc62497ec3d6c77e973abe1e72aa6ad2b72be5a9eac3732a4fc4c1bea8cec11047840242971067eac4270122dfb3b6cb2d799c2ca345a818e1fd9c8db57776e78787ae90981e051ce74fa0d88584e0d5df90919900f092b364a8321bb22d7be421590a2b52061e232f8a4bcf973290284d6c33b3c64ba34004fd9e605e98fc2d2f9a9767013f49a5a24698b2d935b7b32d27e207fb5faa780e1ef173ba457e6ba4afa34a4a30f5c33043c2fbd76922036b92b45823b8fe979d76ab4c08c773a9b431adccf9f928744095e8ef1b7960a1932d8f627ccaba5151d203e65119adc0d133c9adea0905b8e7a2545906335986cff93e9042ccff496709660f6c0ccff44463a13b3718aaa32b0eb96aa0bd85e48e46526c467acc1b1de2a0210252180607e2dcb0dc3343641bf00d2d60e997e2fdbffe3b520e03452a499e0a51be62bd3c31a350c345fb774d00814b1ca803afa895ff6af8e6f806a370307cc9a00435b3279d0ebfe8b60b2d3f9f08f9ad8070ac4887140f5c31390b918826a0a90176b37bd29fae3f00584ea100427144d508e9fe12e136e14a6db234510dd1de4d35ab7b98603ca57adad812a235ad603622e46f68b755b1e8f4469ed3a537626fdf8134ba975f2196efc5e4b7e7832e94372fc7eb19af4ea3cabf9a2a6ab174c19624133bfd2144a81dce2ec29f278388c2ddd47fa117a45318a6a600bb65cc2c1a76976469d5c420e0108e09c84399cb665905c05dce38c49ea18dacafa7ae6af01b9b9c87448aadfd6c474c505d25a5297b9b1cfadcd913b61e69ffb36f2184cc4e56516e55892da63cec10980ce81dd8e5990f4f8d0bb8b3e4d09ddd36165bbdd2ee3e264630ed829e164a8b914cd799de611a0656388b5eb1d56e27f8541ef5a4b902ac09fb839b065f5b94436f1b56d6c2cb111bbfb9d44f27d4682331c4e9de4b36e1059827787d6e2379b15774e7dacd49f34ab059b05d9688af3e22a9cab41b78028aa9bdb2a0ba20130cac40308e4f46468e8bdcd41cde8c001e5f6963fa9da9d5e387077a5c04e247396ec935301396f617429a5b36f3d3d24eb14a0f3b1a4887216b052966bd36a3fb549048eb2bcf764059140f13b9ee047daad3636fc6baebe141698a41ed69e7e51de1fd8c1b6dc022175a0e4352c447c585325b9a91d1a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h852d73fa10f4371bb402748bc00b5ed10601020acf2f2bfc2328ddc44c404c0bfec6506d53a64d5133b44d237b3609629bfe23bc4def3efa1535e02833a55887571d14d3a7381be939a4ee17317df795243729b2014aeaca8e47ae68a19180e6b4273eead87f7582d0c576764ab41312953ee2d837f584784479c3e11aa04d0a9da7e5c65a64f8d2492e9308e98fdb60ac0a2de433d6b46900a5f7be1cb12ce2f05d90c8c00305c4bd1f7864c394b9afcf17201dfa8ead442b93fb75d55e9f2ca48d75f3d6a6f62d9534849739b0259b0ba1cebf90deb853665216ef8639e868ec8b90db4fbecd2c56f9c7259dbd9cb46a80ab7b1d921c71419c098a1f41546de548b450158a0054143c3cdac21bc76dbf34a47712b1ea3d40f93cc1a7543c41e767b4000d21c0c296c0f981803e276868e9a70179ae4b17f29ebd73b8697efacf9c8f7348ea4eb2b4a85901c4e829ae8857877ee940a8b89c53cb9c9d78b2413f875eaa91b5e1e074ecd711783fb8db24a64fe6bb50679cff282acc24b96cb75468d9955b00c978daaab1407ec2ad2feabb42d65de59fd7533d19018910fe615fb05b04b3f05a264b85d30f87266acc5607c06a5a9a5817706233217d01e41024727304083079ff55f1fe7657c38c1923bb3c72883784b022457ea934cf11bb075c23bd01b9a2feacd188eadcc6ebf688b9cf36092963bcd68e343454672af81ba76318fb0c4f4d372a5b3e082963c8c5bffe70ba9642c30e7c8336c8e4bebeb1e5e6660bde918febef5889d9626445659f748b23a99b7a13fc42440af4854b0d2ff526a9ed4b7715c0d9eca1c3e02a04486557e20046b2aa11b11d410d5f1d7993bf7ead507677cc237bca502b149f1c88c21df76cf5216bc10d0c60385a7d652e4a42cda6c4df036caa9f7bc6d522c460981d56a8664a7f0edac454c6817daa493eaddfe4ece2ef9ccf57b16014cc35fdf403abe755d5e3feeb795791fd24d05881a78e1d00cb27f6961c750aedb3ea62ddf1b3d8a4327ceb8dafbd4746a58595b280c7a1d3d186424e560f14142116ff097e0159289a87956515e9e1c0ac277c825744233f3434bbbf91c6212c41da6bdc955df25c5310d43e247370b1fd8dcda55766f79a3b0c5606f877dcce16b176b07242873fc70b47616ed3f3437aa2ad270ca62183e2a9e02e4b00367bc173ea83825ce0fd4facbdd5667c12fbb3a8a8d5b941c22034377cb898f431f4209c65168371de7ce13897ad387f787f732450ff30985e7be6296458946b197f894dd26260b82a183d4a69cfaae8375c3ca6533bfd75aeac99be0e81eb70d24cecd9ca6fb1e6e7ee95e087e8f68a149cf2a2403e7c6b0d0bc6a87653ed4ff5a9c0b142093f4bb98b5eb67b389154d840c5a23b3b60f64742fc870ca6ecf3daf085a0a7ae0c8fc056d128e21860712775fdc71be2c61ba974759f972c1be551e3d86d91ea33a70fd7b320a1dc887e2d0bf96636ded81f5a7b7fb1c2a2990ae038dccf61f9a9b7b2be3ae92d1e9d222960bb22216ee4a3ca64ed1673e7eab4925dbf1f9aa059492d84346920dca57e0e7bf9e6dd1c6ebaefed009698df0e2f4bf9cc6549cfea9ca99b24246edbc55c2069964a98cd11d6a3ab3b1b0e8a0c0867f518969d2df511337f8a93d20a818c5df3a44c062490e98f3fcce86e6bb18a474646459d43f36a2c003a66b5cab0862d6c4f03bd3c5fd98c87eda7d7c9851700a9b545409a31eeab11d227851f3691c9ac4df23147000cc6307db1c305328c4a4d4b09fdcfe310d679ce5b7b4404a358b8929f3e233ca292e950e78d025f6553ae05;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h61a4bf4cc8864e9c968ecc8fddc292dfbb741939fd2c297fb305a914d19859a0d6caabb2dac8fd89cb5c7ca342611f1e5bb7ee280109c0f65bd2de0ce628a5d9490cbb1886b147fb80f869d264babf60a933b4cd082bd08a30a4110b7dc4d0f3716860f1da300cd302fadb933dc1b926ab7d4e9517c457730a1e097620b7efdd6f873192a522b2303398801b122e0049939fa12230ca679e1f26ec8697d6156bea7099305ef0e8c91833313c2fe4bd8c223f07e334186d64587c70d79e2958fded1ac2d0830710d7617572652e7c16bf390ab218fb7c8b0a3ef6958261bbc501be2ef3463995b4045d45da9d3e9b12543b901892f5f786f21cd34fc30e8845db9c0557abdb054838c8f8008eb5b18dc31ca1aab045721ea26c77e961a30f663232dd52fdbeacd060f2e5c96446561eb65d6b34cfc13b1e82709d814b9997048e36754a6685e53c526c84ca050d7e030027cf4cb10b01b8ed21d05ffd7de8fc08a894710de5840ccd2d4467bb50c1db5b4d182f1d99b5727bb5205a6a6c501c367a6c380f8048d1f411284f5ec74bf146a18374caabbb670c83187922fe30e9419520eae4a6da4a0405d7f8b338e9e392ce522e7e1b6302db5052c0d699d2e0e2d8e4e5860b5a35318921e7c1b585e4b20df7179281c14fbe43c997457c58617b191d8fa6b16fc7ad4c09d425050f43cc22b5287faa5e73d68d03a34cc17c4efc973c509b4aca52eb6e37a2116527332a350c53d6e74324521d6793cf97c9fc8f72a40e19a0961ba4098edf9cd4e6334e11e44905e6f5eaee7475c4c052564c40c229890c9532dc400f7ad070db2db63291ade2fe948fb7b445b929f388e3ccc8268e530bef9a7965860fe120c53aa2a0750300829f463d69a5a7da792a972d52211ab516f7dcf3c27879e6e2772e69b3598e58f97e765be8bc057199849dd78611e15f4c20bb86ec738741a54c1a10610c92c4036cd7af897519463db82ccefa1a9011d062cdaf807cbcadb5109d5bad09b1178ed96c30d96f680345fdb41166ca959e37167a78c7506814b6eb5973b6fd2d7300f141babe04ce8305734e5a063e2ba0623203449ac051047314636454a975080d494aac2f90719044a81277995d6d85ff29c5cf4752e936f24b4351cca0a07abce8939adf33858e1d51cce7170ee733ff96ce7fa8f5740afa2776d484b0f04af492d8eb79a5a35086ea0711111089a4d96de1f2e89451c380d75c61d96aea0852443d21d2f1231e0724f43170c76562d92609f915fcde9b0201db8523df9fc5ba5e0c90c95731758cdefa7c9df73cb8857fe59e82f5346f38a9b1fa295c65406bce39267281809aaec7454f866880e585c225e9e4b23e5b0967329c23063dc107b469b84f4a89d3e81654a0e93aa7dec888cf4db4f3236c0f52688b3784f96c4e0789ae69c615956b5e5e2334d432a8faf14f3cef0c0153e3263a572d46b3e447403dd3eec7082f6b557c8f7c8310055bd6dff1699f830dac6a66ad81d616f86d6b26c93a1c66cd856386ceca07bdd7a221668e0e56940d434f7312ee622f841f1cc578927c5e45f2cdd2cb33f7e696574c3b273776e135569e1672d5982aa3dfc78bae34c5689af68efda0692bc1770f947d3062b7a42e85faa27256d2da002d947f9763d74cb165e8b4e3b1afee1c863186b868c63632e277f80cb8704370ef0672c29ce5ee93a149012da4a82042d1714dd6715bf8c1d891c13badea79522c38b0e5acdf4a06581b80accd5dcc3647c7b08068cd1142ae6829d0e46c806381e4953d8d7482d58484044dc06bc242ec3e013d0b53d1bb4d58966174;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'ha99329146d5adcdbc9a02efdd4a07a260fa5fdcb851293a780107cc18d137634f72753c43343c82e8573145b6800388122134c08a8849c11b3209478a10e7d1893d9a802446095ff6a62a480a7cf002ea52a3eafa46b7ba1fcdafb4153acdd71a765eda612f3d60561ee2ab9ef1d40a597241eb717d0bfb803ab5be2c0a83808391da29a2f8c2f5ae2a743d8d02b11ab565e52d81065841025fdc46c51ccb9e5f4aa240c8120d2e465393431aa80b5efacd51b8b567cca52d8373b04340aa34814ca311cbcdc62ed8db738f45242ce0f0d9739fb64ef763db29452c7cfae088fddfed6a7d23e1b5606caa8b88a06e2401faf51a2297a38f75ab07e80c71dd89398111d2ee2e99c688bcc7718d41f679cd23f3c8edb4484e959671796ad0f4f61cf3ed961e1097a7639eeef00e368b8b4ef78183fbbe0f40ece4e2d8942c6abb81e8d978712bb297ffcab02ece6e4e1a9931a7199d84cdf2a86b1f91b8fc988e1e67389fdd7bbfb1439085ed04779a0bb2a44179883956eeb715cc6014012ab7d73b382ab5957825ebdbfdcef2143028dd3aee5f0121c83c484496553a7dec4183eb236d3d630affbe7502995fe45371e76b603fc5e489ec8552de0d5c80654f577f530ef9e7badf4bf37ad5d90a3cc5107045439317031e233cc1cc2ad1290e0e836dc8008e2bf8318cff3f90c11136e2db629a611a5ae0579722f3d92b106a0a6fb13da447556020f13806ab0656c763c5112c800e01211827735ca08c7081683456b9bd576e28b42e5540025d8c079fe2b6c47aba0e456469f628b8b9e1aa30b5875fd67efc9620d091777acfb65b4a45b12c6e28b82ac24837433296f2f8cad937fc8ca97c70cc1579dd7caa3d748da8fdbfb7ac3a5cdb04f2e9b9322cc03b575adc03a40f30a7d1974a13701e43db87dd76e5430ff8df4c9f33ebe3f1870784b68d8b4bbc189b99a3b20101f4492e0011d865e5b31d13508b711590c584e7671dacb66fbe515e62ef793eed1ccf019ef26a61da2f2d14012cf060847a21dfe5238ea2fccff04326fa16d5a608967a2622d2ce11350f70eae71ebc5776881d052ff8443de66dea18c68f18d883b4081f848742c15c9fa1aa21bdbff26bbb3ed9899ba5e97ad60ff43e5575a6b1174eebb1f8309be7aa1c9e22ee78c169d4cc05b30b2da699cae074e0f518d01dfdd3a58d6952c398213a727796089f9953cc7ca8e36213e24dd76c9781c9de06434334bd2eb7e439224f49106fc8385b9b3e71b5b240fba0936a403d8f066d12bb8b653b945965bd73da71e06a73de8eddd136ed157f7db06f35b272527e9c1cdbc96b0eb8336b15b538106fb0e9dcd3d12c1152ee2cbf6b44fd5ac49f8e313512b120e2a11b11f5cedb355e8b50fbea985d261fd404c0b35ef6ac0132748f175f641ceae74ffdef322d1a70f82f27f0858c8129fd8787f7b242083badf995959b392f1a78e33cedf8aa9ec0097a446b72e764ff8fd9a7e53dd69e5e710a162105c48b270e4752ff83998797bef62ab4ad9e67363eeb8c69fcf96d8a2ed9ea1e949ab533ce37ab4192e9f5efdfba1e81a69688b1a76a1ded064bd4df8dca10e91c9199c2f2ebe3eb26badf580577e87557487d38262ef7c4d32623b128f74e9301b368ae1050a117162546fb47e9aca35a13f720db6097b5fc9de6be42ddabecba257e6d947a6c1cca1c23ba0179a6dcd0beb46d9d81704470593b78331028b28178d2838d4aa3f57abd2b91599b863e3c55c7a80aa710b4119238ab9e9f79e2a5600ecb108572193076de1c038af2d2a5f9e49deae90fc15e4cc45b3fcd0c2e69;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1a59288d6c5df4f1933043adb559de28c4e945ce3edb86800258d8233e94089aefeb59ddefb9ae7934ce375ca99ff51745236dc8d06f7bc2db4db20a257b28a130b9b20f9f442fa899f7fae66ac4437c1795544660718e47460cb757131552dd4eb83529b34ab8a037a69bf1cc923b979ab921f5225aaec4364257ee314c9f2031a4049ac87dfab164cd6ba5c29d64a35c3526c82d0638f4de2afa99dda03b137eeb460e98a37064eed2e26cfa4407ba3ca6d07e46f96959750c5d2e75aa592a276744557f0db25117223b7376b80b39d3cb02d16a56c2526ffd443a8dad16eeaf8dada2e74a1e1d4334181b36a9a2556c1ec6cc54c0f0409947ff4f7f29db6432c69fc0c63f6eccfe7cc92aca051706590e9452d336ad8aa3074c8d540f99de57fa342531ff64e367febc4c418938fc06d2176892f271900d9f5f30d27319ba85c0f10b7629503e9ce06f5d7f36faedf4dc6d6e692974e21b8273a70a533ec89bb522b2294857c5355da8dc0c2630b143d17eda3e131fbcc0f8447e50f1b301454da6af607363cfe62ecfbd78d3084052fd762b468c302f66a96b7ef73806518a9876235d2284104ec045c65709934724126e848d2e9eabf85805044c867a7ef7ba483e8c426e4a9adad79c8699adc7b7aae0d76bf8df5ac7e8d0cb913e53113465c72ba438c4b3d97fb46d0c6a0f03049c778764cc0da56a8508475d116589158b6111d180ff9765e0ae2b6555730b4ac8cda23a0adfd8391a857ef79722193a4815e80b8a3809ed84e196babe4f4359e709e38141ca8925b2f2629ec831798a47d94af63cc50da1e06b14b074b284cd72a3928f4512991febacfa6b6a07327d05a1c662c8b2dbed8819ff7307979801bab683d36ff897b4a210660da4c0fde083f8a37851148f4c2973749dc08abcd9a9cf7e383a75ea0c0992e3faa0a1948ffbc94dd079fec3eef0aa37ab1a76d1f068494ebd4edb16a86347e49f572e8d2da87302317e56a02143bb9e6ceb5c35d5a197510c2de45d0dc517b3aa49b323aa7a63891046c8d7c5ac2aac804154c1190419dd19198339a42cb576d20392d741068da77244cba9d9dfec736cafbd157da8aa8f25ad4ce959307d0f7561065de2a98dcc32dabd39181207790ac5b9cee16c4ea6128b8f7ac85c3382bd0ce79f441a7567c7c5e91d2094856d4562541567c93d618f1917da690ca2714bba5d39c9a32e3055de9931e38ef316075192b37630ddf5fdf467383c5a852a2efaedc76e719cc694e7267dd1c79de564d53b7910668d30e0bc27d3135945aafd7261b0ccd4887674bada7d158c5335611058f17073226a79f65cdfacd2810d6302367f7a762de5d64f22fa99462f58ecd12c58e369484b7b78343404c9a56575c14224183772132a3e76260a77cfe818b4e444dd12da8801e8e833365cb39f91a722cefb8caa3f405ddc24cb674fa731c58188f23c11914b5a1552ea788db3e767a861414f8136c07d018c4291008d961c3dd09eec556d0cc8c11a42fb58807a5457fd7e720f94c98fe17e5ce0c4ce9d96079bdacc454ae2b84aaaa4badc07ec47a89b45c6573873c7d48fbc4ba750c675139439a899d9b7cffe8dfe64ec1974dbfac00488b457da058bc285e7762021d63a1711587456086d079b43501c088f806296940c399e0f34fb7c5bc73105e7d32e46764c94309e804a66ac5a293f68ac9ee0425b943a7e8ef19a23808b334ef39748ca1f7fafb800e55c9fc80d5544a5eda8d34cbf36da971cfb58f814d5f110d0e0a27772c36f05ee6c631e78c6e445226efce4f94e762ea99a489859e6049348fb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h5defc4c13f92043f06575be75b8111dd6842390044d2a39667d196ab7b990d8d13ff272b61485912ef46fbccb65db6701cd866ce5797f5047b008150ffd755ab4e2ac9697a8d050ce90b8db85f1d599c6ced31428d7a620a3108f58657a7d99ba3ae909f0c191937fd919df320c62db08af14f9fb9e50514de019c2723944482543a1c988da7b652729010b75362221ccfef82f0d462571587febad0693f1aecd8cc5bd7e07c8d7b51c8f22ef1980a2c74282339db49052223183e59b65e575f64e72e59748ba16d764833de00f9dcf44a694ece3f42c13560fd400eaef6dbfdcee43a8097a8b011be018aa9ac346ebe5fcb15fe4d58015e591ebce1c998b0fa098d80c67f8dc0c0b21312e13f25e0d4a2e9e057bd3d2d9d52a4ef12a2de4626030b7495acbf0f31fffbe1de92f46bcea26546dd6dbce451caeae3fac97104b32a703bf26ae5bc557f7c02f2b35d18e4a58620f5a0c0e76b5ed0e85d94e50d7e7817c823110f282049f6e44ef3d1f86994895d3a536e799566c785e5f1ed3a46d7a6cedc2487b4811701a78a38aebc7df2a1ff600ca4a341ae795a0fc0aa7ad324b286d57996dc9d652f9e7dd7cbb095c810e3f26538147eb3d875ee47f811b4c1db9cf2ce41727e09f327e4027e946960f2613faa33ae17c82dbdfa284d1813016553ee9b394a98a8f477d921b823ae1708bb8c66e5dc21d5861288ebe710e95a557fe77f009a5bb6ab88719cf19220405221c8d646d3509f3688353bcfb8ac714d429a41759f3476fd3d79efe67e0677ea8974aa3597db1f59d4361f9234f70a2f6f10286f686158042f8b4986730d4523db053d08a942439e8014703eda5f371bed92abfffa5276528bf94d6eae1142ea6d78bd97d21b50d82be1fa211050554af619dc18a534f68eccd1a178b45b9da191b37bcdc039465d8cd810dcecca385662232477b68c382ccace0d5e0022946a7abcc573389bc49660d94e69c404bd97abc2f4827c1fd67a33a8c73f23e32ae18e2133737aba062291e0ec42226416702f61694e0814a83747feec8d3c7c637cbdaa532862e34b8a0df9e830ef04dbef1dd80044655825bc6852b27fd263f21177fc52d3a72b56ea86be30f4b93d77004b24f8f243595ebf19117c44bcfbba96fc4fffb57b3131e84a1dd2890e88a04c88aa9477b3a9915abdf19ef036d7c32b60c7c457a3b1940c434142cec82120df60753bb8ecbf6b9f44e85590d25669ed27b77a700ffe28b820880b33348ed949c8483434e6ed6b0e5e1055b1282cee87d7239933702fb1a26c36eff731b9aecccbb4076565d0db707eebfc7309e14aa4ac93814cdb93eaf544bd5a5f6bfc4540daf83aad8d89afc41449d1a122770d0e47be71e7132c808eddeeb87dc16ffa905ac6421fb7b8599b7115ecc0d6a4da3008dbe7f2df185a85bd9ea7f67961b415451296f534902ea861583f86434762716dc9389b49a27ee30d5885e19486a1e3c51487d17e335cbbaecaffc2a10c3c034e6b80d36b16121deca3768ab00d7b8e238e7fe14f9a1e251da8e2499cd011383adf7578f2dec5bcef2d53511318843044dec1f427eb5b58ecb802a693caf0de2c5c90ca3eb735681f8ceb26d1be36de582a18e8596ada513ec7da4c6b837a7c25a9931e932ec10e35fd4694c20c2c32cd495647f202975a6bea17ff9f24853d685fa4e0b6bbf5f4175d65167e889429e4e7ddd9a762e9caab597ce4425c80574a8fcba6a9a91446af98ee0e3cbd6792433cb78d6d7157c15d5f8a2970c7b550c35987e868628deb78a496d6789aa359cb44b66f11bdd72625c9c371f847;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'ha50705f7fca98f128fe50b933dea449168aa128c3cd77387e756a6ffe09a2fc24e7a639b1e65a5dbc943f0c609340dccac8380b2c21a3277a68a860d9ca7bc50873ca1470a8a21a4c05d3f8777bff254e7261bda9dc7edb7955c3e50a63e1134352f978208d9713d0e9bf7c8f1f3725540734fc59cb6f4bd63496f8b3b96a9eb9e15c4845e9b45eef16b25e2d220379a51a2c7121e6d62bbb67a0f87869c1c07c4deedff36ae39ffc1379ac3b2fa83b7b847a3a29ae265751629485944d28f288908231ffacc68fb4da2e0fb333106ebc2afc2db2514470ce37ea37f13dd86bd4b54385561165a99cb33e3d52cbbf9177204f470a195c977926a684653fb52a3767c9dbe4a8278944a36a391c30556c1dd0032125e59f56aedb986ed038c30d85ad3132fae5ab090cc34b6bcc2b0087fdfa071887345a460ecdac80ac3828acd15e4fd0aee8ba51864c8077ada68f1fa86142356e26c0e449d70a9784d351e18d39ddff44dbb4a0f7fad19ab748ec1ef5b8635abd7025ef5865822f0b1781f7e50ea1cfe5d0755e554f0c0e1cb14a87ab99030117d2dd326d0f9a6e10e0e8f4fb1a615e9a791a164450ded846ccc0e8e3375071ac9b961b2d8f36d5427fdf572c3be302b7e48ebe61f84562c439569ecced8ef47516c1d4c2ad5805962c9e7712d8d76bb4954214ef2e33a120eaabf65385e45a90e2c5091d2821af089b69d4a79e91152a8723f58ab5eae074cd2ad0df1ad2dd404c0d406366a7e93545cf193b3fb91216e5d423d89480ed983920e217d3f8b3e2d9ad8703a56ced6f63b05a0a2e515f47f8e79f3daad6fe42acf5f65f0d4fcae4535d557e25d93c60cb30bd011ee73813c5a9aec675db8c8313ec204c501791b2eb86174ea36982e0b0a3b423fef9970892c7c0209f972259eefa9a55ba3f8713d2f45a4e1806c320eaf3f7d001a1a91746b9ac5fb98845d9c4aaa2148a790c8d382d66c3b592b9e04dc87eec5dffddabd2e8c244fe0812bb4b3800a20bdad3f1cb42710f7b38594739c918a7cd417fa92e8969363571f70e596f58737b87a504690788640ed9a8c3e1a0e0b1d71dffac9e9a4f7f246107378ac5a12a3227aac56097a98f4ebf539e81a208d317736aedea363e614975a7083c71374246fbe92a0bb052e1da414d8b84b0b37c0bbcf1d8a6a983175f131608024f5e56784bed3665c040b0a7100fed786dbb4514bf19573647da7d40e551647694aff4d7dbc6e4de4d4bbefb25b3d6e38dda4daa70648f63552fc29695aa3ac352da5f89857b307f21c57c8d076de485207a2eaed24af045b278aa6cc26148d6f730bf68b1d5bec11bd16f8d2f95c2f2af55c97d0691adde581baf892f4ddfea712b6a808442b2c49878d3afa748021ab275f49f04aa47cbc9161a7ca86da5d3c8586bb37bd4bb185f5a81e1e2f2abc812bc31db14a45220f0eac0dcf2307369f67bd4ea820f8b4e38f96291c9186d033687dad46bfcf60945ccdebaf990bd1571b31a9931d554af0a044659c413ed464559f83c789b11c703769aa6854976044e6a1f248d9f910345892ca0c2a27f9794fdeba6b2fdfea4e7ce38d4a833c700aa462f0e84e59aae9ceda96981a6f3deeff14089e7ffe663dfe518ec8ac4d5f52c36fd4715d61acb8a0cfb7405f430ec8bcc6eb291593d356284aa130021c2ed4ab9df64a6aabec718c8d5e373dd1dc70c3351ca5794c01ebfdcd30b705d1ba1cab57214668491b37c3073c01ee496cc78e8c9d892056cefce2eda877cc24e75e293560efe8557fe707275259fda2c453cd3fcbb6fa8b1a33d6e9e6d4ba94978a1045;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h484d140dfbeea5cdaed3788e8d7c5154b9df2a9a9a1a45fc5eb86fab53405ac8eb0c13c29e6b0eeac854f886d4db961eb2a6f61d37957f2303acd5fe1d4e4efeb1a43184919dddf8c6dade5922f38b98e87c7d3009ee2fce8423bdddfd98c7061ad241132e61f4643294b14f2877dcf20a893add090557e33e4c382ba0adaa433b9270bf754b986b648c6f93b4e2743c49af7bb9dabdff1a00aa17cf4920571ff6058af34b300aaee635b2840ded5ae4ef02f72cb8645ec66957f58ee02023284289399f0302f4e71d9f9f81fca2c8c8f7e1967636462b10f4fd8fc46b2f145203db1aabf2e09391ba25f461317a15780915d7993e80b05562db822963dbdf6a18132f79404633ce841d485d8e114c6cf4d789e8841eb772ba3c17fa3f24ccbd4d67c519d34110f2fcd571cd40d8a6ae3328006ccbaae5f4dad9b2d7aa099c7d94bb7297be9138e201a70c5bdd4bc9cdf67306c88d1842bbf42981add2c48c42291a0db2473076a240c69fb3d38a3949453101c4082fc71ce260d66a5492f9673b6f86217f9ac90b28de15895176fec7157fbabac1ad9c90b301aa56a9f6f0ed16687de657c0effd913c03b48083161c3e2027683b06b3dfec792655e26e5ba0a613400fc7d58d38a78ad9c0a778e84bcc00926158a0ae4af34c2c877702ba43df304bec8dfac0ef1bcc326499ad45ba244a4bac7b1b914a1fc91480b679baa3633327a16c0995cdca693deecadbae0bffb3ae6147529cdd02be68a62ebfaebdd97f8b97796e4b77c2f52999634f0e8cd97645a4d9b76fa8f0a5c661bfc6e53490f4af63645dc9fa32b951baf39c5bfd6ff69e8ce5ffb1e3a541bec0106cd1bca60034ec4bbedb116429a282e86290fd87f7f6e98622559cffce9dc5e409b5fed24ece26adf646dc79667097eb16efd56f21c069bb02e9236c99b402247d8024a65bca77b2208d4387598c4df82c8249e440c45591c060e68dfa0ca80d7f6f887876be21ff89d176344f824861b363fc19312c5bf8f88b28d54139a6cc649eee8edbdbe4023e47f1fcb37753c0fe683b55c556a83e3df77aa096b1644c96b7bd18630fd2d1ba6d60cb93531e89fb5b416e4555c4d81bdf9b80aa42a57a6441eedba37114bc77236625d7beba2e9b48b5b01648d4afa3e5879263af49215a48cf3b042253694cb6eace1062fa715fe01d76fa7490c9ef74026e5ce440d7ef1316a6d66544a5dabdf8eaa56df5e2e623ba52c950fc18e63261ca796e1731ad7384a8b94d38e8fd58d36024d8e8a144fa2ec8332467707208faa9d712bfefd46a7f790a2f6c00e9fe4dea62c79bcee0e34740eedaeae8f411eb8f17c7c1631997df59e436682b6d11546bdbba3bad3be9ffedc2f21e4acbc9a32a60e51aea67c42c9db209458594154ad6bfc9f49e8849d55f45bb3e8d4ddbb1b64c7e219131985740f0f427080e0e2cd097368c95232ac2064be38d088750ad1ca0bac6a984e65a6fbb971575c79ea7346804b19e5e78d547a622431a012d269fb5de8a1bb0db5e47aa13011b977ad37fdf78e29236ad53fe85c6641025b31f974d4640f0f336ea92c3d6ba37a938d8bb822b6112ad27495c3cf17c35acc8702a9072c997a58321049e9c1b49d3a2893cd470ec7fa326d34addc076616af99168cbef61495f7071135021c643b8223e8c66d3b4c0f7038519a03cc548c784e4b9b48e0ccd9ed026268dd89bf878b1d3442a1cdfd0811dab30764e4aaffb9aa5b5b06e66c0e31d5147bf1f8f0747d36fd43fd8b3e021e3b1776406640b883c674645d4284c9584fc50b5774842d56c891dfd160ac61ad9dc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h5269bfb334264c0652739394bc17b820660f677eac0e946ab03b68182bf45a4105f041ea63bf5512104695ab2bfb13d5e8991dff365772e78be3eebc7cfe12d4c12e0d127d588ee1661cfe00b3a673486a49874ae4bd227240c5fc056e11de6384a69d1da659ec02a7d1777877360f1fdab632668c654b8ffd06d47d7134ac70f4959d1e70b7c3b8287036a4b7298648b72672feae9187c28714d4ca579e1d84e6954fe8016578745389b5299bdd9df0f6423651a516f39df64b0f8e01e4ba1f917f0644bb8f9b5c3e9aae76122d7fd5850130194cba958260bb279b56748cd2ebac6bc00152f8595a2104f8e1765bc989f02e84d3a260eb15d92c0ebcd181bb9b753fc58dc7b8fa0a5771c33117078f0403c5265f86e4d54af4b72b1415d92387690cee2107bd94fffdfdedf7a37f8f7c063576eb9472fb08accb330f7312b641685a65238e4375f19d583f60cd006d336a8a752f2592e26778a5cbf94b8e25170a9aa02864c8442bbd9dbdba2db1414e0f96bfd60ebc7d30742832da3e050a85566c2b7d619f7e3f48e858cbf4ba8f4c154c3c5e626b0bb77ef4d2afd273bea9148258f20f934c06765cca6868a6da6fcf32bd7ab5a2a14d352700ebf35d934a681c6940dd1788f921d04f043569db5f852cfe522d048f1fb01fa544e57da9522dd0847c626a02c6f9f2c0b7383219e521d9b9c1850c69c6d39c1d5ed2706c59f1feb2bd03a4ce630e11fe9722dc31e656ab6568a879c4a173d359ef6c264d35cc1331cdc3839338e8464e4bc1eeb9a7b31096281e2a3e71ca0c5a861623624b29491340c6222e02b786b1f6ea03710169e5f102235cbd5ae027d8a319935101bfdf997f77c725ebfb16f07a167e38aa0a7e81a949451ccf55401cb63b5764bc5147d9156e9b03693460727b74b62dbece57f544d768585a22713e0daab62eda0c23fd2fe7986c022e96158fbf3d621a8e7f5354cd7ecc1daad4a71b0b60186e3f7963d58ef73d8e55cd52c28a6099725e26d8d6987e76b50e41f2b5dedc67231bb58cfc1fde6515257e7d22987104d95aa6b0d032b54a1fa9d5ed55fff62d4b9b95eab80efce92ec728a096ef2e9441b14cb40a6b6cd4963365797a7e6b54e9d639ec7dcdd20e2295f2bce0bc2d3451cdceb6d1a08ab4710d7ef982740b0b94a1d074618e6e2d76e64bc474d4b45f75ce9c054fe5cdb7b009d392148e3e57d5c18c7c953b4a5637943043e896c92e84a60af1d8e3ae513487948af213833af60c08b5f179baeb3d43e8f1b25c23e1bee99b6938174852af66b79f837ae31a83f64b3d1749e55839c3486a60d5de40890a6ef307b084bd0bf2b7ba831166189a236247de21b1b5ad90e25040b6b6aa95c9c0103a89a9bb91deb09dc7e0d7f57efb9b4f6509e8cdc46c47e27345551f2f357bbd1b7dcd4fbd428659edc6eba61cdde3145b0980cb509289ca4a87f50af6fee53f581b8d05189db4e797eb6e25d8f55e90cd3b5488fe0986a8dd345c38d07c876cb26c3cacb0cc223919ce5db19f91cbbddcdd6b7fc73c6b2939c82dc3ffe5334ccefc57bb2faf78d8ac2de3175c0e7218a0574dbd4efb715dfae4b71357f2221d2b0b0ab5a9c30d6dfb258b15f1365ddbda855ad06bf4814f47cc2732cf669d1e332b094cf46dbdfc1cd9cc3a62ce1f4057a452f268f84c018936aa96fdf2adc90d338b50a0adcaebf3eff8e161916d73566770527b98eab4cae06fe38e3c9880d88c569733caf4a5f7d37a7cc187f0cf5616a985fec832b43cbc2444876125a24fcd12cf502be3900c4e6b7c5bb8829e48ee85141af26310bd77ae5d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8332435619d12e9db12a804127dde7a502ec85735ef7fa21b96594c3825a4eb67718319130da00407672def8f5fcd2d205218d8b100fcb10a29aa7452311a1529167e40a5fc30d0803bae3f3887aea90aa80831b471a9e0a6aa166246cdf7d30b842a00b2127bb5560d207d64401323808a734e9f345e658538fe15e4f4eaeb3587f1b897de2e7279c08b0be83343ef57d3d00b112f5b9882b21a67f0759082038ffbaea1ce1921bd8e7312513c6daf3d70ae64c2f2c0637201abecc8e2fe3772be047c53718f3beb7d6addaf7b8c6b40d6485313ca3ca3b7380f72558ee2f63061aa6701099b3e04176357a40c66b721ad3ac1a2756e835f9144e0a1d73aa36a633f63e631ef189a8afab591659f5ecca724d859811472bf1d8f4c1f1e23f3674a46941c617cd5091625380ec8189212bf9cc1f750efa2fa9281bfb1906e5ac93bc112955f3cdb3638a6322df5dcbefa7f0c623bdb2c4fb180694e4bb6f9773167b0a6491cb01bc192670e8048d6cf68fdbeeb3f81ed5882aae881f44799765e11cd1f2593ddcfc923790b143052836fa7a86f085fc870885513d01d1010a8de3c34a0ae0e115962161e1a768855afbc8d1c74e2fc0b210340c5520771bce8829129a4393c2051c2f6ca104b4776fcb45d9ce892999d03bc78bfe580451bc31633f621b1460f010b51000e3f154b6dbbb1116a4dad576ca0a9353f424bbba9c638c38e91389b29a61c886a53b5a0f5780dd33ad76833ff28f34581980e0560276241d5dca7eba58ac0d1b0314c59e9240cc6c117012dcd0d5a48e0cb4d57401f8be4e24942ec3ce3d56eec45ab8061a042081e39dc4c1e97fb5435f05e1b63c3cb6d7d76f05632dd4bbd275e1c70be0ae57a650bc263a9984732fbcda9e0ec67db42bf4cb8376d37502028f43a1ca81104dd4f32d4996a824c719b6bde0236ed442c5b2ebb8b105edca0feffd5e2c5421ed67bcafa4ff936a0e558b471d77d93ce1510d976341d121c0d9f96dc3199b5db9aff479a45987446382650b6624b10c4c9e25cd89ca098363cb11d7de758f56bb50eb12e2261c2568910d5f0e63c37ccff1af9af7ef24eb5b97b28c7e0a5a3c27c1590ae7d65977ef8e648825bbe11066ed9743a5b8f590ed1c861381f313f383ce66db277a0b2f5991dbc71a8e939e89ab1c164f5d1a6596515ee8c66e6ca5f5fcac67e5062e48f3cbdd6ffcc7a5090115e78ea858703e34c1dbf69ce476d3554abc2258157ed7be204b90c71b9990ba02c6a3f57be3c3517b706cae085161296ac7b3f00b1bdfb9395db92e36d60025a34eaacee231dc35a9465c0a9be35d7816e9b1f76362be684d42297d09bbc3f53558ecbb8787b1b91a790913edc79ea23077942304bd4e589e8b9bdcf687a6bffc635c64cc362c7b20328d08ed66c58bddc4cef6439f6f98504398ea84f4954ba91652aa968c8369eacd6dca3110b52a729e9fd7b51713a91f1999ca177bfc02a668f699a00d8239eed4850a76ae10a366298b7a7bf714c7b1dfb3742f01b77b122127e40dea2b82a5b9f2a989795b4513b32a8731bdc5d34c7dae4d2a3143ff8ee3ab7029b9a95d01aa64d0fa40e93a605f09468761c86760ce3c88da4f43c716045dd2d27a7027f338c887f76920622f588fb29e6f4d85bc34fd5400530695e0af3adaaf0be7696f34aba107ec9828939845fb22157ce218f40af35342e4482fdf6df617aacc05f949daefbc62229ed7bb895cb1b9e65450b1576d720b1aae78041718c3e9893e74d257f5c58fed29d6380b0da2e5b8318b556ef25bfce27fea728fdf5426948148c8356ad075;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hbcdd81673b97e0cdc7ac7835a203a7fe5269e84c06a05d910870cc667bdf325eb90ca9c069b2ddc5ccae900a2ca08de659e30f21e467339fd7f9299bda76887e05614be498b7381951b1557d7b11bbac3eb9401e0fafdc1b11f8400512740e9c977fef4d31b03436e9dd6d329b36efcd5335c158bc44f3ddbb0c53eccd771d2eba1182980cff93c8b39b139aa47ac823588372faae4bb9c1ca9c61199c296d7ea412d82f399b2c1dd1c5c46bb7253e74945993e4daabd6325824d844846667f62c8f69ab85d5e712c804c188be06fca65b74b22ba523ccceeb8861cb61d4d54e962127a91fd5353776af8146164402cd1cd075b8a024873f32a8e10b074e05899efdae0d21a8a8a729eeafceb5e4dacdde150a0553cdc058fc28d7d22c8682e8fb8228638c8b684b4f50ed2a3b0fa14200fea40fce4aba31959a629cf45250d156269ef23f2f4d6b7aeee109119f8b505203c20b38f120026fc5d2d865f77fd7257629d9e675e75570c499ffe0584daa1798cf648273059b5c7ae1f3f28f806fbb6c290c7fd864dbadcc1a8b9299379dec056927e624ceab12ec985480631c1dbe959491eec76f07a93790f29284930aa5dae4dc4806d4985b61c06b5298caeeae32a731bdb8396a851767f9da1490d257953b00ccc653b3a504cef292a4c2b3bc6f5ba535f45413edd74e1d36826b5a2536fc7069e63c7c7566c927bdadb83725417b143372c3324f568303d0cf3dd2e1e76fa9edbaa0d3123a81d8a7d5733e2aa2213b2973c0c506df907f4c16b1b81b17f0cd867347cbf5f55a7cf8a1c25aed097d92ddbada73f14e31dd2c104fc0c18afbeab89dcb28be0c59876382872067e20e9216de36d6c87b72d3be68a67cd7c77866f851bac6c017681da7d9476287f256c9d8e3cf386ed3b5999f23b1b2a2414a6ce2abb273a3711657b9343d6667a9dc2d260d6da2de1b97887a5278fa28dc5e9b26e0422b8a5ee8672b0035d13bea0db58455928fc4f6d514def4a5a9f9c7c716d00a1c7c67ab03acc793e402640362d0b91029544e3a324fe472803e48a64a316e518f3d982aafce8b3d73bb9752e0db7f3ea352fc60d01cb61f650ec49eb58b6f10bb706511b36798eeeaf0f4d395413d36af80d4d6c7c71343e0c6804a3387b7f667271e7af56281cb34eee85c69d9a5458196f0a8afe9595483f2e3eed954cb016491855c9c42476c4f07bc3b65e2596743972e7b0df93e72c844940064f44d247dfa396cd5b79311879c86fe017cb664afca6e2160b1a8d4ec7c19c171520a16903b97a4cefce642e32810d3f865b057f54228dad98015a62c35cde04cbfeb9ddc0fd5326505976d125d3a060b065ba72daaeeefe49af3a815c4ea7be2ec973638781826ab63abc997146f5f6b8788a0ebd034d51ebc3013b040281dd7b643730394acc4c9aa4d16e24dba40c81c3e2f975850925fea464001e9a375224c329704b7820e43c8861de778c2fe53485c3eee1eeb705728b7bc844cfc09be2b22c1899559d7638707d97968e0199c5a77c9a147f3485466a481d75420e187d2db920f4ade1d9dbe70b9108411c2d8ff3c0cd4565637d707a0cdb67fde213eeffc1b2c8462ac52726d01bac6de8d5bde9f800f163e6315dbec6c2effba1df24878198c4afab424dd8e88850b9206afd0e39ae8502a8c2caa35f9b660ebdc03040ee0b8d4a53bbb407f838a77220588c675a57906aa35096db87c8653064009bc698d7f08482e8215483df23846a09cb81019c90fee74777c1a62837d67edafae9d6354bf24785f88fa542bb28b46ebc65179d2b8dc782f221d7f80ab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc757b53e431ac99abcf092fa1cc370f27dc1b505f9a1a6fc9bd450b45cb95361c2314daf1ca09332d8b0f569b69506b564b113074c4cb0696995c45780c8afb9dadfeeddcb92a01e470ffb02c774d16db64c85586bb55255b384c1611e55bbdfec86b3d0966f605d1f5fde1401cb9c6ddd3825e5e7fae73f6f9fede09343ea8780873b84e629ff4bca4115c51789c32919acf936b3975364d6c64851ef3740435e8d84df28b71fffe4ede057c5daefbdc70931ab510a8f7b7b04bca1b327a0e924a2f916640bb6fad0e996a492294c1753371aee5d1a287ce8611dd2e71d131cecaab5062447d1a5677f0fc9d057e93ca002ee4fb734f745a593ded9dcaac59e120faba57a400fb296144836ad71b9e2ccdf69cbc11d75b0dcc0960cc218e53ecf0d007dca12aeee2dadcf07386b3bacb05de11b7dd93c5ad6d4a1291bf113f9733d745b35803f4f86c1423e5512c22f98442125195cbea55a675e6e46900c0c3af8bb6a70ffc7250e7c1a1d9cff4f138b87a4059000dd18047ed68b53bb6d7cda87c0f1b704b8251c83a2e4ea9aa654c03a05386ca4d6763fdd941c30e885dd35a76fb817941de3f57b5fbc03776dedb9d1aef1d8f304b3f0a7a8f591887df8bb81a24bb27268b4a3d3b0ab3261f06ca7ab52ca14c9c78f0710ab9e39861a756c64574f8d03d26a74aeca1e456f9954092732ece5774221f4aeeaee7abbf3b06be4fd215e577ef333b49a12bd9206c7479316af5e0a3912822e622b6209cd7d4b20a943f00d800191552fd65f8ea619e72e1f55a85dceb6d95e1271f8ecc15c4c444ba9ebdb32c2c886ed7c8c373791fbb126711265e517ac1a2a00eea2d2ceeebe48407e108db84ff2f529e6c05c8e8d91710a5d8b455b6e093190013b58a3f7eea5241b0240b09f6c59975d5a139028ae5a5aca21bf243c3b5fd1b1bdd52d9ab64bf0e4cc5ddc64befa5841844975ad51ba6fc4606739151e1795192aa8d34f4a3b02c78337ebd4b4ff16648b0753048c37691001630bca89b2869d690355ab68cc27e426e973462d3f4d5f344c53dd2088efc7cbb9d9059c5ec90a094f89922ae30fbc87204610f73f180189eab1c0d316630f1a651c03dccea8ca3e7317e0b3c91674d55e6631201ab59bc4b75bc5ed5f14febe73bc34b487faf2ed64d72c6d51721b83e8d13edceeee7a6a990eecc1a4d9506d34b1bb1bb5fc04796e22c1a12f3ffdc64e3d6f4cc5cd454be4669c90866cce32db3040e55778b5bbeaddef2bab828ce99f963c2b3f8ac1a124983fea2090833a577de6b3c879b0e7ef6ae976bada5113d197756c40bd4b465b4ca1c429ef8da519400fa4700f658af540776b357fb86fb9fedfda99ec32f22e86105c5dd8a0c66946c3e073bae8183a32cc8066bafae25ca9a18a589494662482fe066e76e39f9ea8cb836dd7a5d61183ad4ba4fce8e6834897aff51ed1d92d8f2e67b6e57a04a7c0f84ffbd94ae5c670c2e7a3a16358c29885c7775ad6d2d74266c76e5849148c98a9d2a9a8f74a6ae8f541b7e821a420bdcb5d752f8bfb4138a3b399e9f7566f4277c761ecf536ee8a40f5f5e56bdfccf42b9a8fb7531410c6c68abe41ab8d4245b9e7f5171127c2f470e9d1459c0bcd614d90b2741bd6543a81f4a049b9802ea0fc0768a3ad51091c1f146bf6f17759ff4c68215b514b26e9ff23f5c40bf0296e5a13673ff9de298873c3065882a1612ef71e473937f22362f6464a6aadda97ec2685a2d314d6abe087179b4815d7ce6597d92018fc1a4580ba261e4a6b88c0848b4037ec4c52d4d6d1e507b22181c92e068b86f01faec667;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he9b654c85c552bfd7f8c4e04bbff6b7d37a24401a5f4068a04ce4eee15904208880209614b24ba0075e01877e9b537b5e8883810240a7a149857c776489681ef23bbe7162ac54dd36c1912ee833af14e6391e95ae71bc17eb8dcf78b82f78d2a7125e6ff108bd74a0e485f2cf250bcbc2f31b4328d5ad0515e63e0aecc03ce5c59fa774be2627c01b13b2a57034117f41afe60006ff65d60b029c29ffd3435175adf87d8fb45b34fb995d05a8e4074fa5dba6fbb2589f405951698a885049e34677adabc4032e5ff02a3ef60d850c551704618e773f83aad1719624430799b057175fc8e13168d919cddeb10ff6cfc626fe64998f0716a4d33f01fea2acc18c2b5b34e7f2a31ad38a23f33df999d0cba13950af01809d34a4de84ae4e65608ba8a784c602c29dd9c1d2d64181c946305e78fa11d4b3232d1bda6882fa8aeba682080c81f5579aa1c4b2af9c11afc20059b58549c3da1a0b858e7fe9aa2e5c94adc969565b301cf322a57fbaac7e9dc1355baba2eb20986017702b1a4b734459c0d46e80f3fcf0a1d0ca660dcfc400dcfbbbe73f39dd78c8d6862bef30869ecb279ce1d95f93cada64fed509c1d98e81857993be59f4ccb9e44b543b4272b1b3fd6099c7b4b4b9053643efa3ae59d4e3fe32485aa7adc1654d1a28039a6a45491173420fee1629de27278649e7b8c70f93b7787e65f39eef6fe7603d89a8f28f2f6ce5b536afae579a5848df55a718b87ff33ec7672b87b748dc766cf0e9410ee83304c87a26a159b82c0b4e1b9ee90d8dd185414bc49f0e0502ef1ae25876844cfb2b1b9c8fd6fd3d2efcf527bcc9890ef178bebbcf1b1e6b54b14a7ec6b4b6f50a8b37f58539422513992d5da96310a2a69182deeb8c0a13b084128f8ede8f83c5a24aab210d4e1e4571fa575c9884df677711ab85da6bea30fa3bb96645fb05a5c2a954601d47af36aea574cf9d28a48ac9861b16ba5f16c43caded81696fe27dd0da1c762a9f84f804323e6e325ba7c162a720be01755e578c163f175e30f1f7f3cb69284ff5c3628f50ae583ad439a9b5d011e9842a553285d6a09586fd192844389f7df6bb79534a06c7a311015519ebc19857005a3dba674fdb0ac517c045909fc2bdc60acf04e4f163752ffb3d337d2bce787dc6d4359f6b72fc8c28f05124213769508acde5c44d6c0322ac7abd7fd813ff392c99e0107c939d67fc100f844fe35bcd8e4389519dd3b9519d8d1d45bde1e4dabab65955a3928a302a90960af3763129a230307377ddb927121478b6dde6e397b26ebeedb79315fb1a3cf619f59c3020f00ca3661eb326a2704e0bd776046a8a6d10f19a19aa53b770ca8e61b05bec0c79ca0cb1a70c52625c61d235ce926ea08f3171a75bc2bab6983f9f2d5a548d9d7e62b461661da845b3e034a0735f0d8bf051ab61cd1db87eb2f98f5c492d2bff6ad9bd67fb818ca9e955277822d73ce5f73f8a62ee43d21a7d8cbd66a6fa709ed9174075c9158067ba1811fabc37f37f7212cdc3d18625b3e511d9d768f20abb9aa2f0f2b7495cb9bba02cbcf8b032d2c20f92030adfb44c6d1c4a4562e28f1827e217138ef4bba95bb4d4de023b54eea5c31270c8a73c864ab8a7045cc355fda62766f6a700d122aaf44a28c560ec1be401c0dd1e0c3ee353150d8a779f55683d9a983e4c4be181676c0d3ab97a1ad6ca7a05e2c5f3b89277d855c5f1f061da47189fcb36535bcd1a1d8393593363a4e60953e83085f2789a00dbdb417ddf4e9fe88cb9010af99ab64f891ee1b18e6ab6bac942a3117dacb755ce3cd0cc9f601f450db3f0ed5c4ce8c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h361d880f1e9816a39c67292db6e9987a5faaece3f9627d69b3aa9567fb999da9cdc49709413200a2db95482488d3ea9255d2ea98d2499e964089a2ef5b310186e5609a070f01714e9eafdbd1a105f89522d6d34186e2269208d741ba1c658398b085afaf3a3c8ab586b612753dee7101202a50d711d5c6ac53a8a4e2da85b547943aa0eba8e8b1c3400941a97c31e454c5fe92148621da0f459bfab4bbf614f25aca962ee2609f3e1dd492499013922f84bc75178e6f9f4751974cae4db85e870e2d88f309b55126541417103a0c27c1abc099051bac7559cbfe1170c808fc4c7002c3c39ac3240b9b18407d5426afc90700345d1b2d85610f2b0f8d6880588b157921128db54952a0627913ed594b6d2b0c33e181f158b9f5ef0b6734bcdaac23c67f63c809295d4d7e259d298f59eee2e31a43b6b9c6c25c8ff41eff19eb631c3f12befb136521dba39b6635f3b6dfa1d86b281941e008bbc8b8ecfb89139201a8d6935a267a1eef36b96b672ad0d542f2b18f061108a11c3afd487508a1773b2569cc298e2f595329a9fafd3122b26cf8c925b11892f2876a9f68dae1bec939bc4c6dfae7169b37ebcd597a95272618e6e6a8d7b4e8724176d453a3bac02b2e305f5fbd5a052770c9951ed5a45de1b3988c03dae15e30207544b507d6d676367539e4734dbf8e371e2f38a87c165f164cbf96f617cb06c3a2fdef418ab47e1356e08c7caf7742e8c546373b0def72022dde58ad14b590f3d3a0d3098050b62d26a812e36518a43475d43f4a5884d49da3260abdc154bc291a64a0f751e06ab2f8a804be7d040eba3ce2e7785fd84fbdd270a9ad3d0b99ff950b9d2ac2bdf1423d97b3e7b79454ce48b50750e09a80152d245f38f39b3a345ad62fc4ff4142c143100ed4e4fb5169e2ce544b7c7d27acc43ba9f155d389b211d3a5c9fc04b17a496855edafc49e6afaa77aa7b22a6ffb4fd49a81705e92cfb6d114d85a4a4c88d51434dc62e6585ab52ee8c4dfee427307b3d4d10fa19abffaf7e2e23027eb5d31affaa2388dbd6c2fd9344739ab93bf4ae1d50d4cc09cb1e6b0da854d4ae1e4013ab2a2dcfd49db75a4eb051347449026b902036deb3691f4c5a2f80331a58a5a852d27850fe9974aa07165b87fa65763203366acbf08684a8769194ae1ba0f62574d4246cb7683e43ac73775342b8cd1b4bc54f0c487e9d1cf589790ee5d1c2a8ac7c3090bad647afa688eeea48386e0a7cbb5f362fdc47a8cc5ed8d64b0c680df41e899b3d149eae51fa157638fb0a25dd559cc9d561289f74def9a0782225e4fe034169bacf15de52a05c97c4e52af5ba242a4aae680b865b6262b41cc74604068e27b0defe391402f857286db740a5a04cb15de299b90f419d391aa9a1ad5661e6111bbd128a90266626e4289e3c99c76a6a4430f6a1a6b00418fa45996691d692b2971a3cfcd8d263df563d2a202b819cb8325e5206325110ec2ee56accf151f4e40fc838bf4b527f41765edfa43afe6fbfaacc7f6867f3f4036e48111e588ccab292e59d1dc3d3bfed13c907c755a960c5ccfa76e5ebfa49f1e475168d9d5a5a37335d5f5fcf2a49e65877a0e7a0eaf63c179e99e518c8f7a0cd83e881847460fbffc0d17794d9b1c9709a0ecebc2bc381a834aaa32ce09fc3c2d0d58bcdb5c8bd86b4f64bfa391abfd7cb172a34ec76cd836ad602b3e18a270a19b13981b45e73bbeb454586e62a0ebbbdf2a53b214c7d4c89f3d9a2f9a5beb41b7c7ac8c710cdec6b4c8f698e39d38bcf3a772f3d533790f6bfc51bd51710d28289ff281898dd73decf45fc41574de8509;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h28aac545e019a529486987142460430a6876d8291f4371c7f1b2759d2475699d05dd7d3d255c1ef4a5ecb1386aeb4f27bd8a3c823bdc115bbe7585d3da3567ae214cac0040abfdb7ad2a71b57f43f0efd2773061b0a687a300ad2c5ce3679e5231ae6d355f06d699be2892065ded2c4a0d48c2a41c273e11a896f34c30225dd47851804357b61656575b489594f8b757e92f17628a7f5aa26df38d8fbebeecd6561b5f2dc0ff65e8d4072db47996c93d0dc8dac644cab0ba28164ce37c7510c1e3b8de716a072b8e1880f9403c95e7fe28a4cbd86a3bb7b1cedd2b8a78e9ae99e85ce8ce5d7372bddd4e5143140866f3204a23e5f3d0e5064b54e31b1d2cc256ee86343d7658fde749f3ff24b8a3291689b8fafe1698edecdcecfe79bd5ab5e261cbfc599d2dc691694f8ec8e0a1edb527f533bf8162205a5df59761eeb7780d38a941e196c9748b3ca8852533a297a3ff94ec68e72a45e675885dd4a658c3a63e2d8a64a4f15ad4c90f8334f8a3779a95f53671382568e345c89cd804ed9e13ba3f19c29478a9f718e8dc3109c59a74baff2a1d6428fec6e31bc32d42d862e07dcd6d729c7e9e595310363368607fd44af7c5ed4e5d496b79dc6b6efc995cd3ea559a2e6e88a64c194f95f5cd7677db16499fb06341d0d35fc6b91ff6599817994ae6159b6dc248ca8daa7f54848d13de77eb19aa87d59de85e4904515ebe8d2544d9763ce456b9c21a4fe44b8ffa00c1dec99bf5b8d8d8c9f093e22877c50e34abf360a34c8fab39c7bd338b0654cb8e206cfe7029fbae779169cfe0a81ff11644c1f2cb8a035567a2c7109c05fb478b723d5d7012c9333515a87235b487b57a3fa243eeccb95e09a0c5c822dc0e37dc32f76d8cad4ae649637912ede0bafe5c9bfd0ade171d33c1ad02f4cf6e752accc70d2a7f59c96bd2c883738a5004d3768f9f02059a03a7a723eb189eaf73a33e7f07bebcea67f9f739c1a4c1ac0ba6331b581534ea9c6869b34a8892be62a608b49a93f3e9ea72a6b7f211469629de35d1f0f367308cc1cc74a085c5a99d629084df29dd499e02384f72c2c9cbd8b5ba9f8005a6708082a43718de3b8bb164d530b660d92d0253119050d3b73e980266b4031a7435c2ffc9c241579bd13cd890eac00351c93168301cba5480984f0f44d34fa9396831bc75047a17185f1c177e2e2eb43a8f249bfc577331b812f80537589df8293b991cb25963c1663b3f64d032a0959f20920fe3b1534375e121fd555d38da8132ac34737fcbb90795d7aba15124a8a80c16d14df4854f024034c72dc40cfd10f3af4e4aa460a034036040080a22979340de1c033cb588864ef5efa7d5633578c9e240f1d284dbd54b01759b29ee103bb30fc5063de712d1265ef25a84a410898d26e880e4480381f2ae60c04f10cab25827af8a646e259c825a5dc29b83a497f25675235544cde064eb964c77d869f37114b19ca92e362ed8c2211b180492c0cebe5ade4b2754601c86ae71b2819d96d7e625f85bcd21fbbeaad564fc8f434b0e5c066d0ed12cad9653a6a4022d412d2de3622a11975177d69299e74b2c48d1fc0fffd8d46af10435f3b1f987038435c2065aa69c51e45c302d47b0ac15ccfbe5b3d28b2bcea2785a78c0f1535d4c354c0985505b766612d9e675d0c00ead2382e73e2f18b76e9ffcfdf3c083b816193e3929b20eb5eba3f01e92d6eac4bb1c2e167f23cd9aa0228cc778a748fda5f84017f1dee6469a0d8e883ae1d27bc5cd011e9658fda3813d74f6aeacbfef24ba3fb66d1f81183d4a689949cfdc1d587e2806fd45be0f1f69fc8010;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1a34e34085395202b0ff6a20c5552488ef93f42c3e980894a9edf414643de23f3c5b261d0e5eda4f2ae381c518997905fe07b717eb083aceadcaca86bf244d2195357711650a8f341629f928eef4a75a0b3698157f85dc32d54421a74f2ee4cd16c07f5f417350b539f1322119c1e26ebedb20cd82529d19e8319fb87bc39820031c541b5ae5d4a231f0e33bd36c8061d9fbaf3f11f17856de24ac28415fd2e8caf234b6958d53e6507cd3c7a7f6862b584e99d6aec3787070fe1dd88726f6a5674a3d9e7613f6f889e876d7baad51a1ab1d8ce1b595d41379c84a7173744840fc25f1a482a883692bbfb4002d6c9f33118f5179c02614a040430b74ab054d8b1a9606c2190370a31ac6086eefbc2ea62342150a894b406e481bff3f06c683cb702d8ad3e94827d9f1b0ee65440f9f7dbe9c6818e18828fa73b03a8fe05491588da93b1c06717a0f811723496be10aad61a71f54bf87e67494b3f91d2c49e696a832f1b14c6e608a639fc3bd8a8fe06d9e576a4a192df0ddf1a4f4a47acbfe12fab9fc8475e736b43606fc0e23d3a4e7657e256605ce40a4fc786e953a23549d0da75a0812b85ffb87c1c4390274675698c03402ad4d4c08ade921db10fb4c4e1a7c26934f1c96a7717f32fc8cdd105c131026eac67b54065a2b5647dc58812200b1c11a2fb1575074c93f8a41b87df8fe798c0d5d43c026bb97225f7a88d371a5a1b9d43647f748edafbfae70bda37bd8c571f57963bfca526e4d3954a36c3cbd8aba3745886c18b0bfcbf8ce1e02b2e9b970ddf7f516da60018a15df58662a8e0e65faebd0b2dde0c92560454c9930a4e500fb4504c905a67a5fff3ef59e33d8363c2469bd9a0a72457c40878e7a258c876db801bc5535c898d41595dcc8d6ab24e11a669eb5e8402c473985aa6228096c15038d4777ea131feeacc8de7530b5fc71a8e71c94d2862412837b093239c99a14bca09141c977f0d737e4d083e850f7ed8e3b787c9eacee0600026830aa8c751d2539b23785480fade659735ce6b3d14ef3a8575545adfe84272d1091bccda03b41004f25cf4a005ec5f0ac0e807d92f74fa810617020c28bb0b6894be8f447a58e46dbca77a38b5ad9234cdbc47f88fb4ba88b9849d0d254690fc1db864cbeeb0ff09eac766b0334725c5dcb6d113285306759e09ef2c5eeb588a168343edbb5b050045fa6520b858978ec6a5870070230dc10344642c986d134ca269b3f772c18f43157e1894aced4d0d529a18a6eceef3c8f953404b963cf8157792f9be72510348451a8bc5570cae64e5e76c6ed18d9131dba3686c2d5c25177bcafec43ca7e56304bd8db7896772293a9afc2562bd280f4af56426ac2824e9a272c91eec903609aff98866852f7301f3e557058471cc4348f5efc01182dc587a8bcef973310b25cf94d9e54c20749f97fe3d4831ca599f003014c2a22f554b02412f84dbfcf706ffbce05d0995a127ba60839bc3de88992e4aa8d139d8a8372d846b62cc62b76b1ad85a96260642de9ef71680df215be3ed4c68942ea83f7a63038e1503b788ae3bf90cab33b9e85b3b900a69ea21f04f2b5100222f0aa44d0889a9e62b00d324a5a01983aa42ddc00fe0cd119c44a71da451c0ffaafe2128b735efe1761c1dd62b6e62c178905290e73e57c4d5f927454e40e9107902b137c6c81cd0078d4d4d9e6340136c0a8981e13a64b26e597d3384f2e214d719c418f8c4ce0e0ec11419636a0ccb5b08488a4ecd9bb0b09c759558b5dad4a9f8434f1d5d7418cf25a94d83eebc311f3a8083e666b689b82a4e5c925176977ef1d707e7576;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hec02ed9f9bf5af998e292e621f14a6b2d420cac76c37de805f8d1b8f90972d7a4e1addc6b21784b344559bf03e4ae86c17b9195b1b5b7f769f6f3c8cefbb7c4d6084fd0198b4e64d095caa76cc28601b082a3040a777945d83667a31a744638f7e2c1f4c83220239e7128db6ec49fde98d80e92cb1cfc6791e44b8462bc6a67279bd715747ac0d9135594e6d2351d9f5db81f64eca18f0165b1839316a753d7de9dff1d1eb4008d571a03a97a6a2e5cf2c09f07c6ed757660273fa3c7a57afe8102dab0eb6319ea4cb587e9b23a3388fa15413d4f8e0ce7f76ead6d91bfa364d9618a406bc8610f3fa69adabc32645dfed1bf71a267c9eddfd04ed85fbd3cb9f78faa8c997c9ed55ec1667e354fbd3f4c1390202da537c6d3fe6df8015db45530e52e32dd549373ebe7775a5ee17bea1774791062c1aad4abedae6363c00f2e8354971f5b6198e68896abc5eb430306bfcb5c423780e7fd02544b6c3d9d37a6356f62bd6d74064f75c7fa4df606ac27f93976c892902712f5aa2b5fddb619195d9de524ff5aff7e4602c63121b2318df6abee1bdb466a0aebaace19e8d3e9b47fe743d5c4974007714d5d6eeadceb1cbe955cd9d1e8291abdc334c0aa9c2b16917521e075c37dbb5e17e1ab33cea705ef8eb7af5350354d0b6f5c48ec174e01f377b55d54a393d4fd4318fb5d8f157c91699f503eb0c397a6dd47baf29bbc2f07d1bd418e9c8378bdf5c0542b28a49a0c684c53a571bafeb7cc4ae271de1274cc1247e3f5cc6c66a82bc542ffb420cbc7427dffb97a8e404c34fbc0e1cf72b951147869414eb5b21c82f240bb9819838c55f1d71a86ba04b79960b0c7b7f5e18291dcc7e5a363da524ce4005331c8b4e0c2013b77230aa3b0d1ae36ff74f398058d305b54d7f245bdca8ef4c20f54fcd8d6b9509c98036277383aef448a32000858b4cd3f81a67342b0397819e27e4a23d9c2f1803b18e1f740df951cca51ce066689d30b144df47cfdf4630d8e3365278e867bacb75a6ed622ad94c88daa7cdc062d888f37bde1e7bd2f59be6d0423d9cd3da85a9a7de546d3beb73515c5e355e77cf6a8df2f4fd0faf501d5f01c36dd6690c7d9157d45f6c407b4b2ae1d03f95442aa873a89276c35197c80d54665ec88a509c45be9da8443c563db86fba4e39d14241a8099f964b82ff3b7530c102b5221c2b4541ab10eacafdbbbd5b9481c8d08a851620da04e953caeb61f131ac230b342b103ad381147dc9d32387208577dfabe80cc7c91a6b5ab384061241a7258d27baba90aee81dc1c18dbcc4acb7a82f3cd7bf0a095629cb5a7a01b4c251190d82a2c618ab9ac5e1add2e8306abb9cc4e17b1efbc0f37a05945d1f44a8645ae35eda5e12484e5dab26dbba929828adce813cb0ec942dda5e80e83e7a997c20ffdf2849434db0014ae50f3e052d6b6d7d779aee548ea5b48d164400b5200ce6a6266d85ee06917d39ef631db70a66dd499875a81ed2a1c3a9f6c1db52fc748f201c37568def6170256c40d661985d2e8191a2fd429243265ac18784bb3b0297eea128d536430378b00afce0ca6ece0a908cc4cbe8db5f40de0eb0fdbaa1680e1c56c60d1c671eb61a92b746051810e5707d34d8ee9222d00ba8c0bc582f74b64635ef24fb6c0e5ed507b3c2c6b8ff0a695f8fb0550b4e9777735a639321bd7a489084c15558db34a45e62026ef1bb814870416441fadce0ef1f406363100d0eb5aa82de7253df33a62ad10ba1f8c7848d530e13453c3ea7c88be8684d3e6c8ae2a72d39a55e8c1c6731c69fe6cc242b8e6323bbfb22069ca12f416c711673;
        #1
        $finish();
    end
endmodule
