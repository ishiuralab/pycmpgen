module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    compressor_CLA128_12 compressor_CLA128_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA128_12(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [0:0] comp_out17;
    wire [1:0] comp_out18;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], 1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [0:0] dst17,
      output wire [1:0] dst18);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [23:0] stage1_0;
   wire [40:0] stage1_1;
   wire [41:0] stage1_2;
   wire [57:0] stage1_3;
   wire [63:0] stage1_4;
   wire [61:0] stage1_5;
   wire [44:0] stage1_6;
   wire [43:0] stage1_7;
   wire [62:0] stage1_8;
   wire [63:0] stage1_9;
   wire [42:0] stage1_10;
   wire [43:0] stage1_11;
   wire [41:0] stage1_12;
   wire [20:0] stage1_13;
   wire [11:0] stage2_0;
   wire [8:0] stage2_1;
   wire [13:0] stage2_2;
   wire [20:0] stage2_3;
   wire [25:0] stage2_4;
   wire [22:0] stage2_5;
   wire [27:0] stage2_6;
   wire [21:0] stage2_7;
   wire [26:0] stage2_8;
   wire [24:0] stage2_9;
   wire [23:0] stage2_10;
   wire [19:0] stage2_11;
   wire [16:0] stage2_12;
   wire [15:0] stage2_13;
   wire [8:0] stage2_14;
   wire [3:0] stage2_15;
   wire [6:0] stage3_0;
   wire [4:0] stage3_1;
   wire [5:0] stage3_2;
   wire [5:0] stage3_3;
   wire [8:0] stage3_4;
   wire [11:0] stage3_5;
   wire [8:0] stage3_6;
   wire [11:0] stage3_7;
   wire [10:0] stage3_8;
   wire [7:0] stage3_9;
   wire [11:0] stage3_10;
   wire [10:0] stage3_11;
   wire [7:0] stage3_12;
   wire [5:0] stage3_13;
   wire [8:0] stage3_14;
   wire [7:0] stage3_15;
   wire [0:0] stage3_16;
   wire [6:0] stage4_0;
   wire [0:0] stage4_1;
   wire [6:0] stage4_2;
   wire [0:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [5:0] stage4_6;
   wire [2:0] stage4_7;
   wire [5:0] stage4_8;
   wire [4:0] stage4_9;
   wire [2:0] stage4_10;
   wire [3:0] stage4_11;
   wire [5:0] stage4_12;
   wire [2:0] stage4_13;
   wire [2:0] stage4_14;
   wire [4:0] stage4_15;
   wire [1:0] stage4_16;
   wire [0:0] stage4_17;
   wire [0:0] stage4_18;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [0:0] stage5_17;
   wire [1:0] stage5_18;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc615_5 gpc21 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_1[18]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc615_5 gpc22 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[19]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[5],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[6],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[7],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[8],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[9],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[10],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[11],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[12],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[13],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[14],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[15],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[16],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[17],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc615_5 gpc41 (
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127]},
      {stage0_3[111]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[18],stage1_4[41],stage1_3[41],stage1_2[41]}
   );
   gpc606_5 gpc42 (
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[1],stage1_5[19],stage1_4[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[2],stage1_5[20],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[3],stage1_5[21],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[4],stage1_5[22],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[5],stage1_5[23],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[6],stage1_5[24],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[7],stage1_5[25],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[8],stage1_5[26],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[9],stage1_5[27],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[10],stage1_5[28],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[11],stage1_5[29],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[12],stage1_5[30],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[13],stage1_5[31],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[14],stage1_5[32],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[15],stage1_5[33],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[16],stage1_5[34],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[17],stage1_5[35],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[18],stage1_5[36],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[19],stage1_5[37],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[20],stage1_5[38],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[20],stage1_7[20],stage1_6[21],stage1_5[39]}
   );
   gpc606_5 gpc63 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[21],stage1_7[21],stage1_6[22],stage1_5[40]}
   );
   gpc606_5 gpc64 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[22],stage1_7[22],stage1_6[23],stage1_5[41]}
   );
   gpc606_5 gpc65 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[23],stage1_7[23],stage1_6[24],stage1_5[42]}
   );
   gpc606_5 gpc66 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[24],stage1_7[24],stage1_6[25],stage1_5[43]}
   );
   gpc606_5 gpc67 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[25],stage1_7[25],stage1_6[26],stage1_5[44]}
   );
   gpc606_5 gpc68 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[26],stage1_7[26],stage1_6[27],stage1_5[45]}
   );
   gpc606_5 gpc69 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[27],stage1_7[27],stage1_6[28],stage1_5[46]}
   );
   gpc606_5 gpc70 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[28],stage1_7[28],stage1_6[29],stage1_5[47]}
   );
   gpc606_5 gpc71 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[29],stage1_7[29],stage1_6[30],stage1_5[48]}
   );
   gpc606_5 gpc72 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[30],stage1_7[30],stage1_6[31],stage1_5[49]}
   );
   gpc606_5 gpc73 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[31],stage1_7[31],stage1_6[32],stage1_5[50]}
   );
   gpc606_5 gpc74 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[32],stage1_7[32],stage1_6[33],stage1_5[51]}
   );
   gpc606_5 gpc75 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[33],stage1_7[33],stage1_6[34],stage1_5[52]}
   );
   gpc606_5 gpc76 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[34],stage1_7[34],stage1_6[35],stage1_5[53]}
   );
   gpc606_5 gpc77 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[35],stage1_7[35],stage1_6[36],stage1_5[54]}
   );
   gpc606_5 gpc78 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[36],stage1_7[36],stage1_6[37],stage1_5[55]}
   );
   gpc606_5 gpc79 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[37],stage1_7[37],stage1_6[38],stage1_5[56]}
   );
   gpc606_5 gpc80 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[38],stage1_7[38],stage1_6[39],stage1_5[57]}
   );
   gpc606_5 gpc81 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[39],stage1_7[39],stage1_6[40],stage1_5[58]}
   );
   gpc606_5 gpc82 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[40],stage1_7[40],stage1_6[41],stage1_5[59]}
   );
   gpc606_5 gpc83 (
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[21],stage1_8[41],stage1_7[41],stage1_6[42]}
   );
   gpc606_5 gpc84 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[22],stage1_8[42]}
   );
   gpc606_5 gpc85 (
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[23],stage1_8[43]}
   );
   gpc606_5 gpc86 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[3],stage1_9[24],stage1_8[44]}
   );
   gpc606_5 gpc87 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[4],stage1_9[25],stage1_8[45]}
   );
   gpc606_5 gpc88 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[5],stage1_9[26],stage1_8[46]}
   );
   gpc606_5 gpc89 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[6],stage1_9[27],stage1_8[47]}
   );
   gpc606_5 gpc90 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[7],stage1_9[28],stage1_8[48]}
   );
   gpc606_5 gpc91 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[8],stage1_9[29],stage1_8[49]}
   );
   gpc606_5 gpc92 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[9],stage1_9[30],stage1_8[50]}
   );
   gpc606_5 gpc93 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[10],stage1_9[31],stage1_8[51]}
   );
   gpc606_5 gpc94 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[11],stage1_9[32],stage1_8[52]}
   );
   gpc606_5 gpc95 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[12],stage1_9[33],stage1_8[53]}
   );
   gpc606_5 gpc96 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[13],stage1_9[34],stage1_8[54]}
   );
   gpc606_5 gpc97 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[14],stage1_9[35],stage1_8[55]}
   );
   gpc606_5 gpc98 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[15],stage1_9[36],stage1_8[56]}
   );
   gpc606_5 gpc99 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[16],stage1_9[37],stage1_8[57]}
   );
   gpc606_5 gpc100 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[17],stage1_9[38],stage1_8[58]}
   );
   gpc615_5 gpc101 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112]},
      {stage0_9[0]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[18],stage1_9[39],stage1_8[59]}
   );
   gpc615_5 gpc102 (
      {stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_9[1]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[19],stage1_9[40],stage1_8[60]}
   );
   gpc615_5 gpc103 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122]},
      {stage0_9[2]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[20],stage1_9[41],stage1_8[61]}
   );
   gpc615_5 gpc104 (
      {stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_9[3]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[21],stage1_9[42],stage1_8[62]}
   );
   gpc606_5 gpc105 (
      {stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[21],stage1_11[21],stage1_10[22],stage1_9[43]}
   );
   gpc606_5 gpc106 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[22],stage1_11[22],stage1_10[23],stage1_9[44]}
   );
   gpc606_5 gpc107 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[23],stage1_11[23],stage1_10[24],stage1_9[45]}
   );
   gpc606_5 gpc108 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[24],stage1_11[24],stage1_10[25],stage1_9[46]}
   );
   gpc606_5 gpc109 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[25],stage1_11[25],stage1_10[26],stage1_9[47]}
   );
   gpc606_5 gpc110 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[26],stage1_11[26],stage1_10[27],stage1_9[48]}
   );
   gpc606_5 gpc111 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[27],stage1_11[27],stage1_10[28],stage1_9[49]}
   );
   gpc606_5 gpc112 (
      {stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[28],stage1_11[28],stage1_10[29],stage1_9[50]}
   );
   gpc606_5 gpc113 (
      {stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[29],stage1_11[29],stage1_10[30],stage1_9[51]}
   );
   gpc606_5 gpc114 (
      {stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[30],stage1_11[30],stage1_10[31],stage1_9[52]}
   );
   gpc606_5 gpc115 (
      {stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[31],stage1_11[31],stage1_10[32],stage1_9[53]}
   );
   gpc606_5 gpc116 (
      {stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[32],stage1_11[32],stage1_10[33],stage1_9[54]}
   );
   gpc606_5 gpc117 (
      {stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[33],stage1_11[33],stage1_10[34],stage1_9[55]}
   );
   gpc606_5 gpc118 (
      {stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[34],stage1_11[34],stage1_10[35],stage1_9[56]}
   );
   gpc606_5 gpc119 (
      {stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[35],stage1_11[35],stage1_10[36],stage1_9[57]}
   );
   gpc606_5 gpc120 (
      {stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[36],stage1_11[36],stage1_10[37],stage1_9[58]}
   );
   gpc606_5 gpc121 (
      {stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[37],stage1_11[37],stage1_10[38],stage1_9[59]}
   );
   gpc606_5 gpc122 (
      {stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[38],stage1_11[38],stage1_10[39],stage1_9[60]}
   );
   gpc606_5 gpc123 (
      {stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[39],stage1_11[39],stage1_10[40],stage1_9[61]}
   );
   gpc615_5 gpc124 (
      {stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122]},
      {stage0_10[126]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[40],stage1_11[40],stage1_10[41],stage1_9[62]}
   );
   gpc615_5 gpc125 (
      {stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127]},
      {stage0_10[127]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[41],stage1_11[41],stage1_10[42],stage1_9[63]}
   );
   gpc1_1 gpc126 (
      {stage0_0[127]},
      {stage1_0[23]}
   );
   gpc1_1 gpc127 (
      {stage0_3[112]},
      {stage1_3[42]}
   );
   gpc1_1 gpc128 (
      {stage0_3[113]},
      {stage1_3[43]}
   );
   gpc1_1 gpc129 (
      {stage0_3[114]},
      {stage1_3[44]}
   );
   gpc1_1 gpc130 (
      {stage0_3[115]},
      {stage1_3[45]}
   );
   gpc1_1 gpc131 (
      {stage0_3[116]},
      {stage1_3[46]}
   );
   gpc1_1 gpc132 (
      {stage0_3[117]},
      {stage1_3[47]}
   );
   gpc1_1 gpc133 (
      {stage0_3[118]},
      {stage1_3[48]}
   );
   gpc1_1 gpc134 (
      {stage0_3[119]},
      {stage1_3[49]}
   );
   gpc1_1 gpc135 (
      {stage0_3[120]},
      {stage1_3[50]}
   );
   gpc1_1 gpc136 (
      {stage0_3[121]},
      {stage1_3[51]}
   );
   gpc1_1 gpc137 (
      {stage0_3[122]},
      {stage1_3[52]}
   );
   gpc1_1 gpc138 (
      {stage0_3[123]},
      {stage1_3[53]}
   );
   gpc1_1 gpc139 (
      {stage0_3[124]},
      {stage1_3[54]}
   );
   gpc1_1 gpc140 (
      {stage0_3[125]},
      {stage1_3[55]}
   );
   gpc1_1 gpc141 (
      {stage0_3[126]},
      {stage1_3[56]}
   );
   gpc1_1 gpc142 (
      {stage0_3[127]},
      {stage1_3[57]}
   );
   gpc1_1 gpc143 (
      {stage0_4[126]},
      {stage1_4[62]}
   );
   gpc1_1 gpc144 (
      {stage0_4[127]},
      {stage1_4[63]}
   );
   gpc1_1 gpc145 (
      {stage0_5[126]},
      {stage1_5[60]}
   );
   gpc1_1 gpc146 (
      {stage0_5[127]},
      {stage1_5[61]}
   );
   gpc1_1 gpc147 (
      {stage0_6[126]},
      {stage1_6[43]}
   );
   gpc1_1 gpc148 (
      {stage0_6[127]},
      {stage1_6[44]}
   );
   gpc1_1 gpc149 (
      {stage0_7[126]},
      {stage1_7[42]}
   );
   gpc1_1 gpc150 (
      {stage0_7[127]},
      {stage1_7[43]}
   );
   gpc1_1 gpc151 (
      {stage0_11[126]},
      {stage1_11[42]}
   );
   gpc1_1 gpc152 (
      {stage0_11[127]},
      {stage1_11[43]}
   );
   gpc2135_5 gpc153 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc154 (
      {stage1_0[5], stage1_0[6], stage1_0[7]},
      {stage1_1[3], stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[1]},
      {stage1_3[2]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc155 (
      {stage1_0[8], stage1_0[9], stage1_0[10]},
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13], stage1_1[14]},
      {stage1_2[2]},
      {stage1_3[3]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc156 (
      {stage1_0[11], stage1_0[12], stage1_0[13]},
      {stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19], stage1_1[20]},
      {stage1_2[3]},
      {stage1_3[4]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc157 (
      {stage1_0[14], stage1_0[15], stage1_0[16]},
      {stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25], stage1_1[26]},
      {stage1_2[4]},
      {stage1_3[5]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc158 (
      {stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31], stage1_1[32]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[0],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc159 (
      {stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37], stage1_1[38]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[1],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc160 (
      {stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[2],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc161 (
      {stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[3],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc615_5 gpc162 (
      {stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage1_3[18]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[4],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc163 (
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage1_3[19]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[5],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc164 (
      {stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31]},
      {stage1_3[20]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[6],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc165 (
      {stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36]},
      {stage1_3[21]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[7],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc166 (
      {stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_3[22]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[8],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc167 (
      {stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_4[42]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[7],stage2_5[9],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc168 (
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32]},
      {stage1_4[43]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[8],stage2_5[10],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc169 (
      {stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage1_4[44]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[9],stage2_5[11],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc170 (
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42]},
      {stage1_4[45]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[10],stage2_5[12],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc171 (
      {stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage1_4[46]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[11],stage2_5[13],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc172 (
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52]},
      {stage1_4[47]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[12],stage2_5[14],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc173 (
      {stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage1_4[48]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[13],stage2_5[15],stage2_4[20],stage2_3[20]}
   );
   gpc606_5 gpc174 (
      {stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[7],stage2_6[14],stage2_5[16],stage2_4[21]}
   );
   gpc606_5 gpc175 (
      {stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[8],stage2_6[15],stage2_5[17],stage2_4[22]}
   );
   gpc606_5 gpc176 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[9],stage2_6[16],stage2_5[18]}
   );
   gpc606_5 gpc177 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[3],stage2_7[10],stage2_6[17],stage2_5[19]}
   );
   gpc606_5 gpc178 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[4],stage2_7[11],stage2_6[18],stage2_5[20]}
   );
   gpc615_5 gpc179 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[18]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[5],stage2_7[12],stage2_6[19]}
   );
   gpc615_5 gpc180 (
      {stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21]},
      {stage1_7[19]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[6],stage2_7[13],stage2_6[20]}
   );
   gpc615_5 gpc181 (
      {stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25], stage1_6[26]},
      {stage1_7[20]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[7],stage2_7[14],stage2_6[21]}
   );
   gpc615_5 gpc182 (
      {stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30], stage1_6[31]},
      {stage1_7[21]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[8],stage2_7[15],stage2_6[22]}
   );
   gpc615_5 gpc183 (
      {stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage1_7[22]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[7],stage2_8[9],stage2_7[16],stage2_6[23]}
   );
   gpc615_5 gpc184 (
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_7[23]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[8],stage2_8[10],stage2_7[17],stage2_6[24]}
   );
   gpc615_5 gpc185 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28]},
      {stage1_8[36]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[6],stage2_9[9],stage2_8[11],stage2_7[18]}
   );
   gpc615_5 gpc186 (
      {stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[37]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[7],stage2_9[10],stage2_8[12],stage2_7[19]}
   );
   gpc615_5 gpc187 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38]},
      {stage1_8[38]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[8],stage2_9[11],stage2_8[13],stage2_7[20]}
   );
   gpc615_5 gpc188 (
      {stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_8[39]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[9],stage2_9[12],stage2_8[14],stage2_7[21]}
   );
   gpc1163_5 gpc189 (
      {stage1_8[40], stage1_8[41], stage1_8[42]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_10[0]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[4],stage2_10[10],stage2_9[13],stage2_8[15]}
   );
   gpc606_5 gpc190 (
      {stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48]},
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage2_12[1],stage2_11[5],stage2_10[11],stage2_9[14],stage2_8[16]}
   );
   gpc615_5 gpc191 (
      {stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_9[30]},
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage2_12[2],stage2_11[6],stage2_10[12],stage2_9[15],stage2_8[17]}
   );
   gpc2135_5 gpc192 (
      {stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_10[13], stage1_10[14], stage1_10[15]},
      {stage1_11[1]},
      {stage1_12[0], stage1_12[1]},
      {stage2_13[0],stage2_12[3],stage2_11[7],stage2_10[13],stage2_9[16]}
   );
   gpc606_5 gpc193 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6], stage1_11[7]},
      {stage2_13[1],stage2_12[4],stage2_11[8],stage2_10[14],stage2_9[17]}
   );
   gpc606_5 gpc194 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13]},
      {stage2_13[2],stage2_12[5],stage2_11[9],stage2_10[15],stage2_9[18]}
   );
   gpc606_5 gpc195 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19]},
      {stage2_13[3],stage2_12[6],stage2_11[10],stage2_10[16],stage2_9[19]}
   );
   gpc606_5 gpc196 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25]},
      {stage2_13[4],stage2_12[7],stage2_11[11],stage2_10[17],stage2_9[20]}
   );
   gpc606_5 gpc197 (
      {stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21]},
      {stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage2_14[0],stage2_13[5],stage2_12[8],stage2_11[12],stage2_10[18]}
   );
   gpc615_5 gpc198 (
      {stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25], stage1_10[26]},
      {stage1_11[26]},
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage2_14[1],stage2_13[6],stage2_12[9],stage2_11[13],stage2_10[19]}
   );
   gpc615_5 gpc199 (
      {stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30], stage1_10[31]},
      {stage1_11[27]},
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage2_14[2],stage2_13[7],stage2_12[10],stage2_11[14],stage2_10[20]}
   );
   gpc615_5 gpc200 (
      {stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_11[28]},
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage2_14[3],stage2_13[8],stage2_12[11],stage2_11[15],stage2_10[21]}
   );
   gpc615_5 gpc201 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_11[29]},
      {stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31]},
      {stage2_14[4],stage2_13[9],stage2_12[12],stage2_11[16],stage2_10[22]}
   );
   gpc615_5 gpc202 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[32]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[10],stage2_12[13],stage2_11[17]}
   );
   gpc615_5 gpc203 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[33]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[11],stage2_12[14],stage2_11[18]}
   );
   gpc615_5 gpc204 (
      {stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43], 1'b0},
      {stage1_12[34]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[7],stage2_13[12],stage2_12[15],stage2_11[19]}
   );
   gpc117_4 gpc205 (
      {stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[18]},
      {1'b0},
      {stage2_15[3],stage2_14[8],stage2_13[13],stage2_12[16]}
   );
   gpc1_1 gpc206 (
      {stage1_0[17]},
      {stage2_0[5]}
   );
   gpc1_1 gpc207 (
      {stage1_0[18]},
      {stage2_0[6]}
   );
   gpc1_1 gpc208 (
      {stage1_0[19]},
      {stage2_0[7]}
   );
   gpc1_1 gpc209 (
      {stage1_0[20]},
      {stage2_0[8]}
   );
   gpc1_1 gpc210 (
      {stage1_0[21]},
      {stage2_0[9]}
   );
   gpc1_1 gpc211 (
      {stage1_0[22]},
      {stage2_0[10]}
   );
   gpc1_1 gpc212 (
      {stage1_0[23]},
      {stage2_0[11]}
   );
   gpc1_1 gpc213 (
      {stage1_1[39]},
      {stage2_1[7]}
   );
   gpc1_1 gpc214 (
      {stage1_1[40]},
      {stage2_1[8]}
   );
   gpc1_1 gpc215 (
      {stage1_4[61]},
      {stage2_4[23]}
   );
   gpc1_1 gpc216 (
      {stage1_4[62]},
      {stage2_4[24]}
   );
   gpc1_1 gpc217 (
      {stage1_4[63]},
      {stage2_4[25]}
   );
   gpc1_1 gpc218 (
      {stage1_5[60]},
      {stage2_5[21]}
   );
   gpc1_1 gpc219 (
      {stage1_5[61]},
      {stage2_5[22]}
   );
   gpc1_1 gpc220 (
      {stage1_6[42]},
      {stage2_6[25]}
   );
   gpc1_1 gpc221 (
      {stage1_6[43]},
      {stage2_6[26]}
   );
   gpc1_1 gpc222 (
      {stage1_6[44]},
      {stage2_6[27]}
   );
   gpc1_1 gpc223 (
      {stage1_8[54]},
      {stage2_8[18]}
   );
   gpc1_1 gpc224 (
      {stage1_8[55]},
      {stage2_8[19]}
   );
   gpc1_1 gpc225 (
      {stage1_8[56]},
      {stage2_8[20]}
   );
   gpc1_1 gpc226 (
      {stage1_8[57]},
      {stage2_8[21]}
   );
   gpc1_1 gpc227 (
      {stage1_8[58]},
      {stage2_8[22]}
   );
   gpc1_1 gpc228 (
      {stage1_8[59]},
      {stage2_8[23]}
   );
   gpc1_1 gpc229 (
      {stage1_8[60]},
      {stage2_8[24]}
   );
   gpc1_1 gpc230 (
      {stage1_8[61]},
      {stage2_8[25]}
   );
   gpc1_1 gpc231 (
      {stage1_8[62]},
      {stage2_8[26]}
   );
   gpc1_1 gpc232 (
      {stage1_9[60]},
      {stage2_9[21]}
   );
   gpc1_1 gpc233 (
      {stage1_9[61]},
      {stage2_9[22]}
   );
   gpc1_1 gpc234 (
      {stage1_9[62]},
      {stage2_9[23]}
   );
   gpc1_1 gpc235 (
      {stage1_9[63]},
      {stage2_9[24]}
   );
   gpc1_1 gpc236 (
      {stage1_10[42]},
      {stage2_10[23]}
   );
   gpc1_1 gpc237 (
      {stage1_13[19]},
      {stage2_13[14]}
   );
   gpc1_1 gpc238 (
      {stage1_13[20]},
      {stage2_13[15]}
   );
   gpc606_5 gpc239 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc240 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc241 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc242 (
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage2_4[6]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[3],stage3_3[3]}
   );
   gpc615_5 gpc243 (
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[7]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[4],stage3_3[4]}
   );
   gpc615_5 gpc244 (
      {stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20], 1'b0},
      {stage2_4[8]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[4],stage3_4[5],stage3_3[5]}
   );
   gpc606_5 gpc245 (
      {stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[4],stage3_5[5],stage3_4[6]}
   );
   gpc606_5 gpc246 (
      {stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[5],stage3_5[6],stage3_4[7]}
   );
   gpc615_5 gpc247 (
      {stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_5[18]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[6],stage3_5[7],stage3_4[8]}
   );
   gpc615_5 gpc248 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[3],stage3_7[6],stage3_6[7]}
   );
   gpc615_5 gpc249 (
      {stage2_6[23], stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27]},
      {stage2_7[1]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[4],stage3_7[7],stage3_6[8]}
   );
   gpc615_5 gpc250 (
      {stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[2],stage3_8[5],stage3_7[8]}
   );
   gpc615_5 gpc251 (
      {stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage2_8[13]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[3],stage3_9[3],stage3_8[6],stage3_7[9]}
   );
   gpc615_5 gpc252 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16]},
      {stage2_8[14]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[4],stage3_9[4],stage3_8[7],stage3_7[10]}
   );
   gpc615_5 gpc253 (
      {stage2_7[17], stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21]},
      {stage2_8[15]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[5],stage3_9[5],stage3_8[8],stage3_7[11]}
   );
   gpc606_5 gpc254 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[6],stage3_9[6],stage3_8[9]}
   );
   gpc615_5 gpc255 (
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26]},
      {stage2_9[24]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[7],stage3_9[7],stage3_8[10]}
   );
   gpc615_5 gpc256 (
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[6],stage3_10[8]}
   );
   gpc615_5 gpc257 (
      {stage2_10[17], stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21]},
      {stage2_11[1]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[7],stage3_10[9]}
   );
   gpc606_5 gpc258 (
      {stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[2],stage3_12[4],stage3_11[8]}
   );
   gpc606_5 gpc259 (
      {stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[3],stage3_12[5],stage3_11[9]}
   );
   gpc606_5 gpc260 (
      {stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], 1'b0, 1'b0},
      {stage3_15[2],stage3_14[4],stage3_13[4],stage3_12[6],stage3_11[10]}
   );
   gpc606_5 gpc261 (
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[3],stage3_14[5],stage3_13[5],stage3_12[7]}
   );
   gpc1_1 gpc262 (
      {stage2_0[6]},
      {stage3_0[1]}
   );
   gpc1_1 gpc263 (
      {stage2_0[7]},
      {stage3_0[2]}
   );
   gpc1_1 gpc264 (
      {stage2_0[8]},
      {stage3_0[3]}
   );
   gpc1_1 gpc265 (
      {stage2_0[9]},
      {stage3_0[4]}
   );
   gpc1_1 gpc266 (
      {stage2_0[10]},
      {stage3_0[5]}
   );
   gpc1_1 gpc267 (
      {stage2_0[11]},
      {stage3_0[6]}
   );
   gpc1_1 gpc268 (
      {stage2_1[6]},
      {stage3_1[2]}
   );
   gpc1_1 gpc269 (
      {stage2_1[7]},
      {stage3_1[3]}
   );
   gpc1_1 gpc270 (
      {stage2_1[8]},
      {stage3_1[4]}
   );
   gpc1_1 gpc271 (
      {stage2_2[11]},
      {stage3_2[3]}
   );
   gpc1_1 gpc272 (
      {stage2_2[12]},
      {stage3_2[4]}
   );
   gpc1_1 gpc273 (
      {stage2_2[13]},
      {stage3_2[5]}
   );
   gpc1_1 gpc274 (
      {stage2_5[19]},
      {stage3_5[8]}
   );
   gpc1_1 gpc275 (
      {stage2_5[20]},
      {stage3_5[9]}
   );
   gpc1_1 gpc276 (
      {stage2_5[21]},
      {stage3_5[10]}
   );
   gpc1_1 gpc277 (
      {stage2_5[22]},
      {stage3_5[11]}
   );
   gpc1_1 gpc278 (
      {stage2_10[22]},
      {stage3_10[10]}
   );
   gpc1_1 gpc279 (
      {stage2_10[23]},
      {stage3_10[11]}
   );
   gpc1_1 gpc280 (
      {stage2_14[6]},
      {stage3_14[6]}
   );
   gpc1_1 gpc281 (
      {stage2_14[7]},
      {stage3_14[7]}
   );
   gpc1_1 gpc282 (
      {stage2_14[8]},
      {stage3_14[8]}
   );
   gpc1_1 gpc283 (
      {stage2_15[0]},
      {stage3_15[4]}
   );
   gpc1_1 gpc284 (
      {stage2_15[1]},
      {stage3_15[5]}
   );
   gpc1_1 gpc285 (
      {stage2_15[2]},
      {stage3_15[6]}
   );
   gpc1_1 gpc286 (
      {stage2_15[3]},
      {stage3_15[7]}
   );
   gpc606_5 gpc287 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], 1'b0},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc288 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[1]}
   );
   gpc606_5 gpc289 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[1],stage4_5[2]}
   );
   gpc606_5 gpc290 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[2],stage4_6[2],stage4_5[3]}
   );
   gpc615_5 gpc291 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[2],stage4_8[3]}
   );
   gpc615_5 gpc292 (
      {stage3_8[5], stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9]},
      {stage3_9[1]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[3],stage4_8[4]}
   );
   gpc606_5 gpc293 (
      {stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[4]}
   );
   gpc615_5 gpc294 (
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc295 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[2],stage4_12[4]}
   );
   gpc1163_5 gpc296 (
      {stage3_14[6], stage3_14[7], stage3_14[8]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage3_16[0]},
      {1'b0},
      {stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[2]}
   );
   gpc1_1 gpc297 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc298 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc299 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc300 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc301 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc302 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc303 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc304 (
      {stage3_2[0]},
      {stage4_2[1]}
   );
   gpc1_1 gpc305 (
      {stage3_2[1]},
      {stage4_2[2]}
   );
   gpc1_1 gpc306 (
      {stage3_2[2]},
      {stage4_2[3]}
   );
   gpc1_1 gpc307 (
      {stage3_2[3]},
      {stage4_2[4]}
   );
   gpc1_1 gpc308 (
      {stage3_2[4]},
      {stage4_2[5]}
   );
   gpc1_1 gpc309 (
      {stage3_2[5]},
      {stage4_2[6]}
   );
   gpc1_1 gpc310 (
      {stage3_4[6]},
      {stage4_4[2]}
   );
   gpc1_1 gpc311 (
      {stage3_4[7]},
      {stage4_4[3]}
   );
   gpc1_1 gpc312 (
      {stage3_4[8]},
      {stage4_4[4]}
   );
   gpc1_1 gpc313 (
      {stage3_6[6]},
      {stage4_6[3]}
   );
   gpc1_1 gpc314 (
      {stage3_6[7]},
      {stage4_6[4]}
   );
   gpc1_1 gpc315 (
      {stage3_6[8]},
      {stage4_6[5]}
   );
   gpc1_1 gpc316 (
      {stage3_8[10]},
      {stage4_8[5]}
   );
   gpc1_1 gpc317 (
      {stage3_12[7]},
      {stage4_12[5]}
   );
   gpc1_1 gpc318 (
      {stage3_15[6]},
      {stage4_15[3]}
   );
   gpc1_1 gpc319 (
      {stage3_15[7]},
      {stage4_15[4]}
   );
   gpc606_5 gpc320 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc2135_5 gpc321 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4]},
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[1]}
   );
   gpc615_5 gpc322 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[2]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc2135_5 gpc323 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[1]}
   );
   gpc1343_5 gpc324 (
      {stage4_11[1], stage4_11[2], stage4_11[3]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1]}
   );
   gpc1163_5 gpc325 (
      {stage4_14[1], stage4_14[2], 1'b0},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], 1'b0},
      {stage4_16[0]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[1]}
   );
   gpc1_1 gpc326 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc327 (
      {stage4_1[0]},
      {stage5_1[1]}
   );
   gpc1_1 gpc328 (
      {stage4_2[6]},
      {stage5_2[1]}
   );
   gpc1_1 gpc329 (
      {stage4_3[0]},
      {stage5_3[1]}
   );
   gpc1_1 gpc330 (
      {stage4_5[3]},
      {stage5_5[1]}
   );
   gpc1_1 gpc331 (
      {stage4_16[1]},
      {stage5_16[1]}
   );
   gpc1_1 gpc332 (
      {stage4_18[0]},
      {stage5_18[1]}
   );
endmodule

module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [18:0] srcsum;
    wire [18:0] dstsum;
    wire test;
    compressor_CLA128_12 compressor_CLA128_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf82cfeba6212a6b8b191891f71ec2e0a87fb6b9d9ed2093da4fbda34804cf92132311ff66bf17ea1a19900c36b2f704769486d66e22290d2d0066164bd673d9c2eb431a836b06e1ae5ce3be351b02621dadd1bdf943aa0100c2d77eb40999aa19237534fdad898b73c5811c7c7d3123c1fe434fa01758d88e7fae9cfbf5eb6974ac8342c65d33b44e59e0b8fb195ca2a1dd28e3b19ee27353962206c4ed220502c7532f7a4e62714e8194a85468f018e1e2f3e63922de53894e674a8fee66aab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h6fb3bf484d12297e2d2d417f887fb5fbfb630c873c10e6b78bb1656c51574fb08209fcf606d5ae5f8110e47d223107d6b460ee1d07f20285422ecb5a57b86ed50b69ef1bd48efa606959189ab5b555989da12af15522855c146f8abbdfd5799829a99a53298e739e3a35f51fda37465bd263ccd941db8036055f51c401c91d4e407c656466d9f96323a97acdcf3cb88dc60a0e1551430419570868d3555669c9ef23f26a886d26dc1edac40653368242368caad6168b41247b7dd44086d60ac3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h185592573b4292c29c0cfb2d2197c72061a38c4a8fb85ab1a3b662132a3d1973fc8828f345224bba815a6e163b3617363f5956e0252d905bb64155c59be815680f7a0d8fcb75c94b869701a6b4cb233b3ff178b73b93d6e217a8a75790744d7fcc26316150d996205d113cd6cc4ac52c61f74a1e8d5e8f9a9c70a50115d5947edf91130b8f47f9536449149f35f4caf742facb2d1c2268b06ad4007d8f10579ed948b8298447feb45958180ed1438d73dd0e2d8d91e6301621fe12cf45e78435;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hacf2b59b515cf745a70dc647ff08ea05b3b448f5095e1d09d619842efd1893510f241452acbe0e9d2145bfc6d976c2993f63478cad295464cf83082b515641aa7f7c8c418088d0aace55b2cbe7d536f43aab09d3767117835328880f7d3aefe7e2428b0daa032e7e71b5ab56c68bd39605352cdeefbc12a29865b200dbb2f302e8c5aaa2becdb70d77b5d5531748ee4454e91a7a49a5d8e384e701a7dad829a8f72347ead657728c356a26e6a3fdc648fc431a3cd7b7c2e016e81c093e883fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h23d447cd9e96db5c5b95bdd277a8a5470323dc50a56af01a009a54152fabf20bdca8b9f54d8f2e1c4a2a050b7606eab8d599a97fbc6c18608bad8ba2a19b6e0b9916a61a3375cbe87e10814bd3686ea7e199a36b10c142b6d98adfa362960489579fa377dea16a4b6d4a44671a6dbd1d94ab78a95354bda5d8fcbc3660c6b383ecd4b254885e70bdb50183188ee48319033113d7333310eac64ec0f20d3b333df952a2035dc50b4e83d199df57ba0147a494d3c500ffa9f3ccfaa0f43e7696b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h60994dd7bee2d2faa6fdfa38aac056050c5d4755fe6f83f22e53a3fea59b2d9cfd12cd5a7492f143a9dd52ce1f2bb608b56660117ecf7c0ad772eac3d20f3a34111b3cf3226fbd44fdaef9f9da4a9f3487a8482ccf26af291b6822c6f5563fa5e41da1243480996e2c42771724fb0b16ff32c7a45b94fae26f71a101e936b168a5b9c02b5f5cd684f872d2a9113690440cac2f5228940bca6b8a49b13021141afdc70ed611b69b0bb5eabd1377c5814d40bfe97bceb03aacfd28a62d6a42a09;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'haa7898813a07b1e8d1b3b72d7c9631af4871c1385ea2a8f2bb8193bb1a48851bf6d94eb72bd21bff634a459f0ae67cf29a923c45c625c35703414f3ab47274363f68a91b89fc7a54287c74edf95bc7c0288c8ec46cf84bf60a422294241b5a3a649554c69aa91f4541d188e662b7ccdee4d1c3a9d69f197ccb63894d90d88c09a1575d41554d3f2ed5aebeddfb74ac278094b6dbe8dce01fe512734d84e8167fbbae47abd422e787c834c71c3665433785925e6f7dace5bc5996b057f7ab37cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8e5b7ca9562f969083fa93a88a101feedfd6a7ffc958e455e1c925215f3b8e3e6c1d1b6a2b017b00e5414a4f75b4c9227fab7678a60bc3bcfe1bb953fe71c031340904b12a97ac13a482e6d22b7d0ab218c79048c53fc44816002ff85aed6d7d0a154f769bc22b920ab11f4999ded3054b7a0cda79d4afd2465bdc84800c8b8ce393e4726fa33dc50b36e3c37ecaed7986933d93fa6d7130bd66c31569fdc6ba0918b5d60ba9152b19d44e2c73e1a9cad1687d6d2b327bf0fd803a5736c4f668;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb1282906cbab98d904fbbe354fc49b1a6810936f55504f1dd95b6324cb1b3cfbbb8f18e9d746b635b9aa18bf8a942c25b82e5ffa60f0700b1fce1d538bc290b277715e5e21945f05b3ff7089f5196f95b8aed84de934dadd4aea097ba32efe25108f35f03854294707a7cdb63fa0929656b5d6a36573b49cb2a1bd8a9882d7daa0bd5b422edc39d80cfd5eb5f60214f5ac6b6b28c50188db3cbea817ed049fd788e50d53ab17bddb6c5e91020f7383d98e670b952baa9cc80bb6adc27ad8796f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7b4fe3074317c7b123be50b1fdfabb7717e2f4279948bbbdcc7f7acb372528e9bf683f346eb984d8e4ad2b252da0b69689bb8ea2982bbae2bccc7530fe88b1e2f71f4234c82e505e19b6ec258d6ed6da6a392c696372677dc37df8cbf1e23e47daeead589e8a7d59c7495e2c33951e9171d1bd041eb303ea6c2356d1afbab89dab0eb0d72b1d097ec874ff2f168287c6f68cac828394bcc2d25c69585b492bb0c856a7ab36b7b8db1007a8b9028485d05cca5189c0b70a5afca33be587db2b3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h62771f4af1052a5de57213a9ff4028918e5c55f496d7f3e2833576e71ac94b98c58c4e66005b792f8631063c1a1c6d6e1347d3eda2f69b932358ca3a87c795007f83d10885ebf021e1541c784e2432c1444db035e1b2b4e29cc3e2f2126f2d102f5647b2115eab976f82742102f95373a8c778d09a2c79618175436511d9aaa5841508f039378ba0d12c79aa431d86f09efadaa40a659072970a9c7fef82e1ee61bb900d52024eaf8c3b71c5eb455aa398e11c299276a5465292a9ef4abd17c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7857412c75fb0c11e17c60f81d17d87467708e01bca654fd3416eca1508ed2643e54567464072a5b1731cd0075ef713e91c7653d7d4f77eafeb6c1d31b7a05e54e078a9b20af37cff1bd9da392f92acf5f7d4a56fb5e674191f12c4674c483aef8c90f15103f9eaa181091b5095417ffd23ca04f5206ab745be31374441119d16fc7887b095beb2184d2be91d85240dcb3cae60338b2948fbd6b2f3689e7b7150f21282a7332beec6f5c3327c95303f6c216f8e2a2af074735913a78fc4fd318;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h9f2708eca43ecea554fe54a88b719d3317011283ec71e0e68990f984e74140d1b9c74e0deb51d449ca598b07b82e7fe7d95a30c5a008112644a547add2596062cc3fc8d0b6e45692fe59f4d44719657d865c508f72653d03b47f4536eabc24210505e09ae1a2b5f84e2d07794331076ec44f5553e69eedca7339c7d73ea73cc88cff8cc1b52fc5e1e4a9db239cc05307ff361485cc01ddf1cc44f5566ee44077a0f6b80e9e32b60f9888ac4f3ff45ee765dae779022802dfe046b1c17cf3f9e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc1f322438483ab0e757b77a60a2c284c2bf863eb9af53126379144af6a79660612819dfe50df0046b80601b02839e2d70139499061ee243564f90a31875b9764490fad1c45228a11a5b2cdbc3132f9cdc67124722c8232f6dcbbcd96c8cf9b772d27f01fd0a7369598fe9884eb035435d3d7fb5d1a7099718851332babe7a437604892db32f37467c12f13b3b314179989f615c9f7ed7aebff5a1712ece3212085ecf1590f74c580eb3d684b166a0132a4c56b60e6374d6debbb0434eb0bdc89;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hbc1c5af4ad73fa27557ca95bcbcf592ab210e50d0a94650735074ca5c259304d4631246e852dc5beaa2bf2970014942117fe9e1724d2c5e27fd2270ec0e57721f1c8091bccac2409e1eba26115c958af905721c0a9438de98ad438e9dbe0fd065cd09d5180ede3bfd3b79ba173364822e5b1c8f69d37fa3284baeb4250ff8c835cdfcea28e682e1d6d5422c1e00aa753d0cdcc6badae130993a6aabf5799c759de27f0b0c1e3ea831b6844bf7e6a7400e951f79c0723934b98c9bf185cf327c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf50b0d4fd4f7c4b13a214fd91e4e6cb3280ec57ed5e9d7d6c21c616da820885776b5081f9fa64c5ace1454d88962e4e97258bf60f01c04f372ceab6c121e51338047fcb9fb747b1b4ff79e981bacb3ecf48a9c1bb1a8a1ce71e33fdb69598cc4db64eec52c9b08a1b354af008d5455c04ff9e1a630682fd802237a89cb6fe5b3a956528e76724cce873da2eb581f6e7992ab2f786946da49bc4491a08e5ffa348bd7c45428d3e2cfc9c32d1296e50f3acd64de682f09097f59cd9a7c00ad8d92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8e20067d302e8fd2d0917ae3c6635c280e8de06eb36cc3c0688979e5110578e828b77295f0379f2a61aecde21818fbe31af27aade05150da708b4b8b79330a2b69c9875252ef451192f276e6e1dc8b0ba5fdaf3e98698a259ad030a2e71c1cc76aed86aa7feccd772c335ca0111b146f1cd2e558e1d699c372f23dcb049ea13f53a9e7f37e87705f660129634a2e03ee13ce6bba459bc7e78da1a8a6b7b16316077f644dea7a8c986d69545f70e377fc8c89bdd5bedad6c1e814af861995a3dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h955fe5587e3e33830fd969a2fd0979f1feec66db1233db8bd5108a1dc63b4584857818505d292aa7a36f52dbfc98ee65f32cc377a450980174b6dc08b2e24c4b98e37cc194b72ba7db8918a85abe54accb957b6d2d3e8bd6bef7dd2d5ec738d8bde168197f014418ef22c62e537fcc3c4bcccd5b85af555acee9bb25883c6df135d9adc2f7a336f3c2a1ed4484233b50ed6d822bd4fb470179d2c7b3797bb5e8848f0874c3e75fcb360c56d2791b6f5365ce27d9be199047cb17e8d25f4fa8c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb3b5687733aad566c4a7aaea3f029e53c2e66c1e5d874360a3ca03dd32dd2841f52266af7b676a7da303a90401c185afb2415e096f8827ae5e58ab35f39068fd2859bd36c06241cb3117e88048b83fdc8360b6d2d8eae44b3a91c9b828faf72a0738e24035fe2845ae62a3150851826e90ecf981bfed505911e66d40a99c6a7b7a9c686590c34cdd6ebf52b97abbf03c3df9327bc268f413b0459eb28139249f125f449585a954ab795989c39b3d12bd421183c70282d4a4a6edd265346a107e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hbdb902a8632ea8b83204dbb36809da5f34e15d4179596df3df133a526e46472fe489333d82266fef2740ec89b74da52735cf5daf9f0a84fa3a81cac23b7b15947e4c9e9259a3bfcb9caca8fbdca89a0c9fe54328c968c1b70a00e7f81125d179da9bd0cf33f28c8803969bef18247cb1ce6274a34833ddd81a81fe805adafb7f6f133aa478d41d192d40f37eff96fdb851c8573086121364a542b3e0e0f089208fae21f5653990cf3d078adcd4f9ebecce02a7505cd9cea50384c1591ff75842;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb627567d55cc8b9dbe4996879714eb3114220f055cd170a47c4f2a27b5f887af3c7d8fca246a0ab5d4f8897e475702550976665cf44cffc631a67cb218d0e43426ee48ea42bab3a156d77fb3ada92f3c31f090b85e92fa8f53face859d5594722dedddb959b31927033dd49d0441d8f37700a9d44c2eff65f7ab7f713da8d0bc85cf2b9c943e5a1209a27c351ec20ce5a14cd34b29feede2b585ae15408b13442c6524b5dd8d5d54a66e345cc33fa854ab102f2f3835108ece190959281577f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc1f3136d744d59f05697aa22124be3f7909d12bea3d3a07aa12cc87a14836aca0e2d07c830f036a5bab4ef8ff27ae658d3d5e70b47ba5f38ebbdc056e7a2db786ee76cb8395261f5b4389859e3176f514f1284bc6dd5cb026f197059180cbd382070ea7d77f67a192bd0b1ae0c5ef111208b7c523938b9543dbd1f02aa9655f802cc8094874b8e657148a99107d83af02972f6b7a798c922ccac0c1a2b9d5854c87ea6ec5d90d9c7e23b9204c08a86670a132376db2e82a6c81c46371bba3e4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h4da080db8757ab82b38ec7214e9850d8b73f4b8887dc3b84a4d335b0108ddebfbc1424e0afefe6cb4914229b5302c1cc1776064be2bcc1d4922351d84935e01758a934d5e811aee4b47006a26eba1d191fc36f5db7d240808bebfb72d732ff6deff828452d2dfc060937c9dec62e38e12ef430d99beaca4ec08736fedd7ce11d195676c27eb28290436b51263d9ee62944d8122ef38ed73fc747cc30c69486b682825f9e8cdd8ecb9c72bebe59e5592c96e218af0cea946ae7be42c836fbaa66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h9a68e1324f1c58c15c01f6e6cf819a28dc2b83518ebf2b22780a5ed97fe2c69a09f2be7a565dbc3cd4d2b814d252144723eb844209b5731d7eaaa81c1ad3edfa79f3e03197c8ddfa17f0c23e59928da2f322d8fa7f8068b1a0de65742d0817e2092a42cf0fb496b41be8a81d8c50dce73aab314e1a244c55409e53ffec42505bfbfe92853c559fa35995b4f7b4c4ea74c62565619aa4801cd3f8bff7970b8d6710aba7f76775abe61111e32fa891f7a64cce9aa537122c786641f92259986154;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h87987e86d744c183a99021f08eae06e39e23093834e2fd331ffbacd3013cfadfeff0c54918501e2f4a3b61d6cb9ceec07e8089d3942ff2bb20879416270be1a375f71be01a70e43ccb14611137166318047703b011d27b2a2e381f1a0be0a10f4c8e5514d4c4c06049b03304327cb8a893ea536bb72dd03debf5968520313024c8eab664a37309c8dfa2bac4faf2334b27cce08da63414d3b158d659444bee303c609a176e3416718fd72c2d842226bb750592ff53a7cdbe6fa2ecbc6ed8ccb5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb20210a7c953263d8c5abceea1c1cd9bbc5ebb223d076eafff7f8ad1e7f526e249ddc2e536c34afae11d0be6a3da6c761a15a09fe80b3b4f18a3db9abdfe265f5617a7a2f0beefff0245e67a56bc428cfd394744e2d404912ea5d9ff71928f8be8af571819b704426d5782a8a0d23465b769c61e4bc72be9792e6bc54a3e0a2562eea91be1fb4d930ace71e0874a488ee6672459d2c77ffb0f0e87abe49abaf09ccf27f3f61ffc21a37e0ff9bd8a31646ec95c362ecccb5174bf724c9aab2271;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb249308a0f5af311754511593aaec140dc72531d89692c9ac27db77aa64e71f5771544ced33b9170a1585d3c154df7e41ace32bffa6776c2bf49c34c736f5aa91fbc2aee7a1d766067653814506a99ce8f3c0b6db76c29d78c8a5c273dfbe4f0aa3465d1636a5738c3751337eec189c5430afa91b81b4ecb86a06da75dd73a17b20b2c1a5de2253483040122d5835807e879479854200570b40102fb2f03a0f9f9639e5803370e511b5fc1c8ee147786ce70a3f884dbd6de77905d93998e8ebb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8933b4be62b9b2790fab34add51de1830cec4e908386292c644d085245e5837d50c5090d33460beff1775eb249a2f7ef1d81cac614c332860b1023aaedcc91c8e134c711c5b5440fa489879e497b654043b1e276bf65c44ef795effcf708c31a4bd252d8795465558b107aeb35270e36bf770a2188202d4956fc00ad173a56901cb5166e73c005e988d60fd0e20c63994ce2f87d8400bac7697798b1e6e7d460c01ba45283aa4a097fda40aa5badbdd066fb73597501419ff98c06f2f4e8c219;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hfbc7df2a443a73c533d0aadffdfeffaf55e82656038686ba2e5d6678bfd917a1b704b709556b6c92eebaecaed59b9292f4cfb283a552e679093d554416ce8c68863e82963a52bd0e303d6d033e51ed149a8083d61ac88a46cdaf9343ab6b81ba171b1e9ae68a0a8098032594876bd9817813a6476571a859ea994ac02cbb05e8ed85919e03e109fd69ce723130ec2e2baa1d3af71afef4fd69a321b5f3d500541d96a4554452f3a21d8dc9bc06d2bb606714570d83dd7828d01826713c7219e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hce39a266f41426fa52a23998a865ab1b3da29a2ad7ee094bc01810b0624518068efeb072812904c376c72bf94afe03fa5de694c09c1405f2ddc2e6e904591c0bf3a0ebfb07e39544a84cab2ce6d5a2d8cc1fbbd6d29de35f07558a85ab8c1b48bf922a43f3eb19572b0658d60be875c47a942ff54f37ddaa7eb5b675b10afb6a922928f9a55dd95af86a834bbdfbe3586d086c35304c820acb6293b491df54aa21d72fe1caa096fdd9f205133e40e32e9ce34d5681e04adc7fd2aac8833d937f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc9e010c0e5c01605127ea5b3e2547cfc2d501d675d4592b93471768ced5bedd6ecd5821d06dbd06a12a9910b89f988196d39027a1418165a1503a0b5d3bbcaaf10b0429b00ecc3d9a54e72ededfec03bf61cc07368b8c1151c3cf406b5028e94366d33d0cc1505376b3a0b088b33f138e9ef1ab8b38501ee04d658724aad3ca4bec41cbd5bdaa10648d0582fd6584555be57e7d3759e864095ba7bcec96253dd1a525fb432779351b27bf589fcb502b3e3c2240f02b2ccb5e91699687da7974c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5123f591c5799b19d6a579fcd02f95ec8121010744e73801115caadf01fb4345b6a150ea171f4435b9b385725ff8f4c0d00d2d18ef493607289908b8826474163154baf2adb7d0906065cbef781d78399ed5ca1b915a3ea781c1ef3dccec8935da1e8e7220e0e1bc06bbba532689cb012b1d19d0159c6052181aa3785653f6fd407fb0fecbefe80122aee4357b1938e8080f675037b604ad29612f35d589e83a30941d726d57fb0544675e5693ec626f482075b6324c4f69736c166bdac97b4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h382d5bf6d91cb5874f2384ab4396f1293d339a4dc75c0ae0d0d3bd883b6913a2c12843f252431dff95665e845ee9f7cf15d6b4e0b86bca35b2284d2a67bc8b1135a97d5e8a87ffb2111dfdef1a832f1d46a2b607a74b8c2bbbda8d39767bb128e5d4a9328e8081868229077b2c073980958c178789ac2bd7f1e34c465b683836b4d479ba90f53adfeeca3839cea3c80428f9dbc19199c39448fb449a8ac46287cdd028e0de94db3630506263f9be0062eacef6006e777d0c11e53d442bf4743a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5638a308b1370b97e5ec3c53734dfbb60dfc2e7bacd7ec22541dc70459833856b04e8704e09add70048efd87d767c9c7aaf150afed914adc47a1d9b5ab9b243a24c2da4ab930e3f06d6041db95a31f663a09c136f76ea443fd0f7e75a3675b1638dc8e744c746c997caf275380670b40780e2ad8d3b45f69b206f076326a9ae7fb05e069f06d42a73c33f14ad66cec2e0b8399efa17b13ac95955b81d186b67d8e7fcb032b20d6735ac5a72c5d5ba70fb8d7e79d65eea07d7b14246074daacf0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h63a78a410d9986429721f240d4e0cec50a465b91c2513e416b2105c219892a684c64ea726f5eacf056fc97cae82f993d9237d8989547bfdd95e713f52e3d7a156f932c4764b4073d8db8a0eba8f0b3c87cf4288e7b8ffee5d3748b923a48645269d8ed16abd17e97de16da6a97cdede0adf2392d79d7eb31afbcad59ab83226453228bfa172bea8505effa3a69d8cb093f38bf70e6d67e8cc160b5e9e2600efd1bc54283aafdbd412b742ecdb3dd81ea778e4cdea9e20e1e90a0aea27e5135e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hcf60c17c545728d36ffa8c4ee0b39f5c0d4d019c5baf5f442a7cb40965c1a9dcad58d29c1a5187660d6eeb247d0e0f3e4a9acaefb14269988134bbfba5900623e949b4bec46c95898b291922dbe335d7001d6f844cd2efb362564e0a14ada54a040ef541f76113a3aca3d7c3b6dfd283f3af0e016349a13aaeec65c96be11ce6ba7bb560164bbc2a63aa605aeb6257c0406cf1b663097a131e455c61f5f3e505ea119c9cbeaaaa2a9ada590f2382dd266484a590d84778bf4e110c48becd9b8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5066dcdc8b2829c0a1337bebff06d9675c185069dc5f9a31dc3a2cec3c6ead4c9a09adc4216d5b4db46c034a75b2d8cee618a366809cfed337d47ea78d512bd43a6dc0236d38927f0e45501559c6dd47d70e15dee18e76e38f2672870fe09c2a9ab72b2f05c55e309a5a714b321e46622821e6cb9ca731abfba4c1065ea98651f015caaa15cb25759295a97d60a9dbfac23d7c0b0a5acf8839d40e1a5cbe8ab00a57d0b6326149b6e1125fbe9b9c043ceb31e4e6029d8bd37ced1c025dabf806;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf0efd5b60625094565c416cc4b2db6840fa71696bf3238ab7efbcf4c47652a5ec80b64eda6b323039bee6a606001a56e659fac301f5d38ea69ef25b1eff40594fc55f0f9b05047f048cd05447c31388c757425e222cc8feccad616d1a6d93ecee8c40ebb3b4e596aaa0aad7865c375c81cb59b548a8e91b8430b0c52a1b28fad77e0daf2e91d9a9d82b618351c58b73523cf536288ef367f2369328e2602b897575f9b1b85845605d2232f092350e575b90b621e1e6b796af0e8339df3abf925;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h74c146487ea3d96a15801835a793dc179682fee2bb3fe5233bd027485258fcd04d1f23fb8ab329b253e80b514cb06c1aa791b282694af64d7a506a9b4a0b7d83bde05a9f586bfa784a2a8126ab31c4717a47c19ac23ea719c5b9460a2c6cb09d90f3600a2db1704c702c46bebc6af9867a99dc619d4dd1aa8b00af8b37374c50e17001acd3922d7156ff131f190bef0e45602f9604763ea04a6b913ef39f8c36e4ae5c62b663ed52279ae5f7aa28323f9816c6154b4aeb759e743d8feebffc7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h917b2173e7abaf3305dc7b40604917989e091c80ff7dced8d5d15faa9e2cf856edf298a5edee83c160713f73a86869775c1d1b7ff0f9124489900dbc33bd3e7ca8f6563bafc8868f258ba465c4bc1729307019626d4f25fd2a8e275a039be283b39992f09a5469218941fcf318e4df58f727fb726159089ab2ced1f98acff08e408ff4a844c2f6f6ee3cd20435f7d6cf95e885cbf5fafe53e74bc619a7a0aee2c5711137bdfd48ffec08a02472458eb85d54efce27862d4e7d9e2e57cbc01502;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hfa9bb8fdd0d25f79a2c9bc588c579dff3236f8a047e04e6e61b6bbfddc9945b59b137bbf0221d7d9cf985981091dd89d39e4cabb98bf336f2a4083de1de9ec7482558362625c6e2fd6d082f86a4eb48b135a2be6dabc02b5ef37fc37b53aa856e33e4b83113f6b6243f05379b4b9a5efbfc78c39e4ae5d3f60d137ce713148f11458e290c22834dd22fddc10238eda270ef6855793b3c1483e95565ba8a73c3ab81eb0f1c6433742bdd7d7ccf6240b1653e123f3610ea9999aa534a4e6384db4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h89257dc1956e9d31fdd2e0a1722b4b0ab141538da975e1a353eedd4d88712d8a2978eed6a149b84a1261f69a2ccd5319d6fe4832437432c2903057262515b372c1afcf18c7770afc88129c0bf7a3b36fa4353a3850bcffb295e0d5053b8a3eaeb63faa2f6529d942aaaa30c541c01b4ae611a4712d7b045e62954d8623ca3c114c2d0140157172fb465654a316e693d80597fb0961ec0295726a54c4c04a3cc6cf9842f7efeb1827c2270aae7eb71cd6034921da654b0394643542201100f04c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hae1e0db636e006e13798ac992d6edb456d4ecca274da4cd084e93317cf4619b36938c277aecd321483147d8964e41f66f176fc9e04c7c8fcbed2aa73fc40a68f343727ba8dd9686bb2c2451d49ac1698a8914a5f58505a5263c6f2cff72bfe9ea5923fc0c1de73b1bc4657825a499727e433a425af856188d334eba4b83ade353d4d2009324ddab3c37fce8949f64e8305d5575cb02dda24183be58974e7b1669cc9f0b53284fb443df48c03bb911fbbb35549e49c965b06c7c7211a1c2f91a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h74586ddb8004307f91056e105bd546f7b6a6e80df541d049b4471fdb0c5cbfa522666364292a1cda7d4c6724b5fe60b363fdb9395202fd3f978c480d3a3f182a853c69a8413de458fa867f6f1ad10f36b3450c0c061f97d51206b9ea5efba9c92f6fd9e0a9e4e7dae5b36da326907fd5540baf9dfabe99e1367c31e7387199aad67117b7558bba95b68e41ad542bb421a81bcbcc975305e825a701917452308c636e416ceb60dbac97dfd58838d07701defee20898e72df242b2516c0287fb00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h2adbc9106816b17f0ad7a59435f1ce57269bab88d9f37f43368dfe5f4e5fca35dd48fb9e149a241ce242c2734094b4c23d44191db95f765dc0b3a9b51bcc5005f30486ca348b75ba6ef49bc6b1e5df69c701a6f71b600021c6c833ed4aa2436a577ca498af1fbfbef203d5022a9b96cbf32aa55c5a6a9b30af0eea884793db102624768eb1fad34c6a1796bd7bb5b6e20c9433e759de4c232564b3c4bbdd092a38af6f5fff9273cd7bbafc05dafc86992893a868754cfdb315f0ad3cd7068673;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h188e97a056d0d13b572ef4f623d4e3ebccde1f3bedd4817d468e36a2a78b8ad05ec9e3d1c4c0c6fa389d9ac72e6e7a83535cab6b7e8c56c0eb1ff42265df7104bf6697d62cc1f6d3688962a792dbad8bd7152a32054bbeb7994c3312f0ff74b2b326f474f569d91e7df93bf68718bceb8bba3975374cdd96bd5db112094615592abad003532810ec1cd6cda406f69634e6f8e785712208f1df7118c3458d18a2c3f46a07c4344ec3902819ac547161d919267ca3e35a8af97a9c56bd2816af28;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h27b0fcd90423c63aeb2691d4dc3b4dda0a0efd9db63a2a62ee69288034fecc3a627ed8922bac14a6da18b8b5927f6040bcb950c6206930db5f41fc23cbac2a1f766a55bcedce4e8120648ea4896f13be0083ef3f1e5bd22ab06e9a483f76f8dc9d67a1a2c57c61e709923a4170e7867a124ad11c5e6cd53068299e34aa41ab55258d19253e1e6fd521df72fb3e0ce348b05a6d6f6773bc9944391a11411bfc5f5d3c46fe5f5956f32a707ccf448daebff8088b01cb71db14fc5734d934cdde0b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h27fa571d49460bd23675713285678d7b3816fb89a0abf12b929e5fca74d36bf741d009c965363f2d1a0ce556cb1faa42b649b1ca893cabbbb4d3cc00a9d020c3735ee13ae123ed71f47cdc01444e0ff5604eed8eec45f73386c9c22b211394e86bdb3a9b2941666a79d6d9979830da2290df40d957ae840b62e60763f20c2fbe9aa594843a4744c0d09bb4edd2d188b5cff5e71a101013babc138460d696ffe465fa243e2c854ce481ed8990b1f938c9621886f4815bf5f8e45aad77c3089c4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h3547338c9cd4ef64f89a1f26ab5f4bb3760eac4a2e150b1a612f06f5e90194c06d7904f01e6c02b7c2ef91e633903e7f917e31c9a280810e60997c6af88764379221be71627d9f06800dc38a32adfb1852218d77cf7d3023ec1997c7b264ad182cbfcd87a33c8419fb6dd2008e84dc5304300cd39d32168502252085e18d348d6758a1e6bd1b995c656d7a8e78213cc0b76443031ce6e062d1b795554d9f2e89250ccdd5281823cdcf24d14c9442f13f23806e66acf12a6a11852a630bc896d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he2d993224c656f4455cbad291c1dba3deea531db0151c537eebf2888cd5c06e45e9bb14ddcb6369f38986121e7a073c8fd3c0dc46f4e103851761d0a152b9d86206554a448e130f1da1e7f62608e5ca40435db2bb84e1f2855122239758bcf06ef576781f7efe2fd3ffef1d5e632439dd98ffecdc5a1f45d889e16f16e0e3446b73ba4b1ec954d051824fc960005538a41ca8b8c2f82b00000dd41fd6a5fe0de37055c1c80a49b53a27794b47fce2aab81dcccbe108466c2f98eebd2fa7ba4ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hda7b1d6c53609127548eefcce05a432d524aee8cf30c480a0f84d7d3917f5a8d9d31976a932a87167b0fa36dee5cfc6643d4174c2a6792bb08567088f7848a1447d6a1f400b4761dec89695e1dec30887b786c6e6aca60e92aa20cbb4d2dc0f7b3e61872faa0d4e6d055f2d9f98443932778f49b44613b2f15ae18613d470873dd02187f6baf18156fa258bdec948406bdc72ab156a43409f0f6707507ed4edfbb8cbefc5ca0a6406b05cf99c650f97705a540b76856c099dc01682882e5b065;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hbfa8d52df353a3f0f83aecb01cd62d30df713fc7a3063960cf8f038e515fffbd706ea590a3b42a499399f283d0227fb028216bfb22096ffa6afce17b19489686ea7ec06aef04ca719eb72dd52b11ced8e9ad42eff7b536784805dfbfc24b082057c89c94267314a57ffae7d78d6df64df40ce68dea5d92cd071d349f5f02c98f7f6ccc72dd5e24985429d208f0cdbfba018d1a8faab823ca0fe448c9ca68c983c7903f27cd2cece63b42a76067b7837366ac2810f905d7171d0755e490564e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h2a54d410b86bab556d36428f29d68fa91d73373ff36a11344bc00eb225e5dfced10cf860b4d96edd1a1e581ab27eaf2459d3a4b7f3620d3809fa307a124aec642836145d248a685b047d8617de52bfe9eeeb344eec57aef5e7a71a763b98ed23dd3261a465b1c25f7c4cafc025207435be6435d9ef016eb92f0b19a85985fed3c8b96416c59e2373836f9302e373a339467276525414c88d62d2f1213eba00fcec60a56e9920aaba83942e15fb5e57a01ee42d3d516b6afc31c2a5d08fcc12fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc3b5ef0ebfea8b22af639455b286a95c409e6550a35ef79f5f6ccae76b6c4de2c2c04353ba40b0c0001f15fae71105e9b631b995dd43879af78f26c6ec60cc9fc9403efcb09abdc423cc21caaf7596322b5bd19d7068bfa6a0b5fcd72874d82141556becd028d0e23590fc8741028613c68b44184fad9edea9656732bfee8c6efcb4fef2002f06a3a3b2d80852d39ab9de04779b2fbc46d6b9f5e12eaeb24b33e4fe86ea6518e95398b622a8c6ded5548f22b288b0e2e69f60545da8f11a5783;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hfbeb5248afb6f568cd59914b3f333873dcdc53517d91c1a5c60d88e6a361f208482516e36c058b2b2ba656c0775bdd34c4b37712df369a6d073a7f0f36c7e64cd90d26a577f1ace68d86856bc5dd9e1c3d80303b8918f93a9b8ac712b1fdf036099ca972d34808942a555c63b100ab3afc1788df3eb18aad2588c3e1682c1cf3e2abbe9047476b5789a62961edb686b06d6f6ed3a65ef07dc367f0e13be32af6978cd41aa13489f1d53ab90d6041aeb1a9ce01ecf6dc5e927c3a7f11febc0360;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h700ba1503d57b48af1b2c6dd3fb9af75b03f90c9d4db46ac00427eed36112d0c723e08166531a3a6cc53b936742d4b104f11f21af3eccc29bf5a1de402dc1c9286aac0c6b12a1231871fae796a2f98f314a0cb82974de66e9945ef109cc4045ae043593bf79af58f96569be3af3466c7e685168cabbed89512410edf2f156b629dff6e404c6b15386a6b768e308b7cebae5c36bc2c81b85b5e5c95f6d93deb8cb2e45edefe7c51611e45fefaa824a6444970754358199d649e59c813795f4c88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd4533a38433ae1775b1285c7fdb962637cd74d99b6115e43fe4ab4cf85270dd1fb89a1d74fde81eeb7d3dcb5c9274de38751135eda3b922afa56ceb2c8872131bc1e83e0acdc7f34082f780453d629a5c00491d336e760a4707f81691420fab67e4231c1b7f3aad7960524dbde8d1d2c44d19154beee68d5ade28327516a736078c92f2b1b065e89edd6a1747fa3619d59fef8086524cd0f7815da9a2a4f2b949693824dad8557ec17088bd6edf02dffabd59bef476a8c1e109fb56d59944557;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5c930f3024b6a792c9bba44ee2e76f34fab15b0694e56166e5cd01d2bf1e60e338677a59477e617d469966ae0c2b34fdca59c6c9538dc81236919d079e320cfa46c326cb32e9173b955b32e73f0890982e394a174255aac8b8885ff89f11490ae452a82cb9538e18a0db87ea638db2047b828da92da6b584be8cbfa1a33a8fb79a02f42c884fe32c77c42db0d0ed7d98e2aaf2570c0accf338c14c6ab2af0cf5d1ee1eaa09214010396710515a27002bdec4989c6a67de04022939e89b9b38f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hafa406e8b3cad1f455a8c2862232281c92159c52bc115de03a7d96bb2ae11f6f79f5382f0cf48d7ec69a091fa7a63267812fc8cceaaeeea5d05187218a46eee4e203d77c60216e691714748e8887af0e165e29a0d8a9e93f939f1bf85149dba61e7a800fe7a94cd2b3092cc42059c8baf414e49f2320587e5e19dd5a8e863b64e40079b10f86fbfd9e7a0d05318c1a2ed9e0b857e1b684d3fdb87bdcdf0cccaf419e406039df0c6f141765b5e1c4c670d28214d87da6651d1cb1aa6b87c0b337;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h4dc338ba195662692b56b815d2795825a920098a491096c1f388085f644a5ea2d324705d68a7528e72757216ae9ff1c0006d4ff172acefdbfc80d524a4f21647697fb3c995db0912f4f87f5268d5bc7b8b628daae0d303b26c5671d2018e014f838079777b0c6d102e5514ca02683ac7b8982c7a14cc5460a85621089fc8b19637b03e52a6b3cb9b09520430d96638585b1752d40eab2e9c0478bbc6620274d46c590d136fa347333be96458c49ec18a791a5960921a3254557d4de13548b7db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h394816012b85b7d0accbf9fd25e4ca0f2c34abe1cfdaad7e316014c32e95f191b002fc4d5b6a1888797bcd841e68c9f153d353ecdd5c05406dfcb8c322dc72bd8d213e37008ddb42c4b18e1f0bd7c057df29c3b833806bacf99a32c9fc1f16cbc2df7f2dd57297dddd4e2a04e18d5ec55fc6cb9a1558f192592304d0f6ac0c9d84363fad78b7556f61dbbfa6f708777d379d7f18a017147d09cadfd9cb2272e0ed0f246dc7ab54be6e449f146648c770f66e36a16cbc1a402413e5b18d180ded;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h58852c5a5e0b788ba71dee31d98af6ea6b399b3fb00a893fbaeba881b959b9fa87a9ce879fc5127a5457c568bfcd9d8a135c7b095dff02949a7f55d6fb717c2620a639a1f608491ebcce9175d90f31c341506f4f8bf145864f194b09d1e3061189639b21ccd48c08390eeb09f1563538b8cf798511e8eeb0f3943e9d93b3e272420f4808af91edfb52b360c534f835618e5780ef2d1bca65a60e718895cf3a4795003424d5a1758f283b76b4060c9561076aff435ab0fcfb65dbbf2056b0f273;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc2685ceed76faffc5d079ab35fa81e19cfb09e49cb3131267a9313ce76dbdc1c04dc15a245d7e04c1f3e727a2ef307358eeb8e77f9f87ac4519e14e35050faa243cddc2f12e12ccfb8b666cf025ee2522140450e911236ee7aa886c2949a9ebdc16af49b588a01d8adb1c882c1d4987f7a6c1cc064e8eb4334b73677695c63f289fde32f92b6c7cc38a372e6006161070a86b6a5ea2aa5b3be9362cd98102597068283aa40c49bf675380cadcdad555d51ae81742a4a7d5d8250f587a6fa04f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb138fdf82fca1da352f712a4312441f3ac5ab56ec983c49cbe5302bab9b0c87ff86ae5221d4158360411abb3c7af85793371c09638c40cf14ab8caea1d746b7fc0ae76aafb79e299dc8de272360dc7f03a1fad8f2e2ba1049d3c64ef5daa62dc4bcb072b0a175b95e85306c0273e25a337c75a05a2ae2eb818d39d954ffd8786581233ee543fda7b1bfab5db8f7b96715cccdc2fb7a53dbcbc75a6ba79f8715bad0a119ade09b92abbd454676af1b7733894b74a108d53bc4904ecda3519b524;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h11a2ba9c3346c0a38ad4b262bb4e2b06b028bba1643b29d942b17a38861860d8c23f7251317e98d134c88379f7a7385cfb93f77be7c7d75e642179165cabde320a7b10f9a25703a8af60b7a7d51065ea4764b1b8a33dee17f2d232478a79349506d4139a25ad9a4ed149094222601842e8cd2b39f3dca48ca56582d17b4838c9fda7a6aa0a57f95ecac72d935558e0ae2ea6e640ec0f6e942b8fe9f4a20b63eefcccac2c36fe045a28c5dc797d611e50f38822bee5dfeae6f96e980785858367;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha5b5523b9c06b975fb3b82655dd57fc02d594f06975d324185596146c14df0e539afeb4781c7169508d279efd4f7e8ccd9cf1656b4471e13c1d43ba978076f4c17647eab87cea5cc2ac769d9d758381e61cb01908e2b91a26e8cc96ff7662ee220c7fedfc02b379be695e2df9a98f0eed43e802b3eba9e555e5e5d2745a69853c5082317df2d1719f5e51529dc6322483909df84c9b5564f1e529b1f62851e6470c5f3fe4b88b0832d84230d614d9cd6379fa688896270e70c7b945a42226fae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf57efe1e966d5111306c8bb10b963064a52be48bc18b13b7eae895c2b66311330b73f5c059e62c6de44d955a5c9e8d771d63720e542bea2ee632b041bfb535420b7b65efc3dd43af12e2c9ec0b7c41b519eac57176ae5a73fd7bf3c6ad147f113b2fe6b059909c300cb1f8de3cef3bda960c3bee70bc268e62f75e0966434d6909e54711fec4fcc42bc9a2e1a40a7f8fbe9d00b99f39a20e2f397a0764eb4528c6f9f39ddc8f8bc3548f08b7a77da05dcf58df6c0449e51541f36b9082458ac5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha9677d4e0471eef107edc2ff651b9465b86ab7277c0c6741596b2e8f5f053f22a4cbe542221dc80e952da682129b373fe1a47f4bc965a8cde3c1e63f56e5fd519cad70196651622db27f85324a65697bfa5d8477d9527c202088d67517ad8c55ac7f5f1f79e35fd842d32e93bcadbc4661fa1fe268dfbec179e583a2efa852a73f1b17d86d9c274dbd70d3ae62a5fe6ead8b33804d8b292983aa1c4938fc1bae98c53387bb23f37c948c52b22eb57b8d1f871c05a18b615fdc04e3aca7640865;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc3184bf58590603009202cc80f5897a34462f22b1f347c49880529c7605bcc054a5b6545bc91aaf866e6517828c276ca73e3c5799eecc554f180a59c445e5632665e4c26dd3818956fd4f7350c350a9edc4d185f5497aa2455998257a70ff55dcbe66776524477f11de7d356f828618a5e364e92c6c506c4c83e5ff2f06fec8f39d557a56b083768401edb22a9a15e7dd86f3af3abe0434e3162d60180dae058b5a2dd95a85e194087529cf7736c6655411eea87712a3c4c8ebe047fece40a1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha5278066125ee54053de80f75df6997b92035a19d54609118c714176278dee61f61ae32c8a08a9bcf8172edb358e3ea4c704729f4b44c8d878cdca187f528e6f907ee72b6c4a2ba37bc2d18eec87e6575bdabd431d5c203a3979980d1f626894a111dfd10ce9177f7e64f0894dad0037113ededf0acf69763f304beb2b21b6f8c82ed4a8e69b5f05e333488762cbb5874c1754ceb31e6899bbe38b5854d9ca377a6ee3715ed2f9a8b186cea1e10963ba3fbe6112b1c27d434e0c07b10b919a8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h9d14b2aef6437dfa756e7c69bfb5dfdad8cd126e0f024a90a92aa9b2db5998a89e3595a405e66fc3c11cad188c134777e2b86ea1cad74ee65ce6b3a4e3f05e89564719c35a316b0d8fe25c868b8dec6468ba9509fc7428cf181c47e971f02c00699928734faaa5fd3f99ca3fa81d2cd83cae9fbcc0a297fd75a49b406e4771452f1c3153a996f91b30938dac6f0c0a3d445b069c46c8b73e37f4d8f22a08c913d394565f2a24114767b972294335d1fb0f0380376efc7a45c0a509144eaa0963;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h62848e6bb68454ff8350655df867782f42c9ef3c185c239390f6a2df4e79054711e143314c93c6aec665ecc1d41926e194154e732dc15048d7013efcc9652413feb1b4f6d341f1a20480e1311c1230e6893364231e01e2de9df1163bb8a58beb3d9c88922fe406969867f5c67f5bdebd09151c7c7eb002d368901cc85a0834b669e8f7f102a0c418e45b51630ab07715986bcba1ca29040b87af13b47c9c43f9d34b57a3474bca7887ca1f0e1d091bd109a5eca5a661a4e140082bef625e6bf5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hbb94f4ee9dbec89e85f540c8a6e47898a86bd77abe14a7b1287bf1455ea707050c97bf84928130cb06ae6d7711014e304a4a416b7dad1d229768c74b2ec50f58a4551687f53e754a76488b6cd6b3f86d1b11f7bcc1e4b5618fa04613d76c174c97ab04bed52f54afbbb4e88269de8a5a285122c4ac673aaf7d5cf9ab98f477f96bb618c6f28e8e48e6c55d93b93451e97b6d7a1cdbe953b87f81b010b30c4e8acfbea889e9b436fcd3281b9315a516cabaa68bfd8ce5122b4220c977b25b2666;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb22a055f23baa94fb922506929b02c9ca2d3cf2fd55a7eca9542afe8acf9c11eb1ac66fe6d7fd459ae9001d8c3c941e5bf54901c895cdccf98d88c9579173a7b73310d66bee792192acc8626fecbf1e70571b1f409dc910cb809ec40e3702dfdef765f156f9bf5e1c3fea842dc81154daa48aa519dee9bec282c1edca0987a819576ef7c1dd3efdf158538ffa6f4961b434966f5b8b16c26dae4ae842e70b7290f6c15036da9dd80cf65e03b4fc8d18808a20d607eb5e529f776bbc1a3364840;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h710c38796ebf0a14a25ebfce3551444615569c05de1aef008476fe07063d37bd4eec6f3dde551ff03c9d5d0416d82916b554b1f6730d12cdff0a362c16b510ab5327616c9afd65e06a3f4031e5f90823b773a150f84880ca2a76cb1dd06b0b76069f7d55a94b2c46497e73e53efcd39f7274536600c174b39f904317cdb2bd15e6520587264a97edb399cac9bfc3299c5505c6a117556e24d9997fe0ab82078ab527fe7e8d1e4d2f82aaa6d09751b0f5f79181006f91d811b1bf1dc3ecd636c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5d500b5825f5f03c16361a247a464a4bf67bb4d5a6c938d56e2286e67efe2f584e5a12e33c2518b60802514cc8d20b3522cccf638e1b28da34f672a0360334309d332b6ee04cc868b1e067cdcdd95b865b158940ffa197dc2f364c2809c8f90741b86441d8d95b22d600495f226e5d82511ef13be55fa4d677eabd542318a3b2914a96d9900ca3251b6338b8aa7167af193f3945d7d458bc26b330c66a0b8914b9ff6da9db8fec2d69c82a10ba2c11413b4701fdfbc1e939b463e24ffe6d610a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h3217270fae8ca7d6becb1c21ae2a91988a7a4b948e5aac49612ebcbfbcbcddc4929a223d4d35d30fff65a812fa9eb63a3583192a0aceea143d9bf03f320b7bcb6803653bf772d2b563fa8041b58115e15776a0822159912421deca4e1b56dd14c58a5bf825d02f9a5cadaa6680fab0e0fe7ba23637dbec6b3794fb49ff347f28dbbecda0e553653241dff11c3dc5797354c8e365ec3b0ef24455ad427fe0d62a9bae01c25f839e1f70ecb23fa46061b2e62e6f4dce73c165a3a4bd41014d555e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h56da0d124a64b3858bdb464f3b05bf7a51f707255e050498db4b18b3da204dadb03a5935ef6960621ff5d094c711508740eaa211724a375b703e1627bea08492c5ef93bff471d9cd2a26b149049d6690e658cc9d3301e094f5348318bb29f9ec007f82dd539d81348d975a28edba21c642e90d12c331969174c5c2ac78bb35b51e42e2e2765f201564b2a1a55a2d197bf7a6d0b907beb7308f5bb366ccb74302bfe04e1eb0406a329d12aa16ae639c185fe0e59a5466a6753aeb2fae45cd1cda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h92742fdfd69f6c693871fb7ce6f00c9b5f617f634606e61ff9b52f43cc8b3b227ee4213446b3ce411e959116a28de91f7b4ce974d4b11fae82a14a36f20603b4b8b5eff5d819af847c30b30aeec2e08bb5d2a8fd254c63ca9c9a1166841d45d9922e21dc5b4d9193cd39b4a9c1facef5fdc72886a7976a7bfe40978927260078cee69d18f7483af073585f16b318a205c4633b5a757decec47ea9bb815e935f5b3a35b7855dd4e2fee789d19ad486b9113d92477b3cef260dae035d69fb99337;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h6427fd03694aa435fc962b884e09b54aeb5497af954d31bd69398a3b30db5d8c8e271694f2e73b948550f01e86a571cc40a50a723030863938b1eee02dcaf3266ab1e6f1a77165492523b22ae775657d07a8f6f6c185ae048bce8fa50743de2325dbaf7792ac4ffc50d0cacf231f40d8526bc5917d272832972170b176ae3d3e55d808d44f0119ba08952054330a83d0eb10fd4f9cbb9fa95b53e0522c1e08b159eee73245a37cb24c2a2aae4a05793f9475e7df7d7d1f651cafda1dcb699b64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h21776c205806a28be3a129c024b891b06135abb98b320dd80d84ff012d991dc13acc64c6318ee258002449ab9f2f3aee2093f0dd2671ac72a14b4abc7a2f42a7dd740f8ede47bd684689618579c008b051b1170e28d7dfc084394858f65d7e938184f6fba1b72d62f0e70d4c6891ffa8ca492b6c007175be89924e19856a78b3d584bdf7706b12cf4e585a7e285612276011f1f83c91de9e84eeb7fb8156374d716a879b12da3935a6daefb0d750e7c23e17a4d09880a7e009788437eae9413;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he129be099c3ad7385a9e7a73e96fe424a7b29bb061e20c8280bc330a8be06ff35dc38933041df51a80d819f3759283f7088347233756e9c5d89ea476e51a0a7b39e92466818359ff46fd2efccc3cf9e73bc3146740692c250d7ae20228cb8c99019e3bd37d3fa583936204939f060e4420f77c3b05ec824930743af91ac7683d61605018a2af6a59463cc1ca123fd03de7bedb4e4b7793a40b4ec5c4a9919cdde1d80808561d25b5c1d456e8ca9624f3a1be0a96626dcf00fcb5a61b1ac29ad7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h9afaf34729e7f894915ca4bbbc448db04f35d8025e5fcaae18afacb4641c15fefca8037fa414a7530d8bb3eab59a59406caf410b236ec94773c9afc0a5c960d3e85efa46b2017dca97f14d4d44a0cd43d2313f83ecb93c0e6ea03405619191e36d6e72a9217016ece483fe3710f63cc7eb16f35c1cd040837e35639e3ec9b1f58837d1939803b9cec114ef2ef9af9443b2a5d90f00b239c0ce1f8ae87d6f5bbc9faa3c9b0ab90793d3b4d4d66fd6320e88c00bd7dd84dbbf5c68c34de598c0b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb773c28a15510f364a318cd63c2f89379cacbb8829d9a674ae585afb8e1ba4e846d8855b137756cb3f1fb06ac5307eb12dd2cd93b4910d1b35230a528ed0f27b7a8807c759837edc4bce86e2d716c9400e04e48785dce83a50021382cb977e5e02083517883a5c4769c5e19162cadd775c7569fc6f50e1715f73e2bc2b66e6d81336b3ea6794505ee63030c212c048109ebf4cb15be2de992df5acaa274ab259759ad63865de4258a67cf099e02ca09c4f8c7b25d73c1ab92b6fe13103f7593d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf04774eb93a4f9c048cd431d33c88760b3dd9012a1e96ab5bde754d7300e916898d1b7da3fdbeefc5105a1e9735f62e24ae49b322b3e47bb4b5c9954686474c99b658e3f3e88a9b2df0093e6e6262ffe3afbfca5e45ffad9ab27a1ee759cf866fb53a470086010c46a549abfaa4b5d9a869c56cefe8f885acceffe1f5ebc999df2ec87a38df82bc62996844c426e19f5223eed664ad31e7eb383b35f314536d032639bac4cdb8ec1b28343ee2f4042a065afd9eb6223ae25090a9dc7f7d8f36;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h823f6d5bff722298bfbaee401e6c14ab2ba235806603a7cefd7b73b91c57e78abfd7e0d5661771f1354340d30bc16c2b3c449cc20db53b61286d857ea33155d8344d3402c71d3812d85ccc0917130ede070dd39819cb9283c12aad6b613c1804aea7e221aff336d9a94a8b815c1c8f179545a47493c54c8dd8082c056e35588d228fbcbc28046f3a0328ab68fc3a87f6530762e66aa70013965ce9d19f18bb4f122c890976d7f516bab65ea4ef07a88217709539bdc031a875bfca65309990a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h45f04f1cd40434609aeda07764beff93ce2ffe4b2406bb05d6d9cac7b8ca13e7a2b878de59e98ddd71277e90714855b43f97208b6a18cee3648fa75e8a48c5043769df273256a78c09201ba6e7ff55b1eae51c6c355c494d7bba2702af9b5cc7f17fea3252167854d54c03f828190899d2311fb8e6dd687bc53e0d7127c7e191eae207c309bfc57e1f4cb028666d10e65fcc8d499e20267dec9728013ca5036d5a26c71083f817aac5e8753eee61b341193f05a2ac392b3969c1d62b15bdf66f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8215160197f9053166a3f94006c60c500d7970238afa2e3cb88b6ee7eecb9bc8121241603a86222b1ca92dfda37e356cc6e61c5e48fa945724c97add5a797afcd52541fdab26ebb30380cb0997e33baf14bb2407ce3d1d60271439dcf37f995186316a2944a1c3cf03b3d4051a0dc4f7bbf7aa4a7e13c203ede1ea3ce95c0120381e4961fa263ff11d59480cd333b352bbdb50186c6c0908e7982ac6ae8e097f4656a489de3a4de0856cfd20aeecd46274ac2ef2c761070d346f520d604320a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb45e1061ce382bfac75498e9ab7011abf60b6ea900ff7e3822a0e430eb8db0709af64ed310b13b076d57f9b40778f04b957f682b15557ed454fdf332fbe3396181cc86670240f822d298b9e8fbaa9041b53b3af87ba0a2e01424ea3804a51bd5cca62faa6773c65f3f88dd9304bb01d8cc2fda8851afe1b114fe1a655b227d8b3dc47e62fbd74330e188f27ac6fb04c0311f53408a14982fa39cb6bde042265d0fbb756ff752fd8e62589fb15e1012698203c035ff542dc7b181ab02643f530f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb292800fc852af0787dfda7c7d63f95e69e6ddb24cc73c606eafb0dd2355bf7b29f9ed05bfc3b85a9620707ef2008139e4f8afefc756fc7a65ca22c22f2f56b0a48ff42afc0dd4a6eee2ea0b57419acba8b1b6df7936d75f3abc3d819e46839e1732fd4fbe957e0b93b33ac9ce0e6d15598a50f4643345e1fb74b3c9267152e0d8427d9d8b54cffb1ab54125a500d98b52e3ec7f9814177e3038f3498586090fcab5d6440edfcf0dddec54c8b7622c82a4e9d600cea69c41e8db5dc288608ce1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h666eed607d398cba1136512f530b7fb51549f3dbff0e1f261a0f40bb14457aef34848d4ad063a1e7c8a084fbace456ea561067b691cd811b7e6e7f90e0326316c2f7183dac6493dd618311ddd74c9aaedc22dba011403502cbc4e93292550158a5c3ec380620a6a6c0c594bee5f769c70a96c6f5a97b46495fe90f8d6b6869024b433212a259778c0af3d68879b85a57898d4ec768c92fc43f42f762df8e05f9682f5200bdf65031af5a41402cc32ece227e4ee86d24d7a79ef6719d5fa367fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd357e09c50bf3ce7d08252b76bef90e12cb8425c6d2f4c2293e25367d6decd578ba35ad32193e75fa962a6a84df5697dd6d12c0e906a108950e1613b0c25c7ea7b4b8882c6a5168d1e31259a5bf90e058bf50ed8cc0aaa7d069b7b722ec6e5c808469149f3379f160060696a6ea84b2f8dc791e7b21888cd4a3517195e51740be09f8640fbb02886e9019ebc88727bf6e7276275151dc94dc9afdf32de5181109ef05c41801aa85e5b10adbeec375fd02655df62c0a6ebbfad8a9c51c9a10c39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h49da616442320be0be6018a04615e946ae409cd256e5515bbe49134bcbe7ca087a6e284595969721450b68d91a1d45abe3cb178ee2aadd182b7913c522c3f7fda7a5dff867afe90e662223b77d20df7da09da05d8f3e87cf04dd388cc97e29315c5bf65f60793eb9f88a14c83735f1b172a4ed316e5c4884463911906b3caa7e0e1156ec765e77f1e97a6132addf5502437346be748557020f45f9e602e9034949a4c9ba8f741329d5e381721bd937e7d55cb17b3ea7e476d1afd47ac822aacf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h1585de2c820577daddbfecad910391c1d464425653642d0ad5838e563396f789e0b515bf52bda6588a286fb378fb076c26e5a131cf7cffc066308faef5a1a1fad2d79254ec3de63a2577c42ad913f60a45cc76ee2068962f5a3a1a4a46edd18ca119d50d99a01129c823aa11e5b57813f1770a55abe8374bdab1068c6ba20149ebf8db5e2b42a27cc3854b20ab3c9bca8670792ad2718439af6c8225490dd3edb65cbe7f835bc30fdb0aee35c3f691fa3d8ee487fef04b78018815a7707a29d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h3e727c9851521857fb8b277aeaf24f1e50a37dd3e5328bceb8478120007101b2d7ef7531085622e05392d8c91dc2117d43c8fac9693bcefcaf938728bef522c49debc7daeea24ede052248cc7d41cfda02b3e25733a04298fe220bcbec6632f1a6912d36b93537cf8a9452e4e7b5a7d3ab9dc48c5f45fd60aa0a750d4f253afcf349e2665fc1a4c6de2849f8721e0dc8a7339dd30ee31e0b0a46dd5d33daf1034312fe631e52f617e5b47a8088e946973409ea2403365aea963778a67709614d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h4de7905f4c5d71a9b557bf4a3b6cd5bc84a3c3fd8432d464593e12a240a2a27d0f1c28c86baaccaf0dbf52eb556a0d2da28d70968cf77ebc250dc1a9f3dcb12b6cdb31e66d8eecdca73114ed2c676ae3f290ba1428f80de867f4e1cfad5db1d1ca690b9ece070f38a65a8e6502cd9d53abe4c351d2aaff854108360ee3f69d39dd0a503056e8ff2ce75e98c69cc70f44526889facac18139ff10f191a1dca25c1670af0a630dd23fb7a60320d99d635907be9a7c9c9296e4a9ed78f5053123ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb3f3ff7151f91a824ffef8ad9bcbb1076e6ea7090d9fd93f75e893a097648e608cfd221bebbd46fada519a5e6abd5c6d46da1720021c75f687ace97ffa2b03918ad5246d0abea3fdd7ca473ff5c4f83811043ae20a20a6304ce7c493723648fc027231b5d29b32d07944056a44f56c31701c15f920bbfcb27d8c08b44a7eb293a81692ce65a49e1e0ec3c25cc9bc4113d09a7b7afc55e9649810491a9518c774297d7256c8bd03eb672857ebe11aedee7b48a2fbcd9245a03b0c12a331bb311f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h6689ee9dbbe8f0c909a408cfb999ea18d83b4d026681ba9cf8dacd3d179e653526e01742ed6ddd0dcaa6760b2ccc4413605f4555f553fe772e99a706c0e9883e93072f3bd8e2f45e304d17b9da034f02ae2f3c35eee3b14076c41f078a30ff0d24cfe87935b17ba220ae2695bcd7b0cd75d67d85c55854920cd0670d9c9d1989d566d7666b68fe7f9537262d7112e25dd68048e3eea476adb9862e8d4352532b08a096f2966ac3263278e0423da2c9fbe7f9da971c62c7348eefb1c549af5709;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h1ebb9567deffed7a3a06b13545de634c04e90859d55910faa379f57c06cb9500cde534bcf455df711a3b633b04affe0e0ba39241fde50359b5d392f1d837aff62a64e7f274c4a1902c2406ec21e39c7512f465c3acae5ce611a4961444fd83450304a35fea7379b3cb97f97f8ab395a9c32ca105e7e02495f2b3303bb25ab8d53e6af7d1ae098e8a6f6210f4c689c2f0f8ca9ce2eab0abd298899865c8e2d95aa458d349440c730529b3f2c042f95b815f158971ac67020d4a04e9cbdf4feffc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8e0c7fd3fbc5dd46cc23ec345f1d83dc6e0cb84cd503aaaaa62fefcffe0e5a18525f1add2908e8ea4df8e08ef4202f009364c112d38865d05c9647c9a28ceccb01bd2883d7272e8ff18a0ca2683d73fdb5b48b6a76f5283a78306e55ffe3ca3cbdf1ff4fa6e4c9eefe242bf57d52bd86fb590b69844325ace6c863d92f5f30d99646fec12461750d8e684c0ce82947bbdee8122090a7f851d5d13563d968240f9532ace7c276a858b7f0dc81e3f0b00decf41d8ec901d83e7ba7f87d0787f751;
        #1
        $finish();
    end
endmodule
