module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [6:0] src8;
    reg [5:0] src9;
    reg [4:0] src10;
    reg [3:0] src11;
    reg [2:0] src12;
    reg [1:0] src13;
    reg [0:0] src14;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3])<<11) + ((src12[0] + src12[1] + src12[2])<<12) + ((src13[0] + src13[1])<<13) + ((src14[0])<<14);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bc3454e8306eaef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b24fe93bad58033;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb2fa79d2b65510f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ea66e9531dcc65b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha859a40817e9d25e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90960ccb334fc1f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb74d2bef6c3cbac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78f1e268ba589439;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37e2902cf7be79b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44823fd942de2848;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf558c9a5b79ffac7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h911c55f4fbfcefba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h814645cda3357912;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31bed02f37599e20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b222af939efa3b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha341b0812d652864;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he35dafa7f7c42867;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83512bf36467ed69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd49c244279f92d79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc99144d724edf501;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a5c64f2880bd2bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4639c0928c3e188;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8fbbc0c78767f56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c1dab0635a5289d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b5caf44b0c3742b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b0f8d0077d9e218;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97e89271a0996cda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h304d4c32fdc2b596;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h803e8c8155d2db33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e8c84ed95929055;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc46e7e9adad856c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha17eee1b61c19013;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf0a8658ec228da3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he387d7c0fb5422b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11401f449f508715;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17bf3fdf2bf36405;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddb306a1eaea4a08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc94887c40905c614;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e5d2800a60d3a1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc9e5b375783e3f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17c0e533d4637964;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e736a5fc414aeb7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0552db9750c4d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58fd0aa37d6f1197;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c393a3af32cbf48;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f062341628bcfc4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1d8157a421e0aec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f0b6e4bbe97a5c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dbc2d2b8638a1f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5070eae884bf9ec4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c5db2eab7b6ce5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63d5ec9627702790;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2564c12bd57c5cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c3f365645093386;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b6efb256d396a2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e57f328398de6cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4ff7a0930be74a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde3fa58d10763e94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5daa09a2fa429919;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd38b293d8416f6be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7bac6604f76ee8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1952d6785e54198c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h398ed16558132987;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h693a42a84000f517;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10d3e65825cf8667;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h609eb5aed096ff77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfcbcc17bbdd71e32;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55839ebf881bf9ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcc0716975cb5c6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f4af5885bac1afa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had7a1abafa0cfabf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9bf6de5e8e163377;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h870936a1fb46e6cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcba4046f8b5a968;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3c6fe8e524d19b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h737baca3e1a58559;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9d895100d5da026;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1653729abca4a70e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33057a1dfc702490;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52408ef95fe7f1b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h416bc28a613428dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1abf211ae5f93ce4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb95e073443a0e020;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6979b9169a3834d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he718dd90214fede5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f438e77779d9e1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf00997aa5a2c609;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc6a2043a438537e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26c8ed6a4e791365;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84d586db07a1fe18;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49141249438d8fee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h594cbb24fc74aecf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2db9f41b8e05279d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57bd619f898af40c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcc2588c91672836;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h206cbac65c2ab1f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b8f76948d50b602;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f8cf9fb58b8db74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a6bdbb5e64713de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfeecc93ce55c5be8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66bb56d7896866f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12f5d1a8900b8f76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9091e77e1ce4f19b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18ac00e6f49710db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f92d2b035dd31b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha808b373e8721343;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb315e124b2349e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h309c4a1b49ce146b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d5da664a424ea38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4199bde2dcce3053;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd764ddde794c98f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h878a02e0ac3b163e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8865a4fcad95aa4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha20ded7bad1de18b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b8d39159500f6cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38ffde25b06c150c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d259c083f0dd4ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2609b9fa49dbd04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44bd6a8f125290e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h567e3063257e7caa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12c8468b3f02e457;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5e96769b354655e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77c4e83e4e37b04f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc7f5d1bcb08849f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70c7bc17c318db5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67a0cba052e5757;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd15e422ceef2abfa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c13ddce7126eb5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h254689c69639d3e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heef14fb2befaf51d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7ee24e07286c4ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b1d3fe83f9efc7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h250328cc5b240426;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e7e179caf59c450;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b5b929a92e13af9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39dde4546601adec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd95b10924ba3ef9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8b6969ed8d04e90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4f0e042421d90f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ca666c05f63456d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d06e6ce1a6f6ce5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66d3384fcfe46192;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8eecd93a2c03d639;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7fdfead1f1005871;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ac2ce6916f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8997f59d58675382;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98aa7cdfcc1c462f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5d21a375511fe77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2bdc7d1cc8ea8752;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedfae8f363440722;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4b5b42174cc9fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2911b2016ea5deb0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h638dc1c2dccc5597;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42dbba3088481541;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h809d14b4910ab274;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8f04230fdf25e1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5da84e4470cc9265;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d1b8d541c2712b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5a59710363e05fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5dc8aef56c64dd1b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f136f3b3ba54dd6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf79ce35b0ebc6459;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bddca9404d72c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5af5f51aa8e635b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50bf36fcb1926f06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9adec82c55da97b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdcd183444459c01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha93dbd61c04e4dcd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74b5bdf881dc1e3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a7c5be18599323b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd457199f97395cb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdf7eec6524d9a98;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h784a1b85cff0ee72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe952ddd89e966ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48c0a54af03b9e68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47e189a9f425a391;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dbe6029efb931e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae6d51bbbf3b4a9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1e1865c2b88e70f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf082d875f79dfc3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h119f7df7e29989b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61d916b915296b19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40b2e625718ac4f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h196c971bbacc452a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc37d5c5011ed997a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95c6ec66b7a0759;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h118bfec4b96a6e3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4690c5b48ec3ef7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24bf8438e9674746;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha499578e80cb5412;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22ff39b29000dbb5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7137f823934c367e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6306e3f2d353079d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9b6a4af7953549e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8ee2b9615cf1228;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43017f43a805b54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9d54df1bc819b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce4da2fd612ebf34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h148d0c305c2d40eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95fa6e296ea22239;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfa64bd97d570fd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h387b0e8b04d36d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9e0063e6a759e76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9313131c69832d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30859803bb11ba43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha88a6b9b5e507242;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcff1f5d221993b58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0dd554880412c15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72f9df69a3b0f24c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a7848da1fa36159;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b434d63f3b6f1be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdaaca198b0e66ce3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h918dd9b3b945a8af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc56e56139775bc9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd89cef6749a3e10a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha232362a8dedb83b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafd7ca62e7f3f5b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34fbf1aa551851d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14862df789d346be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcea1f50b8af721cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha927d9380a57f975;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80529b0cabc03873;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had179fc0ac514604;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82ca632e0d81ee9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42495b5259778dcc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc81fb0839e2bf1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9b437bb3a50aa3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea30204fb4fb977b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ef41a50ef81d3ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccb44127c52a1cd6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24a2faa6611571d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3826a885812fb25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed925ffca48c81e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a347e8a128956d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fc0fd59a99b380d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5f3998d2fbaba80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc483b89578ece7cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b977d0f2fedabb1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b5480c11d3c3e7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefacfc638afb273c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfa5318243be5741;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1297f983f533e175;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb700ecf28a04bd6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65767ccb223d6053;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4d54980ecfd592c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef975dde7e5c18b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5d16b9bb23d4d1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h165ef8d491bac3c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed213d4ead7a1d8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fbe6afc107676e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27cb0fe8ae9c7258;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd66a1269ee5ac77f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h795f87c01600d6bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81725e9abe647312;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3411a2a0126127b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6a0900b7175581;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4512ae700a70975;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89cf4b45ba826e59;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95ba77f859e26e6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he56bc079b1985692;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc72a8dc1a4c98cea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebf089e0aab35fe5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ba0383ae3c0b915;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5bebaed7286370f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdddf500a27272a3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc17ed06404ebd9c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h851fef17a25171d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40715d37c79cff65;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb76082028bc2139;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h920cd0d9eb65d282;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a3c3901c8a8d2b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6fe6fd0499f668c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5cb89992dacf5e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac1dcef5a418233b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12f832c98cd1d5e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f6af0882d0b8e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab56c4980bfc9fd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h626e58714759cd08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4442169a11018cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e576a1a0ef4a89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd57e7c3e09febc8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h701a8270805f266b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h694a5264b4ec02b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41a8ffd873fc6507;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h987e058aedbc21f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94d995081d0c51c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41cb1df232d4c0f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h128c3668d0b9547f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c6d4fa6f108eb5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a3553e9fe1bce9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb1e041adba98d6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c0c1367e5efbc4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebc9f46738508a8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7107c769a081fb3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h798b013dd321ef21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b1bcc704b5d8f07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5956beccb1504e32;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb22b11a7511f8ed6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf91717494b5b73f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddb1ae45f826f367;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c6297f5bc04c0c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0a0d2082fb0ba54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2d72e4057018b89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h576b8cd3a068cc4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ef3d4d0f2aa9a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4661dbc93c8f5942;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcfe88ff881ae982;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55a83ab64291e3e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h746e3dc3141fd7f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68a0a35d8f718f6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ee01bbfb767886d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5278bd953a39078;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37fd6dfbaf81eb32;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee200ce21ac1baf9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96874c2a1a7c5904;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14ad7827e8c8133;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ec54a15a346c635;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8774f29f5e1e170b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6cc11f2e6ddf0bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h513e742a2cb6aab4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h477545c1df5e2332;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26786af4a0df865;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d92b963ea0b11c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87d2c8a1b2861c21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf1fa7c9533fbaa9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec9ff7ca76290b7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ef0a97002482e7d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea16c9ef489d1aea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf1c1bbe15a6872c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefe7dd8e3d9dfd67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he075749ff830fd76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2bf36f1f556b9cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h468dd3c3faf2259a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha23e82133b448694;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f3d224b002bdea1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b710d7561a1c4c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac5b5d5b03a604c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f8608cf0a96e418;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h271ab99c13e69c3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17c5ea548a59f95c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fa4f141738f3752;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8f1461465f67331;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d5b86c68d254942;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1ade0f6e47d44a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d8d81351da9930;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h140d5bc1d6e140fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e8bcec6b1504574;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dfcbefee9080c5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a8d9f70fd8ceebb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1706c28d55547903;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32e1ef5401a9e0e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h918eabe53d21cd3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h520cd7d130add484;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd11d290aab12244;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h112f06169ea78312;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h934ee87cb34aa07b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he33ea61a6be79830;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56ff32ba9ca317b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he94a44b3d948f8fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c5f02b75c28def9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19da687a355fc0ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6f4e5ae433de08d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7326001be7918003;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ac6f0fea6dffd08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6c848b37971abc8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf66e14985e63b9df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b9ae1d4e749dc8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ebfb72686d8e067;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6e99d0231982cf4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h236e39e3aa85d46d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf7cd7e6a3c7fb84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b10ff4f0656cb7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8af59893aa5233d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24bcc9517f876f7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0241cbe7cf16823;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecb813e61c9eef7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4ff5c80f9888e09;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb007e2c658bda97;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6b3215d2cfeb845;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3eeb980af2edba9c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c9f20a27f202e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5bdad41d05bc187;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24d5c4e9ca5f82f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf21e01d1dadaa31e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b76ac37b24cd794;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96e911c35a85507e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e7241d6dc264b8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h633dc1b39243943d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15a06ba9b3013d43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he164f2f3cf2af93d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6e9f12e581ae197;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec5d1836c7f12034;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7430353037c835a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91d98305526dfbe5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefcee195a0411e3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h666bffd3560f3f9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb921d76ad449f722;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a8f673b0ab7539d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67ba16cf8c5927c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b2a5d210b11e119;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he330991241ed3176;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac7210a881e0fead;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d511ba445aa36ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48fa8f81110e2a2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc5b86ce0886dfb0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35dbee14d10e7e6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf12640a540712af6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf1af807e15f1c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd2dc8e900f8db05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd537b6965d628b64;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7a861887635d9d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19fd11f30aaf0670;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20d0260556dd4979;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfaa39621e517756;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc773b44a3e68e5d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda8894b8cfafe00b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd883fa2413c32d38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58db235709bc8674;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4847e0300f98de9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97f3be1a3e6824c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h309b8c6f2a9f0df9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h349f72823d4c8a29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4aba13a2f7e855bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcafc42bb6c542617;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbad4b7ecb7ddb48a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h840a42309c56312b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f553921668eda11;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbc508d7233c044a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h200ea0f331c2b8dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b11f7a97139ba20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h208e51c4f041bc96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c11b6d88d74e1f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h909970648c2ec9c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6bac1c206b359cc3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4231dbe98383239;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f9ebe66de24ad56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9afa635cab7bf01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76d28ee49422a34e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb9f05a9199186e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccbf4c7bb27e6213;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21234e6cb84cc6bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8029ebf01136f1ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc1ad58cf44e537a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae6d430c88986d2a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h621fd33c51f3fc86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2638e7c3ee18ce9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4a524459515caa7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa59c020c7d7a5c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98facf974fb74b3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d08e9b4916c9487;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3acef7e6d568c323;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he99392498ff6912f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7aeb5729307051db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7e2d08dc7493359;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha25614a0fab26936;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5cf6878c0bbd48f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c54749bf4d21b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36907daea4c18070;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3aa626f5aea1e05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc87426b10bb4628;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82720689b5fe9c6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf54d446765585ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91cb87d9f253c421;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd9892dd1b7bf9b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha009f35024165e4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46d37294a1a7d5aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd725ec06c0904b68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb81838be5a6e10e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h677d7835efa35aae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc0558208020c272;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h958810131047e0b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ca8d23bd928a48f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbfde400784397ba4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ffc05cd7873c0d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb19e9d6042838f62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc441c3e1ec43edfa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3edeaafcf4f671fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h196aec7a1a03130b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1326bda692d530f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b4a75e7706ea373;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65a371cc2a278b10;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f0ea8b23946f494;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e645d84643e8317;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h888043690454166e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb99c289bf95e350;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha938d1d1e14117f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8dfb74039617a6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd208fa83844fe164;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80b61022c5459b89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h783efa3ab5bdc75d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50387b2f42bbc7c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h784113e7760c59e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe031199ffd4e03b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae7537896642a98f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h574aaabaf5eedb72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8beba5ecc7ad12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h575e7db0f4649e2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he70955ac08cc347c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha62d4eb23e44af6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h523840c77d5d8895;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19c42091aba00eae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbba087f0199d3af6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h581a2f652cf0dd4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4dea411efdc8b9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h465f3230b041172;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heae5ef6746336a83;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58be23cae75700a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda7cd7a01a91728f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45eaa0df1c24321;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd993cf40f8af494;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ef3b5e34e421361;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e9ddde229dacf21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee5811b7264c1a2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h650e30385414d0d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha590c40b934cbad7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd948da3119e89022;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd562d5fba65d1145;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f84c0a8ee2eb5cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6213dd32e177c7a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57581508ef511988;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd7006f288cd7da0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h479203ef5ef9e5d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd34b3cae5754eb54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd83338ac689282d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21af33ea9756337c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3646e49f01bd664d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b80cdf44f13524;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20516c75fe8a9cdc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8982b35af9b31050;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56f165dc9a8d9a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc9459ff66c31f75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19e1e44f9b3801d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5e8a2a4628e3dfa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd283725d3693fee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33985bf1e8c8b41c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c4d0a92308479a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28cc5a41e55751d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2291b65264eef43a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2de1d68d26c9d7cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cc0f4a3f8eeb4a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69160fcaa11573bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dfe1b400b086b6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde7e367b3c92dcee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf85dbe193f8b0680;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45215a252afbb5ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcdafdfe2bd3eb6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7aba57c568e6d96f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2bc7d6707265461c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b3353301186fb6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h652d5edd27262017;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c0af9eececde382;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3385ab802aef8242;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c208faf68e6f7c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbfac0e0e7772614;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56265e65430a85fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a7d696b8e1b257a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59753bbfbfbc41e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4357f80d2e69eca2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h228df556ccbb8a54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70a36b324b57c14d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb668794245d2111;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3760cac05a5dd5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heeac590c908bc70c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48d21873d255b376;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd1f5e0e5ed95bc7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43c6e08b42ba0860;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6457608183099ce9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9870e3e10e3b48;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h184852f73a749d88;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53647a5c33e12b33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8458a64ad906432;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ba704e9f724fcb2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49414a06f42b3053;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee1df864bf51a4d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c0bd78c7e3bde77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38c8a01e5da0def9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5f84c6df37c2d33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he18e795f18f691a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66790780f1139925;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10b0fe93a564c5a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1bceb450edb3a9c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5334934c7d5ebe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43a50d66ebf4f3a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf061076eb9664d39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3fced83653214118;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h581ae27d31ed5c6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8a57cdda59467b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccfffde2d1c7aa64;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11ec7c7d3438fbe6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1cc5e7e21b4570b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3ff5cd12a2a0dcb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d7d857745ec888d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17c78e317978f19b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3075db5251b3cad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18747a22806cb5e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0577067823ffb87;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb64909910d18338;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ac7c84ded1cef6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd054567608fe6c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6109d967a9cf26e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h413317820e926078;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha37cf5d6e0d9b557;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h443c159cea8a1acc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb11d5feea7f0c644;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57dfc1fc2d3eb71e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed98f5b782473765;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f4b4ebbc16b358b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6812687e3aad636;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf90eeff5e1bd763e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdc3f26316fff1b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha581cd3c845e8e95;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43b667593f5a4390;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c786abac7a6f238;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9752bdb73401858;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b61f3364c079b5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h368de5fd36d398c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54ecde0085e9b3b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd51d304a5e19df58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fbdecfc82b30a4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb23ac1647b1ab4e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he50d02f224923d0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h712ebca9be4f71ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h302af1783a2ff551;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he629956545290d7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23dcf51849c13260;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b778f82269b920b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62af3793622ff6ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb474ba55d46172d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb419317ecd8bb718;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4af977000ac9698a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a178657ee7b32ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a86bf21240dfbb5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bcd85040d6ae467;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf6c30de5dce46c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12b1b8bebfdb35bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1668521862052646;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24996242d54c2e5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b17f0a0316ed16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f18293b71df417f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfcf880b50707c104;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h168b0bafe0c16df7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55170573a12cd55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha17daa83fdbef45e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8021a904ab23dbf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14626500b604afd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heac90e78352afba1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f13f8adae85e9ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcae2c4ea076ce942;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h130b88457162a79e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6534dce256ca0462;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90cccc2bddab84b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefb30ac221196ff7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfae92d47c45a5f79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14a2cf8a851cde9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h528429a50189b6af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h597792dc31ea2008;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbede1e29ea27683f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcb075dc18b801bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac8aeb674d1d4aa0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81ad69c64ec7e774;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35132b64c9c627a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1056d514aa505ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8551a2d7ac5337f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d7da37bf672c143;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff0cf7fa3938e7e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39df6591d5462e2a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3958e440eebd9f31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10c59eea6544a83c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h159387e8c6324965;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h651482abcd6164a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha15c7ffa32411334;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ac432ed6063f55a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c22e66df0ead46a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0eefe5185892503;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h300dec323de30aa9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f75debd896ef094;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h195651d2f4c43a2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha91f1285b2701938;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha98db2890c6bff00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8389b519440e1950;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0f750e97092a162;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf3e175d6475cd40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h722f9ae537f30cb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33ea4068eed5be24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11d5c88a61e798e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he19725832af37c78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a6be344fd1c6c36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ffc9af63752d311;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1cbce4e6f8b7de6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b731aa2f76443ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6211baa2d9c657e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h967559c09dd29e76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf514cc8644a31152;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbede491c1fceaa0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafa05d105c1127a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h691a92cd0b5a83ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2194381a185d7d33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda8917a068b89398;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f6008acee4bf410;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3d091373a5d4f38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe4ff831492ac315;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27df2e39bb5552aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7136f3e28020325d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86687973355c6b2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h433786f5d597a562;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9a2438269ad034a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e3057ffa67544da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd89764b6b42c0a30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbdf767225cfca257;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd44882140ef0a401;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefe8313f2d6f405f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd628c4a9356f102;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he052a487b9d4af2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6499033d8971d2f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8781205fd2d11d2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6789e9e35a9fd685;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf82b3754c5a44af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf04c1971db625b44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heeee1abb3b3d2ece;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b0adec4167969ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb0ac139bd10ec64;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he79de71d244dc429;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93a053611db10b48;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ff9583462605fc8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h532590eaf46b3209;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h916fd2bc998db1d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd54f1f0515ed13fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3717b481a3b4d346;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd5ad5c041f4e690;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7706657c04faead;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9df51a9761a3de12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38c5328e6ca3a2ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba9ad236755dc805;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb70b11ae8f89b54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0c43f6cafb39994;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20fe7db28b44ef62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde6e4a066b8a1f60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b43f0a07fe4ff48;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heceb7405af7d57f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf56634b2518f61fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb667b7924b8f3cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff278d41b8a98f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae7070ea530b62e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84a3bf432e8ff07c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7070a1667d0b2e0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7fba857176c3714e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb82a7ff430e8dd6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84a0a2b83cf167c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7be6fd68f5260f1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h802fbe9bb79586bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f088cee4413cadf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15b656dd513fbaf3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1aaec85b29906434;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f05a88574feed28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5c65bc836ca7e63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7349a5d2c8e7465a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64bf197c9676e486;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h399618db0d4565e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc565cc9e156385d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7bac51c180a84b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64e8ee1a581f7ec2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46df764926b779bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haafa03911895cd4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb81b3f394817aec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f401c7ae2745d6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34b9518b50d6126a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b74fd1e55eb5bcb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b0fd1b948265f68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d77cb94fbbe1bd2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h906ea360a79c0e8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ff50cbbe88ce226;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h682b4010b65c5c5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6450344147968eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d9156a9f780fe39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he16022273a533d74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28fafd8c90fc4f25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0434187489014;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h698bcf2d8feeee9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b1abb3b9e3173d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35afd1b0a0866128;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haac24451c3f106d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7313e9e12f3012f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedd7f1f48d648b1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7904e966281569bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c30b5359c93e2f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51684ddcf2efda3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e764762921800c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h958a8468c32e469;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d78e88c63329cfc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5227f20c46a45af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5aaee46c8da3e365;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed9903be429f1c98;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78b2645f4665ff63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfaaf87c12a01496e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b9d30cbeda2c89e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h789ba7db4c7bf3d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5381778f7fd69813;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h758d7adc1584729c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93dbcb553d0afbd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2916db13167f36c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf58d32e29392128b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a83d0145e19b263;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90e4a15681d6af53;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f6c78c41b489980;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8022491c959b55f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14248ccd0cc1df75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0a4b5bbcac90ac5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd130e4db7a0c2815;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h923ee636b2e641d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53e40caaacc19cbd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20813b0247839656;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6dd1aeba2e97f63a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee309bec7a4bc71e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc962b21dad412ba7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc33ce1f14f505fc3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfaf3173464fbff05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf06e28ceca9b13c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2663218ae6ecd574;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb9f777a3d55dd4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e18b4341f1eb50f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3fcb9076be89081;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62135b0bb126c249;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67eb458dec9e245c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd10a99466bffb5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd79f64b8831b4f26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39a44c28992db3c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb67f6f941a50a835;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52a06a84aa4c334b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha295a144902c9d12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h145e4c8a1dfbdbea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c52484a209608a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64b9350b8ccfce92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f50dc3876b284e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa97cd8aff79e99;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe3d3104d34f36c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39febf9f414f4b0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he61a701b2dc17d56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haab2abe1e69756d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f16812dc9619fe0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6dc14771153a465;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc28c73b80cfc459f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ff32186de37f499;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e7d0501ba538b97;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c9a440d61f64952;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dce373be45cd813;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f49f5f613a09fe0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19b9f716bd9bb888;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9e9415ca6c6b372;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a7dd157ed0daa4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97ba8afba0b9a0be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d2fb13f1e43be5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb13d51c677a1f418;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfff28c1bd647c69a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7681aea73bf5342;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cc16d10d8109e04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha976020b041492e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha39cabaf812d9c26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5aa21705eb578b1d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae74f279b9b94728;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had710cd6d068c510;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90f6d51de3fdb48b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9320a1ecb0bc7283;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71b77f92b1becc8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b5a140804e3622e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h380a0edb371fdc85;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5edef4ebbe4f478;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc36f2a0e38f3887;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77a165f07d2fa037;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d365e4e60cbc3f5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcebaf5d0109e8800;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70b4bee20742ebfc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37d8b703a7089f01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92814751b5bbfdd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bea9349e39edce8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba4e9fa8c4e0848d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f887bf5434bdf74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e1759cb7ea7a194;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef321e7b55b9fe89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0c7e7f3319fdc07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e478f088b9669c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71471ec38eaa65a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8e670d33490ed4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he68277694f9ccfae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7da8bdca43184a3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2d81e21bfe919b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1703f8fbf209e5ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70e87b0feb5b09c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a66e9e94cd23603;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc046dd3880fb2c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f22d0a406adf095;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5be95f97e08680;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ae0882c26ec5dbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ba45a5ab6c5a0a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he37bbb01fa4a3d3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fcb8100224ac2fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5584daaa589cb1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd568db153d0375e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d442f886e4e1c28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbfc6f33b23c7b968;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61ef8c0d3aa382ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83fabed9455f81c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbaac9744cd8521;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ca7bb849fe9dd86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf95735f466dfe355;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3352aa9dd7370f17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ad1b91a988dcf8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1a45bb63b1332d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8473553b21a4e4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b40bfff6e0a5992;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h901aacc73c696e2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he007afc2d8d001ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc55e9c7900f5a265;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6363f377eab8d08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb730650ccc1166f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb159b11834a4eec7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6725462426d07e24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9f21e71df852fa4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb198f1caf753b71e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a1256790236db45;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h385efd963f1fa205;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6da36289a09f62e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3abf2c9936f54c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5245a595396dd10e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d82e3d03dcd90f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91fd5090253f2783;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5bdf2f54f7de4e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd14be435c6ae9eed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e9395f352988baa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d531b00c3d602b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf56976e349d244c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha315af70092d143c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8af42987be467b3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6d3f0feea3e413;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2c3e2b2ed05014b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c106c43dbb0637a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf46fa281b27d49f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49d611a4c5e2e95f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h293743ea1e190d00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h933394c39a7c3479;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f7746aca049c5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32073e2e94054262;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d89c5e62cd1a26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h997dd9c0433103de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6dd4bc623e54f39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0adfdc08a8dd410;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he90b0d2ca06b5592;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb166b158c1ddf346;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc97d40a7fdd7d090;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92ea75c32c71aa51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30800f7a657626a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb41ad514b6b06702;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1955554f1b561d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bac91800fdd7215;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee98b1c2d344837b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdba9af7526c3055c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6cb40d541fa50cfe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a4de84f35f12cb6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6ec74bf4fbca3a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66c500859ee8a5b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha913d1a5b0122113;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95292aaac13e6771;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8be65c4c09115699;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5f77bf86233d3ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0fd79893b30b8c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h203d3bfe7e124d28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3b5a29b601cd7b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7cfa3c86c1d17c54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7987818a641c0d56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe91188406a1f22b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9217e00d405011e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a1d6eea1e6e72d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88def602e03d2378;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5cfc9f9e3d4521da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4525f3dcafbbee67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he09c0bffa3f35a40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h201af15ed5c0fa02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86fa8d4aeb586881;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6a333800573c281;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f741c0e9668c9f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb3bd427edeeb2dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ee7128e00be7af3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce9928ceca5d5877;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf22ba7cf7907627a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7afc915e6c5b8ca9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc29806f9439fd615;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb52589a4148b16f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec14f28d0b4c2e74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3678853f9c855c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb68c023086e86e01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0d100f2bce9fb84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2f527cac5e9df1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he191bd070d7e3253;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f1bd1f24f002fec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h748e1e6b4a890c46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9da6e5f5c7b092a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31a0797156978951;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23c4a37179a7807;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45c8f2951f5a436;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h752fc9b48371a30f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1b4e4062e98add5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h928d7379385d3320;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2397412cc24a041;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8575b7e5f6aa4bac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcfea40bb196d0ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73217c98aa466907;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h240f2dd9ca182cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h248043b85a2a9cb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha93bcd405f913589;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he64070706d98c62a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h313542225db1478a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef38e67980372319;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f75af7021ad6e9c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b33909f2c4b24a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d9ea55963cfeb0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1767d38fd6688456;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd3f5853efb3b8ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc57115ced4b795df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha28f9b75c255c489;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6146edaf12a90636;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0cd1b895b567d02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c63c2c961c739b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he501b7d86f5aa7c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6faab6caaa7123e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10bcb2b5d74b9fd1;
        #1
        $finish();
    end
endmodule
