module testbench();
    reg [18:0] src0;
    reg [18:0] src1;
    reg [18:0] src2;
    reg [18:0] src3;
    reg [18:0] src4;
    reg [18:0] src5;
    reg [18:0] src6;
    reg [18:0] src7;
    reg [18:0] src8;
    reg [18:0] src9;
    reg [18:0] src10;
    reg [18:0] src11;
    reg [18:0] src12;
    reg [18:0] src13;
    reg [18:0] src14;
    reg [18:0] src15;
    reg [18:0] src16;
    reg [18:0] src17;
    reg [18:0] src18;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7f23fe1a57862b70349bb557691be7b2069737b69575d4dc31ed6ed89d421c35a24dd3cc5a4cf53a58fef1dfe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7413856404bea5f9ff0a3a1a0a076d258035b75c3336319afccc61351f75d184f8f462f3e6945035c088c8724;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h247228597f87bf3e6cc78929dd928d40b845b574325751bfb08095eb2fcec786b5dc9a337db39497788f306072;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f391ac5cf4df58248d3e3fb6c3e9fcf483c173e374d9effcb21150c44a55b79d9a74a79f57fbfab48abc5c74e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha42c9984584ea3b8afc45a7f7b5636de2fd974ea97943434a72669b4ffed0f7760bf3a7f2c429c54c3999a1a9e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106bf9f9cd30f55cadd1f75c070428fcbce35917184a4df4abc191e39f0655962f1e4d1620221bb5b3b53557e52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184ac395bb30ab0ef0d86eb731ffd34849a49bc97b3c5bb0ce1010aef6ffd6d8fff413837b4823959337b715be4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb8aedbe632e79789db4a802769a8b32a03dc54b941a2b1e2c13e8601c662ec29171ba97ae8d7b90ba32ddb813;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1898a65e8ddbcb874dfa594230b24c42de53e7ae3b674e2bae9f662741e769d942a5a6286d2272fb89331f49a81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1947f435cd022d89173cc3f010eb1dab142459e36b00ddf1f2d47e3e97962c2dd0ea89cfe7314d9bb4f0d911f47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b444aad9a21957df4b91330a04ba5f9b67121c6b28bce485ae6265a2dd2f66024c0e554b957251c0dd3d19c9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9f83e5512fd841946a5dc8a23fad7fa6dba9ebabe2f49e7c26653944bb654b8123e2615eaaf98b6b5711bd9e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5689edac76a01837cddd3df97ed11e115daeaa460806d178b0337f4d95bbaf4127bfaa52fbaaa9c770e07092a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d819aab41d55747f31c608556f017353dfa2332e83a72b92d71f5e15312c95b28d9281f6ef86875e7e61cf66c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16789b0959f8c4c9612fa4079abaa39ea9e7c80d592d55ffc739a882d9e8eb144fbbbeffcb4e413d2d6bb416;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147b75300a1b30f69d66f4f966d1f66170ed10bddeb75ac9c193a7b8a1541ac4102f1ee7d4d55758645141dd721;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f50583a26ddbcc6b3e1ebb848f0cdd8c3e74aef42e2bebb00c04dc55b8839444e90a79945e17b5d28c4884fde;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h581942d264633fa297f583e976d225a72a155e56de3a78631e0c81b3b4829246f13788b0b0c162a34b066da51e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8af2d5a3e3efb660582fa723c14a94c7974bc5126c06172f45f12e1421d353e07fb578f8bd9dcbaf11d7fed695;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f386e4ba60101c9f7ddc72c518fdced299ac5b2b5aeedb379074ffb0770a735089964b52f587a154ddb23f2e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2774cdd48f3e0f89aa033fc19bea831531e7d90cdc1783e3b3bd7579ba52ba875d9260558627a59ffa643b66a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha77fad07c4b1fc3bdfd6d9e2ffe16745e051b36cc3de50a4122ff95d2b933729a92c4d82f5c9416723291f8927;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7d6200ca7d309c00c23c05bd651bd3e7937449ac296e9e02bd602367786d353519c34663b2bb10a6cc7070096;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h412870547bb81a1469b4674ad552826d587b279642db26f36c4acb723c866b7fe67ca3abcce49d3a3f814d8a40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h84867a1f9bf2c550528a5a76a5d1eae2fdab657e01d6f782bcc13918b4fec03de1e9f1758e046f36931831eb20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3da4673ab6adac696f13275ceb695db27062b77fd8779dc40ee71f8fd5f0311bd181c3c0e24ec888b8ce79a21a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1260b5a2440765dcbe7e30a0aa2127a4efb7e84870833a2dc04bee4b0333b97a9f09e8958905d5e0e7a31ca2ae8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de27648aaf906df7c3c9b0059a85c1687e1195f6482b17db9b6e5b1f767e2def65d43edc8d26e92005c6baaceb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbd5c2da3286cf66d6851956d4e0559fc7849ba4d594bf4bd65ff88cbeea6c1dc2fb884a51130c1fdd59b8c63d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h85e2cc3768b0d541be34f159bc3f6646aa4c402aa16873b0cf1ea24bf73421dd7d4245491815704386f51cb16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h275da6d259a6c88b826d6edfe3984fba645cada97a1ab18c0eebf45065c571ec9df30f5e4bd8cd9a30c56ad18a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149ed45bcf4b031437f21b5b7d9c15ed717e85d8a566449717306589490159ce5a583134e228ad2885de9032c44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f32fa9f32ff4abcbd3c221b3ce928da52ba11b9688a1a855863909454e8f9aaad28c8d582bbc65f45b66156491;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a6f586b3411871bb123c67a3b45635b02aa2507c2a3c41555df7b4ae2dc9ddd6c33f73178fe0c3ab99b4c0a30;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132dfb65d6ca5ed32d365e8670f6d0be6a0bdba9c535c645fc0f18d0e89dd76e9d3d149b07bd07c6a9e52972caa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70a73396373e875fe3df748ca58b2afdabe9e0665fa4dae89ecda4ecf7c2493f7178b0204dbb572b5e6d2d9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb76b506e03aac43ba076b09380e45e95e45f5b637f76401eb71fd3774d50530621a026f8a4d349458e18c23e1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1db24c8977418b799145dcd708d6608b50f0e41b27487cf89c0f7a3708fce8c5b3317fa8778c6b1d894a81b01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h610e2406877b4eb8623d71a6813c7c2266191f7302c4e3b4ea5734c66a5b31be08019ed6e8acbc7189d9748980;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3c114235b949cb3d8c96833d7afbf7cc1cdb3f5d54228229bc89d39f1a60779c30b0e7c04e32c739303d6f78d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a88b634beb306cd790baa8746d94093e994d1fb70f53b1d7348996d631239b6fa6eec813b4f4f336a533c921d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1701bc73dbe8e0c5c7372fb94ee227593a7d143e0a8d61acfe00eda000f93c7b1af341af7446976e98592f6f532;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h183527bd246583683f369c457db743208577ba854f13dc10a24002378a2b612d433838d2368e0ce6f4ae477af77;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10da4a2c84a064041a3e6a2d019fd8cfa25ea7748383920808a6c9819f8c408a291b2472115125fa9aca833e3a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f44de0faa19d925848b496fa2f3fee97b31f32ac8e70e2e664f8ebac4ab66063817e5d0f387f51a5b7ee09c0a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf54a035e956d3725cc6c47081dc423939e78e7cc3afda4b6bbde4731140c3da948e26fc1bdd79a59af8a04d3bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c50aa2d3520f1757f7377004f78f0723a211c23170c33aea2e4dde479795ef005d393f557c74f4214634750b59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a6cdaa2981821bbd15641f7564139b233dcd1e37fb5ea6945a76efddb755a07fb225f8d0a16432b4baa8a1174;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12432e340c703fa3a5747e87bc21ef5c4336a8e58ad409832f4eb50a80c36503d96efafca6859e9eb913d855408;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf5f15a579a6bfbea893c33260c731d3eccc1f4df1bea45bfc4541bf5aa35d12552dc515df725ca20d84c05391;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9f9b496062342964871c2005034bf1e9b6d7872f80ffeb7d9df6be5ff798c76b90e409c3574f08f44a79a0c47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c1c81b7839ea02b4ada67bbdc580289adc99e61eee64d01e808c34423ca8ef2c27af188aab801dc45c62909ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1f890abc1daa11327386e9685d2067c1a8b4073f869f9e1f2d2f9832006edd61104e3f7d4a5135159bbd235a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha0630cafde20880308690bceefd645ad8b0133ed03b5feab2ababd2234b7e2c1a88234ea4f891e4205c89a249e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41828d3131385405e1bd03f625c36a55252887e2d18324899cc6acd0beeaa17bd86c8881f2d9d2714d4744fffe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164c4dba7507957de9e54851f964daf15be7b994a7056f4158e57e283bde720640c3c128986ce522fb17ea2dc98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fdce6d2fa1fb259603db48f5b812036742d6f69f7e8437ff75da7c61bb807954eee376161b8e654c40536079e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189ba3fede7c3f01708dd5dfa0a19de45b433f225c8c13059de0b39527c2f51850dc19148ee065887864d67b755;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f6d164d6f52c6342d16e435ae945c7aef951ceaf568c409ba4297d3ac98e4de7ac7edd737f74f5f530828bbcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc174501809913a06e3dfd650b36afa406965e2746c1564188d2fb1cd9061b9229579cc091d8c1619796c18387b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1233fbd0e281a05e89ecab7ffcdcf20a3c5cdab81b6c9b28a9cc922f4d88dc413aaadec03df9c2d1fefbaacac0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30133ff595b65538b9ebf1b07eaab83dd68bf405aa8002bd57167835c487f7e0f3274db0f4a7d61a64731d0686;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2264d8e0c442d669f989521fae6d6166af7eb5d18a1f5f1f131e9ed75a49dd7ddaf2be63d7e1339f9ee5cfc9b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d7c27be87cdda1d8ecc3f9f493bc713456bbafef8f43d685c046a357988e25d8865579eb054c211020760fad0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10eedbd69c9f13a30a8c2f5e7ce120208e513cab7639289143615223469c071631f7e667d34ec2b9c25a7002bc2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a1147d98e10ca3fe777077a783f20caea507f1700565b23d07b76de39a24e0ffdd1e4cc0cb081edec0c26bc72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e927deffb2f3ab6203d93ed28881db62a72db9c93a9f62f92e69dd36c9ceb2ed43a1b47ae6a4f84b61932bf0be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h83e43993e45c9ed081ad80969d9ba358414b6193ef52d1b12f45c0789abcff4d944b11eb71f3bcffe155837cbc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f43ed2fe723e7fc1b2eeffebdc5a5df47efd2934a6726d77b392a73a81a09fabde92ba7988ddd708950ef581f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1030de2d6ee33b15de09bcc2fb6de9e0580ae0b5873d46033cfc5c15e76473c9c574a451478cbcfd12355dc181c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c6b020acfcbadf30e17a27f618a75a6133ff9e93328f52cf66d3842ab3f1d167d4a5f366974db03743a82959a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1094ecdb4259ce35aaec716a15a67596d696be424b9838bf349334d26c2a4ac713df99cc00812bc7ebcca6a7d64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a80490eeaec2969078e9144e8a25e1c92c2ebaa180eff28fcfce69e29858f383ba5b77bddd8baadcf3b0a480c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72eda22835243c5d036d54767af4f2fb9e32dd60bfa65893d18700e7fd192e6508169aff89279e707afa1b1b02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c296b146241df6f7a37ffba1afddef90b2e2d86a5f52c84da97e19ccbd594533e10cf48dd853ef671040458f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199e5643f02c47357628965da173758e1ffa5d2f48e2b8c362fabb65c26781ecd500c88bf8e2ce784e7491eaf32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17922171392a66038a7c04ebe513b49fec8784613591757105eef7e09617d8b3784cb19728b93dbe45c2bb09e0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd3f3b700139d4a716011eb4570f10a3d236eb2c03019264f34a926c80a8e2cade4ebbc3a4a5e3cf1a26f8bba1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h102b6ca981059b11c9a862848c0fbdc9496694cca8f472bc521b0e271b8c0327d68af7ebec856eb3cba862e0bf8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf532a1a27d6e57c528c45663a18ae13f23c83763df77504436acd6877bc00a4a1f144f81cabe00203e3ff43588;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28343e5481069aab8fe003fc8c2ee9137fa546c12402dd19534025ff89f6cc03c3ab268d582062ed624b1dd71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1381b132b0227fc2c83db5f4f1c0c2487784b686649e3b86e8692839f769f4b616fb80bcc8994adc7858b71e025;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156a319b891e0638d06760ce60b6a9aa53315e6e309a5ca87089b62064e0039946e66d2225421e0eee5e00fc2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c19d8dee7d91b3a024b396972a0c4fd1d1d56a82c9d67ebb77e3a9d834ce1063226d157c83b70670927f8fd81f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4869dd99207b81931c5efd61180bc579a9035691fe3052ad7af55c4b74bc397d56fb4d5d554324b9468cec5052;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103a0a971d5bac1474d978cb20c1edcdadd3e75e5e38bbeafb62a7172868acf207f00a1dac4d6852a18dc42b55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18e10a48911ae6fbd72083e6fd94868944d21cca6131382943c22c3013234b1ef88003ad9cda8415ca89f7381dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dfcad0d15c90bcb2cf2c5dfcd456e29d8ad2a3b5e290ed91bb403a68fe9b71d48b983e0aa079e6f9c8d4c0aa24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149590f13b0494cb1655eeca4e400e57e79b8d0c4bf2d8f20003472e9e043c53a2e306f35edecb21962b6675eb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf14acd8254c777fed2b1fea8cf9383f01c955d7f1209bc71a66efd41867a382dd981beb9c56656af449b12c02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd678d65229017c91006a31002d81ad9b87d52cd9be907023f2dd2e15acdcb9d12764c5fc6e9f98f8fc010c1b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd79fd989d39dac60e4f081c1b288a2326908eeb2b5bb2b896e6cc0f06ec0c6f49f900b3430bdabafe216925179;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2ea3fb98c445da9e37bd61f7b726f06d262e67c50c583b18c8f7332717ab77e37b57144f4ca46303c1694a5b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1edcae6dcecf03913da52a518342e3ebb7ed5a3aa68b01749821eae426b59807de0163a11609fa740b0da706eae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c516d5362c87e9f0f2396190ddae208e8c03e980e12321cdd890273fc33d749d36e0ff49b096cea9082ab47d5e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164099fcd143f5e0283c3174b204af430c1da75b33ff789d685ce08d4bee8ba5866bf4f3d94b68785dc94ea348f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16477a5b8bbaeb7a6e7e06e9f072c471afcf1888de6ee69e6ba8f638a3628656ec7776f045da535d445a678c9f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c977816fa9c25b72e00b405f271c60f183fd69d886804edfcd4ef8a23f10d1781145794486769a0a8c54fae26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53d2ed28654104fa9ed52ad79bdd746a0a65d59935effc0fdc151d52c57372a67f175004f2aae7b04f78d4a62a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef07623af32236dc888dc7ce67af9c3183fff33cd30413477a14109fe293117791220c33f684697ae33edd8f20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c215e01c6e8481f270a5fa9a6d74961756ad79764866f30beb52f42edea72631eb4480aaac5b4475ab6d64d4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2ee74ef6dd88b32778a45e453821f6d6b096fbe702330cb8b86f4385154d898258c9de82e3c097d5e6e4eced0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175e51a4438713ffbdf50056f46f90e7477a17ef0aa613a68731ddb67bb51ec504167d1c6d61279f9e59ba866a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f3cb31de47a77ef4c7923461129513067a8087af34bef1764e28e65a05fed62206eb5f45e0d300cd6123ef21c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be843ab1d19f818f97c2690543f326383c89beb2287730809af69ba058e2a7a8e2143abbc9c73337d9e6560b21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3278beffcd38c366a98fc826bea4a53590e5d0b843016762938ed31635759c98921df893846078d6c5947370ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15eece0596bcc38f20f41344f4ef4f66685188be32807f5c52c42efdd478c794ac79f3fec3f9d0816422115ed61;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1559ad01e8d3eb0f007a8c4b027be2d65a0f00cd2e09f50605fd19fc342d8de2c33aec6d0ac6811ba935343d32c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1605a3d3f653201f4f11d8298a9420265d2fc408cad204d9730864f705641f88644a5bf72894efedb16bd90cf74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e18616d43ac374068ad78af302b44a348297957bc0bf0738129df374ca206096ecc66590572a3eb627bb0f47d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16409c2efe78903dd8414acf09fbacbeb925ad8e1062ac57477e14973153de96081c8f9ebedfdbf81a0479e75cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28c33b8383207875c9ed39cc5f1ec875ed0ca68e6fd031739dda5d8d8f3b2171c8378c80fb593426df26f125e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1914d6a9d2e67e77962595ca9fcc4d5902d62ebbcfa3c349373b66f32a2731216f951d0244bce5a28dcda478483;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf4fe447fdf86b131c8f6939d58fcd49f50662a1c7488cb75d84b688e726effc55fa178cdaf1fc005e967349bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h531eb9dd9eab7a5c73eed925c8d7f1e09d1b5c8e315f4b31ad667f2c644aa583275716de38eedb11090a096482;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c2edafef7653a51c27cb9dbf1a99f571adabc0b1d517dd9ecf0c1528c9f5668020ab9b33ccf7cfb7bb90888c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a455f3e8b4df3fbe8bc2d2016f1c95bf7c4c91d97dd8886792e7b9da5a06b460b4e589c0cbf0df6dc0a8a73c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f5ec5ba01b7b3af91732679735f24a5e380b0f58909fd57343c9248880aede5917b9bf6c43156a6457ccb3bcea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1134203734cec888d9f82429cbd53f3069f48f24de6b224cf80f5ccbf69bccf31cc5ead3f724f9a189ea562c9f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4230b8688a4325f7e7bd0185a01e4fe237928a10675c6ba619e5fadc439a16d6a6ce452a2263c535f6e9eac6ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha95a71681bd7566756c0a55b9295b48fb8c0c05f3d63a706baa99ee1b2da551bc736bf54a5d3947b696491827c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ae8497bdcbc7a1bb9ff103208ced69a88463964d852db34a2a1323740db994aac837195698ffc24e9f314bda9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35f446c0571e950acfb5ca2e296c43c215af91b7a5ddaf6dd8de8ae67aa0b5b43f8cb46843d9db82f52aa92460;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h263a19767f54cf9ebfb0047e555150caef9151a9a5aa2ca3a83b72f5136a99c641104fdc1bf54569c19cfdac8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c95191e4ef95ef2a3636bff1d853cd3eebb86129446497cacb78eb2e9e9e45f2c390ef4a6ad079d9e70f49612;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a2535c1a1b04b8fa2ae1c11c46cbee2643c00bde9a9af7ec452c4a29db28bedaba919db1733b8a94ad1e3daf2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda7255491d7ae05671889402c480da5544f67f7db32d7a41d39fdc3f00e44affcc182f2fc457f0fcf6694da0b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128d8e1ebe74da5501d86501673dc8ccf09321ca11a093623298803cbd88ce78fa899b7a733224ebe6664b62f72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d01281c576c759cf8efdc1c8250484d9b9d6a2bf8c8e91c7acad4de7ad819caad2103cb9909f63f7d91873b85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11dd222ea97ff0749e5fc7e78dc4b5b4bad17f565fefa7a2f786e68a2639f1e9ef8bbcc227be6c472515680a4c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f38658da71454108c0dc48289a87e4cec43f417fc2e2aaf861ee16f3f53f3ede0e081ebafa72e3dc7abbaae67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f785b96cb1d78620414ccd440865985a0ed0e289b1734946803b3cf82b51a0ed9340347dc58fc9d960ba3a42d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h699413ba6d1c673d1d7574bcd589de085ad49b0d2d18e69304a95e68bd0f19f4e9786bff95f6d26745ee86f3cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9fd0e0b4587564eee22cc4e188cc7cbdaf9e43604fec5fc291c6cc16264b3390c85487520c94edd99daace074;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h566332f10f6c220a3b90bbe93c3f1ec671bd9e984bc4236c9ec56c19f0da8bcb91ebba3428b480b23def3ee358;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7eb641d10aefa27d4fde15905a514cb9158915dc0bafa9d5f5cc65b9af218e0ee531f943e2bd79027e627e47c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4db2bd861fd82fa4dd23dbca822df82628ca6f8a156542bcd0424dc2ca42f290050f95eab25aa4d227285ff296;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heef97454f82821a1cbf916a18f61e44116c96ff3aa22bb2d6d2b594f6468552687c1f475d41f4617b84b8b18f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0e68175548fe3e6aa8a1b3e81e007ec1fe971d0d4db24df02775e5c6d6e8c3562dc28d114bb61a9ca930354bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62ddf51910974eb4916e6a416339ea46493c5c5319234032a34d616a5f836ec4a005d64d942e08e5b4ab718aa2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0a3b1a896ebadd3537ce66d1ec77794d0b71153747cb2e03d455de9b5a8a9740e7c3ae0304629eb06ce2df124;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12f66f1141cc06cca2a8c5d11224bfbe29988bb5d081cb599c5b2ad0f7c97eed5115f3cff83ecc740a8c612744e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb06b015a8e109645256d56ad412dd7b4cd67062eaa6000176c3bee956bb50f47590bf684d9764e56cfc1195ffe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f0ea79ca34730af2e32edd7b0894b8c65b9d295d0749ac202c0c58baa502b0f28177ec7deabb5a3e6f79ada7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b9151a223f3ea146551c682acba0ae8a050e7db8ead3e700310e66b410048ec9b09e3212e12618a08d60dd19cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170cf7e42d0f5d5ef03b34501f3d41fce4ac5dc821dbcfe80e9841334b928d544e6f74577fb352cf6642e193c84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a05d736b0ad30baf4b9783b5836847b130403e6de67ebee0fd353c3c85a82849dfb68698a623c9442720cb92d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c6f77cd12f7d1001456d83dabeff732a6b60df2eb4280e63f9dcac35206c52a0a3f209465e1e1cdc28058138a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h56e7b67f73a9dc7dffa4b0d8a0cbed3fb86da946ef6dc4a59e6a4ce2d530d660fc0799758f8a7b412247d02b7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb1ab99f6ceabe868efb520c4694b185c8208babef2d1eee3ba50a5368cb9d7d151ca5715eb6c515ab590183d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5c35e1711093d22ab8448d4f3e32c51c2a195415197d97e1553180475121dab17051db1952fdfc0d1cc2f53c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65184d3585ea97d204b204e705ab2593a9c1000228e26d89c67d16403082f05e48a1991497fde88e8cf83a6802;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd3e7daa75f2cf45a20c5ee1e19bb5d2b16a73c60552258990d33c5b3a349d071592fa02e206d18a6ab4a0d7b4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5f38bf7be1a7d7b374214ec9f87934461d30c38178a71502be64492186031ca78016da00889caeccf470bb6db4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f433c6ba1770e7f3cc31a0c60c1f19f6afc3da763f1d9b22a63d7dd6007fee5be62299c4ec0615fa2e04c0aa51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha372c46449d37613f170337f68f98cdba8fd2e6d7d1c6d27910f6c137e7eafe86fec43a0b744843e55f82a3d85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac4d47504845358d1ba16e9d1c05bebbc42f05083310eb7988b0f55147a8e91d5f08731887b80c8e418c251971;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf294837ec56850f29518e630bc891bd5183b22a968b5d816784e0dfbd1fd2259f450ad09fde89c2d5a8a311b61;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2854b0195a13d459f0a781aed2443966697f3443bd87990039eb21e63de7da87e2c174410fc8cfee6b40a103e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1392145af46234fdbdeccac3d18400a84f82745ac01a6311a80badabab93630771a69ed64d6fce6ba43c51281e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d3d607f3900f8adabd7fe87d49f6c0f0aebe1fe7311c75f47acd7b696c9f44b3c7399028c2656c126e2399869;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h420200cfc3713eecb959ee3f938edae0144a8362b985d1f75d2262950b28efafb2edae5ae0e9d67ab2079375b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17eec1dc7843b5d2cc5c6db6b5450ff71e2bf55717adf290a0978f93533ab4e76b51a7aee7a9f559bbd39d57c3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1367af4314303096f9b980b6bd491fbf39cc18de7ca9e0245f44652f570549aebe94011558438249411626a225b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1a31f2e76ca378bef45cfd415ece7777241dce63d2abc7788d428ca05218fecae024fb304f0dde7faa5a30c53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1de207d3b27c232510855426b6a5cc5f1b75a0350b5e9f105320e1d8e13b9a84dfcf8ee2db733f9ba1a8cc442;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha82f594d945f55b2fc22e4ed16f057a6117ee1509b191d9ec8c223ff065067d0d3bd8504d85b6015cccc55b84f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122df89e193bdf954d4b99765b4bf1631251f0020fc73e32a70a1c600b530a9899dcfe83a3755988c9d93f17dc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2de7f8998a617d20bedbe34e7c29f3fdc49a21a861b69b6796237e50da756e51b1c24e2cc1169a22b19d1e72d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha0c45244f611b1c5aabd2be25f866f18f35c8659658625533eb55bfd9f2d216a6af0322189db5cb7e6b0ee9426;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170ac7184dd6e6e5d6e55bfe5eea6f9bad93164e65ba1b515b5cbb09bdf6fae49b0569266fad87d0c742e6fe498;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11be4e138d9eec538321a485c828bd05272edcea8207b0e3db183db9a6ad28aadc51bb763b4698ab63bc3918322;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118881815719074ee418e1e7a73515f9bdfa1aca2d77f543996d59f6aae9542bf035f5d178c6ee2f32c8d93ebba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h102b705dd99273febf0d7ef5e42fd5ed0590bf7036fd0fd0758758e8563056e1b12c7f971afa906145cb6e08bdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112837b2fb7215a0f7049f94ec7f9f81586738524fa0112fb4deb64f8787e7a23421050b5d02e50266b67362757;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac5a0f6e869d2d1897083130e4b75a91696595abf73da43c8ab3357bc8a85ada92575f185963feaf67a86e605;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b37b012ac9c760fcd48f255a646f6a63ae0c0b392a5182b13057f28118bee376f62a907c117b5ed5e042f796e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h979c6928631c6ceace04179acf8f3bc5a82c04bfe718deb7e9270d13613e35ab8ebc452a0f8daaac894a895eb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h31ca7c60df2eee9ade0f8e3587eba23e08330715c8adf84c0f7b14f109884a81fffb48e3b3139fba87ab8861e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b174d1c9a11959d57bdbd16d7167a64f50fec0dccadac21827411746df3b69dd6c5938fc60711a2c576b62bd24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ba0c502a101fdd39710848d2f872668ec52f041220dda9129a46ae92dd9973cd3cf99ee6ff375cb644c458b65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ce35518f2cd35dd9f614bc14814ea2bde0b194c37c17ffa145a490f22546da3bc09fa8b4ac38f4bef2aaef481;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda9fcf7f0a921dd32d38070425a49d1281722f9204a89a9c14a7053e31f0b816d1377f7de424b2469856d16d4e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf12937ef8753c47c48b775ec82e1679cf800e964ab863654f0d876c070ae6b6c5e1c3b37ce6567d389c0b03d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7384837166c6d13ebd3117f21a3110e65b44abf764f633bea636ea5c7f51ac88d8825a1d3c755c5ab5ca57d5ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6464005ccb3a3885e204dfa5642d8c4bee3436483fbf93e142803fe7aaa478850da7fd6dae0bfb8dc7e563a8f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194c31538638eb75a251093d581c99e44bb8df7157ab9de91e94d916f7d47ecdfb8933eb091d9617302091f7a13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca1107df82ed3545f26728d47ed3ba54a8ecc9c891c11e7b3ad4f127b924f7dff14ebf3f95192979c219df955c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122d3012425c2880fcca1b07250ff7cb0eb43318bed5c9c216428a6cce0573be83a7e7dbda652d86ec8f66d4d74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf8f64c04eb5d77645bc2a2482ad65180b4cb99fe81d70d8d844eb6a5467aa2f45aed3efb0b6cf9fb3e9fb2ab5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114c8736c881a8619de0284b17500329132531a66cdefd011807c7d542fcf7dc3456a91392d10ef79e04243071c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7324380c5f25b03a4b3dc4d921c668c96d74a594a30f6d534fc634a85f5f47ae52137d66a433bdbf3bfaf0074;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3eab1197935c76744c62bb52918427b2a7d7eb01cb0eb9e9b83930fc9d3cda9cd9b37eab1d1d47ff4c428c03dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h101cf8f346838ac303a87876c9f29bbee14ca1dc5239082b0b7cbc09c0ce2dfa900804bd808ee0c476d8590ff13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hacf8d4756e3ce60f31c1535997a071bf9a8995c26e016419ed85cf2fae0e875548c46c61f0a7dc57ed656d8d8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dce55b6daddbc0672689f4e4b18e1a3857a487a016be24a43785086fcdd616c423ba1118568ec88b1c3cd6a4e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3c41094ae25da0c29e6225448dea1cf05d2175b9a44ec1a55a79ddb403c7c5e01815adb6696f6a246a9120d72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c691200977befd1df495e291c771d9468aef2581ecddf660bf7013a899668bffa5402cb9c1c8314cffa053c7c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e47b4089233b45a4b86fd60d8943ec7e4cf6158a1b558c605a4ef7deaba7929f9f9b4b24537b74400c34eee79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12eac3cfa634da29b8c5755fc008f867c7cbe992b89f3972fb7d3befc249644da8a0691e1be6716b51fd6035b15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec39bcd812bdfd16754f89dadfa02c9a946610ef39c4b91b014c6976cc9c4cb95703c6bf8f316e64e50441d89e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcee382b3abb03ca41212f8237f6699b32c86c23dabcca343bef2ea74d124e575f85182b637d7b20b40e456df32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d28bb9074f5036e865f6177ed0f9bf7c6066687416ebb6f5f7e6eefaaefdc0263531fcdb3b02bc2d0961c9bfb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3209d4e57469b5a75c599b50f612718da40f99182d49dd8d8541a130c313e31e5f615a13f21fcd7f2f917976c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f05c1ed6171b172d47445cc11972f0f853f753310c00c414098aabf1f1bf012f7fbef4b06f069a316c24e713c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1569e2e64a283fc1dfe8b4b9eecb61a9b56f3d2b8899b8478a51f46db7aa8450cb3774d9aec02d2f644a4ed727;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cceed4da780f18999640bdeaacdea94c5a4f838ad29dfe1de38022ac4ba970219c13c8a225d138bbc294d786d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3448d5beb7bef6b9b7730136fb88d4c22c7963b825ccc1817b13b54500ae8ce49aee0333a5c9c22182dea66cf5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d94da541a565b17a45095f8e2e7084cc572f0279127caf929c36d92995bacb2d90c8191578b2339e1d2be911a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1d44430650d3a1e1a98c829ecce2102e8b6e402f871f3509b3164ce5e5c3c92c6d906fe6571bd42cfbfc46639;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6a5edeec1574f7a7d1d21fdabddda564691756df9923dbc4391730edf3aec5efc47a488773494bbc117a54498;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf89d13b7df77088962cf6c75c9745b6934afe3db3c429c5e91115f4fbe225f85aca13794aa4642b12ac008c25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcac2adbc304c5f13840849a37dab3ba0da1985a1f462e7830372d6172b7d5874c4facbfe62856f3620a248e667;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3ad3e75c610c953b69f9e1270a5848cdd294069594daf10fef7b43c244360795fc8158cc06f0e5aef4b6841e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146b536e6934adcc2cabc7d17b49a54c244723d64d215bd6201d1a444e9d426cd5ef6bd437fef19cac0296916ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he19ffecd4f136cef786a6a8d8de9411fab3ddad4c2d9d30d0b993224b5aadcb6f1e63d868db167ef4c1c87fbc8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18094f3be45d0f933af2cb35dce0d6e2ef682311e5c9de6ae2db0c1f7e8e64e7e7d30afaafa9e1105110df44ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4c52f7487bc3d51eb1cdbf42194ed46845c53afae71776ffbd627ca81a16aaa4ff9c442c599d6142f8fcbd45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7bb8d5eccdf7d47207288158c38e501ed133875a4cb290e28c877f6299ce1d85fe762b1e2f2ca6739b8038133;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eaddba2053687241a592892e151c9f647a3d5d5d50770a9a90162e26cd96b2eb854315d4bfb589842d472c3ace;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71378667f17a9aaabc6819473ba17bf11e485e7f1d71b0c59cfa96fe15d0f56b362a9c8d550b966c052941c1cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f8bff8d9d1394ee3ec80c49f931499fecc7effbb0e978fd3d3032505f6faf4609df6ce8ec58c21d6d244854f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbbd704ba8cc2a30d8796992964b50d42df1472780bc164fe3081de4a621fcbb68f3c5379f17c3583e4eee8cb76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d78b20021f74318fb5e21c42ec3697321a52ad2ade96687c0c5f6eefa6d4d5d31db2fb2cb8250ba4e154ddd01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b28b30bb511a7897daf81cf8beb35d905187004f2214f7793681b0aec9ff75d4f1dfa94ef5cb978d8d0f99a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc50c2f236ea2b38a807665e953f7cf9b89ec4329e47e11ff7c8a9319e65e92dddcde6cfca1ebf74bf7ce4285e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hffb9637dd646d99e85f3af18a35a7bafe9f281987778aef362558ce50bf84bb75dda459e1e1915dc444d60afd3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc13e33cc1bc392aa2bc5cb3dbbcd9fec1349d08836b16133e02ee67f385a5d303ec281f0a0f268d53a84f2372;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12f772eec025d920ac760539eb83b2469a923f12fbe14f7a617854f90b8f7c8a68afc3c8e6e44e8c883bbfb2f61;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1baa3a32cd9dba16d4e03d8c99e71ace0fc399868e12cd418a161bf1cb6220469dd48268306f6a04ed7efcb37ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ca95f45c7ed09f40235bab11585c8b86debc657719f2181d50526a20b256006616c4d533d82415271cee34dbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45ed2bfa2dce3789a51f825b8147528bff5c1b8d5f79529cc7514f92b80ef6a014db8b29bfacf0ec7b4f5fb968;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hea1aee514a6fcf6955d16b4dfe19408e6b196f33747bc663737e62a80f72be20b8717e1d0f38ff1c83f05882ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1532cf5c8c1204e8492a407a1e86bb4595fa865a2410c3a1ba727c3378983bbd7558a1adbe4a6ae8a28ea0e6ef7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6de47dba60fac55ad0846968274f8a0a14ce3eb514240b28d1b1331e7418b8b092f8611df312e10007de70fae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134be5dd2650c8121832bbbd4a0cc4443221a43d61ae069e4061a22826fa2422f820624e5e3d1c5324ae0486a2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17fac3641e5955d32b94540529e6dac6082574de82b6d479c863cf734c317ccf69e134e4c7ad5ffc0c2dbaae001;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b9b2b0ae06c664108ebe483149babd1bc6bd6ff7933ad1d6c96ecc6a41b4834464c2cc4900ca93ccd2565039e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d7ae9a36cc52000636c6aaaf5d15368d1d09504b90bfe26e8f5d0e4b085ac87bbdccd2f44f651d56524eef0ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99bdac8caab38bf1936ea93d92717c12d726b2fde1116ba73222ab122566c39cb05048b7967d0c4b0dc8e2069f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8deb5eb415241def49dd481019c17d3679a3017335fb1ce96d6bf75bce862ccfbe325c8e4c6f2731465cac7d18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18091b8beb7c9a83344c3e6c10f80e81b4241ce59ffed61a0e670fe5f0ed71fc2dbecafba35a2ae3490501eb5c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99652d0b47a272fca43912d305555a34c8411946b79ba2383ae40855bf47c09a8f3ee67c02affb06f498cd72cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1637ea9a089f9ac091c157bf30a1937e819e9378e35925dd6babe3e7ca5bca187c706b873d39213a3e3c5a04ba6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h44aa22fad3af1bd79e22ef0b831d1a074090512aea26f278bb3cc7471b8276dab73b77dc5d52fe85e97edbbafe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h135007174f551bb658dfd6520eb6c7beb1be7175282cfbe36f644c8f8188b1fbb1c6b474260a7cf87d1aad3a845;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1180c2aa7c8531e2669bcf5675cbdd51f3da01ade25ea14a8990fcf38621498a1a3c135f266e7806965c79d0146;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94fff47a817bc7667afb3472ab78e5b7716e91acbd5277c34271835d42f234ac4af909426fb92344cf22705f80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde0cdb5439b5eb901e27e03770c00afc17dc61c525fc833f0fee808eed50423fa7a151897353a6f0b7680da2a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70c55dd3bedd5d4795cf9d479c3f181c923d3f10f8427131fe42e3015614d332f0af3835c18d08b930eda35c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9b5a2f7b889881b01896048f13870d8763fdacbae920dfbd7b2e09db47fe421ebf4426823bcca1c882cd938d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e68ccd188348529afb7b13cc3a37f0b3705b1b3544f03cba24d19c6122043036d2cbcdb467e073b865705f7f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d0ad19a6fcf8d7b55b31b5458ae2f6425ba45794afb5837cd44bbc3af3ce34142709e2081b644aab29d477bc50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d04717edea0a7dd8d408ffa81786457ef4330f596fea14abdfd45f2d21dcfe3bb6bb89c5b31a8fa09fb153cc1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c55c8135ceeef532ef41ab626254459790e61689190c0d9d916d56482e5953405526c6a30c3689f623c5c5ec94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2494e94a05e9892b9ec0097f7e50c7a1ac74dd8d4076ff48633944863c19b059ab99bd5e01975b6f67738ad10d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6e2bb9eb2cb13c9150309770cbedee0a21ed765d9e3cb0c4038e11d69b84c7c3485dde1c7153ec02eebfd5924;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fca404b4f50ff84c8c70697eea3bea606201be62c6d854da1a400a61f3d65d36030198eaebe8dfbf94f87b6bb8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b9979464e10dad7ee5f50d07bcebdc9e2966bd6e537633d374e0bb229c25609da4a4a94fda71e04084975c6e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d6590809906097d5d45db6ea9b570ee8021b804cfd1bd3ec3b9b19772094dc00f52cd0404755f1d56041228fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe082ef1c8d74608cf88ff49d53d6219d1f4f64238cc0acf229662470383ae11e54060b335a53d189f2eccbff2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae0927aa9dc2b367e966207b0680af3879cd5688ad0ead61bf2523007732f9afdfc84a8e72a4d40824169830a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc991d94e1f924a40e04c8c5258a44125051bc0142d670732cc8d415449afc909ad918f1470620c1096318c553c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c2b6a2d497ca89fe4dc084e1bae7c321f0d8dc9784060fa17927a364888a73f03e7f31ea051ff320848b7c2c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc872cbce8437884d511212ab841dbdb6ea0394683d0aad5e2a47cc849e565549da0dbb3f0c669182ecd6aea465;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194e5c7b274b4553c0818d6b2d56b6a81d8ebdd20683a3df6ff2add68a00638414834ede0dd911338983d65add0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a13d2003f42c1529be29bc9a7a6baa5225301e265ab33a99a07a93ca6e0eb941742f0c8467daa4f6657d6b2512;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5582ab683562555316a7385432e3058e3f1ae49de3176e77d72bcf8d7cfb8b32732a25dafd0a181e637a259d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha120fb7ce89c9be59e10ad355482ac846105d5a4e2564bc31e923ac27d5e347a7f1f6f64ce65b71fe6f7f151fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2181f58e001c4f2b541b23f9d0f80226af4d6cadaa0f3f23df1fb81e6069a46566630784a3cb774f2967b2d3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af051baf0a46356be52db60bf1ec169214d1044715925f9c3e672b0aa09992d25d29cbb2716d2239631bc1f62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1915e4ff457fbb01e3eaaa9ceba05037d2ec3ff5de225e605b99a8a7f5fa387cf89d7f17bab175219e00debf46e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha0befdb7890c75d5fc82e1fb90aa5401ad60256d578758d3b942cd7f9168a1eea5e1aa33b5a82fe41ba4ef181e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcdfc22b23efa4e23875867925a2ed77cdededde2e09c88f19c1ad39e3c835f6bdb6b1f75fcb29abcada909fdc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h478bb9eed739cdbd48de55b662df96c451c18d7adf9cfc328bb9bd9fa370e9198b5bf7b803ab18b0de373de05e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18aba40e4ac6e5145e9fdffcf171b360a64e693c74aa45b25cfd47998d8086d06f8e184c2f343cd23efc6da3a05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e037c6181fe250655d8f87caeba1bbc266cefd19f4d3174e066c9797b26032aa5443956ba889a667bd99debb68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1533acec2bcb7dcb3e31b328a530f9aef545e7e4ea9960f0883cd08bf7ae72032be804a1416a4f0dcd2338c85d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b2d31f9b2e1240e720fc593be3863e9a2e2a5c7551b00fecc11a0768156780e8b828cb719b0dd8d22da8057f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8b1563751508b389ba7ebca6b5eed4bc801cebf588e7213bddfdec8ee3434407caa64abc6b3204bf0b90b7dbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hafca8eba012032e3f42d7c9726a65e099a0270fbca985e5fd0213c55912895f73357f5ac9a3a484f3da1393ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12070539343668e9b83cd280ee9bceb848e14a638857dce3fdfd95a3f0623dd38405e6bf7fc0a051d44ae8112b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b23bd834b82e5f9d6366c5e74718576aa9f6f625ee3b7222f71962d590874dd1bb51927c1d1fd1938c4b974a2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca059eaac62e6c5291033b074a147f17a2381d5cf47bb3e20f3beb8de42ceba0e617d670bdc1c57ea923a81a8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9559224911459ec07e99b405425b9d15c2440eefe5f594cc772af2dc2966b7d97c523687b295090edd2099edb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13bec7400019663ec79d91194aa7ab9225bd777495b2b8074f81a407319d68251a7076c706b3305af57f17212a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f46eb7f9f7f00b4e92f1f7f8a5094abc4fdd3251618f2a464195d428601096ae2fbb333eb3f6890118e05abe9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had2b8fed740a40741a3bfdf48f7121e8c73390361ecdab49f52d5566c22b035f39aa06b7ebdbe0e563777ccc2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6573e2bc6b298b5e24b199ad1f3e187a55776f02752666a7fd8be8780181ec5f5af3a75e3508f869b0c02cac3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a22cca5007dcf47091fff3a35f4bb3f01a8874d4e99bf3c06f4f8647ae324254ed9b87de28da23acced21cc34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a0ad6be38929a270d20638bd5f7bdabc3bf4b994d791f99391f3807269c247a503370bbba20c655bbf76cff47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf317f66ee889cdcfbccb15cc284db7ee5f8bc989a222fbda80a791743c579acc5d03fc0128ac998ee9a3b8225;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51341d705a13ac63c32f4806a981d8db753d5ebd2a02a14804e5444d3dbf0ebfcdb01fd9562e0ad469aa19a3b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148240a747f9d949c421200d80fbaae5459b5f4684b7e515c5a78c47a381c5114a909014e5fc371cc3bcd434c47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1902483cf8809faadc01eb58afdce55e24cf8b0d851bd9cda2a1c37e5a25461aed83a489f34091e8a26855e88dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b1dd0fa0544c4e56492020899b7e1ed9dcd304982b49f4083792d07778ee6eeb978d9c61579897ff93dba0193;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cf19ac8bcb89384caf9513370fad47d93b8a4ba4d7a58608f0e02e4f786424a556d9d7b909ec627e46511fe7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4415e028c5d8ed140761a7477c76bc9f94bf6ea69c2509f58179c36471e50d7fd88a57d62c70802f31f3a4decd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5ea541189a8f5b0ae348748238ff620e942f445f6666162f87139e705442ed3b80392cbb50c950b118d06a4b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9b324d9765ffce1294b2d25dfcd5effd4f9ae99c20228cfb75748dda40e9f77becebfad3dba9cbfb2409f94bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9d74edce6abee1f5420e1db8670ee2567921d58ffd78f51a1c0fa0e5b9fb9f74287b4527a8fbf8003582971fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b5cb00a5a8999f8efa5ecf443a9d29c169b48b0b7e98a3f1c56b8c1df7cd37e8d734b1918bdbacdc8e11269a97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bccf210cf9dc2af8fb412670b86a2bc5b18e55da7f5cee3b9e9104e24febb6717932c519745f915e84bc2ae757;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b3708d54d2bfaaf1f238097ed72289b6fa8143455231624c74c5c5adb6e91e83e67e2d0bc39c64aa9c65f954a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125f40c2035e029bd56dc151e78901299331f3d5a1929eb59895c4191f07de15ef2cc8c7b031af6a9523cab7ee4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d176ae74eb2b22659baf8c29dc4ef287dacaeb5c06d216eea7188d1d5224205ac82a20497dd303fa408af8dfe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f67e6043f3fb3115e2df3dcd340aaa4b819ae57c755ec88c63053f2cc2834810ac790a7623fc223c4eaaa065b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc8da45d404f0741608df786296aad55e87e2b2e764ce0b1780a0b41a01760f51811e9fb788f07ad212e756dad2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7814ce2c2f71a1ca5c7d782adc70f8372eae8271e3b3d096e4e16a9ae4759e5c9330a21e436cf5268f99f2c46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c31dc23c671a3d23abae65cee36ca6242e588eeff3f2c7eac2c22b5537452d346cddadc9e3b9c2edb1c178119;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64e7730ef70de164a0d460fa0e3c4d094570325fa6f387ca10c98857dacd43a1535baa0b5c7714ca2c74c652aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb006b3a400f284cd48bce3bb4e783aa0ac1f1a42b7a618129e311a2b729143b2702dec38d7720802cd8f276662;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76b792fe2806415aa7a155df1a6a0cf026e6e6e7857c011824a02fb0bf76a7ef7be6664e657b32a7a0dfeb2654;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ac1fd7ac75ba2478fc59bac0287442bd55a3dcc0e63b54adf8b92bb183c91fd05902e7e86910554bf94889b52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d5c029517cb980c93b35805bb3b67c0facc2885cf24211d015f98c723f162f19b7288fa318465566c935dd541;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29d80922d25e7f776fab03c869ea965c7baeba134a2cb79cb472f4b819f513d81893dd346d306fdf9525297f1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he563233e375df4e1c88a24c60ed3a2b85a9a321daec92de49c2dc4b27678ef51eb704036c26711d018bae02576;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h173c5bf0f94d538d1e40624abd76ec537a7bfe33b9d06200affd47b982cc57ee7ed472cf353ac373bf6583aae96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfa0ad77c2570fc6c6d33f05d4e51a5988ad315341b786b9b57caf5de0a23a8af25cbf8e1403c4cc7095a881303;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b5f8fddaffadb6c3a14ce69f23e29e2526e257c7986ca8e229c74b6342d2e25a430bea3b489f77f6dc329e1ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8cd149d920268df1a356e4948139794e45631bae44417bcb248dc08dc50f2ca947979bcd344c4bed626e24cfb8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba911da6eb8a4db37a4089d59f778b8321a610a6f11624bbce36fc8592f7dfbfcfd8796547ab67e3bf0efb9707;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a8302e27c45fc6c1e1510baa60a702cd194171123c1e1eb70e464d4262438f800ce15dbd815600cdf8dd24229;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha22fda7c58f8874d36e1d450967b90c243c1ddf759966c6741bfb4eee4639e30476021aa624bbf1fececb7c08e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26db1d330b5063fa8ffde7a49f3c3b9e71134155d539d1301cf7cb43a07f48a9b655538b21b9e531db6dfdaff2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8da063d65a8d2a5860e7533062026baa06538048b72d63b12b8d25bbb0fa0e5e8509d2200a4d8dfc3168d69cec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194f1775e8c028d90933b26898e34599e99fea1f4189894d695630444ea136202b69edfbe8680fc53d6fa88d3dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdd73a6b8b041f52161e60a48eb36cf9622ae355816f95ab07a09d2fb1865ac150d8c203e6e19dde5a44091b08;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a06a8389f4d36093e5892fce82caf7f35693d4d748bcc36f8863754b12b0dd62bd19bce95943a02557e3ce6261;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156374a24ddcd4bbbfd8a8c92b711f9946541d91d7abed27e3685c5a888b9d45d6f360f8f6a88457f4a63577665;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc8d971211d8a946b810c658602a25214ccb04ac9ec79a2cb6b97f2afea14b0325f08f20a247626616f677fffec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cbc46a6fb044ae1f3c07daaace5c3313e199eb64ebb790b6af72a077068d35e6b1649bf3cec63f68d35e32f67b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he78afa63d8e37a6e33a03dbe1b19efc1759b3999b91a06de4b3ba1deb327efd8e430d4575d5b088036bd315449;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b015451ad82d63089b0da3200f88f3e417f89621ba6f8cbde9b30b3e43a94ecb7a557ad6a2b9cc6ced1d792136;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13318cb2a4bdca42b759b095ffbc047886d3a2362a9fa4f7bf84341fcd00fcbc8598caa1f661340aae978afc785;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a5f5c2edd7b19489fac6d618ad6cda244bf9724d425416d88697c0d33c2d923c095ff7e3039019c403562391e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdaf63c847124e86a2e9f56e7dd4d15c4981bf4ae551680740e2585ff7aa75021c572427fd487ec23aaa3924377;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2b2b27feb9a81d676c7fc63328de8888cd72032d34bf68d5d468d4a669e37375fbb44eaf75dbd879092bc835e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19995f26ea7fd847dac5b9b82bef99b0dae2bfd0491b906ca2073c5d7eededc6b4a6d9b1f2cfc7c21b2bd04fc5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h775fa1136a0e777530ca787569ebbca4293fba53962a25d985a35c4d14a055ec04d1d6eeb3ba8329e246ebf50c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b299805d51425d3a7aefd9e4123da359a3b00f17dd621bdc3c81d0f362ab02f5b1c2c13599f66856bfd86ee283;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff322429b9711a384ed470e44fac89e5e9dbf1bde2de149d13604f9d70ca6b533174eba3e82a1dc0d74d35035;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he89bf94fb8069219f860624013ab7e9d58fa9633a626e4f82c30a79c601e4ac8180ea3b1149483997284df9a88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb13c75c1a75b3be34e85a2a17ddc0b8dcca2bb25c8745e90517e5bd4b9e4108d1ea7aeea5ee7b6f8260cb2681a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c882f22defd03cb0ee31592abfd8075997158dd856a1c3ba22dbe129b5955f6b53748c0d67757aa3f678a4a14b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17de9be3de678762d50340068706f3b35c49b2344fb62956d6f153ec49721af08b0b389c4ca4f7997b549e73d0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1dfb2ba7fd691f82b42b18c459436369fc4fbf1f67808097673578b3059706a653044f164ce1e09a402235116;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5f28f1ad503cbe3e496aabc692275e00123b7d1ac06af724b01488ff2392e9d88b1b299fdf23dfd75f9dc7aaa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc1d63dbfd27beccc35454f5ba0e6922deb93c1da7b80323605a1adbb87ce9a66a2b34ac554de31ecb36060ca8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89b8a0157d67e8e51d06803061757b0cc8570ce9bbea385174a8f05ff1eb6d10eab7c64fd2c86fe2e285ab8e18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8dbfaff2c8990e96bdeaa24fbd256607ff08481ae1e64d99ab6154cadfdea11fd91efe801f2ce734129632dd7c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a69f569b5ceccbe56ff17f7788e32c50d4e5487573cb58c9e144601bf019e06a9286873fff54c173e99152d7d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4cb4769b8470d9ff7aa96c25b66324513a0712ee910ddbf1e3787a8d0d95bae3ad48ab39b496dfb8587704f0d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h145ee3e62095f738d7a39291e876f12a75f3abff8e924f3391414f9279f907f88bbaa05f6a849eac122fc7508d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143cfa09034da31506709b3b55b2f8a81372af7044bb40bae540f35f5cbd685419502e73835340f847d4e1b16f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5bcec83189740fbe90305532b2f55496c5d6e109c981731c7ecef4a3caed31469bb8b80bded0751cf1cd1a8837;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12acb0aea1f560abcbdc14b684689784927870120261fe9a239f3fc4c71482bf70a057ee414f629cae432a77f8d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hadd0ae842234a13aa494cd7ed5573ca47b57f0770f0d5f8b998f24e757bce5f562b98549812c47d8747106c847;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9900bba25748a73f1b340856992a167fff5bfeaa1d757d8369468e0c7e4b776932dc8a4ab51253b6a70115fb26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1476267c8ea381bccff2d6df5a855a690ac2d9ac4c1537c37b6973408181077fc3597b2b63186d134ad53ed7237;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8be9f835bc3b3172b18c118016da5cdc091889155a5bdaec78a8a35e99827fa83266eb88efc715c45cd0147bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c6316f06d887d554f21912eeb43123fc7b20b1eaaab665385f4d797101e932c752fb6b53dc6bde86236590f7d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16345195d816956245dc19ee12370b2012cb14e30fcfdfbbfffd313e9b342a393c84334c0b61d9c952d01ff7424;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc23197ae7f739e962e8e1b83cfc71c2be74265ca08cec67791b0dc472e11b330c7807db058e414163bf792939;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9fdcd2d89b70cd2ee56d049f64caf3e255a5ec85269b29e861cd22bf4bdb694c09d2355e6ee00452427f4a0e37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c0be5c5f47ec76ca786f4b208963cc504c2bea7925a54b45370c7bf2a6ae6dfc81b60483185b59638ed6015a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ee16a7f544a3dbddab717e3a5a09ddb4124f51ca7bed5c9267cc212752fbdcc09df2d1483cdc95f9347a035a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c20da6587a360c90910a4bf93a6bd31f246151b943800849c0501921ad12e099716c2cc13abfda7cbc0e76ac7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12fdd6c9bc52a196603c3713563c2f9dd11165d7dd20d89ab78026a775b7889907e585e54ab6610ee119f9dcc02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5f66f4f365993027268075863ad22423b3095e9b12c85f97c049327bd7c30e3d37e78d9b70934f4f635d0aa9cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16287946e7c443f887d32cbdc78a1c153f3b6cb7a5650d30b93353fb223e3daf43858061d0caad2a65628614560;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a96a910278f85d9f5900178bfe68ed3785655bd533a570525148d22ab6184c019a7c4ea7de9d02b30ef7a6db00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12af2e62c3908c081877706910980cd0eeb40e58a4fe39767e473704491a5aaed4a54ab171aa4dd0b7f732e13e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6949858d3cb67503e1731e16507a1f28b9e6cee17cdca678e2d745e367066e60469a2bb20767fb45c0c680b01b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16e667593a7eb981f23d914fddc705aaecd84acd0ddda9d25938321a3df1fe4bd246cccf58b2b85fd1eea82e783;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fffaf9bd9fc6a6638429dfc8999791010fa4d10ed96e1d20661086daeffad4404ea56b989eb89aff240ab3cd07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7e3ed203697ab8ae5d7adcdc1a75b1cc0ef89a9836beefcfdbbbb744d01ae699c2279f9d702c6ed7f17c0a9d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h863933cd43f34291c0f210536794c977aca2434cea5ffeb43072a4d37220a81d1b32bf0bc9906b517a2fa8094c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156dbd3db0e68a913c1fa3a72588491bd15ecd28701af65c7fbf15717755629c71e14f5307baf274b0b0cfe2c1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b0acc3a3da2d59c699f6d299684357701fef53948406f52477a037e45dba7b74fe703ef885796f89094843cf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ebbe8ce93ebd6d7ac4aca0bbfcc1aa22b7393dac3529fd2cb994161b55f01148df227f250d78666080acd4579e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he36a26131a2de447878d4f6a64e8734cb96b00a9e2e9717e03a2769b042c81716c39e4f38b014e562b64599d22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfa5e57c2075fa2c3f6dadf8d6ad3ce76117874eb90903f0cbfb5b3c921f5eb195be41c014f0148432cf2d77296;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175fd6981ab3bba68daf39396d504501bb28cf3c478acbbdd34e70a6a947a9a82b961f07901c6175398ef48ddbc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155d067c40208a6354bccff90ded0e5074acd858bc3cdd736ce930780fc246ba043d97021b48c81a421c1ede122;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1accdaa98095caa49e97801c6f95bfc3edfe70098b9c92538e503337a0cc00b25f69e6d6952da98c4b059f90f4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4128f9c2beb22944d59796b5eb4836a6f22553ceab7af7db42324c49ef02847043b10d9c7d49e99e74e1a62c87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161b958ddb831bd97505dc23c7d5380f3df0ea28e30cf4af36222257ead954e887a2e9f07664fa12e7e148a4620;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5cc3ff92da941f95301f279daa57025462bda13deeb7ad77fdeaa7fcb19ad46a03be5078b9e55e7b96b86dd737;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h105efc48128b97a061bf676c59b666a806b8477fd4e59ef3891a4cc7bd1e84d4e994c95185afcda5e315ad0302;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb0c1936b28d7f2c41ca3a76525a98cbc7aa1c3e2d7094e1fcf50afdb33b614806e51591f31040a0ac044b47ef3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e4c9d38df73a47e35da834054e579a8fa70f1feedca7a295e2e9601d5ccd675d3f1e357636d8ae28ef69ed0e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142cc110e0822ced887388588612aeaf144494c4d2d83ed9d060506ef2768afd18ef3ba997370a4732d57b0adae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h321ceb639f0d1155d928065f28b2bd951809ca8e167837fe847dea1f0598153cd1ee9f9599e7f2224a539cad6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b2a9d9043151a1847bdda59796ccb92a0e51a6b355fd549af3856eb1d1caa2818674ad6389312d68e9bd178f24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149f643159eab5a9867456babf2c997d897e8093bb096f99dce16c90605d9bf42549b61a2f341bd2b8c4b6001d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h618d28e181302d2e91e479c7fa4bbf7c39f9cd88cf4e5cd4ce8206c31597af38bffdcd40dea8c5417b1488f255;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47e79e83c7e3b35f271265c7930281d17e18dea615c821573bf43fafdd52d5c7d58a7ef44c801df94fc237018a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1044e86b8f9f2c4074621d4282d80be9b57e285bab3aca4bd81769b82c028d20f75077e2d7df23a88eb155f271d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2aa3dc9b89dda1d82a9c02b5f96b49a1f4bbb79afaeb29c948d90fc6825c5b986525a0cb47f8a8c2b8dabde46d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18280dd0539cbbf67e6f306d073eb18ec85e47eede137fc800d763bce6840b2d86b99b00553860f4a786ffc478f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153cf6389b0fe9168cc759c784442026adb2529bdcc9a73aa3c5ebf7f60db06b7981923ab04a6c0239a86080486;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c542ee423af5e29366587199a699a8fce9c2883226ba9e552e8f5dfc4694e78e1aad96bc99c58ec00bfb86f3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172a2035c228c66c2bb19c77daff458a5189c4627974b77a5ddb07893eea84023d3fb0923ce0dcdc3123728a597;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d400e4aa5d3292993dbf9e38e9aaab9832656a8eb53231fa1c8f47517789169dd5880f0ceafb0896f8b707e83e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12111b655ad53ff87cc6e4771e241b2e3269bbbd95d01c77741d764377af64ed88f3368b3c4d2ef7a8fd9f16653;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f83b0fac565e61106feb60a1a64b1a7cedea406ad1be7d8530731838c7fa6c6103c26598cf8a51a44f7ee093f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcaf7a37f31f070e0e9f90d86d93fee9a28f280562b2078acb30461cf0ffc876f86689b6751a20cf779b27b3fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb8d2a37900e96696c82f6f8dabc58d6e2a821492ef37c5f071378fc2be4b58e3df05d406b9717b6c08f40ef271;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ec5a5435f213cf3a10401ba8d042bf728398d322b6b3d2bf2439c96c1d58f0b5d68606c2acc87c3afa253474e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h340e3a4a9cacd8357a78dc3f3ad015787f6305d2f8ac668910afb791b3459b1c9e02d78188c91bcf3de0791919;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42e41e171b5584214080b518cabf74c250320d6f299d9d7d2e0cd237cc6f506534f963055194b0510df3ae9fb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haaf7e10569b10164c0993e9cbcf255d616827f845d194344232f8db7118bb378078bd5fc961daeabf400f31214;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf78a3c0019aadf4b15e24b832ca7872d846a36962faf0c3002d79d84b7b939d46443b80f735ec19b2331aa6a35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heba6ab098b46d4b9daadfd89ec60af3f0ceb7647aae2d6cce2b3e780ad0fd99611f05440733a816058552aa3a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185df7622b379127199c6bfa895b890ea435458d034012c37c4a7e0dab21964b8ca94c497eb8e71f3232045d471;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c3f01d99ea0f3f3adbeda069adab33f271d80e67b055658689ea186ba88199291ac8ed0a0c2f0dc6510716114;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c9acef93cc2ee5be43500398036c0e68827273decdf022f3e884dba174d0681c4b68ca35a9bbf56be762fb8c81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d70d483b5459a4ddac731ff7e9aa875d447e7901fd149a6680cb6a1ba4328f79dd9a1ac426dbefc03e8cc7ade;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1169859848cd29bbe48beedfa5622724cfdbeb92a7c4a9928ae5802abbc29aefa61e95a971ffdfc910d2565adb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e86195f035725a4c7a1f295514357b284828b98feb3d13c6b8e8e872f9c7f790096a732cf60b536e8ff1accf1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc8f7bebbe3ca02771c09ae1d773217456b8aaff7967cfe76e4bf58a82bd7225f6176a862b43e818e9e417165d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd6a2a02f8be72c9c9b321888633615c3fd480afd9fe405ce23bdc964468271df0174d5acec279f1f191940f90c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e0895d1356d6ba5165c7ef3ea219178c449da061e464a32a540a2e22e8b7f11f35c6a381d89519610aff410a4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda77a6abc150139832529fd1e5a8da89b8ec602ed4c8d29216f306583cb75d61fda9115c3b5ab0f2cb801ca028;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcc032adc08fc26d407a5335d0302a0703767919030a0ed576613976cf60eb151aac06d4404ed0bb44ea467afc2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107b0b03d8d9f97df5024526e02a807c30d7ac8ec1ac44104fdd21e17cd25cd7f296d7251689cee2982d6c2af35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12f5ef7d78b43cf4a4747c2bef8ba286f20ef6f6148b3bd8383a575807e5e85c5d8be802952cb0cfa06e89cd0de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b6123b9ce0245a757055293096d321fb79544f079c0b1ef2793a5c5aee9a70e2556eeac6c6c8524a8f9ec4fe2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f331f1e8d1652fc26ccf06223bf51c204d3a8a6bb800700a8e0ba399b5d620ae656aa7d0335c1f593508c3060;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c4f1da938d3a3fb5c6bc8d7485cdb5e0603aa137d930febb1e6f9d8a5d582723536fce5fc785ad86607e5388;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ec2cbbcd581539d1796fbce9d881b78d7e0c82419a1b52d48a3d828624018c88d3bc27d9c7c37288f5d8bcec8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha04d1904ee9e5681fd6487b2f33285b2036451375cd23562b64680eff74ed4b17b85a7d079752e02e235f2811d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17105ffeab11ed47743e52a9bf7d4da561c8db13e2a80085400018c328896d6693281fe59fd7071cece24c37916;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h570478a104ca293039a7c6a1b01403898df03f6c108b336c6d2fc68b4453a13a86eaca314ee9e2aed7c8addac2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h57d1463379b68e01e5004cb387584a4382d0b2ed9c5f5456b6b99f329e8253c58a77cfeeda7d15fb32876a34f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc70bf14b5defc5c9a1a7ad18f994d01774e2f701e1eaef549f145b0bcc560d9e87ba92bdaff072b3f5fd5d3f60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c92b2ede9d3fd0d715fef347d279c0f4acc42c26a53ab232300d442c7943526b35a134234a5f99211450aa80d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a1df77d1925ab8fdc43b4b4a86799a5fda6d4923cc9d11d7fa9b6ad7115335c774e6a65956f1ee6f0dae321a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aecb13a6803450b7828ca7912f46999a38091d570ba6c3f93264f3bd5834a22311658376724a4db98f95e13b2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a38bcdfc900394a85f0426d1dc7558f13a668f4e7844a0a011e5c3de899678a6557a2ad705caf63149c33aab6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4570272d13e94b75def8fe628b4835eaa50e797cfa27e9c021778a88f5d8d296ba4c9440e35bc565217b2f9a5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9aaaaee2145ba9c0f9eb703ac90d744e4ee932fd6e57cceed385a668a2209af3998d6174b7dd249554b41701e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170180e2649ea77052603998f8ad3d44c590a923eadc871853c443253c3642baa3b811dc817830321c25fb12fb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91be72dd1d9454654071ffe46cb1761b2304d8e38b557e794cc1b2a679695a90420be2cfddeeab17bc78d160ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23227c02d10e81bfcc5a5b1831f85d69fa0f612be87b4804aef93e182686c51cb59e2ad40b0212602218e2c268;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf386589f5bec9fa52f58db0ab7a71a7221adb7413c5bbd2665518aee81a8280c3b62e13eaa453d07c68edd2647;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe8d3544071fcf082b6889a729ff1420f039b3bc3937d2afce4a4bc8b299cc1786c6033de7aab70b244a833a4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97feef7094f2731a3fef39b1d124d8ff46b961277497e9a52e557460da1f931da5f437e2ab1bdf0b40df63870a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd361fa28890595abd5700cb357c5eced59bf963dd46459c720197a8e25737c7cb712207faef6e4c44a9b278a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2c77d04824ca585a27027fe3f6ae39ec59a0b0f4110d51155834cc3850396c2da9b0827f0825ae498dd54118e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ada0305683f5606f98e665bb04c142985085684da12f9a2ef12b31f55d26daa29adea5ffc6d669acdf59207fac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc7dbc168a94141ef4512b9b815ae4542c7ce5eec4779e6ca2bb91bc66a85a70600646eb01901ffd8251956492a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185b8ab1cd83f8c7652fecc5c6f5a3f5c0e96a702ec9bbfc0492ed191b801f092f5d9a2fd7abd0dc1199109608c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7cf26685a7ef652d91135998ff079ca76b01a7a26a2bc9cebe7a3beea643cb45697c64a20396be668a49d3504;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdf59e7c33e0ec742b0b94d4fbd0aaf89797a841adc318e867f8baf665a3d330c3765dbb073cab245c5d922065;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c00ac97b7314c1252aa7409c58221f68959f24c506e6518df0bbdb8ba07d275c6440b2cc0b6bd7b013fabdfb4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38c2c8a57cf51e2536a5f5b0ed7f347fc1910fa5c07d7052291f477c5eb246573189d3d75874fd6e0bac2287c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148617edecfe761b950835b0058dd197c606a23b6869f8d5965a6bd27c5879932a79236107c226ae9e8b4bbe250;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bac90411931ff98060026f5e70077a4a0fd96914665435a59f0d16072c40046d014584cdffa072cae7e1ad1db1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4478f933b7827cf493dd7627040a07e45359094171e8a67d7785b11de8388bd5aca93d0bb131d45bfc7a73f02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c86329835c060b8b6db9f33a86977cb13958ce221bfe6e082ce50aa0486766a041cecff21b5cc1b9e7f3f44d19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h471cd29b6fc97f3a9ae204156d62fa5dd99a5dd873ec7d9d3a4d051f0e6ef007cc067efb0a01ea57b76ab2f34f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141db9aacaf09eb97221bd9b0ac94ec66fbd4a68b91f6a5870d4cf1fb1b080a79d76dc1970f90228f637dc46bc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35a09e8294c8b5b344c8e23836cd3b244dc3bc771c0fb91a7558db4b7d9ddfa2c50b2fa6e9aa56e6394182afce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93320c775519a91dd2c96b4262a730c74df98ffd93e158169f64715265ea3f320c099113f5b05df522243a98ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h754157ac441c8944dd244e9e00ffc95b4c09b8d3b3c5ed7c84606dc1fd595b87aaac40480b66d6740e75c486df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb316eef6138351a64d481206225136f494c7532328907e3f821fc1ea44b270349eb94ff1e788d8e6d64e3e269d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3945ce3739c155eddbaa2fe4dbb4b0ed6db1d6d522809041bcdc6cbcf749e9b25a87ca8fd348e6a09b49623831;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff07ea1433b9550a0d4c329e81462790cebdddcfbb14350c5761322f7a9e795753cc6795377e9bcb65282b022f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17291bc66a3389876321c3d27a3f19956093aeb7e7c21cbd43ddf49cd8bea7d7fcad83f547ea88b5fd85df9b49b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb731709dcabe21f5979f1c38472b70eeabfa1c2b9d51afa986842ddeb804ab5118466a25b845c48942e70ce5e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf33ebf435f3fb5355a9bcecca117fea38c79736c87b02b0329590fe5a92f6e9a11d579bb79dde8e95e7042c439;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a7f795dab1cd7140e93d6dcc1bc3e2e18f4a3ea8965a25f905e388993e9349d9ff054984b4e9b68ce1bda1ce6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5dcdd56677e157fd740375f155f661e7db79e6de482775bacd7530fd2397c06b131745b110998e3f233e00659f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6337f624b8f1c8f135663d4f8c84e087d6ce23c976f2833e8b85930928c82b6feaee1f03eb2f94d3230f143ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h611471b16f403a1b6814c6bb588620155e760a834a69daee2d1bd127a725328e331750911a6821ffd98132cf9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2b0e09333aa60d0789fe72cf084d8e2ee6f33b8ef1ee23b6c5197da349957bfe4f1394d998942f2cd41078fa8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec86f04c2e0f155483d51afb94cd96e3923997505cca178583b61b9fc3811cf61165f95602c6c05fc500918b88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a0314a0b43b276381c946f397fafbd0c342ac27ded4679ee2c1f4b873e730c73ed7c7fe875cea993a51a0375f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4692cee6cb891aff8bb7760a5ab78673541d1fd90fddb4ea2c347c69ed9b8d45653a4b4d62d435754d6b4effef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1785f65d4541c7bca84b46a2b6006f3862164ee2b20572cfc135519880a3fd151b3800fbcf7a7e28fcc64e1c73c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heca77201ab5d44fffabfe09416856c8641612d23a3d8722090b46261497b213f4807d23f0541b340ddab270897;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178e7e51bdcd5d3d3fb353794d6077fb1e10b13d1caaf49c56e001bbd7ba1586550e68811e0f08cdc6f877a4acd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17defab514f06c782592dc100fc2f0747f2cafbc589ba6b25f13c509eeffe37753ae315f4432d5b2e689c5be216;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b7d79cb9210da21e1edd7afcfc1ae8a4e25c0bcca58194249a4cfa938eda5cb8a8b405564acee84f297af767f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ec5c962ab45ea81522808243c024a1cc8689f2f3ba6668f2e549c28cd6743efad82502ef8e039f42813fe100e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154cdda618e7b8afe676e53f5be8426e9028f7c939bf5c6f89dfbda30e1ead3c50ac4bfba9595c3600b20f46a29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb366b5ebfe3dcbadf33c82b6426ddf9b24cf12ff3546d5860bbe69d7edc97795f49ce162a71d9ad5b2adc46f33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h592132cd7bfffd8f0ee4e8d7ddb3af25c0a83b321839d3643cf8c14eb980d7eb144ce119be2a5f105655c71606;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7eec6767b1d577c1acc0bd97ecc5fdfde16a409986b8b21300f670c5ea9a6346c0b1f54bd7189905ccd08323cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c7e63c6abf5734e542d0712b1186dd2a4c2530e27cf54cddba8d12c061244425da9514e70aa716a37ef118a04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e09a060a9c9ab7f79c3a1f202561c997cb8f44d03c7de06530ebbd69162d871131b736dde53d7d441a15b7e3b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae7647b76d1fa3bb355aa576a45db340695386644e9da167fc7983d159a2a067059eccc002f4388ad9053c3222;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7662642f3ee752bcc9186ef665783639380f0bfe90f827dc25dbe951437786aed83bf75d4b04aacab67982f12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he173b1aefa19c8c19231b6750a8bbe465f54a47cd1f0daa6388049085b59a5d0e60304bf98392c61b1d59eed5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99f1b92adbe4057dd9799b6477c8126344fde089173776885381bc571a7d6fc9ef5d6e586db04ab83a8fdaba6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hade4007776e5b1b9507c15fe50a8e5272a4183c489a95dd6e2703789d3dc9aa23bdb93fae11435b3286c9c893d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c6e4e5d50bb6ebdc18cc64658a7965cf1f6fb6e8556dceb388e6ddc91a1f768ff74371230060054dfc640b48e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heace3fa7207342f54dd36403f3d904e5d99b870bb31b79f9d99fe218de3d9cf782da44744e858f61e1cf97f9eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf57f5d49007251bcb2746d50d84eac137233442011ba24039afc082b016b72a82f8248421aa98057846416d58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3203af7136a64398e52336e33d858eed74144177453284d13f6a05dc25653488814c7ba5faa86d9ed97ccbf84a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d817e67229ae1e7b290e5ac232bef8f235766d48cc0126827bcd489bf3afd29fcee4a9aa60481f5c7f3dca9317;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4de7094d9776ecc92cda4c75a7bd8336a867fe0ba6081f5cb494415e5687e2f598d7ea2ea681fa7a9b03df7aef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hec45723a1bc9d9e1ec99c98ee9112312466495c4923474329111e78b59d6a95efaa55c28091c62101f3b7c89c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa66a05ba95aed445299674228e7b10b63f4885479585e1d14d31a24cb8319fb598dc4b6d14b4faa20b868c769;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bdb25797f435f9d9705a93d34a35048dbd30ee6ed15251b899dc9234c044efd0d9a7f584855ec3e02f79face49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf9398ce1b7dbc1a54cf5c1a19e63513cd81a5f02d372d70a00018e1fa08c47e71ffdf48d39f777200e26562828;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc40be49c1371f51562566f849fb0c1020a5aa513402e571aba1fd79255a84b210d830980a52f85c74ef5762390;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2be9ac52a80ebc8deab1e524bbe3871a811c600a853094882a6301978554b09e6b69938661c30ad4a1772eb9e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111213407b929e56fd4de1043a2ef8cd8fcead1bbbc1a0c5a5bf97f65052d11b5f022213157ab536448cfc14d77;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae0f8d5324d5baa4cfe81614c5608de97e6d3e838016edebe04ac524da77680237af426b611646388f06a6838f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c1bfce03bfe45eb2ec73c23479e7a557f747808e4d83689a48406779f765fcdaac14bbcad7a5d83f0f1778223;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18e94ccee804d8d4d1ae022b36e2adcbdf276bc6791feafd4b6c8859a0e7af399179033910c3ee702f567f8567e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124a721d870b4ef719f9a50737cb8295e8977e49b9297dc891a68db3a05f10edf3bd267e05f8c14ef3e60683594;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c8e412ba3d8a4b3befd20b25760a97fbea053a3ae4595cc975cbb7e852e119736dda38c09a412d2e989822d1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38c9c0487b151096c07e3b5eddfa4734a9eee7a1e8ea2487edb2380b5105ae64fa70e31ba478dead79c133fd09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2fbaa730ceed2d314ed3523e69d42466cee7276a48d0124b79b000a5f73815af74cb399191e35bd98e84fe1b0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114fcff08930009659e9ad43afcb339463d2e0dfd7bce533b43e62979e64ef1e827c7e4a5ce2167d98dcd6b0e4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1754e578ba070a227f6c9048f7566fb925d6ea92f4ca1baf4b17ad918661b4ee82de082c2028f01649008a9ca75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a23974b5f262a553dadac1fb2a9c7496040da9184bed8c9f26b7d717eef1ad70e2dff3fb8faa6b966cb979aa8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15386f3485575de92471cf835f70e4c78b3bbba2e58c40099204cfbe915faa97293b1261d7754b0a41757f720c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7262a8f39c25dc27a37cf6b8d9ce174b1f615b74bde4611146565a3b9c35500418254eca754642dd4e573d9609;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ea73d784e5792e66b9616bd18c32ed195a306ad879c02cb2d6219212642cc009167060b0b08fb2cfc1177674;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f232948771d7180b50e2902f5ac759e8f6ef94619e79490847b9c282a78bfb5dc1fcdef38b0ad0892a1cceb22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcaea2b285b1d250c68d55af9a397898acad17d28b6942c63f562fdfcefff333ba0e95795b892e21c90962b1e0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h537fb197cfc168699d62e9781d556f25a0c5ed1aaff7db2eeb46cdb75840a50ce27e4dc13bd2bc930476ef71d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb166bfa84861b59d71d0951876ffe65ae0d3e3fbedc7b14771acecdbd0aa4da3a73581476cb198e6b053dda47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e4f0e5703220697bcb75fb5c3b5326d2f6b25b48ad7c55e9b1d57210fe670bf7666b4ffba67112ffceb47d373;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f80dcd137812ba3853ea66ca9dde6534d98f8277afb5babfa68c658675df40395ac959d0c6ad817a94daa5c04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb306ef07a9ab9930ddc671b6f9fc7306207fddd57bef1a0dad17997e289fee0776a968b7ee71bcf4aa85b5924b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9729e6c780945b3149f5f495abd32bf95e5e0b0f6f437cc9cb7009799f99dbce2e3375cec97a13eca384a7a9df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14461c5716f9bf0eb7264d7a05b83d7a6e10cf447f7963914334d73f79d4b29f0827038226d21a0357fe0a9fc3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e37a7833e391013a3ff1ac7b4a4cff8375b6ffcf4b083311da761505851c9a520ef64628a92ddf37dd1819fb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19238f5144ecedcc2200ed109100a83d352632d27dec4731ae9280208ee41c5a92c1c62980a0bb16a414c4d5de9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b1506dc064b72ed8829e0c70064f5117fd05ee0b85f4a19bddc68f8eed71fdbc54b4848f173db034d00ac3d9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c89841b909b5418b652a84cfb0ce0fbbad79ff47121cc7ba7563963914314499a5614eed2d9906da76af86ecb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d14224267eec3e818bbadd308c603874acbf8a1d0864a1a46e64a4d5f5a124b01e953111a2eff88e96b9382c63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb6e2e428bffc0da9a3573c2a23839cdace31d76f8604989211dd93cc96cdf5bbb0721446794961f8db6d15476;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f4ace22bbb0d22941b71d3b2465f84df76a9dcaa145b40868f668f96ec38a3aadcfb8177f5564dfc73e61d0b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1abc6d53caa8e6b6b395d7694021e1f43e7a51215d74d3b9ae44fd4907d5df4f6de88636046551f5a3f1c3c511f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7ff11f2ae272d7423f3532a566db298138e619fae371fdd04c0f8e15ede42ba507cf2b15bbb7b40aafa32afb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h177426e64dc43453c4590fdf1e58652975a5c6d63be9f55d39caffc073fbfd965ef22f8e9a971fd1243eee4987b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h629ae27fef50b1df7c391bf89811755dbb7113ab1048fa2036330981782c64daa25a9ad2d488d3f487178d687;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5296bf8ab853b30850974008290aee8730c50824a410ce8cd74ecc1af701195dffc74a797d48489ccc1caf2a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb254c7e0792c407e95082e59196c9fb7727c3574913816efd41883c38ad5148045aa43e81f4c114d4eca73ff7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3e9b087757f0dc37ffc9b31cb06decb39c8cc132a5b2a3e5ed609a5dee460fd70a8d8aa25f9e64ff7aed7003f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88bfef778a22d982c98fe5eae06bb081fc2aeb39f0605937c6b58d5742240a6f816c9d91f6662690633e2d735c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2646eeb7c4bfebfa562d16091e700bfc77d9055686096ba96bf484616ee4a2a4c5bdf9088f98453ad67ff148fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h803d65d7590881201ed1f4a81cc5b7b82be8aa5ae72381e1cd360fb79343c7b6bf22d40a21978f8bcbcfabe2d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8de2ce7d0354cfcc6a58627471062bfc66793416ca9c62b4ae4eadcb12421b36608fd7359cfe443a23f38facc3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136a69c5f7db541f0fc1e75513f1b8fb1b22d42272ca330a644a0e95c208750f7f5e0badf448c677e7d167b5421;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1484194fd3d399b83ab06f0b69205716fddb97fb7a0c10a6dd60af26725af11a7747f0447938e4d3d58fe62e793;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154b77674c373ed112e263fa8d9def2491b0f02e9d447f5b3ef9a27f8f8e53fd9f21d7aeface197073cf2fd3e8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6715b0f06a1048c443527ea2a90daddbdde7a02b65f973c11bb843a146804b77b0b6a308a91cde1d607b6b4e3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h537038c019b60e2534dd4a96d00379b88b88643137e3ca1f8eb279758728ddd18a43d540b6b0e439659e28a18d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a180b7399f685a73ce990891b76499da3cb30065a2b21d09ae71a0504c0a9fd924f9b42c23e4101a58b65bd3b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h960a051f254cb6838a87f0eaca09b84b57fdbe6381ea8fd9be09ab777516d5228d9bf82dc9b7fc932306437ae3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18254d5f753cce6ea7fbc963e625fe72e8cad324ef84814099d63b14733d0e73e70a8aca7c5dcceb4722b064180;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf33611ba1dd536024bcc728936e9e9ccbdcd2c402031772e73f5a71793c32642a520e684a06b701ade5c25efc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0fea67b2a5e75369df2630d83e2a623db93399812e6b5cbe09bf47df1fbca0bf569594017f40820624f387e23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3e3d0f23e5f01a4e0a3a94f45c38c2861a5e1a71ca3e4a12c414ef6bbd446edac489cbbe44c72b85e49e7f0e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82dbe792adf5f71ae63178ffd1fece4d64c28156d9e6e1d313bf35027d9e40b5599680f2e773bf066b73fb707c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fad98d10f19cf5fc99cc4f7cf350e5b597d6227892f2f3d23e891d82693667a6a10516ed5f77d4db77a5c809b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b61dc871c6ab49c47b1061a354de4e50a0aa4825d0fc2d7bcbe025ac5910985326f2fad69249cbec11003fbfa4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13779bdb7d02b3c1e4c287c2fa71fadf0e0dd3f9f4f84b215b324fee76533caac1fd686e49d5a13fd22583e022f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cc9ecf0afdd5137d562d59924414393d4dbade4a9b74aa2429ab28f986c5d0901085f9e549a744312606843c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h49f797ccfb3360d366f02883a2d9bc5a6278778dc4768e9e70bce0c5c91d2cbf95e15b812a4a02dcbcda3409ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee346a79cc76a15e35a04a1e1efddeb867e0de02367ec0e4e6fd66495e24e8143c6f9c3b07fae00e7ad1c714b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6eb30e15593023e58ddde4883c4eac9c815f17445766a21a47019ed19b88e28eceb592732895b5bdc8b3372592;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14732a203ad3a2f57ada2c66a491c0e19b157e9366d47f4c7c35d86e7a2378b53bc3438399309e2cbfcc2ab516b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a8af24afc037c74ec7437ab0e428265e9d32d0afee2417a8e992d999c27f43667dd56cf2873bb9d3d6ab780986;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd961e3e7314084ff6ca891abc0dd565f455483fa5689b206010db76d0de051fa8598ff92d630c0f37a6a3331d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e14a34e54a1e1dd68f29fa14d9a8c7e545efe84e6acd1e0c78ce9d4d737ecc7417dabd92679746e0bd130b486a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a110f67c4017094f1541952c85c7f2643bd46e6ab7e76ec8596642151bc260ee62810871a09e0f3bfbae3b8fdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he907ee5fc43a0eacf7ccadc44ca1f57f9f3b5ca5ae75b846a414e7fa0c5ce75930125a7b9eb267853aacb89180;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha39b27ad20fb4a5974f68c880163c0a424490648d1e2beb901352329d146545be979cf7cbf9811b01b97aee6a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4cf5fece649f8598eb73cf0badc93f11a7eebfaee01221afd441daeab07117331a4d8ea99f9832c659d59e05fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7281e3b2990d8de89ae8eebca2a20bfaa3b766be5b804defedf412248c4c732a6c5ae9902e426e0ce0d56dfab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193ab4a3e3fab3817c30bad6807654d840fc64caa3f05cabc0364b59b2f92b8254ebcd2bf6187979911e3207783;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1142e2cc5e07fbe01b9fa618405b209c7856bbb5c5b644fa62652a472acc0c922accf1d78648619a5619c38b2ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cfad6422589ec3bdb4d28da0aa59dbcfff95763d6ddefabf9fd831ed638d3054da03a2a517ce23a7096d981f32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72db4caf8d17332b8dfb420608634e33c99d64eb4797ea5b8b51763e6e3e02aed0073ac174028724352b00b0d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf327722181bdf66bf449982b5e5838ee267ccdade6fe76d0c0bcd04971365d93e0ce9c7a8753bf79bd702bf445;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h611186889110d3daa7b9a61d8d3408007254496e31368f78e80e4d49f360c8ac73655b3641fac990d261bcb4ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dc70fa0ba504c36c9d0010f53a8de72aa05b41c95908ae4b4a3d356b6250fcccb15252c3d1ca6b7fa66892a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb59884eaaca85831e622466cdff0845be342392ebfe4574b01dc624c59225124b2f48492f740377c67beb82ac1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d6af54860bcc3db8144624cf14bbcd6f7e47431f8b15c1895f0b0a50f602ba0eb95f086a744252563387ad023;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89f67c36f734fe135331f0689b6b48afb1193c3417d69cc52f8c9817f4c794f200890d104b0ed9c93e0833f42e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19862aa44d9bd8b2dd5a68eebbacc230e0be1aefa6ee82af6870e6bf9c2d98b6a482eec61db0914ee065e07bdcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe746c84c6672b5af1e8fe8c94ae758cab12e18dac5e13ec902296a0f577a150ec4401524a38dac6c203a9c8e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9d03aab38c1b9b585552b8672dc9cbba5c6ee5309731fc3931e1a71bfe6953fdfbdfe463d40f27d30575f30cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf097c832e0c714e0a01110228f9100a4790def0dd15e8cc097e873a4893bc2cf95ccf19d04d7bd060ae9ab82a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2cb18af1c4cec681eabde95186fbd40065507ea1b6eda7dd34a363e876043e0efa5b6139d6cf20cc9066818be7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e0b2d0d1e001f816ebd0ccef28021a7913f9c1fcbff8fe7e076e9b0aa19274bc9f35f416dda92f79087a303ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf3983ce53e6bb8d58863885294f98a332200231d22bb01fb39fa09af0e17cffb9fe2aaad9716cbcde34cc1f93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16d1d88b4afb8045e73ffd0240849dca5f2a063b0f57e0f9f85f00015254bf0ae8efedfdcb96292b15335bb7524;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda36b22ba17defca5846e6fd759daedc3420b18a42c3ccd2d62ebc94a26ad60778e7bd874b4ac69bb557c5f941;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce63f5cea8aa7f52b47b7b64061a4c712e32eda06a03c696d71e81f1caea27440412359a9caabe4e280f38098d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48f1d20ec35acff01d536ea7aff5505f890c58de6e0be962036b0f1a883903ff6bdf8b925f755585aedfbab57b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2b0b8bd4ae1474b68b9e6859e19e5383f69c027457355158943bc37a7b24bd62b911a20d8ca15c257b7b2c5e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc3cee69d4059a17b40751e082a6bed76be7d847d3cfe1714b9de70386d399c8f7a1dd7a54d57eb6f81cfdebf1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30c1e3fa761f660beb4d8bfd1c1adc517abc60d4d94a8a477a15210c9bb9e7388db73cde463b89be941ba0c790;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147d8eb870c83238c89d8585ea371c5cb1f51673248e848f0417989c9dd8341d05ca9c15572352e85a6518299ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161a4ce5e904b71e3c5eb28431722bf20ae848aa143bcf0e914596e00456a099d97c32844be465ac486b11ad6af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6305de06db5eafc80947c57cd3b2e42c29c1f6373c508647939393ee0ba2f2f9abafa97b8fc3ed055b8e613fd7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb5f88efc9def46756ff77244dd504f2f1a264ced5490da26165924959f81873a091b1fd418833e48caeedc84b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ea0ed748dc595f28ccfe7bfca1bec775ef9caf7ba9f54a3122ca8ad928df19d0829112aec459c86cfb262695c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14af7b4d70ef505b58fa7f7c75878b95d9145f81f89c427019310a9ed6bda951db18b49dd0a946c302e868ebaa0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75e0ea0d4fa1582d9b32eb5ebd487d405d0008816fc2190ae46ebd3f04843e2e32c9c3c0fea64bf0e1e2c96ba5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h584143cec6a6a112e8a3d8b799bb53c97eb716ea27c580dd20526ca359a5052fe6b58ad2c090edfae1eae5239e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb14f83ebd99e31c5280b5ef9bc93cc664c4a90dfb10fe3f4af1633daf65d5a277e63661dd156c47704ebceca5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c9d250dc36e20f113f003117f8ee94d13cde8e0cc476e5fca0a531529b33d87e1dceb4354e9f6413fea8a07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0a7eb2d9f33e07eb93c31d5893ba30be1568c9740ad453a643b9e4b9f4ebdf15740c7c89dbb4ef0464cc379c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1344ee5e01f10cb5c41b7342daa3bd3bab21d9056985561175ebfd89d2652019f315b0dad2190bd42edfce31979;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had7707eff07dd4e0b96ed8e016a8391f643e81b2d7cff3d71a39ed93afb3aa92182ad6399ffa9b6af416d8a487;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a6916bde8744d4118a5be976b90bb15554edba4084c952145d2c10784ea9f269b4172b7e44dddd474ac4b773c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h587a6645003a6ffd10ee731373b598c5913a5daf5ac6022fa2f68db9b6cdf2fbf1db3cc06a8262c924a47b2bde;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f50c51380247c1e5bcd4f8e1e6c24dc663a8b35d0a727241ac99a79ada84f9b64fcef3bca4114ae5375ee9b15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2af286143dc2be18927f683906bc6150462b7559c3fd505731dbc0a1ad997f2591eba65e52e6562deeff98e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1350da12a3c37f97735324d9d8cb04ba7cad16b36a93b621f6837f50aa72698d7117e0941bd96eb09d6fcfc02f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f5960a40b03205d4e281b6d77820f15681a7e37a0cef1f9bf258bc98cdc6566cc155b6008a472fe059836e2b16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15946ded55a929b935758cb0e23fd5bd68d8ab1a30a0b0fd813185ec0b64b4e8140f80529df22a9276c36b751c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbfde93dc80d6cc538418172a1934ab3c66cee8e5e08e3312710d2fb5339fccdda4690e99f3aab8ebfa7a9d4c81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4deff93c63c4061dd2cf46af60ae84bc497245147e8e2c5a93c456de148b89aa59e93b7e7932b0f2a8c401949a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc005c18ff646d38ea1af19ff93da16d52b2accb3a91d4416c3f20244554bc3e94769fae2a38e16f4187b89cc10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133086eea6206b6bdde4048633afd71dfa6c88f9c83c0942a04a283b621c1e157f2a55ab2e9534a55ff4fce222b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10e5e880dc78c09d6600a4b90b39a948a32237ad3b5c2a94a009112d385bf9d7be4f58d0c62bb25cbe453a2be5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h115263ed11cd591a1c66d5f1f1a5f559193bea59135e62f29fe14b5524db5cc87e3d23f97397f5300b057ed5ed0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e66f88d48af0824d52b2a3937660f01799b5c2e732231e6c85fc9dba21a8930bbdad9c578d3e655467f0d7da7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0b3fe6995fd541abac0823f121e4c4d524c0d19c2350e546991c052a4f04214c222df05a137a12fe44dce2d05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he03340b502b176db6397931eb3a3c9e5c8bbcf06fc8c1be3ddd1f7b21729c5ee9ea2af9d53732da9bc8c453cfe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108659d57d5a91b24443ab125ee33b1e2877f3b2260df962368748f892997ccd1199a83e2201f68a0476cb3c9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12dc04de6fe24afd16f0beb252329bfcc4f18b9589ce19c1462dc93870fc52bd20e4d2c774b26e7613c50ff2301;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a7387a2f7aea8a2e787062908f835d7ca9277f76f18c983667c72878e779a6f2e7e9261a567aa81ccb5f590bd8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca12558ce5686c16e5d9cb80984aed5e65b6b962bba1adab6bb4eabcbe2de2909956afc45b56dcb78c4ae3962e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc8ab0a20059149b088518902d3d4b762620b679f794bf662e226658dbdace7813fb5dd9e4185d0b6345ea0309b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae2149e514e00674f6c0d37ce207d9ac4712c40cfd1b8a1c24fad5c2f5a6cd7467ea42aca940aa4c36956436e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d9779a31eff3b21579666844665cce6187d6118063b4799d8f3b96157ba865f5a4f5252dea7cc627dcd5f961b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6254b59e7751886885dfb6e8162678abb2c106d1b48a7504fd8b595a37b02be122e8afe034d75e8b8f43f11fbb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb07374a8ac48447694eebaba978ee7471d87ffb0570ba199cb05f9aa9b0b06bf56840553abde3ea18518d4d840;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2e5aa8ff2a210db886e1a927ef29e8799b1fe586d88fec6247ae0a00430f75af8bf017307e1f9137757ba3161;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a10986b19d0e82c512967ba23a49fac4e5a2ddbd607e8545ab779c1477b036066bcca9ae1f7c5dd867d5f348e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127291249af70dbe73838962cc7cbd5865d6c5051b004d02ebb05e33e845807e56048f435e7c9e376537a3d2685;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc6bfc122918a593992655c0fe545ead542e2326a063398bf48164f1ba12a80c43aaf50152402a9fd9d8225637c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15569492b434be1cba610f87119090bb1e05abdb2d06647749817935e86bfd7a1e4c558dd12d0d5ae60010ccc58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ada0a9ad953712402f0f0550ffdcea8dbf5a0b8c4292aa03a5dd9833e815cfcfe3bbc2c5ad4cc0ef374cc28b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c31fd67ccf86e05b38b18bc70e0d539d6c0e032d88f0d830e5422f42f4c48524d45ab06e85dd4db6282fdbce2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f6fb23478f249f3f80f383853a58a009bc93247f888990bf89f35ade795e51b7ae9435cd8dafa82e67fc1d29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a101e7f15e98db362000e91b0b7c0a731c665b81e78973ab8c5c14607a56cd31fb89352d307a99e6e157aa0d68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16d325b7a11483d4454b5d8b47c27901fa806f281b2b52583ace254ba077fe7101292de36cb0c898840fe7467cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172b055e5dfdd22f61994ec4b18cf97ae16afdd05a1c92020628ec2a2c12265e1ba175c28ce5e72db6ef8eebd7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ccdca0f6620b7d1eb4e33443dc454e746667e5ef3398984ad7192ce886e94925358718f557e380ade8e893a3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d833d76788ee3ae12537cd4ed8d042d0effa64fc375e724bf7e596056375fbc835ba0dd3338b54d892471f3cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h177541c2ed67efd195b34c30b805074e220db4b7a1d88ba4597f75cadc9f54216f5cc15d001c5467c139ea4f274;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc27132cc9905545179faa912449dbb47941e1055915e19c095064f83d9b1f5d1083512e3f150336944b517c225;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142f116229c514fc87d0459169404242e11e13ad6798e6a035916e2a9bcebf6eb9f505067edc882689714c7b6fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f1db46dd8bce74685c35cda59cec32e0a99be4622ba120a2101c62819643c4add2da3513a5a8356fe9d979710;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e4a0c74af459a5b5508b23a9a66ccd0bec3204a5f47adeefa2889cf0893ab185bed531deadc6c146ca8f857e16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ba1d895f503ef5a78db8349e1bda243be94198907b516bd03869c1d39c73b93a1dd0fb8a9c059fed8e34f940a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19567ecc7bc7352e35c91c4e3fd35b80043962e7c1cb55ce7889412e21888dcd08122354f52ba3480986c63ab59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a19ba9a430bf0a9bd24183b39562db94e035eb746d2b12f31faf664b2a23983fa2451a4fc060c758eaa40674d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1acf831e3e2d9922e4442bc9502a1d13e3c5cde376b9a7b43e849688e8c81f0bb145c18ba19ef650a4ee79b1cba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a75897369e15a483cede80a5f179fd5a8cbc9a51a66265fbd3b7f38567baec9de351e079a4ad6d1dfd2e076cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdddc604b0ba21f06566dcf8035bdc6238b3e419f75d8a87bdd56b76f719350a88cb60c058c4e1b811be28233d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h942658c7f1ce41372d9e2162fa655d6bac3417868813630d799e7473d92b6354c4b96a6b0a25cca60e6d3627b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad7708d417aaaae84b335c8bdd07be4f34ab9cb529ceb2089158ba3ac19940772ae26d2153e11bffa50c7320f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1801b84862945ca41fe1727801372089cd55de2dc05dceb36887af4eebd08c8682d5ac80e4f6e5a3880e0cabba8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f21c090938f1dad796420491b00da45d2c32743c2ebef1e212b13c18fe433a43f8fb6da83a7ef7674b3a709e6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111862c4cc8a96c6cf410b2126faf5d713ab077ed884884ea4766892c4dfe45498e604b7764d1849a67162fe489;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc744c63de68e1187ea896e302ad8d0ab41a030a128554d549bcca4e734946518c51bb2f84677a7592db2cfe14f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1965a22d0632ce6f011678d40b08456da916a5d1868f5c0a064880ddec983d07b8d1f87c6872fd4f9243329d93f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h169b5b9d4a8ab18acd5e81c60111ab33274a28bfb421dd2e21d89191430765ecbd482de1f5d899603cb74fb0367;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde7d2035493a68076326006a6b09e544ed92a570ea9ddd4f389c2cec751bc7f71e2a7f438312c3bc36e821ce61;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c45d2b8ba90937d58133813607e65405c4e1494e868c6a1b4d24c7f7dd1e3910730af14a12c22f9c0cfba1b163;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10edec19cdfa5ec4b6a057462ec561bfa0683d334231d6e48feeab7155bce0dc409dc12b68e326b4b47543ff33b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16e8571aa315906c025c4ef9c76593cb5283c91978426ec2f13f3e091847f2768490257b0cf39bda79d2d5450e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1519417de8b4234dba5aeb6076d7f9e1faf7d89310d69940b7cfee6c03197da642aea335ed3b005f24670f767cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9227307a5d1bf615b18e57eaa6981323265a101ed9cca0f5ba5536df5cfe687d088422ff87956b71fef628a1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h269969dc37c3b3f0b31e8e0bd4e45053641a2fde0b990e4c2b45bb0928e7ee5a48e5a68f271ee621ade7deb4d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbbf3385ad817db45b65d15b8e2e2d86f1d69902ca4c6d25da7c087220a3815063c79c1b7db9d0cc081ad966c06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5052d736d1bacdf7ae71866d33d0eac23b3922a1d33f04f99fa9a76ae3b20d59346d6bad80d829cebf376cf343;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he0e1f71a2ab8cd828e7ed2f406398bcaa848d460ae769d6dd27d141c99eb3735e78bdb01e817f8ccbd17f42181;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dcdd3c8991054815744c706b139747fe72d2a9a8f78fd2fa963b4c941c3c006ed92c7a6f898a355969cb9a9abc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2818c94bd8e0022c8bbb7cc2a952c9445361e4fcf9d6daf53cab5be81ecdea1e25878d51b41374d79c825a6282;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e201e30145d56438c2d9e74f0dc9e8deb6bfeb26c2006aaf34cba069dcc0d29e03d51c9d041f54f07db2f8940;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3554fd8fa64c65381637fe415a793d94bc0819b5903cf01c47a819e93adbcddeb24fc5df8257dd31d436b248e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d3b3a7d72479a0695349025bd2dab2942cc877b5328dd7ed8fbd6876a81ec3f25178567f5a7d0cc3b74fa10d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe78eb319aa670b3a432fdf352db72c054a8ae510aeb92c1cd33f383894bf23bb79377b0fd15eab54eb0d4df09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186ef9f763cbca8ec682303d0d6cdd7fa48063dbb76536091afde9a27d670ebc49c051685824144809693c6f256;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1fd05da5dc58098897c3c2dbad30ab7816800edf844ad579078ff86ef34e16f4dd6d8b9b96cdf940fb3977116;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e243b4ed02ceaa20b92aa2c256e0b8ea98b1d337b8b887e8e0675d24f643969d59ed2d85e15ea8f6335642520;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195ccc29fdedf5d9380fa3d4335668afc3a5bfe1134ec227c89e8bf2e8a15a64b85dc93b4fe2ad15e5cb8dc09ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb68b739af03d75d2c2c65be9e05acd8ec2334a723eba8bfe64fb646043bfcc6e7881110dd18f93bfb0b097cd20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d435eacbd3c19c956f89870fa8c303143ce8413b4b0f39973bcc1232a95ef09d8d8ccb1620d3bd0f8883a0ef8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff1d67412fc5c46a8616ef8eb1540ba138327ece0a270ff87c807971bd142dd762c2adcd9e5eb4fc7e16b0940c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7186259b229023e87d27f39fcaade276b20d9d3eb76fd646cc5315252fac34aeb9beb3094721b0c2b318bc8e45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14da51cd4d3aaa50880a63d00d0a56bd20345f229fca96cc1c6429acfcf7423460a7bcf84fd9c8d8f72635475a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc8eaa908941c772cbdff17851c44b8599b292ba6b94f6edab3910bcd7adcc665c9595241da7cd9d09aa395ef58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189a74e2fc1352f429e3b7e3c3d447673aab21a8cf154e1020b60bbe5f77d45d158bb4102130501b6fd543a1cb4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha72b620e544d5e25390761f70eea833adf4fe8134cc3e1c3f75caf99d65fdec962259a5575f52400bd7d2d37ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h402334ffb35a3c99a1f12c4fcb7ccc8bfae8dce0af9e5c9e93faa5188ddd42a8a2526186c17c6f8c64f319c3a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f7d48171ece5f40878c183a3afbec454c5ee4b035886b0a872aaeff6474c4a20519484b2db74f58175dbec2ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11481811d460302afd6cbd8d90e0c092f42fb292473797797fc0357bbf695c822e8e397a0b7711fc703af9a7dc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h92d3c484b968f7db2f2287c07643426077da4a392380d914384487af75fac08a510a1d0d00e05fe08e1184bbd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf28488770ea209d831ef0f17152535a1750404577597cd222051ab66fbb14242fb1422ed80de0a2612affd82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1c3a427a3c2b926325326ffe64c9f3c02ac912cc8fcd08de9f44e9fa3c26df1d36ffd2a56c559958d4877d36c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h86e491dac131d5ea9b0d4c2e9d35faf94f3d0ff77378e7ee3387c4502eaef04da7c8f035ebe49e08c531cdab5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h139001b4edecd87a5b44b16e27b472f6702ad2a6453efa27fdf9bb2bfb7ab236257f40075a41fed513326d80732;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd0f14c25829adf6293dd58ade2aed1280350ffcf3452e9993e2f9c17fb080db60b5ff04abfc7df5e4def5bd22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c9aabcdeb69bf69d86171887dbae5fd05fe02cc9a3b97541c64c93eb388e9e3662f916a2fd3370c19b18a125b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ba3706d7ca8d1970b72768b63d571486673733a0958f15cd4f0c0cf41cfc40a168b21f4acc951094dededcf47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h687d32a5dd8d817bc1b613017e459845af68f4d2ed4789f3ee88f3fff356b0f84dd33a352325a33f33711d01e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h137e683a60f85b8cdd32b27114ffacb508d6b36b342cc4c8d81b5844b255b89dbc46cf74688836f14d9c134c9f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf447597d905c069bb5401ecfe8cc826a2bb1c4d2e26bbdac73911765218592c33926fe9fdecc4e8b4e3293082d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c1fa87d5d7558f83521a533b5f8fb2b48585722b20dee82e03ea63f818722d1c1a10f4e0c8df8fd820cb26695;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163b169df9209716484870ea6e3f6cc25ac26ec189477ca49e1f5d02218a99e5d33fabd023cc30e11218b4e6ffc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34e22d1110be9f6840f8308bcc098d166d47235dfa2f54d91fac1d50deac7fe7604b2b25c96b7bcd826ebc8814;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e46aca6b1eb951a97cab9d218d49be85aa5d3be2dbe7c72842aeae08142edf70fbf69d547664a5071520b293c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8acc0e54c6c00bf2c3b0c4e7d7a4a03e2ed5e5bb4b60d8b119c8f65393ff0aa8996be92446b4676c764726241;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha39f375e0914d2249919f2195c29089a3e07ca6d4022f9d545ba0f05bb4bb84b398efdfabc20ea8e444dabde76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ddac47d531f727e8711d1708454b4b4d8186898f157d0a577b1a3fb482c7f523d64b96c23abb35846906ef0dc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b0c9556e368b7b7e5c91c7a8b69fb3396b9e4043b4247a5a2313799fedb974a29b85a80e14f9cc38ca4201f70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9353eac72edb116f681676309e25e53b7e49916e6da96630e4e4bb9ff153e78442b3f790d43346467c1d734cc2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2f3cc52fe36ab221fe95f6948a7fff8912ca71d8ec1721fc66222ac8ee2d8f9ba83f30836ae8c24b8bf5c55f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f6e0d0e215adc6534e60ce01faf4a4b89297cd20981c6620bbfb6528370758e413d2c155d1fc00538dd39698d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12439e6b6b8f99e1e59af8caea8b66cd2c9cd8fa55a0a0b99a2edaca41772319f46d253e13cff52d07fac6675d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd548e61fd617a76386739e8a4731fafbb362ceb7aeb0b2b1fc510b764e7cb12376da24d48b6a4703cfb3f6021a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b86c26113bb0f4152c77cfc7d7d39b045f9725b31df3c31ae417400c80b2819c5836fc2483973e625a7f63ce3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h171768625b0f43453a864610e80e20d9b41f503c185ec6f61acd4702fc1ada32b672e61ebb5b347030824bfc0c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4823ce796fac7c920d3f7bea82bf902675fd3aab00085ad6d4e7317150bab04c76b826bcb0228ff604321afabb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h655f967d8c0f17b2e64a42f682c6b84d5c922a66a7ca42d4610ebfa28a896c9ee79c28c1d85b7443babb324444;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ee3ad5a08bf6fd2ba8de5d2e6b886fda844d06b7e0ab457c658f9e336070d8da8cf2186027ad83b2efd52ab2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d24ddc4bff47dabbc786a8ff3b13529e7b73f4c92ab54ed63b2b9cd5cd49411d653fb0588f0bddff844b11c86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19365b5679056060527eda771c9ad08b3db2d386b930790c802eb9759a68ac7c86c25374ee1c64f4aa21e141888;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h32f3446d4e6d79333f2d9c56e031abc5964f4d918a6f5af55a0bb3ef50916deaf792c1334a1ef3d11d0f27e32a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51dfdb90736e6d460c00e001baba6dd742f6530b2bd1991172dddfdaef9a3170f2cfbbd44ab7dfa8af60336b6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1183e1ca1195c3201dd442d55fc4fc27f250b6cf3b16257255858e11d08794f5f374835015ea380e6e84f95e3be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d33fb143b0c6f46b174e9b6ff06b0b43d16471f276a97ff152d0e322feb8d69321a0d4a61d1893cdf0461cc04d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1247f2a1beca6831097bd433024ed2233190b853185e4e5bb5a98ad6e5a416c935cef4cfd3558ec1373399414ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd395940e20b0281421a2975dd451b0c7bae1d743627c4735850581f3a72b37fc93e3c5834b06bb200575c5903;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd47440edb98e10e626eb1877e99875f66cb12351cac620c9fb7f83b0ce162c9be3632a4726f225d1050d970d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1adb0b926a14801e519859ab6ac4b8053d03fa66bf60c17028fbeb1e883a9741fa8299d8e10f898364a28afcc22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175fae15962fd3e85eeee733dee5be6b9dc595a7281f480bbe2b118df2fedcfe91a39e6e9334c69d0e50f4c1267;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea7c4238fb7704dd3317cf5960359a23636494a20c0743959cd98f2e269f641ef78802297001f66165a28f775d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he85e345efbfa632ba4b02acd9df7fd4c4792447e022133e7ab00ffe1355d676fa1197a44130f8aa78ad3b0dcdc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8eb7d025b20f7fcb21b13fe7ad3a8911d1901d295480c6e29ff19881cea1a533f50fc86f16529c17b71046b90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178af7111f4ad6c992f5191c763f0c602878669f58cb1a6434731433183fb71f343ece76b8972e32cf66998f878;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d8b6b6a0da65bce4d21f484842d02f455053a6d658076dbd78565749a3960b614e17f863916186b7870e43c4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17daa021bc58a90b4ebcea369be725587f7347adfb763ecf33f50356660a4e6a26c518f8884bb0e0f40c3646682;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd65865700507450d6e9a44674ef0d267c2ea60f9a35ec79e2a1207c902daa3694ce1b0813ade24b81be6c04ca3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h21867210dfa7c548338428f08ce2afcf9a0eb43490ae2da3002839877f3f5a7c91ddf095233e9ebaa724e0be65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c66a5f18c5be2dc8cd4575963de21bba98ddaa3b6be9619d34914daf71ee85fc8aca507a02fbc2a0254aa0afc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14578371b22c364021e86bf3ded12967ca3374938ca782b407e2ed7aaa45caec82a04eb4041358c50424295db65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd7174dc4a8836a7d6747cc6ccb7b079e0f03a70d087c86b1c251d4e12085632620370982c0359461a6bd9e0287;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d0d1737952e832b66b913582e2edb44b6d968b54db969995f3f994154c250a70eb61e437ee54428db3d34e631a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h985264339035582396684b6c750d99180d1dd00b7001fdc9ca272d0bbc5a1bed116f49dc5a2d6a449c4983ecc8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2928c018c95eac8f5f8d1ae6b08a9310f48c8691c71040fb1ce06954e26fee065bae1a5e26ffd8dc3daf5e7c98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3bd958d5f3f2392ee945c717a40584ee46d9b14ddc4a6e4c3446cfa5075623026e57fd90051ef2a5f17a86b11c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd925230a1d31725ae0328f8ef6e3dd7000ac7c4027dc1f96536449979e893e38f4c5facddef159d0c6f1a90c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf383178d96629daf56f316462ea2b1706c6c7f4f8659e6194d625431117f95119b5601ef391d6ddb76f62ed42b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf646c90c83f4f55aa6bf0724620a56e5f7cb3439cad7a3ce08feb18c36f5dc0488066802c502edff7ab203aab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3482c458515ecd0db3600b6d1b3a7faac485c0037bad8f3cfb612c5847504a1b3d51ef680f31940992c127e744;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h109da57ef9b4b58f655694a36827b9061863cf04d8bb543d5226f3de9e26aa9414e1b37d5214c0c4c7325953da2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he40374983bc3c472150625d845a6bf55acb8b6fe87b912588a38ea87c48721c75c8ee34a06b12822aa285014d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e420c7c4eafa8d139ee988a6a42ca2da1e3b73e75f0941c259d4f79b8b7ccdc4066f436e5ac1162d7ebe4fd1ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1b6b187d18f9ca874a0d2702ace76102a8f00e4a8b92b03bcd2d66a1e1acdb54301e99f8cf4705ef42fdabc22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76415ee7020024b9651ee0ee1c423640958e21fc73de1a3fdb5fcfcb02d0a5ade49dbbe974f59ef991084bc141;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e74eb4e11f5f665150e5177e499e32068f45297650300a914159679bedbccf8d743083d483c7563d195874520;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hafad3e4b732192eef8569c8617bd12f0d4ef21a9d19eb830714f100a334578ec3022b3529402f7f038216cac69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd21a0e7785c46ec1f6f3f950d4816b284979266d71f82b118afcd9aa248aadd171620553c02ecc1aead69afb1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c10854b76eae3efb4c44bb5e84b92771cab28f9da3b2072a8e752c10e6b40b370605848e2c90a33b14374ec37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de884e7452f90330dafd3556b3aa4698ab7d2dd291aae2c33a083804d9a383d3997444bb72a7786d6a4b3be8f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h169a38b5ed7d21080a429984dad67c386fa41424398d5320b33239d8d8beac6c39ef536d2db671d1d1d109ee098;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b19e14a160ac531b78373bde39c791e5f260fa9b1c6406be2d4fa53a3046d81e25db3e2e192820fbe0653956cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he646b9ef854870ae3dfe436f32ca0d68287e46a52bb5b5b90a36e3d814198e8952b486185a0681caf2d204ece8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h57371fd296190235b5cc2c4800418aa06e70b6d83d1c911ed90e1c1178d8c1a035c8bdf254d6e70dda0b1488a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a298ab9e52502b74c490154b5a08b43439511583b16cb260612f1a2c1b93aa8b4f499fe0bcdefce373e8a0dd27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1091cde6ecd9e361c493ebe97bec1ae206defadc52821d6a3a7ea5359d2197a618f7a17dab3cc2aa42f45b7c2c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d53602eda47ebeac8ecfe8938854bfee0465b917c0f99b9a49a4f27cb756c2bde5cd0dc61133e599f7eb6fd53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha452939a9b35eb7b32f0a52ee17d65a4b00397799a1d1c34adb57f99e6e952f9aa2edc136e296af8d5bd31a17c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h920036c595f547ee7b9be99068cebbc5c8145f4441aec6f358ed3eddd7aa9ddd97aae289eda6292b36ed2dc950;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb63a5b2b580024b14f02e971d3afee9892c38cbad9bd73f3335d04c6e01fe07cfba52373ec2ed9ffde0c930301;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16da836602ed494faa49284146a044e0a1da7f72a41118c4e4f8b8133176c3f0c52cb8aa8d3ba683157ae6b6660;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5a4eccf9955a7e8aff4ddd89938589981ae6259ca0fd4c49b2575b422de6fd248a5a4dd0f1571ebe56c3902f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ee7bd649d5cc9f930a0ced027e942a7668b0ad6d243b1280e46fde387b717dcfc197f2161e90872630519d2ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66e9a24d4063c8b89f32c3eb45476fe6d95221cc3112dac173fe4fc757860f52e672f26fd0da6f22a42b629e45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc65fcee765e4a0d68925f6cbc1a4efadce28b7b9086d0cee5f3825bc04b9be2d521d5a70033a983c729f12139c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he129ea4abbabb4307251af48d9015216c99855c81a3f56bcc2502c3742954ff49f72a58a866c005875d6f7f154;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142531c356c3bb44cd1806980deab04f53bb5fb8f8a906cff498189dd06a9e0ba8c26ace035c0051afeffa9cdef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f157d0a3df04bd36d53b75ee4a5ca54421c776b2ff5c49a8574f463b214768605c7874989848641fd75251403;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36378598e44318379c16c15542fc01e5e539f39535d4d43541cc7204181a502d16e60faf068d0b86d616d6df87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h295692a823f673e0a4b98b6adf9401cbfce0b8bd03fa696128adf65bc3ea6c9f29fe4af431ff11d4718d6eedc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd2e6f731185912bf2b746ff8a5498aef54c792c65221a989012d9e00bd556e6d481d71c58cd6aeb0fdcd9160c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e918f5e6cdd94494674a93548438d868ba34880f4433d2daa79d0eacf7a6173e3c0f0a985d0477291ebdc0d2d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha6f4e416067adba7e63d43d7ccf46798ca0631cf5a993cebb612277920bd88243f337870bc4902161026b99f05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h843d5db1d6250f587369d21673c8e971b66c0d6bc5370ceb78a13b8e909824a0550fdb950d7bf2f03e655b48ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c269358e15d8735fe4d5173183f3054a038a2fb4a211ba65ddecc612815916230d0ac6ece884c6121a1e884b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141c100c3645b6b6cc9e5ecff3f10cbe94f788766d21c23d7b6b0ecd74ab93403f8e4aa4da4c1fba816a9c4e190;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e047d5fae9de3d345d8a9c6a28ee1314138459b88e4354a73ed310a52cedc3838fb3503d06e6f9bddaf96d1e8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab1464bab7817e750f0974b95da0f7d60f567787262275b8f76d66a63b1a976dcf1274c48c70ef5db84b09a7a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf541af94984b4ed390b7d5213bc1203251ae38c20db420222364df39d85c50cb5958d6f0865c04dec246638600;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h83b7fa8332ba460bbf5ee435a924ae0fe8ceabd1a2ed22a0d175d7cdf8306d3a9c415bf6f3c427787bdb8a0bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb942a390107de92ba633ef51a2f3bb33520e6ac09e875aba32f518e4836f512d82b3f989eddd4fc115398e008;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hafb4d9a0faa0fd7f2974f36fc211d36a4b5241dd51e7dfd0c4be3dc43563a9fdf6f17c33774d243080de1849a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12febe927b040d60823477e74b4ebc3f9a4c8793d60ae08c080e93c7225cf6c1786fc135963b25a5a5d716b33ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6a36221bf09ae4cbb3cf0eab481e8221f8724d95c84ef88fbd732986c0396804927e7ac5962a79809d396a325;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5e49e155747d1ef016bac92313ec6c1502527a033cbc1a6dd7b69373bcb491c989b2920d880d135e234eccbf5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ef9577e7bc780ff879fbffb77cffd8b061ed3c361051f8d743f34298737d121388a3daa4df047b64f0d443073;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h872c82e08a8af135a27844c8de60b1044d41c969c77e027b938c809d38dcf42fadaf932ce43b089462a0c2a3d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18db4d040c9ac10d3a1b3b0a095128aab4da6dc5dc26661dbd19e6f998f22fc95d6b118f69f183de613eabe302b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb83e2c81728fc8e78994fb8bb51fd6b5fbfae9830205f94a304c5e9138b5616d55451aa93c616885b170eedc66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac28d9c20fea771255bd6a608b54ccb74251b8f8fca7d9805b55f69c862c4447dfcd43fa759a523e73a56fe3e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91179b34777c575b87be5153c136b636b30835fb80ef9996ac5127eba0a71683f449cc402adb103e76228f80a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b09f00b080ac47748dca8657626bdf728870836eaf539978aa924e4153ff108a8a76fc084518abb2a644c12a52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8190acb5cdaea7b88023497f4f3b4c9507d5e6c5714fdaf2cee0f1d339979cdf7f75c4832646fc0b699c835cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb310ae2541dd63970c622b0fce40d1d8cfbfa5274813a218d796715eca3088f4ecd20b5c3f13487a6b02f45db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e34c2ecab34887df1d8df2c06c1b454516e85064bfe9483d95c224d186940572262d37ea019e817a0af6fda0ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9666eeef936ffa9275925f4b923cd3c6285bfa7783defa5e6927284c368507b87eb8ac35ff81b5b1dc0d355f9e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ec57e071c6c9707d42e237650d445bdb24734e87f6fee6ec614eb3da40cbb25204467017969e20e4233ae1281;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198cf3fa08d5f378bf362da683827d6de9407e01b38773a10f1db9be5da3ce6f048b4bc3e43eca881edd7cc2582;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41e378d6a2ea0063e3827bb2d325c23a7ef2dff8230f064ede4b680ba8e0262f60f8963049ad47ca6f559e885c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bde5b5b83d556b7075a4b4894d49d341a2b3a4ddf89def1902fac678e94fc8b9d4de9f0b87d7adda7fb45723da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha76926e864d5bdf3bb2fbd25a4725f8ea56bacd9c8fc49dcaff3e4ae04556fa7fb58b85fc6fc6e655c8fa1ad0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107e042b8b685b3dce042061133816c1049e7e192f23d7c09afa7b6936868c8e833075b64acb67f96f4de383a17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1873562d3bde81e63b62840a48af480b24f915fcc6399081871b7a55d19745f0871bdf0ff894e970d679c2f999e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he58b7a73ee71dba062c42a4cbd136b08bc1a2c95de69f37a55fa0c6973dd41b65b763db6d4cf8027c1de31d619;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fd649e5cdaf6359f63989d90ae0adf384c3209e0e9b3c9d812510705151bb3212be1b96a48e98ef24bc45158ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16266ea58862efdc1f30c8959b6f98d61f4f0231cb89f0bd254b118f43fcd5a4f2d26af66f28423184748a9c22d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff34f1b78b35ea294eb3b317f3852d360f0f15e7517a8c563e4711644a477358c5298229ec5213b23f99359b21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12eb2998d91d02d54962f983204c6af4c21926e05b425a0df8c9cb925c91b820775f4c923dab3bd97938cbd27df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc16685ca02a145552354c12e5ea8e4bfc44955e07ea03ccfecdadd6cd7f2869ff1f26726d0e83e153da6a729a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c402a917a0870fbcdde6ba40e4f5c65a2b1abd5579523a7466c253bfa406c3015b8d43eae56684e69504a9cb75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186f5699c30b9d2e8e9f8923b25d99d5b09a6fed41efa3fe9df00376f5c616ff4d09b6adcd5a5d0fff60933d46a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136c2fd3408ed28bf936c8a93d255f64bd428ed8b6fcb66608ebe624b7322318c0d9cfdf15573db1df364c94230;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16b2f51363a9ceed322c65285d82fee24f168c8f8e13583d1cfc6c95d2ed43a2c0dc99c0918e2aa345fe2de7777;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d33ff0cdc7adf5870bdc5015f28955f7edbd3b08e512cf287c1e299e6ebec78db38b76c24e0d6b9e1967e4059;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19040e505cea0ca976cfccc894db82a57fa00f78dc5d7b5b90d1ebf17236ab434a7fa9eeaec3adee891832336d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a2c650fdec52e3902d4a195622d7ed7d4d5d526c8c3032d24a8c7fbb48d817fd13b5ceb7d29f4065962215a73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had6ffb66413e8fbb67dcdef0823f874e9d887282e683ba540f960e5d06c0744719a620766202e590343d6798b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a6f37b2f3ffd44e1c14e81bd840380cb78026eb97afffa4b626a2c854ec04ade1603ad3c71e98ac487aec861a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1045a8a4660eceb062a7bd4c8d30e028a483cd4eff511db356240db8d0172c7960bd284d79884e424a141f8ec6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f154f1fa4b795b2b6e2696612cf824e1fa855161cc068d41df6753fc75c8ef8dfc5253161a365b4b56be89a599;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heca8a42b6022b20a3de2429692e39b15ceb218e7481cce7707d81d108a9e1a55a59abda494fc637206ca44c8a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182f50b973aa02dca2a61e5770feae603adbb489497c9f644b720a5d3b2fd95534abba1b03e81280d28ea2148c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199f83019f7cf51d7df153b6fc3c564186ee86ed4986e487e27baab3f290b9f671b981cde66cf80629d5b516a5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1de55f7a70dda056de989875f165cb0bcbfe01359565be7b0bbc628e442904cc86fc8f105400af05d3366e419;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c83e466f4414801bbe399bd29918bb2caa01e0bfcda1c94083028c9416600880070f05d6886eb299f7e52591d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1563071037778accb7a40312ff62393e5d7178db0285474e051bdfc0f631ef0445d61ac9cf1384a311058639e16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a716ac46d8b678fb93d5e7c8491081f2afe738ad71ff2edc3f83527a10c2e89f6677209719a3be4a7414c4186;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h152f89f861ac5896c08b69c7120096766319c9f8c0559a5135ab68f8fe15c15ca54d30aa4c6ab80292ade1b3cc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f6a6d3651107c660a52550a4a7620401919e8e92addc9fc6b17a3a8805291d62d0831491f506100524bbf68e5a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc8cbd22f2eb551cb2d84d3427c33de9e1e0a4942f8813cb7120dad484947a52c6af51acc014edd1a632fb187ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0d32a33fa18ef32eb06735a34dbc98a0380accacbf3c2d2c7ea369a7d713c5d1ebdd92201a3f4b2f89029b185;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cff68d40f81d397c0bfcb7db0359434b8784a4a64d8fcfab76bdb9123f61c1fb751222f9bd640b3b9424e52878;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4225e2f137c6cb691e586e6bcbb8bf899715e1151f366c9a41fade8e6890adf7003f927f023441b87b882e403;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14acedcd9c101d749931960334ae91a1c1c1f9e9dd8cab638be86d849bc923e156cceafe2a57577aefd5617258b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c3ebc43840b355148cde6099d0709292e23108523b88f0d1126cce8f47b0887472a84e1b00dca6c54edf145cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he64ba3581dea9c1629dd84ee4857670b802a1d517aac3e9a5914320e1de317b9857aa90ff9f212a6b688f78cfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1791242c57e394d7eb55766df533cf7e279c39100a8b0e99385cff24eec4884ef8b025f76331d3653edc1c5c7b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6998d560491fa808230b5f876608d6f3b0dc08a74bedd66c6c6de058d7f6ebb09a9a393bcc3a2ca60581ad70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he81650be2e26decd84e3ec30b60f9dfb9758c333507c8023c179a55277b5b584fb01c6f1530f068321e92445e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88be453409da4da3b21e1ddc66e5a565a31157e349dd7bfbb295d3962c190fe5af41ccbc2790bffa5190633f15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h22c3433d7c232b9cb8f73920f2c7c0ccb4d775dcef11dc4e8bf66bd9b2e458cb05a6ef24c1b101a79e084372e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h100a4959a6cad431813657baa8f21ae4e18900fcd315b2af1cd9780d3c6e6909c07dc44f6a5e92ed9d02e829b2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc6ac0f238b76b53569d0ed0bd19b7875a031f39d88a476b4622812e9e964234da147c6e02d130841c76d9a2303;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af603c13e46c93b16aa2803ed0cc634193945465a694f242c9811428438b0c1a4411e216edec16ca6c310b5c21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c597a1ea743f5638be0c08ca5b2d65cdaa5d56712419277154404537b7936c25470dd736d63c0a4c38d0b9ab0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f9f9c9d093d7b1279db27b6ef64e18bfe2ee37c922e8c3acc188c96f9a5936f22cf7395798753fc1d33dbd508;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h710ad0330dee8419e9c97c80b346e67986d0f35aa3038df1ef8230c9badba5a3fb1ac30723657fddb05fc05928;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159fb792c5f7198ed96b38662688e77ad09a303e867f883447c2bd7f6cc14ff5ed99650ad970ebfdc5b8d22b94e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cb001bd6a06d78fc4a8434b08ca6dd014a36460655d696048fb4c5235b408e8b29fcbf33e82c37e0a29ddfb09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b14ca783c7c3edf4e302a2110cdab59be62dfc1fc981525f6b344f7940764c7bbc97a99fdaebd85bbdc921159d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d3c9e14abf4172e0300d9c53703f897b0359a1a474c97030123590c80c7fc6329342a194dfc98f9910c029917;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6794060c093a514eb2005755fb7c65eec50329f1b15579f66b988a8258684e538babbed326de143c4d529a35f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d9a5294d9d66b72fb4836cf1329ccae7bde3485dae5813a778f03cb23de1ccccc82337d34eff17a94da96339d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hffb59606dc46bb7557e008eacfd0f636e6bae4ba175e8deca0eda376e587d09e5f358e5820aa89fe5dc8d65abd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1955e98ac6b800e4c2e9121e3b8d8e0153aba0220aee6de4e63de33750a036a9cacb48e2df9d1fc500b95f54f8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a42a6385cadc3c94bf75554a95ad0a7abe396397517ba7ba7b244333771c812f89ac6678ab67b206594a53c72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b45289f724c5e7513ade6b2766964584fff0c1b0102d678cfde79d44459b224c37d71b8970d67abad398cf70a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a76c24bf315af16460301228ed0be8cc42194ad8dee44fa94d985b885f5430bd22f3399b354af059dab1517ea9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h84284ec9140be334e6ce7bfac0d847a0f39e1dee9a66f8554bf5af99a6fadada6f2db1ea425dd910f608d8ab5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc9f86d30156048efca5daacb0b4cdfd499627f97137df4acd1d4220617d6638dee857c79df24b4314145e7f85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d4098924d6fcf96dbf2997615bed7b3eff8157bf383775f7d7e51fe8f80e60142f33dcfff995b99a1c74865d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9c94ccd765041ee8e8bdf1a4b1ad5ed037eed6695f8b0d8eabd559c5076b9b19a8a099c9aa90b1ec80b76836a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1735cb0000eeb9a5e22efc585fe2846b656b5e0df95787717a3db7f77993f8c04d4db198b1d720cd6c33f08df17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb8cd34368b27948e92eeee86219592d534d665ab43edf3ce195333665889e608ad207fd224529e560c26de919;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb92eb3a7063e2d838d513ad33fc738b0797cbf27bef181f98ec98e8237fa5890938ce414718e2cead27583828;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6875f8ae62ff9ceb26d3d129405a99ac8c58ef3aa98cb123b778a7bef0140333b8c0d1c2def33e3478406edc9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c90fd6cf1f7481cdb44759059820c2c2154d3615df8298a6ecff2a5f2b7a6a21586db87ccfcde1d4747a457b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be2dd7ac7706bb679e0d90946ef242a08140ab97442d3eb7b70f57a2dabc042895621d5606da4c9736085c982f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9b794cb0868e4eeaf794f0421679ffb8d556b9969f1625488905fe1390b4ce81d3647d380ff5a392cf6bcf49a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb24db65cf40f88b21996787a03ef3ab471330b5550f18d06616506671da52637a7e3fe8330eeb9a17dcea75a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1535ebfa2724e846ef08cc8b3f397b0f50e0e20a85af908993456143d0d852d2a3d251a3dad4e58e6495f6b5114;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hec7d62010d93327beee4306958cc19980f2ae089aeecf77db74b7cc8e5ffd15e2cce63527a1ff14b13ec7ba7c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e66f0a700986527b3bd0bc2f9ef7bccae795eefaf1d84fd51256d2ba8480e8d08144494aa7ed9bb0b9d29bb923;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19fcf5a1ffcbd00ee15426a0cf0c001294e262249eda3696f3ec967514b5e93946469d5230b2c2549b6af97c6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a573d6aebeccc1b54926e7ba1e0853cb7d4f92cdd72f57f062679ce11b7e0b577f38f0125207b1747b9b061e09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f1d9f39928a383a61f02a8ee5bd0318dbe39839fb52dc900ec95672b47fbc2374f7d32523d6aa28eba75fa837f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he52f81c57ce8a3fddf363300c3cf71b8c703a3542447446581bb019bdb44fc35d039db21f6a456f891972a93da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h96ccf5a189b5d20291fa81441e5f64568aaae4f613f1900d38e84c88770fa8b3de21c7e23fd4806d392f48ccca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7785335c792c6515b9463a19522389d10bdaf2299d938ecd7f4f50c47e7e2eba248dbbdac63c58eb22133a0375;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h719319cfc229530703245455dd0166a49e39cab421d12d51ccdbaf50a19d3978676d6e20d459cf51a44be33638;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132e27124edf9ed6c9828a2dd881580b40d5df1cca1b6823dce9dc2e4a91b1275367e797606b2adae719487150c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160fa5732ec06b9b307f8bfe0329ec674681580a291e7056587f7cd0c95de22bf6028a9730ce4d2e0ae68094116;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d63cddecc94717a31485d969319b38459cb0247a747a1d9637e190e1e625f1fe54d8a5a78848dde108cda6806;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac61ecf48a4567ca9128ebb6cef2ae3c138bd46f1f4928c05c6b141069f132a42c8210c94e34c7bd7d19d39df0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75d6d7e9448d284a6cf155e5fc7f710bdd339800cc0bd8e89fb49b8312047faf8da3d4d6c816643a95874c1643;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd2077d87dfeb05866f7deb1079ff45b3ed69d77ae81495a5d6838d6f393fb00263d5801b60f146e419eea2592f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc24de010978ef1f143365ed9f6ab97aeb785df67a744711b9c5a9ca9a2d877fb0afecd596fe93c3b096ab6bb68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18db782aec81698d42fae20bbbc069775a9a5042a05350a1851d008df079f1c6420ca81fb7249195e76d53a5341;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef556fc2e0d57dd44fdbffd8db7c9f425a9590e08d63edbc452ddbdd1e6af0c93ff77a979d3dd30433240ef41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f361360626c614478741699cd3ea4f3876dcf10b46887748351d9380ee53bdefd628303099f2c1137eb061872;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd55574eacf5cddbba4f908310f6d236e373e7673658fe02852b160e37c46e3ddabbe0a0ec9fb720d7c9b6bb8e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159f86dbc5650aa7d9e0cfdabd65f111213c5f8bed195f10a06ee88c2556580d1b352618273d11110f5da96c72e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fed2cb42a6a26aa8fa4335adeadd8c8ef383208521678b252c18dd6e65b5cfe0d0c4cac82715caefe6bf1ba646;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1861a3e6c1feece9b76d4805e55ce3591caa5de080584c43a77b2ebaf2888b458a32073a805ebe7f3a8d6e460ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he88bfe1b7d79ff7209669a2cf994f246ae2168d9d5d9b46124155ef30bb28699e6039e78645e24031324b16b2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4adbf5dab7889472b3adab44397337a52e5207e1d2f92d2ffead3091010618ed8e79b6608aa5759d18128ad0f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b385d5c5ddfc6fe865093b69202c270134e7f0f9d43ca6667b9a0b0b6205670ae32cacd4c49c361e8635e41895;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d0eb0d99271cc3a7e5c0bf22e4c2b5fa844d5afd0f6572337603ca7170cdbee17da327af26e5e54e126f8b559;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a42b4336ef653bf35bde4cc4e50ff769aeabfe94c6d862c56ad5bb02d10e29055a1cdb1933edf6ee762bc084e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d0fd5c0a46fc6cb1d296aa1bd78e08fb4a4d2d847ccb85422ba40cc443f920269dda5338afedc07da8f6740f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he1203e3a37d9f3ebf6fbbb4519d2f124a5394ac9f8a86dfbd0af08d4a083161725468457c6b198d7552fb17876;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ab88d40a8d9ca73bf6f5d4e8ba0d36fa5f31d5192f9950c042608202318448e151bb7bba0f78bbf54291ad773;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a67ab71438a225fb0ab4489b405ddb04b3a65cbbf5a32f7de87e41f55681457aedfe5b2f5f91d45f40ec77e98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127ecee22f7724db3e2ffa02e39b6d1a50d2f97ed18e5462bad4f5cb1d2f6fd2e7df895ae051ce829c8ea2249ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf84fdeacd6b9c147435ce02be9f339a2b9e898dbd974fe90b711d554723fa7517f265453dd48b71cc94c4e4068;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b7f4e55f64304a49b3aee30e034f7477df6d5f02173cff735fba2f947d2b637fb6947090c0902d9dc3068ef4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117ea5f921bbf59a11c5784fb96e3a7c3430ac3f49e1b79b4305d0141a8eb7b2c37c7451e45316b48e4d5a9f477;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45e5b548e1046339db82d9ede156aaa328e3d1f52661b5b31b29a53690f1c62cf5ede3ea1b6a75bf8d362ad601;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c7932644c5f2b7f0d6b0de2c3d5fcd3be75c07c54d871565c06de7495d829e3fa6605330b9e44175b1bbc51ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e3edfe1b24b5228c50cff5d1aa0fb5bfffe4ab0848f26f9a9b3acde9ed01a9fa6ea56c7523a5c21862dc3b248;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h137c20ee25be136b55de1e334934d75a00b9fbc54083e09fc982b4f725226307e0e826083e5e9bc16f0ff6600;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7fefab5c2fc9a168136839ce0fa46ccd69825fb6381ae9d814b525ca0551ae943540e9a7928597f309e1dc6d56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89fcdfa7a9865d10ec86ae34d1ea0c32f8844206a8df3bda8747013598a0008643d0bcf406f6c7f3b98a03fd5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18e0beddebd256ae048f7af6bce2f43f4c2c7d1063dd7429a7616b6135ec910adbd86a5d31bfb72df60d2c267e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e9ba57332d54f693fabdd697a895e2e04de72b6c2221ca55428c12d4f93023002c792a0fc741acc12be1b883e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53b815ada12d6ddb64d8a48d976627d3d2853fd8e770c09cf14caf9ac0fae83d5a62cd1b26f3ad8676d737c476;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h200bb445b2e478c24f5229bdb30c851172715c003411d415be226dbab15382c92f0d73dc79a10cac5bc241108d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf516abd02fc5b9723951a3dffea26408b92c72d07748d39364ea743bf0206fc4cd930c5562560dbfe7de09f8aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb06ee6f863bc0cc52cd6972a5385c5c10cef4bdad4d2ed0fd9074ac8630bc96eacaa1c7c01c8bfb2ebc9f60617;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c026f48f9fb9928beba33012f5f933d51b008f8d1bcbabfc1b7b0fb611787da4876e2c0c29bfaf1056381979c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3dd8c1241e0e53bde0c4dfab8b68b1dd65a2e6bcef32d9b801469fda3405a25fa0b0a032e255ffbdcae52f554;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e4f76b9408b59a452b87da81ef4a38f017f348739a17cb19b015e3cf46a530424fc7fe19b2b3a4dbb36ed7587;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98ddd855f31fa9caf8b9c9dcb64b769077e88e79663d9d66e15323a727a7a86e004c26207eccc8e53db0e0d884;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8f0e501396ad7c2e28e4a62a07afa7898586c7cd10b817aecd4beb2609a83016bcae3adb28aae8ea06017524;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48f164165f203dd11d3895d521148f8ef1fd942aec9ab6024e55fdd539a39d2d9646c8d3c1825fc744966044f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h59e27fc63058ce01fd5e898c0a69930f22a24ba227e795fd8faa6ebc6e4fe40d29b45d529c38e701d1ae8f581a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103a6be6351a004da888687e8b6859d33c82b7a965c1335de9c5492767743c26c1f82dab6e0822a1159f8f4c01e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df2fa005193a9ea737f3ea4e3db102a3d768157947fcae7a2379b4f1cec9a54d45d9418f7c9db7de75c0807f55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122ed6a754918d1986df275eb00f8d10b8983103ad8b025b4ac9a754c960ec2db4516d7c1f0c77eed6533071944;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c548a78b95411f2079404948f92af8c6670aef9e8377436bc025d4c352ce0839430afe81ea0d96cd3340fdf3ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1531947e51213b129e941d7d721c9e2d83777dd1262b0f84337e55b1f73597d1d00aab28e22ed53f24f266b249c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17524a36b7fa8ccbb7a1d9c53f2c3b296d7f74c694a529fdf34b7c2cdfd46e0400f169cbd10209e20f3d2426822;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd9ad991c980f005a964cd800a6f5fcd0384be20b860b03c8a56cc27ac39048bca5c953d78ce1c4d1204b021988;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122786b09a0e4d99fe6b2f7ecd03ae279b02c67cad5e6582c0e1d25bd098c5ae43468b4f167b2ad730f9b41e7f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167e1a76669a4389b1cc776633deff2089e538ec10a2a41c7883e64ad81640216dd77269897bddcc554f367464b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de1e563bf151aa30df46314eae29bfa98924901dea8613f08c7d45ec8323835c76dc494bce62cd70e324d19f74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1649dc58873a728e4715e6cc88fb08a3440588367f3ec91b9d2164dfe6631fac835c78f8cf502a55d2e9eef9598;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1dcc5652c02314d94de7945c6cc1eb781e68330f48dd23b6355932db82c11f03cdb55d3f05127ff2f5cd96d0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ffd7cf5e7fbc1cbb9903f68780e585bb1e498a1463d831bcd2525ca7dcb54721adca7f0614916ecf7dd2280b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c7076585e03fa74f2dd60c2f1947f3e9bcd4b7f5becf9cb19d92a5ab5d633bb06ef877e8d4077ea8dd3dc71979;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c10ce0a47ceb9831b9610b60581aa5eb1b29b1d7ecaa14c02e007fd22c2761fdc4bd278b53b2ef9ce1647e067;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hebd2e07b0a8bc8459231854eb109638fe7799b4ea1e4132bc7f301e76bca916f35a258bd59f42f49a1caf22780;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154f83af045bb9249d995c2f4809e2e0348df6a4f83e1f418f2a62ac443495212903a8e19e7ceccd55b94bf51ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h174f915ab003d6b9bc64f5469a471d564c4cf6b2c72340c2f773e4d976768e4a4a531df213b7131a49d66070029;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ba040cb3a85a2b2cd68424f7571b5982bd54d1d373fecc634ed7a9673c2c396984ff69fb7cadff493fb3ef568;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ba414419a0a4b4bb4f2f42238c1bf0976e25f059e038997331e2a479ba77310bf7b09b12c00bb40cfd7e452b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed7ed88d6fa4dc55a20e549b0d251531cbca778369f1389d5d061d9bc17a4df502409e2c8b3388dc7c99b43c4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b8f7392b1eea2ef3c53bb860891767e1de4fe0fceea95208e60505df027c940f03c3b9ac10339c4c9ab87bb7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4af10eb108d10a7a13b720ac52d19257353e74d5bd94fd130b5f1e7a3fa36ccebae267f71f29a8654e8fe41fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c729c4dee23102bbc0298a4130b013cb5cfa80ad93a504a9bea082dc528ad769631176cb11472dbc2365b152;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121cca76db960fd3240b0b033f74bf2d511ac188f9983cb035cd020328cfcd6ed74b6e4a7a41cfdf4c1f09c0551;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3d9672c7699d13aecae5d5398a69794bfc5c40280e66a761649672caab9b750a3e6ea952425037c386f3426e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20784c6e085d7b03a015622fce2fa3ad32f8a0a56255cd7f89edde568e1e0f4e442d920673818ccc24ecf10a19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15761ae0ae91ccbddfa676d03a6c52c997068b78f875380263d3f4f25edf932f76f891f093293866e5cc0a8a4a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b2d4ae1b102a56375b62d5676e967198551b0a46c489d6d469c15f96e3a82d361e2142f132483d63ad59a8ea78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1896b47b11204c5e9d1024dd5c0e891257a47b58a68c9fbbff408ea3c16f1512acf1c25283d4db0463fdfa8aea5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d41eaf212da2f604796994fb53411e33ebc22f7e21e0b8221f48473fbe8e8435fec42eb9643ef959ff5a38381;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104f23c9d7263039804e6130ce2672f8994ff3d8123f37fbb6a674b13b8e64dc2f48bf7e0bca2401c86de98a79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9ba60cdeb3cb7ba60352a0a786f8a49046517b2e7b80c76ec179c408f807cae54df524aedd2452da8f1a12277;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb76652c79612d657ab613665f129dcf069ee258c45e55093181c4ae371fe3c59b9e107037e66a51071a5a71a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd5733d43ad950f2b6c31a27e95527865178708176805c193ee0ccdacc85453243c8b659b8d4fd7100fa3d4886;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3ac473b9f23644354b18f081fa3a67fecf4252a8756c9dd06556c2e979f27487c1225ca150b742a9125f35d6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14006c73a240123925ee6fdbf860ff19d5f0488c4f14c692a18a701e6d003a49e56e65ccc7f8b6ada07e80617b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd7b0a2c2f7cee9ab102f8def66494f572e13150809220ed522a579909eb819f098dfd422e3a2a20867188af01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2e2cded578b060bc8982604dd8e006e0349e0d28baca48581b96f70c38ab9097343965672e3de9fb2bd4dfed9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e92ce8ce99faf36e9db7ce4d06d7292bb16c96cc5ecd18419c09dd0d0481a19f79270310cd222ff3d82cb0324;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2003ee97f634623627ba9d413f45e1df8cabf59895ccc79c1fc9f6cf2adadd040caa73e1c07dca17b5c20bce1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1559700769ad6c54bcc80effc130449f0fa8ae91c1a7bd34767d56b33ef572bf78a2fac9660fea95c8829aadcd7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ca46ef8ea1df24b737c880592ca797bdf98b9be7a87fddc5b12310675bdf0c1f60bf993eedaead35773f19baa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h810c71f3bfd0ec9bcbfe46fc591f6a0c20f2eb7c04eadefc68b6bcaaaaa281d6baa50ad4e09ce2bee52c022401;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172e15354731cb0490289981286ad7c1cfa623fa5dc3ba826ad3222c436d1b50d54ce8ecea8ae4df8f371511ebe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50ff09acd55ff6cbbad5e34d9d1b8a9ae6a877337554074eddc87bc4df7a3581e933b9165aee5df16071f318ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb9f76c6ae4a38a4d2838e976fb0fa425807a5c874ced4ccfdea79f870a87c7fc6195386bda4a2ddaef93064d84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2dedc89e2be276d6bd5ac05dad03206b1c1d8c2ad93c56fb19a2ee9bb053e65b22ae353bd552391279c705b2cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90ae07a542ac3a768f835732d6a485b6f043f9e0ba8b4647d806db4e1e089d55554f8189b5fc624ed943c02f33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e7b0dd8769eaef6b5ecf8201bace2a0145241e824cd59cf4c9460ea2a4424d032628f573cde12c637a733d1f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac356edc5260353eb53e6e80d07736bfe2c7f4edda99ce55a8c6c83dc71721abd28387f6a47959c011a098a307;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8d8f6b755a8c1d2d0cf08b186d4633c59527ee06c70bb343e47236e701ca7237fd4775170f3cee069b4e6ef48;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c359ac113d997609f59099d2a1fcf20ef2ff2a8697c99ae40901ecad5b877a33baf38e1c0236492ab68d4770f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha4350f698cb5fdf56dcb7b3115de4665dde0b6263a85a84845d3c7953553dde549a2e09398997e0ed30092e779;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h126978e579ba2c4bf172fcf6a3b3542bc7a1b887b88a0796be869c4390b5f3f364655fce1713d6c0455c49981a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16379dc0fdff8821e31812cf81ce038970cdd9fbe5b9b12e3fd0acf6a612c4b7b33059066bae6349088b5328487;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf9880ab49f7360dce1013e116ea1b299db1ffc5e397d1ea33534abce19746f358dee6a7532f0f62a3ac7ce7f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h922b36df3a7d17230e6c076f62d81ae4d2c0a435b814502e91f64c15c94adb1ced10ff033d527836410086d6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108f18b31e1793a2a4d4d4fd68b04d961139b8ec9f9b3bfe5ddc64e347b3bb2e4b4e34013904d3c5f6798654c83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h674b399d709e24ad03ed5dc6d437b24acfc6ac7265f7a646d6f927286869a6e959e0f5cc7c804d73e4ff9ca90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4041dee6138906f930bc085573f69dfed7e0bec6c35ec296b9fe0469798f82db688702176dcbfe680d033d0cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f1ec652498d691a98cf85a930a06ec10a6cc4e91c60b1c3707da76591d202736e3892a3897b5215018f78314;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcf9bf90573ae4355dc26c24a26153f71de3efcdc41e51e7044e3c1e83765fd0534130ef863c911f3edcd6a6818;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4cee5324ff6f805247f0d0ddd260ea8b1c29fb1afd35d3b0b943532b70ead5f5971b4de597d62c3bbd8b5342e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15da3dda0690cc42fcc431d922437b8b93b5079cbde20ec0119040bc9b08f633beadeacde55169b1b45b5458a02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1217742b82c36e95b280710c52df1f1804844b7dc9838bf3724a1143cf309eed5ffa9df84e4e8d59816de7d052f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149e387b8458120519663bc6ea2307f5d123c54fde69cd26ae8a7f48d7984f1e1858039137fee1aaeb048640e8d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf18605feb6fc32d6372f6af10911f051835c1dff2185fea06be753095270a477caafd46f7c090a9c1a7b15a945;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94336de6991faf0a5e259d1f210401bbfc20f42bf32f3561b114e1dc6777f8b4d8397a6eb2c4b2de84a03da768;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf658ddd3da47c926248a1032c3a1d0f3e8ba085314a5b51686e65b3241bebad6fff30647e5ffce0c182fb30212;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e58724cab71c94a8ee5687bc176217d7e5221bc582ecb7d4f1c52076c77cfb93eab9cca90aa57444ffeaa616d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbfd823d7660fdf07f1e7144b3bf49319a6e710f7ab2fd89be7fe535dd6c5c01bbd6c36a5319e83cf5192ae8d9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199aef807fb300897b7b78d4b8db60f81eea279e27328ad561499ab0849d73ff0c365a721a8cb07a3ba8e8adb91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb9310ec379b8617b6865c099850a8e8107a4b6cfa98c326c3f50eeb55a9aab10109a8f329757b460af3d292b73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7bf967e38a620eb8cea58edb5af7e5c05f0b80f208398554f3e632359ddd5b618ccafdbc50409f6b9501a6e1c;
        #1
        $finish();
    end
endmodule
