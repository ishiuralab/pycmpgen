module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    compressor_CLA162_12 compressor_CLA162_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA162_12(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [0:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], 1'h0, comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [0:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [30:0] stage1_0;
   wire [52:0] stage1_1;
   wire [65:0] stage1_2;
   wire [57:0] stage1_3;
   wire [138:0] stage1_4;
   wire [67:0] stage1_5;
   wire [111:0] stage1_6;
   wire [47:0] stage1_7;
   wire [72:0] stage1_8;
   wire [78:0] stage1_9;
   wire [58:0] stage1_10;
   wire [52:0] stage1_11;
   wire [52:0] stage1_12;
   wire [26:0] stage1_13;
   wire [18:0] stage2_0;
   wire [22:0] stage2_1;
   wire [26:0] stage2_2;
   wire [32:0] stage2_3;
   wire [44:0] stage2_4;
   wire [37:0] stage2_5;
   wire [49:0] stage2_6;
   wire [33:0] stage2_7;
   wire [41:0] stage2_8;
   wire [29:0] stage2_9;
   wire [29:0] stage2_10;
   wire [24:0] stage2_11;
   wire [27:0] stage2_12;
   wire [28:0] stage2_13;
   wire [8:0] stage2_14;
   wire [2:0] stage2_15;
   wire [11:0] stage3_0;
   wire [13:0] stage3_1;
   wire [18:0] stage3_2;
   wire [14:0] stage3_3;
   wire [18:0] stage3_4;
   wire [17:0] stage3_5;
   wire [17:0] stage3_6;
   wire [18:0] stage3_7;
   wire [16:0] stage3_8;
   wire [11:0] stage3_9;
   wire [13:0] stage3_10;
   wire [17:0] stage3_11;
   wire [9:0] stage3_12;
   wire [12:0] stage3_13;
   wire [10:0] stage3_14;
   wire [7:0] stage3_15;
   wire [0:0] stage3_16;
   wire [6:0] stage4_0;
   wire [4:0] stage4_1;
   wire [15:0] stage4_2;
   wire [5:0] stage4_3;
   wire [6:0] stage4_4;
   wire [7:0] stage4_5;
   wire [5:0] stage4_6;
   wire [6:0] stage4_7;
   wire [9:0] stage4_8;
   wire [6:0] stage4_9;
   wire [5:0] stage4_10;
   wire [5:0] stage4_11;
   wire [8:0] stage4_12;
   wire [4:0] stage4_13;
   wire [8:0] stage4_14;
   wire [4:0] stage4_15;
   wire [2:0] stage4_16;
   wire [0:0] stage4_17;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [4:0] stage5_2;
   wire [5:0] stage5_3;
   wire [2:0] stage5_4;
   wire [5:0] stage5_5;
   wire [2:0] stage5_6;
   wire [1:0] stage5_7;
   wire [5:0] stage5_8;
   wire [3:0] stage5_9;
   wire [2:0] stage5_10;
   wire [1:0] stage5_11;
   wire [2:0] stage5_12;
   wire [3:0] stage5_13;
   wire [4:0] stage5_14;
   wire [4:0] stage5_15;
   wire [1:0] stage5_16;
   wire [0:0] stage5_17;
   wire [0:0] stage5_18;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [0:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [0:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31]},
      {stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73]},
      {stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85]},
      {stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133]},
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc615_5 gpc23 (
      {stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[12]},
      {stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc615_5 gpc24 (
      {stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143]},
      {stage0_1[13]},
      {stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc615_5 gpc25 (
      {stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147], stage0_0[148]},
      {stage0_1[14]},
      {stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc615_5 gpc26 (
      {stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[15]},
      {stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc615_5 gpc27 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158]},
      {stage0_1[16]},
      {stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[0],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[1],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[2],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[3],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[4],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[5],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[6],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[7],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[8],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[9],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[10],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[11],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85]},
      {stage1_5[12],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100]},
      {stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage1_5[13],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106]},
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97]},
      {stage1_5[14],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112]},
      {stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage1_5[15],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118]},
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage1_5[16],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124]},
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115]},
      {stage1_5[17],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130]},
      {stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage1_5[18],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136]},
      {stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127]},
      {stage1_5[19],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142]},
      {stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage1_5[20],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148]},
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage1_5[21],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154]},
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145]},
      {stage1_5[22],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160]},
      {stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151]},
      {stage1_5[23],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc615_5 gpc52 (
      {stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage0_4[0]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[24],stage1_4[52],stage1_3[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[1],stage1_5[25],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[2],stage1_5[26],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[3],stage1_5[27],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[4],stage1_5[28],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[5],stage1_5[29],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[6],stage1_5[30],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[7],stage1_5[31],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[8],stage1_5[32],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[9],stage1_6[9],stage1_5[33],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[10],stage1_6[10],stage1_5[34],stage1_4[62]}
   );
   gpc606_5 gpc63 (
      {stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[11],stage1_6[11],stage1_5[35],stage1_4[63]}
   );
   gpc606_5 gpc64 (
      {stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[12],stage1_6[12],stage1_5[36],stage1_4[64]}
   );
   gpc606_5 gpc65 (
      {stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[13],stage1_6[13],stage1_5[37],stage1_4[65]}
   );
   gpc606_5 gpc66 (
      {stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[14],stage1_6[14],stage1_5[38],stage1_4[66]}
   );
   gpc606_5 gpc67 (
      {stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[15],stage1_6[15],stage1_5[39],stage1_4[67]}
   );
   gpc606_5 gpc68 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[15],stage1_7[16],stage1_6[16],stage1_5[40]}
   );
   gpc606_5 gpc69 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[16],stage1_7[17],stage1_6[17],stage1_5[41]}
   );
   gpc606_5 gpc70 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[17],stage1_7[18],stage1_6[18],stage1_5[42]}
   );
   gpc606_5 gpc71 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[18],stage1_7[19],stage1_6[19],stage1_5[43]}
   );
   gpc606_5 gpc72 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[19],stage1_7[20],stage1_6[20],stage1_5[44]}
   );
   gpc606_5 gpc73 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[20],stage1_7[21],stage1_6[21],stage1_5[45]}
   );
   gpc606_5 gpc74 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[21],stage1_7[22],stage1_6[22],stage1_5[46]}
   );
   gpc606_5 gpc75 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[22],stage1_7[23],stage1_6[23],stage1_5[47]}
   );
   gpc606_5 gpc76 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[23],stage1_7[24],stage1_6[24],stage1_5[48]}
   );
   gpc606_5 gpc77 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[24],stage1_7[25],stage1_6[25],stage1_5[49]}
   );
   gpc606_5 gpc78 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[25],stage1_7[26],stage1_6[26],stage1_5[50]}
   );
   gpc606_5 gpc79 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[26],stage1_7[27],stage1_6[27],stage1_5[51]}
   );
   gpc606_5 gpc80 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[27],stage1_7[28],stage1_6[28],stage1_5[52]}
   );
   gpc606_5 gpc81 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[28],stage1_7[29],stage1_6[29],stage1_5[53]}
   );
   gpc606_5 gpc82 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[29],stage1_7[30],stage1_6[30],stage1_5[54]}
   );
   gpc606_5 gpc83 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[30],stage1_7[31],stage1_6[31],stage1_5[55]}
   );
   gpc606_5 gpc84 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[31],stage1_7[32],stage1_6[32],stage1_5[56]}
   );
   gpc606_5 gpc85 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[32],stage1_7[33],stage1_6[33],stage1_5[57]}
   );
   gpc606_5 gpc86 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[33],stage1_7[34],stage1_6[34],stage1_5[58]}
   );
   gpc606_5 gpc87 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[34],stage1_7[35],stage1_6[35],stage1_5[59]}
   );
   gpc606_5 gpc88 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[35],stage1_7[36],stage1_6[36],stage1_5[60]}
   );
   gpc606_5 gpc89 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[36],stage1_7[37],stage1_6[37],stage1_5[61]}
   );
   gpc606_5 gpc90 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[37],stage1_7[38],stage1_6[38],stage1_5[62]}
   );
   gpc606_5 gpc91 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[38],stage1_7[39],stage1_6[39],stage1_5[63]}
   );
   gpc615_5 gpc92 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154]},
      {stage0_6[90]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[39],stage1_7[40],stage1_6[40],stage1_5[64]}
   );
   gpc615_5 gpc93 (
      {stage0_5[155], stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159]},
      {stage0_6[91]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[40],stage1_7[41],stage1_6[41],stage1_5[65]}
   );
   gpc606_5 gpc94 (
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[0],stage1_9[26],stage1_8[41]}
   );
   gpc606_5 gpc95 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[1],stage1_9[27],stage1_8[42]}
   );
   gpc606_5 gpc96 (
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[2],stage1_9[28],stage1_8[43]}
   );
   gpc606_5 gpc97 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[3],stage1_9[29],stage1_8[44]}
   );
   gpc606_5 gpc98 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[4],stage1_9[30],stage1_8[45]}
   );
   gpc606_5 gpc99 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[5],stage1_9[31],stage1_8[46]}
   );
   gpc606_5 gpc100 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[6],stage1_9[32],stage1_8[47]}
   );
   gpc606_5 gpc101 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[7],stage1_9[33],stage1_8[48]}
   );
   gpc606_5 gpc102 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[8],stage1_9[34],stage1_8[49]}
   );
   gpc606_5 gpc103 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[9],stage1_9[35],stage1_8[50]}
   );
   gpc606_5 gpc104 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[10],stage1_9[36],stage1_8[51]}
   );
   gpc606_5 gpc105 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[11],stage1_9[37],stage1_8[52]}
   );
   gpc606_5 gpc106 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[12],stage1_9[38],stage1_8[53]}
   );
   gpc606_5 gpc107 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[13],stage1_9[39],stage1_8[54]}
   );
   gpc606_5 gpc108 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[14],stage1_9[40],stage1_8[55]}
   );
   gpc606_5 gpc109 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[15],stage1_9[41],stage1_8[56]}
   );
   gpc606_5 gpc110 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[16],stage1_9[42],stage1_8[57]}
   );
   gpc606_5 gpc111 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[17],stage1_9[43],stage1_8[58]}
   );
   gpc606_5 gpc112 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[18],stage1_9[44],stage1_8[59]}
   );
   gpc606_5 gpc113 (
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[19],stage1_9[45],stage1_8[60]}
   );
   gpc606_5 gpc114 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[20],stage1_9[46],stage1_8[61]}
   );
   gpc606_5 gpc115 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[21],stage1_10[21],stage1_9[47],stage1_8[62]}
   );
   gpc606_5 gpc116 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[22],stage1_10[22],stage1_9[48],stage1_8[63]}
   );
   gpc606_5 gpc117 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[23],stage1_10[23],stage1_9[49],stage1_8[64]}
   );
   gpc606_5 gpc118 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[24],stage1_10[24],stage1_9[50],stage1_8[65]}
   );
   gpc606_5 gpc119 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[25],stage1_10[25],stage1_9[51],stage1_8[66]}
   );
   gpc606_5 gpc120 (
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[26],stage1_11[26],stage1_10[26],stage1_9[52]}
   );
   gpc606_5 gpc121 (
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[27],stage1_11[27],stage1_10[27],stage1_9[53]}
   );
   gpc606_5 gpc122 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[28],stage1_11[28],stage1_10[28],stage1_9[54]}
   );
   gpc606_5 gpc123 (
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[29],stage1_11[29],stage1_10[29],stage1_9[55]}
   );
   gpc606_5 gpc124 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[30],stage1_11[30],stage1_10[30],stage1_9[56]}
   );
   gpc606_5 gpc125 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[31],stage1_11[31],stage1_10[31],stage1_9[57]}
   );
   gpc606_5 gpc126 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[32],stage1_11[32],stage1_10[32],stage1_9[58]}
   );
   gpc606_5 gpc127 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[33],stage1_11[33],stage1_10[33],stage1_9[59]}
   );
   gpc606_5 gpc128 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[34],stage1_11[34],stage1_10[34],stage1_9[60]}
   );
   gpc606_5 gpc129 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[35],stage1_11[35],stage1_10[35],stage1_9[61]}
   );
   gpc606_5 gpc130 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[36],stage1_11[36],stage1_10[36],stage1_9[62]}
   );
   gpc606_5 gpc131 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[37],stage1_11[37],stage1_10[37],stage1_9[63]}
   );
   gpc606_5 gpc132 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[38],stage1_11[38],stage1_10[38],stage1_9[64]}
   );
   gpc606_5 gpc133 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[39],stage1_11[39],stage1_10[39],stage1_9[65]}
   );
   gpc606_5 gpc134 (
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[40],stage1_11[40],stage1_10[40],stage1_9[66]}
   );
   gpc606_5 gpc135 (
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[41],stage1_11[41],stage1_10[41],stage1_9[67]}
   );
   gpc606_5 gpc136 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[42],stage1_11[42],stage1_10[42],stage1_9[68]}
   );
   gpc606_5 gpc137 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[43],stage1_11[43],stage1_10[43],stage1_9[69]}
   );
   gpc606_5 gpc138 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[44],stage1_11[44],stage1_10[44],stage1_9[70]}
   );
   gpc606_5 gpc139 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[45],stage1_11[45],stage1_10[45],stage1_9[71]}
   );
   gpc606_5 gpc140 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[46],stage1_11[46],stage1_10[46],stage1_9[72]}
   );
   gpc606_5 gpc141 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[47],stage1_11[47],stage1_10[47],stage1_9[73]}
   );
   gpc606_5 gpc142 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[48],stage1_11[48],stage1_10[48],stage1_9[74]}
   );
   gpc606_5 gpc143 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[49],stage1_11[49],stage1_10[49],stage1_9[75]}
   );
   gpc606_5 gpc144 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[50],stage1_11[50],stage1_10[50],stage1_9[76]}
   );
   gpc606_5 gpc145 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[51],stage1_11[51],stage1_10[51],stage1_9[77]}
   );
   gpc606_5 gpc146 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[52],stage1_11[52],stage1_10[52],stage1_9[78]}
   );
   gpc1_1 gpc147 (
      {stage0_0[159]},
      {stage1_0[28]}
   );
   gpc1_1 gpc148 (
      {stage0_0[160]},
      {stage1_0[29]}
   );
   gpc1_1 gpc149 (
      {stage0_0[161]},
      {stage1_0[30]}
   );
   gpc1_1 gpc150 (
      {stage0_1[161]},
      {stage1_1[52]}
   );
   gpc1_1 gpc151 (
      {stage0_2[148]},
      {stage1_2[52]}
   );
   gpc1_1 gpc152 (
      {stage0_2[149]},
      {stage1_2[53]}
   );
   gpc1_1 gpc153 (
      {stage0_2[150]},
      {stage1_2[54]}
   );
   gpc1_1 gpc154 (
      {stage0_2[151]},
      {stage1_2[55]}
   );
   gpc1_1 gpc155 (
      {stage0_2[152]},
      {stage1_2[56]}
   );
   gpc1_1 gpc156 (
      {stage0_2[153]},
      {stage1_2[57]}
   );
   gpc1_1 gpc157 (
      {stage0_2[154]},
      {stage1_2[58]}
   );
   gpc1_1 gpc158 (
      {stage0_2[155]},
      {stage1_2[59]}
   );
   gpc1_1 gpc159 (
      {stage0_2[156]},
      {stage1_2[60]}
   );
   gpc1_1 gpc160 (
      {stage0_2[157]},
      {stage1_2[61]}
   );
   gpc1_1 gpc161 (
      {stage0_2[158]},
      {stage1_2[62]}
   );
   gpc1_1 gpc162 (
      {stage0_2[159]},
      {stage1_2[63]}
   );
   gpc1_1 gpc163 (
      {stage0_2[160]},
      {stage1_2[64]}
   );
   gpc1_1 gpc164 (
      {stage0_2[161]},
      {stage1_2[65]}
   );
   gpc1_1 gpc165 (
      {stage0_3[157]},
      {stage1_3[53]}
   );
   gpc1_1 gpc166 (
      {stage0_3[158]},
      {stage1_3[54]}
   );
   gpc1_1 gpc167 (
      {stage0_3[159]},
      {stage1_3[55]}
   );
   gpc1_1 gpc168 (
      {stage0_3[160]},
      {stage1_3[56]}
   );
   gpc1_1 gpc169 (
      {stage0_3[161]},
      {stage1_3[57]}
   );
   gpc1_1 gpc170 (
      {stage0_4[91]},
      {stage1_4[68]}
   );
   gpc1_1 gpc171 (
      {stage0_4[92]},
      {stage1_4[69]}
   );
   gpc1_1 gpc172 (
      {stage0_4[93]},
      {stage1_4[70]}
   );
   gpc1_1 gpc173 (
      {stage0_4[94]},
      {stage1_4[71]}
   );
   gpc1_1 gpc174 (
      {stage0_4[95]},
      {stage1_4[72]}
   );
   gpc1_1 gpc175 (
      {stage0_4[96]},
      {stage1_4[73]}
   );
   gpc1_1 gpc176 (
      {stage0_4[97]},
      {stage1_4[74]}
   );
   gpc1_1 gpc177 (
      {stage0_4[98]},
      {stage1_4[75]}
   );
   gpc1_1 gpc178 (
      {stage0_4[99]},
      {stage1_4[76]}
   );
   gpc1_1 gpc179 (
      {stage0_4[100]},
      {stage1_4[77]}
   );
   gpc1_1 gpc180 (
      {stage0_4[101]},
      {stage1_4[78]}
   );
   gpc1_1 gpc181 (
      {stage0_4[102]},
      {stage1_4[79]}
   );
   gpc1_1 gpc182 (
      {stage0_4[103]},
      {stage1_4[80]}
   );
   gpc1_1 gpc183 (
      {stage0_4[104]},
      {stage1_4[81]}
   );
   gpc1_1 gpc184 (
      {stage0_4[105]},
      {stage1_4[82]}
   );
   gpc1_1 gpc185 (
      {stage0_4[106]},
      {stage1_4[83]}
   );
   gpc1_1 gpc186 (
      {stage0_4[107]},
      {stage1_4[84]}
   );
   gpc1_1 gpc187 (
      {stage0_4[108]},
      {stage1_4[85]}
   );
   gpc1_1 gpc188 (
      {stage0_4[109]},
      {stage1_4[86]}
   );
   gpc1_1 gpc189 (
      {stage0_4[110]},
      {stage1_4[87]}
   );
   gpc1_1 gpc190 (
      {stage0_4[111]},
      {stage1_4[88]}
   );
   gpc1_1 gpc191 (
      {stage0_4[112]},
      {stage1_4[89]}
   );
   gpc1_1 gpc192 (
      {stage0_4[113]},
      {stage1_4[90]}
   );
   gpc1_1 gpc193 (
      {stage0_4[114]},
      {stage1_4[91]}
   );
   gpc1_1 gpc194 (
      {stage0_4[115]},
      {stage1_4[92]}
   );
   gpc1_1 gpc195 (
      {stage0_4[116]},
      {stage1_4[93]}
   );
   gpc1_1 gpc196 (
      {stage0_4[117]},
      {stage1_4[94]}
   );
   gpc1_1 gpc197 (
      {stage0_4[118]},
      {stage1_4[95]}
   );
   gpc1_1 gpc198 (
      {stage0_4[119]},
      {stage1_4[96]}
   );
   gpc1_1 gpc199 (
      {stage0_4[120]},
      {stage1_4[97]}
   );
   gpc1_1 gpc200 (
      {stage0_4[121]},
      {stage1_4[98]}
   );
   gpc1_1 gpc201 (
      {stage0_4[122]},
      {stage1_4[99]}
   );
   gpc1_1 gpc202 (
      {stage0_4[123]},
      {stage1_4[100]}
   );
   gpc1_1 gpc203 (
      {stage0_4[124]},
      {stage1_4[101]}
   );
   gpc1_1 gpc204 (
      {stage0_4[125]},
      {stage1_4[102]}
   );
   gpc1_1 gpc205 (
      {stage0_4[126]},
      {stage1_4[103]}
   );
   gpc1_1 gpc206 (
      {stage0_4[127]},
      {stage1_4[104]}
   );
   gpc1_1 gpc207 (
      {stage0_4[128]},
      {stage1_4[105]}
   );
   gpc1_1 gpc208 (
      {stage0_4[129]},
      {stage1_4[106]}
   );
   gpc1_1 gpc209 (
      {stage0_4[130]},
      {stage1_4[107]}
   );
   gpc1_1 gpc210 (
      {stage0_4[131]},
      {stage1_4[108]}
   );
   gpc1_1 gpc211 (
      {stage0_4[132]},
      {stage1_4[109]}
   );
   gpc1_1 gpc212 (
      {stage0_4[133]},
      {stage1_4[110]}
   );
   gpc1_1 gpc213 (
      {stage0_4[134]},
      {stage1_4[111]}
   );
   gpc1_1 gpc214 (
      {stage0_4[135]},
      {stage1_4[112]}
   );
   gpc1_1 gpc215 (
      {stage0_4[136]},
      {stage1_4[113]}
   );
   gpc1_1 gpc216 (
      {stage0_4[137]},
      {stage1_4[114]}
   );
   gpc1_1 gpc217 (
      {stage0_4[138]},
      {stage1_4[115]}
   );
   gpc1_1 gpc218 (
      {stage0_4[139]},
      {stage1_4[116]}
   );
   gpc1_1 gpc219 (
      {stage0_4[140]},
      {stage1_4[117]}
   );
   gpc1_1 gpc220 (
      {stage0_4[141]},
      {stage1_4[118]}
   );
   gpc1_1 gpc221 (
      {stage0_4[142]},
      {stage1_4[119]}
   );
   gpc1_1 gpc222 (
      {stage0_4[143]},
      {stage1_4[120]}
   );
   gpc1_1 gpc223 (
      {stage0_4[144]},
      {stage1_4[121]}
   );
   gpc1_1 gpc224 (
      {stage0_4[145]},
      {stage1_4[122]}
   );
   gpc1_1 gpc225 (
      {stage0_4[146]},
      {stage1_4[123]}
   );
   gpc1_1 gpc226 (
      {stage0_4[147]},
      {stage1_4[124]}
   );
   gpc1_1 gpc227 (
      {stage0_4[148]},
      {stage1_4[125]}
   );
   gpc1_1 gpc228 (
      {stage0_4[149]},
      {stage1_4[126]}
   );
   gpc1_1 gpc229 (
      {stage0_4[150]},
      {stage1_4[127]}
   );
   gpc1_1 gpc230 (
      {stage0_4[151]},
      {stage1_4[128]}
   );
   gpc1_1 gpc231 (
      {stage0_4[152]},
      {stage1_4[129]}
   );
   gpc1_1 gpc232 (
      {stage0_4[153]},
      {stage1_4[130]}
   );
   gpc1_1 gpc233 (
      {stage0_4[154]},
      {stage1_4[131]}
   );
   gpc1_1 gpc234 (
      {stage0_4[155]},
      {stage1_4[132]}
   );
   gpc1_1 gpc235 (
      {stage0_4[156]},
      {stage1_4[133]}
   );
   gpc1_1 gpc236 (
      {stage0_4[157]},
      {stage1_4[134]}
   );
   gpc1_1 gpc237 (
      {stage0_4[158]},
      {stage1_4[135]}
   );
   gpc1_1 gpc238 (
      {stage0_4[159]},
      {stage1_4[136]}
   );
   gpc1_1 gpc239 (
      {stage0_4[160]},
      {stage1_4[137]}
   );
   gpc1_1 gpc240 (
      {stage0_4[161]},
      {stage1_4[138]}
   );
   gpc1_1 gpc241 (
      {stage0_5[160]},
      {stage1_5[66]}
   );
   gpc1_1 gpc242 (
      {stage0_5[161]},
      {stage1_5[67]}
   );
   gpc1_1 gpc243 (
      {stage0_6[92]},
      {stage1_6[42]}
   );
   gpc1_1 gpc244 (
      {stage0_6[93]},
      {stage1_6[43]}
   );
   gpc1_1 gpc245 (
      {stage0_6[94]},
      {stage1_6[44]}
   );
   gpc1_1 gpc246 (
      {stage0_6[95]},
      {stage1_6[45]}
   );
   gpc1_1 gpc247 (
      {stage0_6[96]},
      {stage1_6[46]}
   );
   gpc1_1 gpc248 (
      {stage0_6[97]},
      {stage1_6[47]}
   );
   gpc1_1 gpc249 (
      {stage0_6[98]},
      {stage1_6[48]}
   );
   gpc1_1 gpc250 (
      {stage0_6[99]},
      {stage1_6[49]}
   );
   gpc1_1 gpc251 (
      {stage0_6[100]},
      {stage1_6[50]}
   );
   gpc1_1 gpc252 (
      {stage0_6[101]},
      {stage1_6[51]}
   );
   gpc1_1 gpc253 (
      {stage0_6[102]},
      {stage1_6[52]}
   );
   gpc1_1 gpc254 (
      {stage0_6[103]},
      {stage1_6[53]}
   );
   gpc1_1 gpc255 (
      {stage0_6[104]},
      {stage1_6[54]}
   );
   gpc1_1 gpc256 (
      {stage0_6[105]},
      {stage1_6[55]}
   );
   gpc1_1 gpc257 (
      {stage0_6[106]},
      {stage1_6[56]}
   );
   gpc1_1 gpc258 (
      {stage0_6[107]},
      {stage1_6[57]}
   );
   gpc1_1 gpc259 (
      {stage0_6[108]},
      {stage1_6[58]}
   );
   gpc1_1 gpc260 (
      {stage0_6[109]},
      {stage1_6[59]}
   );
   gpc1_1 gpc261 (
      {stage0_6[110]},
      {stage1_6[60]}
   );
   gpc1_1 gpc262 (
      {stage0_6[111]},
      {stage1_6[61]}
   );
   gpc1_1 gpc263 (
      {stage0_6[112]},
      {stage1_6[62]}
   );
   gpc1_1 gpc264 (
      {stage0_6[113]},
      {stage1_6[63]}
   );
   gpc1_1 gpc265 (
      {stage0_6[114]},
      {stage1_6[64]}
   );
   gpc1_1 gpc266 (
      {stage0_6[115]},
      {stage1_6[65]}
   );
   gpc1_1 gpc267 (
      {stage0_6[116]},
      {stage1_6[66]}
   );
   gpc1_1 gpc268 (
      {stage0_6[117]},
      {stage1_6[67]}
   );
   gpc1_1 gpc269 (
      {stage0_6[118]},
      {stage1_6[68]}
   );
   gpc1_1 gpc270 (
      {stage0_6[119]},
      {stage1_6[69]}
   );
   gpc1_1 gpc271 (
      {stage0_6[120]},
      {stage1_6[70]}
   );
   gpc1_1 gpc272 (
      {stage0_6[121]},
      {stage1_6[71]}
   );
   gpc1_1 gpc273 (
      {stage0_6[122]},
      {stage1_6[72]}
   );
   gpc1_1 gpc274 (
      {stage0_6[123]},
      {stage1_6[73]}
   );
   gpc1_1 gpc275 (
      {stage0_6[124]},
      {stage1_6[74]}
   );
   gpc1_1 gpc276 (
      {stage0_6[125]},
      {stage1_6[75]}
   );
   gpc1_1 gpc277 (
      {stage0_6[126]},
      {stage1_6[76]}
   );
   gpc1_1 gpc278 (
      {stage0_6[127]},
      {stage1_6[77]}
   );
   gpc1_1 gpc279 (
      {stage0_6[128]},
      {stage1_6[78]}
   );
   gpc1_1 gpc280 (
      {stage0_6[129]},
      {stage1_6[79]}
   );
   gpc1_1 gpc281 (
      {stage0_6[130]},
      {stage1_6[80]}
   );
   gpc1_1 gpc282 (
      {stage0_6[131]},
      {stage1_6[81]}
   );
   gpc1_1 gpc283 (
      {stage0_6[132]},
      {stage1_6[82]}
   );
   gpc1_1 gpc284 (
      {stage0_6[133]},
      {stage1_6[83]}
   );
   gpc1_1 gpc285 (
      {stage0_6[134]},
      {stage1_6[84]}
   );
   gpc1_1 gpc286 (
      {stage0_6[135]},
      {stage1_6[85]}
   );
   gpc1_1 gpc287 (
      {stage0_6[136]},
      {stage1_6[86]}
   );
   gpc1_1 gpc288 (
      {stage0_6[137]},
      {stage1_6[87]}
   );
   gpc1_1 gpc289 (
      {stage0_6[138]},
      {stage1_6[88]}
   );
   gpc1_1 gpc290 (
      {stage0_6[139]},
      {stage1_6[89]}
   );
   gpc1_1 gpc291 (
      {stage0_6[140]},
      {stage1_6[90]}
   );
   gpc1_1 gpc292 (
      {stage0_6[141]},
      {stage1_6[91]}
   );
   gpc1_1 gpc293 (
      {stage0_6[142]},
      {stage1_6[92]}
   );
   gpc1_1 gpc294 (
      {stage0_6[143]},
      {stage1_6[93]}
   );
   gpc1_1 gpc295 (
      {stage0_6[144]},
      {stage1_6[94]}
   );
   gpc1_1 gpc296 (
      {stage0_6[145]},
      {stage1_6[95]}
   );
   gpc1_1 gpc297 (
      {stage0_6[146]},
      {stage1_6[96]}
   );
   gpc1_1 gpc298 (
      {stage0_6[147]},
      {stage1_6[97]}
   );
   gpc1_1 gpc299 (
      {stage0_6[148]},
      {stage1_6[98]}
   );
   gpc1_1 gpc300 (
      {stage0_6[149]},
      {stage1_6[99]}
   );
   gpc1_1 gpc301 (
      {stage0_6[150]},
      {stage1_6[100]}
   );
   gpc1_1 gpc302 (
      {stage0_6[151]},
      {stage1_6[101]}
   );
   gpc1_1 gpc303 (
      {stage0_6[152]},
      {stage1_6[102]}
   );
   gpc1_1 gpc304 (
      {stage0_6[153]},
      {stage1_6[103]}
   );
   gpc1_1 gpc305 (
      {stage0_6[154]},
      {stage1_6[104]}
   );
   gpc1_1 gpc306 (
      {stage0_6[155]},
      {stage1_6[105]}
   );
   gpc1_1 gpc307 (
      {stage0_6[156]},
      {stage1_6[106]}
   );
   gpc1_1 gpc308 (
      {stage0_6[157]},
      {stage1_6[107]}
   );
   gpc1_1 gpc309 (
      {stage0_6[158]},
      {stage1_6[108]}
   );
   gpc1_1 gpc310 (
      {stage0_6[159]},
      {stage1_6[109]}
   );
   gpc1_1 gpc311 (
      {stage0_6[160]},
      {stage1_6[110]}
   );
   gpc1_1 gpc312 (
      {stage0_6[161]},
      {stage1_6[111]}
   );
   gpc1_1 gpc313 (
      {stage0_7[156]},
      {stage1_7[42]}
   );
   gpc1_1 gpc314 (
      {stage0_7[157]},
      {stage1_7[43]}
   );
   gpc1_1 gpc315 (
      {stage0_7[158]},
      {stage1_7[44]}
   );
   gpc1_1 gpc316 (
      {stage0_7[159]},
      {stage1_7[45]}
   );
   gpc1_1 gpc317 (
      {stage0_7[160]},
      {stage1_7[46]}
   );
   gpc1_1 gpc318 (
      {stage0_7[161]},
      {stage1_7[47]}
   );
   gpc1_1 gpc319 (
      {stage0_8[156]},
      {stage1_8[67]}
   );
   gpc1_1 gpc320 (
      {stage0_8[157]},
      {stage1_8[68]}
   );
   gpc1_1 gpc321 (
      {stage0_8[158]},
      {stage1_8[69]}
   );
   gpc1_1 gpc322 (
      {stage0_8[159]},
      {stage1_8[70]}
   );
   gpc1_1 gpc323 (
      {stage0_8[160]},
      {stage1_8[71]}
   );
   gpc1_1 gpc324 (
      {stage0_8[161]},
      {stage1_8[72]}
   );
   gpc1_1 gpc325 (
      {stage0_10[156]},
      {stage1_10[53]}
   );
   gpc1_1 gpc326 (
      {stage0_10[157]},
      {stage1_10[54]}
   );
   gpc1_1 gpc327 (
      {stage0_10[158]},
      {stage1_10[55]}
   );
   gpc1_1 gpc328 (
      {stage0_10[159]},
      {stage1_10[56]}
   );
   gpc1_1 gpc329 (
      {stage0_10[160]},
      {stage1_10[57]}
   );
   gpc1_1 gpc330 (
      {stage0_10[161]},
      {stage1_10[58]}
   );
   gpc1163_5 gpc331 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc332 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc333 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc334 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc335 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc336 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc337 (
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc606_5 gpc338 (
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc339 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc606_5 gpc340 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc606_5 gpc341 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc606_5 gpc342 (
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc606_5 gpc343 (
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc344 (
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52]},
      {stage1_3[6]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc345 (
      {stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage1_4[48]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[8],stage2_5[8],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc346 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[49]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[9],stage2_5[9],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc347 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[50]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[10],stage2_5[10],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc348 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[51]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[11],stage2_5[11],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc349 (
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_4[52]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[12],stage2_5[12],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc350 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[53]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[13],stage2_5[13],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc351 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[54]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[14],stage2_5[14],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc352 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[55]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[15],stage2_5[15],stage2_4[21],stage2_3[21]}
   );
   gpc606_5 gpc353 (
      {stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[8],stage2_6[16],stage2_5[16],stage2_4[22]}
   );
   gpc606_5 gpc354 (
      {stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[9],stage2_6[17],stage2_5[17],stage2_4[23]}
   );
   gpc606_5 gpc355 (
      {stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[10],stage2_6[18],stage2_5[18],stage2_4[24]}
   );
   gpc606_5 gpc356 (
      {stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77], stage1_4[78], stage1_4[79]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[11],stage2_6[19],stage2_5[19],stage2_4[25]}
   );
   gpc606_5 gpc357 (
      {stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[12],stage2_6[20],stage2_5[20],stage2_4[26]}
   );
   gpc606_5 gpc358 (
      {stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[13],stage2_6[21],stage2_5[21],stage2_4[27]}
   );
   gpc606_5 gpc359 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96], stage1_4[97]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[14],stage2_6[22],stage2_5[22],stage2_4[28]}
   );
   gpc606_5 gpc360 (
      {stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101], stage1_4[102], stage1_4[103]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[15],stage2_6[23],stage2_5[23],stage2_4[29]}
   );
   gpc606_5 gpc361 (
      {stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107], stage1_4[108], stage1_4[109]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[16],stage2_6[24],stage2_5[24],stage2_4[30]}
   );
   gpc606_5 gpc362 (
      {stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[17],stage2_6[25],stage2_5[25],stage2_4[31]}
   );
   gpc606_5 gpc363 (
      {stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[18],stage2_6[26],stage2_5[26],stage2_4[32]}
   );
   gpc606_5 gpc364 (
      {stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126], stage1_4[127]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[19],stage2_6[27],stage2_5[27],stage2_4[33]}
   );
   gpc606_5 gpc365 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[12],stage2_7[20],stage2_6[28],stage2_5[28]}
   );
   gpc606_5 gpc366 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[13],stage2_7[21],stage2_6[29],stage2_5[29]}
   );
   gpc615_5 gpc367 (
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76]},
      {stage1_7[12]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[14],stage2_7[22],stage2_6[30]}
   );
   gpc615_5 gpc368 (
      {stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81]},
      {stage1_7[13]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[15],stage2_7[23],stage2_6[31]}
   );
   gpc615_5 gpc369 (
      {stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85], stage1_6[86]},
      {stage1_7[14]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[4],stage2_8[16],stage2_7[24],stage2_6[32]}
   );
   gpc615_5 gpc370 (
      {stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90], stage1_6[91]},
      {stage1_7[15]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[5],stage2_8[17],stage2_7[25],stage2_6[33]}
   );
   gpc615_5 gpc371 (
      {stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage1_7[16]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[6],stage2_8[18],stage2_7[26],stage2_6[34]}
   );
   gpc615_5 gpc372 (
      {stage1_7[17], stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21]},
      {stage1_8[30]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[5],stage2_9[7],stage2_8[19],stage2_7[27]}
   );
   gpc615_5 gpc373 (
      {stage1_7[22], stage1_7[23], stage1_7[24], stage1_7[25], stage1_7[26]},
      {stage1_8[31]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[6],stage2_9[8],stage2_8[20],stage2_7[28]}
   );
   gpc615_5 gpc374 (
      {stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31]},
      {stage1_8[32]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[7],stage2_9[9],stage2_8[21],stage2_7[29]}
   );
   gpc615_5 gpc375 (
      {stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage1_8[33]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[8],stage2_9[10],stage2_8[22],stage2_7[30]}
   );
   gpc615_5 gpc376 (
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage1_8[34]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[9],stage2_9[11],stage2_8[23],stage2_7[31]}
   );
   gpc615_5 gpc377 (
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46]},
      {stage1_8[35]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[10],stage2_9[12],stage2_8[24],stage2_7[32]}
   );
   gpc606_5 gpc378 (
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[6],stage2_10[11],stage2_9[13],stage2_8[25]}
   );
   gpc606_5 gpc379 (
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[7],stage2_10[12],stage2_9[14],stage2_8[26]}
   );
   gpc606_5 gpc380 (
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[8],stage2_10[13],stage2_9[15],stage2_8[27]}
   );
   gpc606_5 gpc381 (
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[9],stage2_10[14],stage2_9[16],stage2_8[28]}
   );
   gpc606_5 gpc382 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[4],stage2_11[10],stage2_10[15],stage2_9[17]}
   );
   gpc606_5 gpc383 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[5],stage2_11[11],stage2_10[16],stage2_9[18]}
   );
   gpc606_5 gpc384 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[6],stage2_11[12],stage2_10[17],stage2_9[19]}
   );
   gpc606_5 gpc385 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[7],stage2_11[13],stage2_10[18],stage2_9[20]}
   );
   gpc606_5 gpc386 (
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[8],stage2_11[14],stage2_10[19],stage2_9[21]}
   );
   gpc606_5 gpc387 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[9],stage2_11[15],stage2_10[20],stage2_9[22]}
   );
   gpc606_5 gpc388 (
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[6],stage2_12[10],stage2_11[16],stage2_10[21]}
   );
   gpc606_5 gpc389 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[7],stage2_12[11],stage2_11[17],stage2_10[22]}
   );
   gpc615_5 gpc390 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40]},
      {stage1_11[36]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[8],stage2_12[12],stage2_11[18],stage2_10[23]}
   );
   gpc615_5 gpc391 (
      {stage1_10[41], stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45]},
      {stage1_11[37]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[9],stage2_12[13],stage2_11[19],stage2_10[24]}
   );
   gpc615_5 gpc392 (
      {stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50]},
      {stage1_11[38]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[10],stage2_12[14],stage2_11[20],stage2_10[25]}
   );
   gpc615_5 gpc393 (
      {stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55]},
      {stage1_11[39]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[11],stage2_12[15],stage2_11[21],stage2_10[26]}
   );
   gpc1163_5 gpc394 (
      {stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[0]},
      {1'b0},
      {stage2_15[0],stage2_14[6],stage2_13[12],stage2_12[16],stage2_11[22]}
   );
   gpc615_5 gpc395 (
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage1_12[42]},
      {stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6]},
      {stage2_15[1],stage2_14[7],stage2_13[13],stage2_12[17],stage2_11[23]}
   );
   gpc615_5 gpc396 (
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52]},
      {stage1_12[43]},
      {stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12]},
      {stage2_15[2],stage2_14[8],stage2_13[14],stage2_12[18],stage2_11[24]}
   );
   gpc1_1 gpc397 (
      {stage1_0[18]},
      {stage2_0[6]}
   );
   gpc1_1 gpc398 (
      {stage1_0[19]},
      {stage2_0[7]}
   );
   gpc1_1 gpc399 (
      {stage1_0[20]},
      {stage2_0[8]}
   );
   gpc1_1 gpc400 (
      {stage1_0[21]},
      {stage2_0[9]}
   );
   gpc1_1 gpc401 (
      {stage1_0[22]},
      {stage2_0[10]}
   );
   gpc1_1 gpc402 (
      {stage1_0[23]},
      {stage2_0[11]}
   );
   gpc1_1 gpc403 (
      {stage1_0[24]},
      {stage2_0[12]}
   );
   gpc1_1 gpc404 (
      {stage1_0[25]},
      {stage2_0[13]}
   );
   gpc1_1 gpc405 (
      {stage1_0[26]},
      {stage2_0[14]}
   );
   gpc1_1 gpc406 (
      {stage1_0[27]},
      {stage2_0[15]}
   );
   gpc1_1 gpc407 (
      {stage1_0[28]},
      {stage2_0[16]}
   );
   gpc1_1 gpc408 (
      {stage1_0[29]},
      {stage2_0[17]}
   );
   gpc1_1 gpc409 (
      {stage1_0[30]},
      {stage2_0[18]}
   );
   gpc1_1 gpc410 (
      {stage1_1[36]},
      {stage2_1[6]}
   );
   gpc1_1 gpc411 (
      {stage1_1[37]},
      {stage2_1[7]}
   );
   gpc1_1 gpc412 (
      {stage1_1[38]},
      {stage2_1[8]}
   );
   gpc1_1 gpc413 (
      {stage1_1[39]},
      {stage2_1[9]}
   );
   gpc1_1 gpc414 (
      {stage1_1[40]},
      {stage2_1[10]}
   );
   gpc1_1 gpc415 (
      {stage1_1[41]},
      {stage2_1[11]}
   );
   gpc1_1 gpc416 (
      {stage1_1[42]},
      {stage2_1[12]}
   );
   gpc1_1 gpc417 (
      {stage1_1[43]},
      {stage2_1[13]}
   );
   gpc1_1 gpc418 (
      {stage1_1[44]},
      {stage2_1[14]}
   );
   gpc1_1 gpc419 (
      {stage1_1[45]},
      {stage2_1[15]}
   );
   gpc1_1 gpc420 (
      {stage1_1[46]},
      {stage2_1[16]}
   );
   gpc1_1 gpc421 (
      {stage1_1[47]},
      {stage2_1[17]}
   );
   gpc1_1 gpc422 (
      {stage1_1[48]},
      {stage2_1[18]}
   );
   gpc1_1 gpc423 (
      {stage1_1[49]},
      {stage2_1[19]}
   );
   gpc1_1 gpc424 (
      {stage1_1[50]},
      {stage2_1[20]}
   );
   gpc1_1 gpc425 (
      {stage1_1[51]},
      {stage2_1[21]}
   );
   gpc1_1 gpc426 (
      {stage1_1[52]},
      {stage2_1[22]}
   );
   gpc1_1 gpc427 (
      {stage1_2[53]},
      {stage2_2[14]}
   );
   gpc1_1 gpc428 (
      {stage1_2[54]},
      {stage2_2[15]}
   );
   gpc1_1 gpc429 (
      {stage1_2[55]},
      {stage2_2[16]}
   );
   gpc1_1 gpc430 (
      {stage1_2[56]},
      {stage2_2[17]}
   );
   gpc1_1 gpc431 (
      {stage1_2[57]},
      {stage2_2[18]}
   );
   gpc1_1 gpc432 (
      {stage1_2[58]},
      {stage2_2[19]}
   );
   gpc1_1 gpc433 (
      {stage1_2[59]},
      {stage2_2[20]}
   );
   gpc1_1 gpc434 (
      {stage1_2[60]},
      {stage2_2[21]}
   );
   gpc1_1 gpc435 (
      {stage1_2[61]},
      {stage2_2[22]}
   );
   gpc1_1 gpc436 (
      {stage1_2[62]},
      {stage2_2[23]}
   );
   gpc1_1 gpc437 (
      {stage1_2[63]},
      {stage2_2[24]}
   );
   gpc1_1 gpc438 (
      {stage1_2[64]},
      {stage2_2[25]}
   );
   gpc1_1 gpc439 (
      {stage1_2[65]},
      {stage2_2[26]}
   );
   gpc1_1 gpc440 (
      {stage1_3[47]},
      {stage2_3[22]}
   );
   gpc1_1 gpc441 (
      {stage1_3[48]},
      {stage2_3[23]}
   );
   gpc1_1 gpc442 (
      {stage1_3[49]},
      {stage2_3[24]}
   );
   gpc1_1 gpc443 (
      {stage1_3[50]},
      {stage2_3[25]}
   );
   gpc1_1 gpc444 (
      {stage1_3[51]},
      {stage2_3[26]}
   );
   gpc1_1 gpc445 (
      {stage1_3[52]},
      {stage2_3[27]}
   );
   gpc1_1 gpc446 (
      {stage1_3[53]},
      {stage2_3[28]}
   );
   gpc1_1 gpc447 (
      {stage1_3[54]},
      {stage2_3[29]}
   );
   gpc1_1 gpc448 (
      {stage1_3[55]},
      {stage2_3[30]}
   );
   gpc1_1 gpc449 (
      {stage1_3[56]},
      {stage2_3[31]}
   );
   gpc1_1 gpc450 (
      {stage1_3[57]},
      {stage2_3[32]}
   );
   gpc1_1 gpc451 (
      {stage1_4[128]},
      {stage2_4[34]}
   );
   gpc1_1 gpc452 (
      {stage1_4[129]},
      {stage2_4[35]}
   );
   gpc1_1 gpc453 (
      {stage1_4[130]},
      {stage2_4[36]}
   );
   gpc1_1 gpc454 (
      {stage1_4[131]},
      {stage2_4[37]}
   );
   gpc1_1 gpc455 (
      {stage1_4[132]},
      {stage2_4[38]}
   );
   gpc1_1 gpc456 (
      {stage1_4[133]},
      {stage2_4[39]}
   );
   gpc1_1 gpc457 (
      {stage1_4[134]},
      {stage2_4[40]}
   );
   gpc1_1 gpc458 (
      {stage1_4[135]},
      {stage2_4[41]}
   );
   gpc1_1 gpc459 (
      {stage1_4[136]},
      {stage2_4[42]}
   );
   gpc1_1 gpc460 (
      {stage1_4[137]},
      {stage2_4[43]}
   );
   gpc1_1 gpc461 (
      {stage1_4[138]},
      {stage2_4[44]}
   );
   gpc1_1 gpc462 (
      {stage1_5[60]},
      {stage2_5[30]}
   );
   gpc1_1 gpc463 (
      {stage1_5[61]},
      {stage2_5[31]}
   );
   gpc1_1 gpc464 (
      {stage1_5[62]},
      {stage2_5[32]}
   );
   gpc1_1 gpc465 (
      {stage1_5[63]},
      {stage2_5[33]}
   );
   gpc1_1 gpc466 (
      {stage1_5[64]},
      {stage2_5[34]}
   );
   gpc1_1 gpc467 (
      {stage1_5[65]},
      {stage2_5[35]}
   );
   gpc1_1 gpc468 (
      {stage1_5[66]},
      {stage2_5[36]}
   );
   gpc1_1 gpc469 (
      {stage1_5[67]},
      {stage2_5[37]}
   );
   gpc1_1 gpc470 (
      {stage1_6[97]},
      {stage2_6[35]}
   );
   gpc1_1 gpc471 (
      {stage1_6[98]},
      {stage2_6[36]}
   );
   gpc1_1 gpc472 (
      {stage1_6[99]},
      {stage2_6[37]}
   );
   gpc1_1 gpc473 (
      {stage1_6[100]},
      {stage2_6[38]}
   );
   gpc1_1 gpc474 (
      {stage1_6[101]},
      {stage2_6[39]}
   );
   gpc1_1 gpc475 (
      {stage1_6[102]},
      {stage2_6[40]}
   );
   gpc1_1 gpc476 (
      {stage1_6[103]},
      {stage2_6[41]}
   );
   gpc1_1 gpc477 (
      {stage1_6[104]},
      {stage2_6[42]}
   );
   gpc1_1 gpc478 (
      {stage1_6[105]},
      {stage2_6[43]}
   );
   gpc1_1 gpc479 (
      {stage1_6[106]},
      {stage2_6[44]}
   );
   gpc1_1 gpc480 (
      {stage1_6[107]},
      {stage2_6[45]}
   );
   gpc1_1 gpc481 (
      {stage1_6[108]},
      {stage2_6[46]}
   );
   gpc1_1 gpc482 (
      {stage1_6[109]},
      {stage2_6[47]}
   );
   gpc1_1 gpc483 (
      {stage1_6[110]},
      {stage2_6[48]}
   );
   gpc1_1 gpc484 (
      {stage1_6[111]},
      {stage2_6[49]}
   );
   gpc1_1 gpc485 (
      {stage1_7[47]},
      {stage2_7[33]}
   );
   gpc1_1 gpc486 (
      {stage1_8[60]},
      {stage2_8[29]}
   );
   gpc1_1 gpc487 (
      {stage1_8[61]},
      {stage2_8[30]}
   );
   gpc1_1 gpc488 (
      {stage1_8[62]},
      {stage2_8[31]}
   );
   gpc1_1 gpc489 (
      {stage1_8[63]},
      {stage2_8[32]}
   );
   gpc1_1 gpc490 (
      {stage1_8[64]},
      {stage2_8[33]}
   );
   gpc1_1 gpc491 (
      {stage1_8[65]},
      {stage2_8[34]}
   );
   gpc1_1 gpc492 (
      {stage1_8[66]},
      {stage2_8[35]}
   );
   gpc1_1 gpc493 (
      {stage1_8[67]},
      {stage2_8[36]}
   );
   gpc1_1 gpc494 (
      {stage1_8[68]},
      {stage2_8[37]}
   );
   gpc1_1 gpc495 (
      {stage1_8[69]},
      {stage2_8[38]}
   );
   gpc1_1 gpc496 (
      {stage1_8[70]},
      {stage2_8[39]}
   );
   gpc1_1 gpc497 (
      {stage1_8[71]},
      {stage2_8[40]}
   );
   gpc1_1 gpc498 (
      {stage1_8[72]},
      {stage2_8[41]}
   );
   gpc1_1 gpc499 (
      {stage1_9[72]},
      {stage2_9[23]}
   );
   gpc1_1 gpc500 (
      {stage1_9[73]},
      {stage2_9[24]}
   );
   gpc1_1 gpc501 (
      {stage1_9[74]},
      {stage2_9[25]}
   );
   gpc1_1 gpc502 (
      {stage1_9[75]},
      {stage2_9[26]}
   );
   gpc1_1 gpc503 (
      {stage1_9[76]},
      {stage2_9[27]}
   );
   gpc1_1 gpc504 (
      {stage1_9[77]},
      {stage2_9[28]}
   );
   gpc1_1 gpc505 (
      {stage1_9[78]},
      {stage2_9[29]}
   );
   gpc1_1 gpc506 (
      {stage1_10[56]},
      {stage2_10[27]}
   );
   gpc1_1 gpc507 (
      {stage1_10[57]},
      {stage2_10[28]}
   );
   gpc1_1 gpc508 (
      {stage1_10[58]},
      {stage2_10[29]}
   );
   gpc1_1 gpc509 (
      {stage1_12[44]},
      {stage2_12[19]}
   );
   gpc1_1 gpc510 (
      {stage1_12[45]},
      {stage2_12[20]}
   );
   gpc1_1 gpc511 (
      {stage1_12[46]},
      {stage2_12[21]}
   );
   gpc1_1 gpc512 (
      {stage1_12[47]},
      {stage2_12[22]}
   );
   gpc1_1 gpc513 (
      {stage1_12[48]},
      {stage2_12[23]}
   );
   gpc1_1 gpc514 (
      {stage1_12[49]},
      {stage2_12[24]}
   );
   gpc1_1 gpc515 (
      {stage1_12[50]},
      {stage2_12[25]}
   );
   gpc1_1 gpc516 (
      {stage1_12[51]},
      {stage2_12[26]}
   );
   gpc1_1 gpc517 (
      {stage1_12[52]},
      {stage2_12[27]}
   );
   gpc1_1 gpc518 (
      {stage1_13[13]},
      {stage2_13[15]}
   );
   gpc1_1 gpc519 (
      {stage1_13[14]},
      {stage2_13[16]}
   );
   gpc1_1 gpc520 (
      {stage1_13[15]},
      {stage2_13[17]}
   );
   gpc1_1 gpc521 (
      {stage1_13[16]},
      {stage2_13[18]}
   );
   gpc1_1 gpc522 (
      {stage1_13[17]},
      {stage2_13[19]}
   );
   gpc1_1 gpc523 (
      {stage1_13[18]},
      {stage2_13[20]}
   );
   gpc1_1 gpc524 (
      {stage1_13[19]},
      {stage2_13[21]}
   );
   gpc1_1 gpc525 (
      {stage1_13[20]},
      {stage2_13[22]}
   );
   gpc1_1 gpc526 (
      {stage1_13[21]},
      {stage2_13[23]}
   );
   gpc1_1 gpc527 (
      {stage1_13[22]},
      {stage2_13[24]}
   );
   gpc1_1 gpc528 (
      {stage1_13[23]},
      {stage2_13[25]}
   );
   gpc1_1 gpc529 (
      {stage1_13[24]},
      {stage2_13[26]}
   );
   gpc1_1 gpc530 (
      {stage1_13[25]},
      {stage2_13[27]}
   );
   gpc1_1 gpc531 (
      {stage1_13[26]},
      {stage2_13[28]}
   );
   gpc1163_5 gpc532 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc533 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1406_5 gpc534 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc615_5 gpc535 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_3[5]},
      {stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage3_6[0],stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc536 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[7]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[4],stage3_3[4]}
   );
   gpc615_5 gpc537 (
      {stage2_3[11], stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15]},
      {stage2_4[8]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[5],stage3_3[5]}
   );
   gpc615_5 gpc538 (
      {stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20]},
      {stage2_4[9]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[4],stage3_4[6],stage3_3[6]}
   );
   gpc615_5 gpc539 (
      {stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25]},
      {stage2_4[10]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[4],stage3_5[5],stage3_4[7],stage3_3[7]}
   );
   gpc606_5 gpc540 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[4],stage3_6[5],stage3_5[6],stage3_4[8]}
   );
   gpc606_5 gpc541 (
      {stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[5],stage3_6[6],stage3_5[7],stage3_4[9]}
   );
   gpc606_5 gpc542 (
      {stage2_4[23], stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[6],stage3_6[7],stage3_5[8],stage3_4[10]}
   );
   gpc615_5 gpc543 (
      {stage2_4[29], stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33]},
      {stage2_5[24]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[7],stage3_6[8],stage3_5[9],stage3_4[11]}
   );
   gpc615_5 gpc544 (
      {stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37], stage2_4[38]},
      {stage2_5[25]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[8],stage3_6[9],stage3_5[10],stage3_4[12]}
   );
   gpc606_5 gpc545 (
      {stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29], stage2_5[30], stage2_5[31]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[5],stage3_7[9],stage3_6[10],stage3_5[11]}
   );
   gpc606_5 gpc546 (
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[1],stage3_8[6],stage3_7[10],stage3_6[11]}
   );
   gpc615_5 gpc547 (
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40]},
      {stage2_7[6]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[2],stage3_8[7],stage3_7[11],stage3_6[12]}
   );
   gpc615_5 gpc548 (
      {stage2_6[41], stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45]},
      {stage2_7[7]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[3],stage3_8[8],stage3_7[12],stage3_6[13]}
   );
   gpc1343_5 gpc549 (
      {stage2_7[8], stage2_7[9], stage2_7[10]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_9[0], stage2_9[1], stage2_9[2]},
      {stage2_10[0]},
      {stage3_11[0],stage3_10[3],stage3_9[4],stage3_8[9],stage3_7[13]}
   );
   gpc1343_5 gpc550 (
      {stage2_7[11], stage2_7[12], stage2_7[13]},
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_10[1]},
      {stage3_11[1],stage3_10[4],stage3_9[5],stage3_8[10],stage3_7[14]}
   );
   gpc615_5 gpc551 (
      {stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18]},
      {stage2_8[26]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[2],stage3_10[5],stage3_9[6],stage3_8[11],stage3_7[15]}
   );
   gpc615_5 gpc552 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage2_8[27]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[3],stage3_10[6],stage3_9[7],stage3_8[12],stage3_7[16]}
   );
   gpc615_5 gpc553 (
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28]},
      {stage2_8[28]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[4],stage3_10[7],stage3_9[8],stage3_8[13],stage3_7[17]}
   );
   gpc615_5 gpc554 (
      {stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33]},
      {stage2_8[29]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[5],stage3_10[8],stage3_9[9],stage3_8[14],stage3_7[18]}
   );
   gpc606_5 gpc555 (
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6], stage2_10[7]},
      {stage3_12[0],stage3_11[6],stage3_10[9],stage3_9[10],stage3_8[15]}
   );
   gpc606_5 gpc556 (
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12], stage2_10[13]},
      {stage3_12[1],stage3_11[7],stage3_10[10],stage3_9[11],stage3_8[16]}
   );
   gpc606_5 gpc557 (
      {stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[8],stage3_10[11]}
   );
   gpc615_5 gpc558 (
      {stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24]},
      {stage2_11[0]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[9],stage3_10[12]}
   );
   gpc615_5 gpc559 (
      {stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage2_11[1]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[2],stage3_12[4],stage3_11[10],stage3_10[13]}
   );
   gpc615_5 gpc560 (
      {stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_12[18]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[3],stage3_12[5],stage3_11[11]}
   );
   gpc615_5 gpc561 (
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[19]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[4],stage3_12[6],stage3_11[12]}
   );
   gpc615_5 gpc562 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16]},
      {stage2_12[20]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[5],stage3_12[7],stage3_11[13]}
   );
   gpc615_5 gpc563 (
      {stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage2_12[21]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[6],stage3_13[6],stage3_12[8],stage3_11[14]}
   );
   gpc606_5 gpc564 (
      {stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[4],stage3_14[7],stage3_13[7],stage3_12[9]}
   );
   gpc1_1 gpc565 (
      {stage2_0[9]},
      {stage3_0[2]}
   );
   gpc1_1 gpc566 (
      {stage2_0[10]},
      {stage3_0[3]}
   );
   gpc1_1 gpc567 (
      {stage2_0[11]},
      {stage3_0[4]}
   );
   gpc1_1 gpc568 (
      {stage2_0[12]},
      {stage3_0[5]}
   );
   gpc1_1 gpc569 (
      {stage2_0[13]},
      {stage3_0[6]}
   );
   gpc1_1 gpc570 (
      {stage2_0[14]},
      {stage3_0[7]}
   );
   gpc1_1 gpc571 (
      {stage2_0[15]},
      {stage3_0[8]}
   );
   gpc1_1 gpc572 (
      {stage2_0[16]},
      {stage3_0[9]}
   );
   gpc1_1 gpc573 (
      {stage2_0[17]},
      {stage3_0[10]}
   );
   gpc1_1 gpc574 (
      {stage2_0[18]},
      {stage3_0[11]}
   );
   gpc1_1 gpc575 (
      {stage2_1[12]},
      {stage3_1[3]}
   );
   gpc1_1 gpc576 (
      {stage2_1[13]},
      {stage3_1[4]}
   );
   gpc1_1 gpc577 (
      {stage2_1[14]},
      {stage3_1[5]}
   );
   gpc1_1 gpc578 (
      {stage2_1[15]},
      {stage3_1[6]}
   );
   gpc1_1 gpc579 (
      {stage2_1[16]},
      {stage3_1[7]}
   );
   gpc1_1 gpc580 (
      {stage2_1[17]},
      {stage3_1[8]}
   );
   gpc1_1 gpc581 (
      {stage2_1[18]},
      {stage3_1[9]}
   );
   gpc1_1 gpc582 (
      {stage2_1[19]},
      {stage3_1[10]}
   );
   gpc1_1 gpc583 (
      {stage2_1[20]},
      {stage3_1[11]}
   );
   gpc1_1 gpc584 (
      {stage2_1[21]},
      {stage3_1[12]}
   );
   gpc1_1 gpc585 (
      {stage2_1[22]},
      {stage3_1[13]}
   );
   gpc1_1 gpc586 (
      {stage2_2[12]},
      {stage3_2[4]}
   );
   gpc1_1 gpc587 (
      {stage2_2[13]},
      {stage3_2[5]}
   );
   gpc1_1 gpc588 (
      {stage2_2[14]},
      {stage3_2[6]}
   );
   gpc1_1 gpc589 (
      {stage2_2[15]},
      {stage3_2[7]}
   );
   gpc1_1 gpc590 (
      {stage2_2[16]},
      {stage3_2[8]}
   );
   gpc1_1 gpc591 (
      {stage2_2[17]},
      {stage3_2[9]}
   );
   gpc1_1 gpc592 (
      {stage2_2[18]},
      {stage3_2[10]}
   );
   gpc1_1 gpc593 (
      {stage2_2[19]},
      {stage3_2[11]}
   );
   gpc1_1 gpc594 (
      {stage2_2[20]},
      {stage3_2[12]}
   );
   gpc1_1 gpc595 (
      {stage2_2[21]},
      {stage3_2[13]}
   );
   gpc1_1 gpc596 (
      {stage2_2[22]},
      {stage3_2[14]}
   );
   gpc1_1 gpc597 (
      {stage2_2[23]},
      {stage3_2[15]}
   );
   gpc1_1 gpc598 (
      {stage2_2[24]},
      {stage3_2[16]}
   );
   gpc1_1 gpc599 (
      {stage2_2[25]},
      {stage3_2[17]}
   );
   gpc1_1 gpc600 (
      {stage2_2[26]},
      {stage3_2[18]}
   );
   gpc1_1 gpc601 (
      {stage2_3[26]},
      {stage3_3[8]}
   );
   gpc1_1 gpc602 (
      {stage2_3[27]},
      {stage3_3[9]}
   );
   gpc1_1 gpc603 (
      {stage2_3[28]},
      {stage3_3[10]}
   );
   gpc1_1 gpc604 (
      {stage2_3[29]},
      {stage3_3[11]}
   );
   gpc1_1 gpc605 (
      {stage2_3[30]},
      {stage3_3[12]}
   );
   gpc1_1 gpc606 (
      {stage2_3[31]},
      {stage3_3[13]}
   );
   gpc1_1 gpc607 (
      {stage2_3[32]},
      {stage3_3[14]}
   );
   gpc1_1 gpc608 (
      {stage2_4[39]},
      {stage3_4[13]}
   );
   gpc1_1 gpc609 (
      {stage2_4[40]},
      {stage3_4[14]}
   );
   gpc1_1 gpc610 (
      {stage2_4[41]},
      {stage3_4[15]}
   );
   gpc1_1 gpc611 (
      {stage2_4[42]},
      {stage3_4[16]}
   );
   gpc1_1 gpc612 (
      {stage2_4[43]},
      {stage3_4[17]}
   );
   gpc1_1 gpc613 (
      {stage2_4[44]},
      {stage3_4[18]}
   );
   gpc1_1 gpc614 (
      {stage2_5[32]},
      {stage3_5[12]}
   );
   gpc1_1 gpc615 (
      {stage2_5[33]},
      {stage3_5[13]}
   );
   gpc1_1 gpc616 (
      {stage2_5[34]},
      {stage3_5[14]}
   );
   gpc1_1 gpc617 (
      {stage2_5[35]},
      {stage3_5[15]}
   );
   gpc1_1 gpc618 (
      {stage2_5[36]},
      {stage3_5[16]}
   );
   gpc1_1 gpc619 (
      {stage2_5[37]},
      {stage3_5[17]}
   );
   gpc1_1 gpc620 (
      {stage2_6[46]},
      {stage3_6[14]}
   );
   gpc1_1 gpc621 (
      {stage2_6[47]},
      {stage3_6[15]}
   );
   gpc1_1 gpc622 (
      {stage2_6[48]},
      {stage3_6[16]}
   );
   gpc1_1 gpc623 (
      {stage2_6[49]},
      {stage3_6[17]}
   );
   gpc1_1 gpc624 (
      {stage2_11[22]},
      {stage3_11[15]}
   );
   gpc1_1 gpc625 (
      {stage2_11[23]},
      {stage3_11[16]}
   );
   gpc1_1 gpc626 (
      {stage2_11[24]},
      {stage3_11[17]}
   );
   gpc1_1 gpc627 (
      {stage2_13[24]},
      {stage3_13[8]}
   );
   gpc1_1 gpc628 (
      {stage2_13[25]},
      {stage3_13[9]}
   );
   gpc1_1 gpc629 (
      {stage2_13[26]},
      {stage3_13[10]}
   );
   gpc1_1 gpc630 (
      {stage2_13[27]},
      {stage3_13[11]}
   );
   gpc1_1 gpc631 (
      {stage2_13[28]},
      {stage3_13[12]}
   );
   gpc1_1 gpc632 (
      {stage2_14[6]},
      {stage3_14[8]}
   );
   gpc1_1 gpc633 (
      {stage2_14[7]},
      {stage3_14[9]}
   );
   gpc1_1 gpc634 (
      {stage2_14[8]},
      {stage3_14[10]}
   );
   gpc1_1 gpc635 (
      {stage2_15[0]},
      {stage3_15[5]}
   );
   gpc1_1 gpc636 (
      {stage2_15[1]},
      {stage3_15[6]}
   );
   gpc1_1 gpc637 (
      {stage2_15[2]},
      {stage3_15[7]}
   );
   gpc606_5 gpc638 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc639 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc640 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc641 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[2],stage4_4[3]}
   );
   gpc606_5 gpc642 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[1],stage4_6[1],stage4_5[3],stage4_4[4]}
   );
   gpc606_5 gpc643 (
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[2],stage4_6[2],stage4_5[4],stage4_4[5]}
   );
   gpc606_5 gpc644 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[3],stage4_7[3],stage4_6[3],stage4_5[5]}
   );
   gpc606_5 gpc645 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[4],stage4_7[4],stage4_6[4],stage4_5[6]}
   );
   gpc606_5 gpc646 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[5],stage4_7[5],stage4_6[5],stage4_5[7]}
   );
   gpc2135_5 gpc647 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[3],stage4_8[6]}
   );
   gpc2135_5 gpc648 (
      {stage3_8[5], stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9]},
      {stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_10[1]},
      {stage3_11[2], stage3_11[3]},
      {stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[4],stage4_8[7]}
   );
   gpc606_5 gpc649 (
      {stage3_8[10], stage3_8[11], stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15]},
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[5],stage4_8[8]}
   );
   gpc606_5 gpc650 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage3_11[4], stage3_11[5], stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9]},
      {stage4_13[0],stage4_12[3],stage4_11[3],stage4_10[3],stage4_9[6]}
   );
   gpc1325_5 gpc651 (
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12]},
      {stage3_11[10], stage3_11[11]},
      {stage3_12[0], stage3_12[1], stage3_12[2]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[1],stage4_12[4],stage4_11[4],stage4_10[4]}
   );
   gpc606_5 gpc652 (
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6]},
      {stage4_15[0],stage4_14[1],stage4_13[2],stage4_12[5],stage4_11[5]}
   );
   gpc615_5 gpc653 (
      {stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7]},
      {stage3_13[7]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[2],stage4_13[3],stage4_12[6]}
   );
   gpc606_5 gpc654 (
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], 1'b0},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[3],stage4_13[4]}
   );
   gpc1_1 gpc655 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc656 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc657 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc658 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc659 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc660 (
      {stage3_0[11]},
      {stage4_0[6]}
   );
   gpc1_1 gpc661 (
      {stage3_1[12]},
      {stage4_1[3]}
   );
   gpc1_1 gpc662 (
      {stage3_1[13]},
      {stage4_1[4]}
   );
   gpc1_1 gpc663 (
      {stage3_2[6]},
      {stage4_2[3]}
   );
   gpc1_1 gpc664 (
      {stage3_2[7]},
      {stage4_2[4]}
   );
   gpc1_1 gpc665 (
      {stage3_2[8]},
      {stage4_2[5]}
   );
   gpc1_1 gpc666 (
      {stage3_2[9]},
      {stage4_2[6]}
   );
   gpc1_1 gpc667 (
      {stage3_2[10]},
      {stage4_2[7]}
   );
   gpc1_1 gpc668 (
      {stage3_2[11]},
      {stage4_2[8]}
   );
   gpc1_1 gpc669 (
      {stage3_2[12]},
      {stage4_2[9]}
   );
   gpc1_1 gpc670 (
      {stage3_2[13]},
      {stage4_2[10]}
   );
   gpc1_1 gpc671 (
      {stage3_2[14]},
      {stage4_2[11]}
   );
   gpc1_1 gpc672 (
      {stage3_2[15]},
      {stage4_2[12]}
   );
   gpc1_1 gpc673 (
      {stage3_2[16]},
      {stage4_2[13]}
   );
   gpc1_1 gpc674 (
      {stage3_2[17]},
      {stage4_2[14]}
   );
   gpc1_1 gpc675 (
      {stage3_2[18]},
      {stage4_2[15]}
   );
   gpc1_1 gpc676 (
      {stage3_3[12]},
      {stage4_3[3]}
   );
   gpc1_1 gpc677 (
      {stage3_3[13]},
      {stage4_3[4]}
   );
   gpc1_1 gpc678 (
      {stage3_3[14]},
      {stage4_3[5]}
   );
   gpc1_1 gpc679 (
      {stage3_4[18]},
      {stage4_4[6]}
   );
   gpc1_1 gpc680 (
      {stage3_7[18]},
      {stage4_7[6]}
   );
   gpc1_1 gpc681 (
      {stage3_8[16]},
      {stage4_8[9]}
   );
   gpc1_1 gpc682 (
      {stage3_10[13]},
      {stage4_10[5]}
   );
   gpc1_1 gpc683 (
      {stage3_12[8]},
      {stage4_12[7]}
   );
   gpc1_1 gpc684 (
      {stage3_12[9]},
      {stage4_12[8]}
   );
   gpc1_1 gpc685 (
      {stage3_14[6]},
      {stage4_14[4]}
   );
   gpc1_1 gpc686 (
      {stage3_14[7]},
      {stage4_14[5]}
   );
   gpc1_1 gpc687 (
      {stage3_14[8]},
      {stage4_14[6]}
   );
   gpc1_1 gpc688 (
      {stage3_14[9]},
      {stage4_14[7]}
   );
   gpc1_1 gpc689 (
      {stage3_14[10]},
      {stage4_14[8]}
   );
   gpc1_1 gpc690 (
      {stage3_15[6]},
      {stage4_15[3]}
   );
   gpc1_1 gpc691 (
      {stage3_15[7]},
      {stage4_15[4]}
   );
   gpc1_1 gpc692 (
      {stage3_16[0]},
      {stage4_16[2]}
   );
   gpc606_5 gpc693 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc1325_5 gpc694 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4]},
      {stage4_2[6], stage4_2[7]},
      {stage4_3[0], stage4_3[1], stage4_3[2]},
      {stage4_4[0]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc606_5 gpc695 (
      {stage4_2[8], stage4_2[9], stage4_2[10], stage4_2[11], stage4_2[12], stage4_2[13]},
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5], stage4_4[6]},
      {stage5_6[0],stage5_5[1],stage5_4[2],stage5_3[2],stage5_2[2]}
   );
   gpc615_5 gpc696 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[2]}
   );
   gpc615_5 gpc697 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[6]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[1],stage5_8[1],stage5_7[1],stage5_6[2]}
   );
   gpc606_5 gpc698 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[2]}
   );
   gpc1406_5 gpc699 (
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[2]}
   );
   gpc2135_5 gpc700 (
      {stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7], stage4_12[8]},
      {stage4_13[1], stage4_13[2], stage4_13[3]},
      {stage4_14[0]},
      {stage4_15[0], stage4_15[1]},
      {stage5_16[0],stage5_15[0],stage5_14[1],stage5_13[2],stage5_12[2]}
   );
   gpc1406_5 gpc701 (
      {stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5], stage4_14[6]},
      {stage4_16[0], stage4_16[1], stage4_16[2], 1'b0},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1],stage5_14[2]}
   );
   gpc1_1 gpc702 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc703 (
      {stage4_2[14]},
      {stage5_2[3]}
   );
   gpc1_1 gpc704 (
      {stage4_2[15]},
      {stage5_2[4]}
   );
   gpc1_1 gpc705 (
      {stage4_3[3]},
      {stage5_3[3]}
   );
   gpc1_1 gpc706 (
      {stage4_3[4]},
      {stage5_3[4]}
   );
   gpc1_1 gpc707 (
      {stage4_3[5]},
      {stage5_3[5]}
   );
   gpc1_1 gpc708 (
      {stage4_5[5]},
      {stage5_5[3]}
   );
   gpc1_1 gpc709 (
      {stage4_5[6]},
      {stage5_5[4]}
   );
   gpc1_1 gpc710 (
      {stage4_5[7]},
      {stage5_5[5]}
   );
   gpc1_1 gpc711 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc712 (
      {stage4_8[7]},
      {stage5_8[3]}
   );
   gpc1_1 gpc713 (
      {stage4_8[8]},
      {stage5_8[4]}
   );
   gpc1_1 gpc714 (
      {stage4_8[9]},
      {stage5_8[5]}
   );
   gpc1_1 gpc715 (
      {stage4_9[6]},
      {stage5_9[3]}
   );
   gpc1_1 gpc716 (
      {stage4_13[4]},
      {stage5_13[3]}
   );
   gpc1_1 gpc717 (
      {stage4_14[7]},
      {stage5_14[3]}
   );
   gpc1_1 gpc718 (
      {stage4_14[8]},
      {stage5_14[4]}
   );
   gpc1_1 gpc719 (
      {stage4_15[2]},
      {stage5_15[2]}
   );
   gpc1_1 gpc720 (
      {stage4_15[3]},
      {stage5_15[3]}
   );
   gpc1_1 gpc721 (
      {stage4_15[4]},
      {stage5_15[4]}
   );
   gpc215_4 gpc722 (
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4]},
      {stage5_3[0]},
      {stage5_4[0], stage5_4[1]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc615_5 gpc723 (
      {stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5]},
      {stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc623_5 gpc724 (
      {stage5_6[0], stage5_6[1], stage5_6[2]},
      {stage5_7[0], stage5_7[1]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc2135_5 gpc725 (
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], 1'b0},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage5_12[0], stage5_12[1]},
      {stage6_13[0],stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[1]}
   );
   gpc615_5 gpc726 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], 1'b0},
      {stage5_14[0]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], 1'b0},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[1]}
   );
   gpc1325_5 gpc727 (
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], 1'b0},
      {1'b0, 1'b0},
      {stage5_16[0], stage5_16[1], 1'b0},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1],stage6_14[1]}
   );
   gpc1_1 gpc728 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc729 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc730 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc731 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc732 (
      {stage5_11[1]},
      {stage6_11[1]}
   );
   gpc1_1 gpc733 (
      {stage5_12[2]},
      {stage6_12[1]}
   );
   gpc1_1 gpc734 (
      {stage5_18[0]},
      {stage6_18[1]}
   );
endmodule

module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor_CLA162_12 compressor_CLA162_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9944525788f0c2ae62e7baf7745a2b4f1d556df011e4ad6ac40fc2026f6c740ecbee65057d07d9d4b1ded1a8abdc79fda25a1798058d739b512e0157000731d50a5ecd16f003afe908a38ed71f53918197f315767f6ac56798f7391313e4156aa89a7b34eddb5931ff5ca24520f276d618786fbbb2c70e44ae7387bd3e580fa607d5398979072cb5f656f7cf6d895c52c0a87dfeea4ea00a1c1943b7fb21699d18017eb7efc66096cee3c1a367a9643724ec1bbd7aefd220cc1275e878a884ec45670aa5604074831671e71876a8f19abc56999de4979235614d2868c9913a25ba28d79d078da1c12d99b6466ae96c753213c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h48e22041f5898e2f0845ac252f486a4cc1c3bccfaa8eeeee0e0a3708ffde1097183af8fe2aefc6a7e546f64c27dec0dbe4162850849c17d44f9ab16bc7466e2861d1d420886bfd6de5d9c571d1d7ea2c76c464c10b2947fd9a748031d9b6aad85f540906ed7acce0a7a17a56b5bc59758e225fb5c296546e5b032e2c78f8e6208187e33b698d8c5c39c4d52a6ae4eaa3ff8ad09856c9abf2c0b06590d5c2cbdd631c62a6b59c8d079adfdbfa15983185a91bae663b645c6fcb6d99087f6af1caf2dbc0056b7d48bd66a3e6f5d0503edc14d3f7493687c87273198ff2511b6586aab508aa38acc3282be6b2f282b296a06b150c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h73f5ba1f3e5c1dfad62b7e73a025ba84fff5bea9c24ff15c4dd9e9defef582336463ef774995d27c461183c4c055e8904c2a7605a44c6a643ed12470e46419262a3d47ed2df372d18ec9a6996f778e2ade6d9cde06936601658356d04fc02f40fb1072c31f3aa5b162ff3d1e3c1389c65f42e184b505c077f3d9da407cea1ab656724214f4f859e5394c9fc7c3c535b367dea31e32ea38a485cc8db7265bf4ec0873a5b3983573613c81ab09acd1863365cd8a9cceb1768480d4882d3fbcd21daa46230422caaf69f51f5cdfbaeb430425ba847d8db33fb80626dca669c5093a9b4df91f9508b1afa3ce854b6b765718b25433;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc5ef6f800a22b514c75475dcdb581352c086feeba4bd756e20d304e35e48056eccad3a8c7b8de154ea061767474c72dc21c13134b9bbfb6e9af980205579ef95e4e9371472c7f084e3c1e0341cbe246b4f1e3dad92eeda76ca36aae380c3614394246a75582e8128e997a04abc491e3e89318f6ffe3d4c04f30b80ebc679f7b5ceaef6b279b6417d27a272b4a81371685944780e5f41534b3b8d8a57189857fe7fab80bd19ce2ff087904159eb4d7b826d134cd31b71f9a6870ad0349bb45f8c03e566a4e0bf3a2b1da0e8a4917fcce50a244e1f1e741a58954b1defce146588e2d5e2201d528ed70d74c9b683643b14db574f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h43f3c68a2a2a4d38b194fb850f1902ab57214ba94644c914877f635e0f1c0102b09b4cd78a3b6fa2700a62c00a30dd0ae6e4d5571530198d772d065a6781e9d04d3d047861a75ecaa2b08757a548ec48c6d1253f7f46038a34755f7a144dbaad62ea6c330d70fdc84b9ea138e976f8cf3ea1caab0c0942240c8668c12d47f9b6c23dd35ee9a97ac0be7449ce0d2c17838babbfe2955685dd2836eeadfb0dbf8cf4b52144f424adae97cc76615ebea418dd8c86f4c04d96cadef4946c960c91013c829e631bcea23a1ada771dec53ce6b13169845b5870b04ea3c709a4b5b2733838d337cc855d829d09dc3e1c43a1addfae9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h432e34313aa8edb873de5a472666ed1a41e749ddbe7e1f326f7f6bd60cf4a9c02aa175eaf0b470c415de4e4b73cbbe461bdd897918f312daec4924ea6e085f9fc6c7a109034724c18674a19d3da5ae9c3b91ee0c1175a31696e625e22296bb91b3ec4aa91d0e7342ff4a62b2592bfdaf7d96708835546373855b27b6389aad38d2a76ea3b8142ff4dbf4e6f5b0529aa8b69d75e5e50bdfb7ce26d845511cd4c04bd8d6c403b6be08c911663eca95480c7d0a7632f90043cf083ca9ae7c93e4d9a9905b9275d5a7ef1fc73f62d69db64426bb702685df5e68a870fe056409b10561d899f14224180153f69e6d8a83805769a03d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h7a1e6f0608d880d6b57f37755105cf6eabe4d87ce6bf2fa216b6c7bdc88c029112ade2ca857fbe13f625032353f0b370e6067514b87cd49f25a32311e8addf77764b9200a61324a47069358b383e3fddbea642f3137ba25cd0ed6b78d7c9eaa15fc035c30dd3f2d32acb060961a03b1e9e0376c0ff264c0d5d21dd4367a78dd04c0eab86431ca1bf8ccc4beb78d57c87e1b0e8ec8ab3ff3449cbaf8048d86aac1aebbc62a59cec1a23024f4ee4ec2db3c1a1d4be96e19580015a545cd373a6b322fca7c20e67a7512793e4d44abca76bcf993b9701514a6a2d6fa6a2c949c87d572217e02661e5faba57e1f0adf65a370c105e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h47f4a1f1e9d8e9a8789c7cb8a59afb1a245f449e17e30d25e8ef26f005f9307b692850346599f5708a55348c6f8e6010a697408b62be85b527884b1a01db5a2743eecf4057a95f6cc583b69182c661acdfcf1ae9e5d27f43686123c46cd894dfde4c35c2f2e2fe31ae7bbb9c01dfa4911b3922b3046a118e5b199a8a5f22bbc17379cd48f313461d7f40e7f0f1e7c09b4e7d69a02ee03b72fbf1fff057b0aeb568c5f19583eb6846c0df65034eaba6e548c554b2119eeee90f6e7d1548cb88238f887b49eb6b223835695356e7ee804c2963e55f17844abf201d5ccf1a243a994520aceb0a120d84afbac9743a79259f5f1ebb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha4c83c2010c06119897a3ee38847599d975c4f9a1798f46baba484b4fde03f0250c2e8c74b66d443cf59be6aaf358dc2c6a95655ca8593e4db59a18ccfd00fcf1ca81c133b3b5989f31d667c3a55b9cf38f03c57dfaf242759e3bbd6e1a456464b023141b021d6f7884374dac707644a1091f574180ea9bd94f22b1e96aaf282bb12353ca026127879b8a7b80f443b92e9591f6bb749bc778078c7bf75bcfea1c80912502cfc0334120708ee8078ccaf4a95954dffdc4b2de069fa7e376b7d6e35be01ba8e695d6dba2c802e3033afcb83b817eb0e43ae1607cd8e0e2042207aa20d8fc1be80a1526d26098010518586f73fd3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h29885ac6e137958f0a4363ec7fad386d87b8a6b585a7f32be549d6d43702de3b6a677d2a131cf2cba29d04b186457ba8a3cf816ff3b6ef61ddb82dc5ffea91633c56fa01be74c34643c61715391853e4f15af3688cd42fd7a8172cd5a1628f7e5972ed1209aa534c2df5aad7c9e243d60dbc94547bdd359ec5e158d05e214bd9e75f22b359ab7aeb0274848c49f4ed2a1fd450330cfbc09c29ba2a0d0b87d8b6830496253d70e719177881ffc433860cead7b2b639297e22ca31fe7504f624abd74a69c5262249e8a407b9477d24f5b05a860fb590db2f8cb52ee5ad8dee3743207c45b694662106e348d54e8b694676a87118;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h13bff150a87e7dd0bb7faab9cab680f1afdd398961c5301638c491073d33df9f83580dc04d4f82d8e050f65962000e78b860a792d7e50a9cf53cbfd8915e6c87f8b71261f1f9ba81199baf3dce040472342bc75ea5a060efcf775c849d7dc162e305453aa73d3ea2e4823e92b933344756b8577fe50179782a19e19b13307ad64a1911966ededf375416739fa799d36ce1f4e39a5d363c1731ee1aa6808f18b60108ba457ae75fedbd550de3133e5a6ffda9e2c32df7fdc31cd3d5e79732d477ca91227f9c95776ad83fac068554381bc5a7fff4eef698462ce54e57c3b5019c6e76f19f2d24cfe8e6d39ebec3a410a09916aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hb8fe66870f29666e3e73892e5356feb9f0bb86eac996f8cf5c156f07c9d195c9d4c1aa47e7f1a7c0580a283966ca5f85b276dd633386efa2e3edd2c209680993aaf3bb17debf429a0cb9e83599c3c98c712418d1e3d950d56be5921912036b0b1f4ca40c18c74165cbf2b1d3a5dec8f0f1a0675f1d09d0af30a5820ba19d2ea5cd7cd058a697765684f2f639759ca4bfbc0063d06fe3594861d9a91f90c4cf3073857c33386a67cfccdf9a2841be82fbe199f2f7911167617d3d9e91661642a4119d4a0df644fbacead71067c169ef65aec59a453b6ea451ba1c0385c4bcbfca2391a36222d23d10d610138a4a47daa892a81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h6e3fe3f0e1ae4e35a6dea077858a6039ae1535eeddd8c9116aec9a3468a6c976c62620cc227420bd6ddb8a5982dbf166bab548699188f2c50f6ecc6bae52f8fcfe97fdd738ed42e61969472066b9de7806e57c713791afb20c4e1a087dc0eb5f54c95426242dcea304d76470cb0e2dc352ee633c07f08d85559427e5b1fd670fc12856f3391bde52225c9a51a9f08b5af1cc4d2c194a66f162d2a6a0b46f10051c5ab9b612afadf9d5b6b74b4ea7a57ff10e0bf10e3143ac21251acf4fa4c6ad61b369761773f416c73e2a4c5ec424f8f3dab6d8fa87a8cfd82b024924f81eee2a7f5e6df14eef43c1d5f73e6de31278c75b8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h92d2c96f1b07224b825dcc28d6977ad988684c9d7836657a44cec471c8fe2f21115f815bc852cec979d899ead9cfd548b7409886ff8f3ca6ae9e7d711451872c8757034632a4c01302877aeaa78afc35f05dcd588e4fbf25888e27601da33f929b769bd1e691aeba55576620b82e8ad81e8b41205fd4f0295d5ea14a1f9fe7080c7fa5649e13591ed86d9bb4df8e71c6afd3271684eeef6edd32658f8d2539a3d1e353806359bd9038bfe0aa9c7de4e16f66c2eee3171c202180d9ab6a0c0f8433593f8bdad67983ee6fefeaa1fb9e7753b76434180da5d5d2f7ef18ab53f6b8206a67e03cd3a4eb22ce997d0b84389154d096;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h45cb419ab9c35625b5904a1ff9c32428bfcec0cc48c15f2b95100692cb4000278639749ac6f2fca565debada6499ba5e347ea9e8dc46e09044496bc83c7518b020c45c5eec49d919e10e155f5b18ccf1291c022b78a5fc62225c751d8f02fcafcbb4a91a3a7b4741bea8c85cf5a372a75b474b57f1bb9d17999c50785c17c82bce843428208a2982e853e96fd1fffc065c4f0bd2deb49c68f5af0f52f36fe22e360335f27cc680d64421a22db0ef07ec16b06dc18b9c9d62dac3b4995518f4959677b5157332a59c5c7b61dcf10616d11f3717177b4cff639a4baedbc681fada22b5897d8d894f57480a145485df1a3bbaeb05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h481c5007bc6e8b65ba78e30618b85cf5b18048acf7ae08fbc9c9a2e218869245b6e97932bfad400f8b3723a1b67c419e5e4134ed39fdbd37423e99a777963e69d505bf69b4e127839ed293b3b99cd30a6111cae8e70b162084105c9df3cca7b8d7b237356fa278000e4fd94a8cb53f784a0d2c941b6d8a4601bf257f4e72db6caecff59fe9996e4ef6e315e6f004c0f0deb85597acdcae6cbbb355479387dc5b2f2e1f3b877589ecc7061384915ba020e6873626dae46853dd4c929f1f712e609e6569b9ca515bfc09c492feb25d454580e09a5d8f0726ffabc12c63ac1bcaa5ba7dfeba3cbecc73534e300d7b472411a19d48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf0219092da537cea2039c5b73f663e8d4ca2dc520da0915943140fb56f8d18a56547469d3ab128823a7d72ef4b957b0f6bfeb2cda8926cfd28fa0bdd31108a842b4e8aa902c3bad4f59b20b8a41a2e427cfbb60344adf292f6ab20f7c2d981a17c5479c5a91660b2db37216500839d2cdd8e5afe49bffe629aa70d79e5c370912f11b418f1a5699a11cf74fc990691ecee62b70efe8a24571361cb15ae4abe2fc731b670f5a964334c66db5ebc4ce2525471a24ea14339f650571204b850faf11022be04906288722c19c01ff91d7822f0c61e8f3ec3f0e3ab9cc5d17ad84b3d2a63d04b41d053c868add1bfc390a3e77fe741;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h149bf68906a3b2ee96d59fcec6ff84b92130b6ecaddec155b6890891e86d3b17e79f60415c0c1b399aa6083e1fb644f2318f8a0b12c4cb11a9a79d054bdf882d445c32e059954a5b988f3546ff702d82a7afc7888053d2de8cadbb17026d23ab89dd70ca1e1d25938fcd88963302db404811fc06feb9b7cb7e373b31242b1410bdd3dc202d69ea0d3613057b7df5ac093399f33fe53754715c903b1fb03735fc388840e1ce48ad2230bcf327929d64aa503fc50652818b60c1cff79acc9105ab0a402465cf901a72b5a13ebf2637087224eb4c3c3af7845ae6c8ffc637a19dad856d5e1e5602a9782d49ddc2ca548443935d2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9da223f23e2896968156f8eadde66b819d2afe0d42b759ade126a6d53e7bd54b5d49d962548dc917b542a5728601bb8bbfe06c2d99f3137884ea3450b2cd0c269b5e07f8440a3f6b1381a8e7b1f0ca418fd11a7734e8f7d332a8beb1269f5386ce06cfa901931c8df7d08699404fba76bc51b3efe1116655039734a3d99408ad30f6fb4667fd2f94b1d17183a5126682b3bbba981825cb8628a2b11654a97a69f5c6b08ca69acdca92678b4f168193fcb2c6dac0e731b3353998f8f5d3bf20709858b7479994ed5f033737c59ba0e6f28e4b6a86ff55ec4f8cc6d2537419ad2ecf2bd9f75c2b5eab8b5baf22565ff246fecdea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h69b214526e4d7ec315de97030ff854c67d65ab183eaa1fdba1d3b6cfac04f8db82f27f60e61c9f14cae1f95188aa362226f322b0b5dcc61acc791441365a5d0f3c8cf6f4219ae8dcae0517f1cddfee0266f7e1c639d2ce1ecc9a60bf9baffeb864b9ccd06d735c7b6232f5434f878c2b6160d592a7c5003dacafb1b81e52815e68fe568d91ac559c093a43fe8547cdef661780cb5d1a38ad34a491fad85d5371f5567aadeb6fa95a2697e1bfbd7dc8b00d4389614216230e2a542bfc7d6852bc807a9acc932b35181fcd4ff816bad7ad093b211ad5adaf676366bf734d899ae8edae1485b47a2372322a164211c70c01331a19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd874dcb1fb59d1b2dd0cd369dcbd0157ef93a40068cd025ffdb39a9bc14b41851dd17e3a15c6b72779efbd16f1aedfeeb0cd46fd61d72ce7ef73a656fb6c9ddc5322e4af9d66b1207f566a6a831834f26aca344d44cd16f02574b5b6b3a984dd0e69b884035549a40213165c3f2f3c41681c8baf6b816b5ab479645e030d8e8d6f22a7ed9a67a49b61dd77dee2eb07ffd32b172ab34e823df0888e0e32864ec1725d020489074261d346255d6d9b1915882739b2eca5fc79c22441e922a51c9dcc8dcf6e71d8de9e83651c3d4e69b3c37ccea401bd23d6055a7c48a991633044c3a7d3615331e84cd8aaec4009239124f4f6d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h199b26097b65c9b95bfec6d97a4b3f01bfadb95ce96b11b269c7c5fbf5b24fa1abc95ec580ab04db44e89b39cc55bb7037e23aac55233655f6c060b16e6a850d959c7648451b4566037b1d908cdddd90a1d7f7be6675548835d5ba32f18e9aeacb79cabbfe9d0c863973cee89dd405a04005f7c51e25d5a0f24c0b239b0ffdc98f3d65ffe128623d738846141024066f41506b54854d900fd5dffb2c21464e28e7d508f8d0d7ab875824132319203cb3b9e8acd3b4e8835c17566f826ef3360d40cc8bee1853ea3fb75c96dd47d3a3ecd181e9fc7aba7ff318e8de184d6415ebe2c91cd8cc18f0dc2b632898913ef76568a1dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h88abe437be673c3d14a94c78e5ed093a72f178fe8ebd88b8fc2488f785a7bbb4f00f8f3d5a830c8e2ee6d261dc7d1579df9d5924034b574931ccacdd787b23d4e41e1d4909b903ddad8ee28a828bded8807927f9718f46810e8bd87422db655d40c7092844a63c897059d73e09e8d8eefa0924dc3870ddf67d7770f7d81f71efaf6a624366a081a0b20e06430560c7ad138c70881427af1b4e80b20bb7cfaa2d727c9dc79e57c22641d970b9b2c00f9ff34d25fa7b8958a07450065c4ad918b156edeb573a47f990fdda882d5b3e7a57e12f4f0ca880a92e1a5988a9802aff7e2bd02cdc63f4287e8ed1509a6484e7d7f58902;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc99c597bb894f6be22f0a391b644495063ea92428061e25c1d24d89bfd49d981a9c6e3946b4c3920e9e8b0f2829eac2f1b75b96cd58ae3760156ad00089e2d45e024d54b47f17a23d748b061cac9409f948a08e02038a11b6d8ab51a85c0b1ec43bb557d6edadf0db945758c94f61c7eabaef1249ba5dfe2efb1a438d99e55683568bae3060ee743769be4ba0024345f8b7e10a340d3137af49a09e6af8a0bf34a2306341aa91cbda6efbb5c8e8b373b1c748dde06c9224bbab1f30e4bd94b9830b9d49486cd75430e3653e4decc4deb51f14d392ac849298d49a7f4742462544b5a2c9e5c2c149bda573adfb8bda8cb887404;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2e8cfcc450417b040a4e3371fd05b50511c887d8e8430a3d691f671fd8fa4792a6f506625c999ad1572823b36d1bd7f3bf204c66e912812e964831b43334844f6fa35b7ddd4d186c342717052116e72337d146adb10e42215d702e0b2a711ad944baee2f7ca465dd7f0ad8a0eb8fdaf582c844e28bf391fe006b459191ae22160aef5491417ac95eab965dc4f5605dc37a44bf7d704baf4a7631da7490700b111c0ef76c7876f8e47b0ceed44a759fe7f2e316683e28cdd19e5ed57a156534fb4661445b5dafafe4e37de9bc748396b834d9320f6bb3f6057aa1bf28b973fc763a01d2935c7991bca4bf7f1bef72eced5b391c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h896f0b03f97c61b33f80d6c544ae2af629a7e73505509ef8935ad009f85a72cb231d2a324cfc70239973b70fe7838d47cbc41e0857eaa50ced863974fc00e3008691eee1b9f159930d0d622c08b9cd0ed2049f34fa70eae5462ffe74ff4afa595840706402f7d6270a6fe753316b957d29b37674474f93923df915db9985d62da9f2c8528740301a749b11135a95db60f66bfa5744954de6be17f1bb1ac00b35d8a33a753eeaff7a3c95d641493b2d026a8bed0f270bc9fceb2900a3efae8374a96811818ebf071c226f712f6ca6ee9c4904213d54fc75e7d5ca29bc63a65f5a841c01e29619c6cb52e8de350fa7d01614a554;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h1a50309de00f0320ac5e6dec6f4f48c8ba2a221eea0098c90c2ee9b36c0f19a9b7fc6ae99ab3671ed6bd89efa2f1a36d34e4fa9e67ef087bed76d20a8f05933cef331af95e41cefda90e250ebcf5dceffbf0efe9c6a9bdac1d3cecc2631970492dae950e9cb0526d5252568746b46d19acf469aa4cafbf05eb862ffe0c87fcf424c2142c3ff7fa400dcd4abf4e326b57e0865e1d117b1120e337de7ad388181cf9ef755e83fef06f10393ca152dd52d28d1132ae26a0ae572be6c3680c3b7e5a0e2030503f1be3d2b22c99142643617ac95d271f4ae59d9dc4cc4436018f6bbf38afe2d51e923f691c7f4c086e1a06fdef89da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h62da13ea876eb01c5ee38c0955986994cdc43d919d19dbf453e7e1be8d069291ff46a86dddbeda94d6e50af5eb92f664f696ea5fde7be4157b7838e8f72a98d56db34e2043acfb4b7054785055559ba13afe4a910e2f01d17bcdf43eecb86c56c9dc2c6e26098ab0164f9c11b80c36fd368cca49698768171ed6cd18231c598550ffabd84bed47e37c5cf13029510decfce230a1128642ee6dd8e0a3368dc51a56d5e6a2cfb735c604210adefec616786e50c6d719d0b7342f3668aae3b3e109a6841911e7ffc48aacbc327718d2a06790422f938fccc4615e8911f22d6911b108875b8bae0ea5081d4ea8eede2daeeaea312d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h982327c03fcc9ef779a6ee157d7b72b341694d0e4c9a9c54a1a969b8f534b209899c48b573f1c160944518510419019f4ecd28c31cc8399228520392210b880a7b5f251c01a6364d2b4552d960aa92735365913d229201e86ed4af20dd52d49c5909cd27d583ae29429bd98d125bb99af6b5232cda70c94a9f6236a82ba5394ab886c099adc89d16249e1c4fa5fe10a209085ddb1d78d0c0e7f1c0fca91a902f6fe625cc0591697805541a366c13868d777711f2f138cc3f53e01daf79d013d5d31701cc173e473aa2fc34f3a5c1b4857f63e9e5d6f62ec955ba52ea8d1819539932fb3393f00570122811511d2066f3d84ad7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hdad1dd076bff4527c31a095847e9a226d0e1f290fcb8265d9d4f05200edbbbe9fd9152338b6331c8dc32b097b6f2eb5139ae167fa9168f1693428e25dbcd29cbe1ccb6c0540ef895bb7095929c80d795cb144241556c606468015f1366dc5ca0d6e2f4451d13f36dd6e18fce66dafe482b27bc727775b29cd5bf69c4d7ccefb387c0ec734c831f49e89240426c3cb5ccddf2057768a8bf467e4c58099338d81867b5916a634e7f1d1cdd2d3b13a33ab44d5a686a01f4ac4b5b182f00ec97dd87b94ce482356a3777b0c1ecb0367131b84d79983becbfd53d716d750bc01f982cf25d30433ecaa4edfb743d32e44c3499b4553b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h8e392bd0d79c514a35543d5d4065c81f7cf596b5e0c4c9932d92cfae69ee4ec84ff34554c3c4efe1ea9284c32444d50318d9598da18232d244babbcd4132773be9515e5eac76519e9728d15c67b74d54f9293af9ff31e0e357bd08587c07f857a89a369a34194a4daf5d9a960d697d7c4e748c22f631501dfd6e57ac1afcee77bffa6d9e4d46abe42f4be22c5975ca1f4545d071375737c037ce50415913de5f205ddae004f08106bc6a492f17e383d4c6a10c02be33a8e0f289c03f6c93913e6b1cab464e8f1f1cf83bbc571fdf7c5277ed7126b2746badc8b74b963c11a25b5ba66735a4e9548b887b4f70a1c20f2cdd0264;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h83ec5e22a37eae08f4be3b0e9e7b27fb631acc7511af53aeb917d6513ac8ce2140968987e7b2c3f20d1603f2fc88209950c28121051344c35d597058d8d0d82b3f96a82f17936e49c9bd4e94c8812b805eb6c96fc6f7e974ac94ea09b786f9772856dec79fa3afb63437bd8fce19f22c5005adf45a2da4e3c6f44c8db8014e1fd138a7d9c880311525bfd500f5b88b86067c4bc1013efa592c6d44c6e85f874c0637e4b6ab119dc8b9f35e0a3e0bc0fea49c932eaded0931c410af310eaeafcaead94bcabe33903e1d3e4e757732caa39a718affc92a597636b2e1bdd1db9a741c4724874390332a37826434ca0b487a0b848;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h3a5b61ca7b0be10c1cb125549b2dafdda7a3e09f8a1dcc098b9f46aba161c07a0bd507ba4c7fe24c4330e4972c4ba5e865aea857c6aa5b0decafcf25339b39efc7aa4f3c2d02630c9261aa642cae4aa7515c20cd06b4342572ab21461c6c54f7099e632980928b0185fa6f1b2f52985f68df70334c79029be6ee1a1a3982c7179b157478ea7faec6579a65a83fc3b7bd411bfd1bf9f14b36905a069fc6ca7123fa52bba99c9b308a4b1579a7254f6ea9723dedea0428dffdadac071d498cf44e6deaadd942a93a3aed46d07cb99fccc74f30ee9516071f3197e970b54f932ea39c3505ee0f7b2b33caa64ad32e29eb947d6ae3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h162a92fc726fbe896b8741aa4e6d4afc19cf76f3a3de5d549869cf10abb7e66761e413eb4e65a68292ae03a3125edb7b3bc2c4e7d50311014721645756d092f0b69b868de92f4d95595637bc751232ff44625858bfb0d932fa989faeff6aa83c8d4cd43f37a5fc241ae426fbbd5b4620b765acfbe53732f454ccc0806e41c19c42c5866da6d1030bba03561d7dfbe2ac567c399567bfecc97d2a51336516afdeebb262d4ebc6d53061573a186fb68432cda620206b87d01c43eb41ce83af8a78ca5d845ba640daf48440065313daa6736192c1cde58f211a44042f15aa0ba7caf76bdbae3960c4cf42081acdd01825510057bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h3854f959b470bffa75e7682771b6c36e395c149ac0579a4db3887715e2bd76ee13c6712a0d2bcb24d84c3db863f74d83dbfd90c26c778ef703f1dc719a8768d12eb18b9a2332f0a92622c19ed95c5dd1763e4d20cf546e9ba85db44f9b3f3805cd4cb39e9845b48593f1ac31434b9d1d95e0f9d184dfd89c87470b0406d946afa74f95d98311b2802cafa939f39a26188f2082dc5b91865dc4198300021d6ee108b1881b94181902dc4d5099e4c6527ccef379bcca42ed91f7dcffe4e0e8acd05cd9cef6b0228e918887fda7c986aa44c024134e46002cd950374e8f583c134853c7506908c215db165772c809e845d171cfec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h114d851885979a9ba843331de8aab65d30688c86407451853c396c95a40eb278b9b26dfef9d44a5a766626af015939d566e0c02769e63a849b94192ad0d15cc5e18965052842be33b43a2e6a9a45cf4d08253219e5b563f2c7a776817e3b333fe2934235a64e7fbfd48b8155672258c6553675fdc95144b482354db1803e959a4a71471991c01005403e70f67cbbd8cdc8fb21dbfc76f80a9661963cb2c21496e416f302b4280b35066b5017894c2ec7c71fdc5e41e6e678ceaba17195c8c08f298d2e095acf4afd078828211aa699ca323f154cd588bf0376ffddab2c4418c078dfed0bebf59d8d263a42f2e8dc0942b17a1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha58b0dba59dfb4dbb257bb99219f71a70a5001273d8f481354738c2747ff000f4c534e72a153e885d3b3a1c3fa35fd02c881ea8a59855ab634be17c8da5f8d70abf381d0367ad45776ed185e381a8bcc59bb44401d15e3116a57b6d715f9c04030b373d39bf0992d8ad1824a9d018ba5c613de58d3e5f566ef41449504b0b2c02a11c43ed68bb4a93acff0c2a87a67627c7a819827e3147c309845ec1dcfb0db0befb385e5b0266627630e64816336c00c42f54183cc7cd037db34a552c055595dc5406005010e1f5c597052bb5f989def91a2263b7f89d2f2bf7e72b6c204b667ffedbea8926420c78715499f343b26c5db5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h53eec2311a90b358994db0cc325dd607625450b4e2b28d027bccd709df696408da740e3f1cdbc78356f8e3ecc15f7bc6528a265d9adaac198a459695c8e6904bc4701c8405a7e59f4c619b040db70e3f68b1c37a89373f63bd2e5841b314b7e556b2c7f4b87ace75a9d8b8b3a7d2fa68a884f983578f0d81c4ad20345f58a631f9bfa7bbb1f7239f1af33b9e8fa548a1787f770266b659d7bdd0819398d753974fecdcbdc934caa08ba7dcb5f629060865e1ac7746724701cf4a0a065d87ef639a6a2b6fd267b73ffab083aaa3108ffe7b9eaaef3534016dd24bb1387d95d1fe2ae265f2167c3ef90d56cce6776525a4f9e12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9a842178b53feb927dd8c5a7c9dbe6f669901f48a9cad586a25d115e2b3238dcf2ba57adfe3f2860405699878d0371a14a037e2f885df5752968fa8be1276df65d3b5e7d062725a85effc1cb4c03c14e5616a5d5c6f324d1e992a5c9119db8d990dda58d440295fd04440edc97f1720832058bec0c0b8b9b0cc1e511bb60d8aaa8936e32f1a380581c462f793464d52a12877d4b0173e355018ca227d6a43772aacdea36b5bdc85b4796a832745dda42b607c07991a1a856a8cf3d7137789eda3b54886342b745169c3cacd244b5fd5fdc2b578a8711f85bfa6c4b2d95fbe8869fbcb0b27e2f44e41bb47c7be3955952606752;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h8020d3fbad3253b6e2e0ceb7fd460595b6aa481f170f8769f5d3222d3cf1ea4f699d57def32f40edc1ca2e9a1c92a20f59393b989bfcf2a3799810ab2b266e02a4e6c86560b62e6b1956dd8fcf8563d83847957464343dcb7ba4e46b3fde541f611e4534faafe20f4c503cb0d94731107333cbbddd09ccccbcc2bcba9c7d5624816065c0df120164b4681ca4ee8fabeb5b0f07dd0832923d78ebdcb5a136bac0c76d1a14b1a69391c949a198db268e57e739825b04ed8a5b4064f8bc63e9f8b2387f66af33ba3079733a9fe3678d6a89884d39730bbc8cac604d1fb6bc43ce9ff60ed38b450ef29f000f9d0f4853c37794c04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hcbf60df16675a50e4ebd328ca54d9b4aef984aaf6c28e6b62bf64daee3fadccb3d3f53be21d778e0169cbd72e3368a81dc498276791663bca9f406ca6013ab4abec791c787482d71a7e34cf26f38192e459a9d51d0828d6c294591845dd4e636d53318647b61912f5bd4578a0ce14044fc3d122e6317281eaa6d2d30af5fb8f7bedbbd333bd28d39e50183c6689e3e598a3421564d465565f9dca0ecab3789c60a269b9724e5bbea19275dfbce311504fa44318646469b46571ba69f99f2c575f7e35f29f40b8e2bdb0b1b7f48a5888b199e8d4f90c30e166fa48616b36fba94a15fac13772eaa5194a5dadabe4e2cac8d54b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h23717d24577768cf17d1011c784cfda42d3f73680b0eb6a21ffd4a97c04a73bb145ff1c08b3f6a638180e20372fd5cf19d67b11ab44ea9059e3d81c97745ff916659a417a4ff547da43ecf645bcf6462f0bc63e8a58d31a14dacdeaf579fd64f0a81249ed156de062e360622daec8f8e5e48369fe5bffcf41ee89aa6ad94be9e57dc98b89704b56f9046e6124f925ec98e0e66eb19ea84ea372e38fe84a94c587c3480a74d81dc256a7cf1849ef1bc3c86eb1ac979c5716ad3132d8416e0bf7c068c25bf5fd6ed0e3afcabce298b7986d01d5ca790b703c39abda13e20ed81630d04d32182b6263c965c95033c46f26d54f7be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h95387810256e372bfe3f23c1eea42527f4eb606ab83452c2c6e6357aea8017c117bbe4ef619d48f5b5f47bb4fb7324e129d3dae27e78bd5f29d3a93820cd4c4541f5aa174d5847c2a5eff1edac6326c65a2afcd9bd1c32b4814f0a81aa3fa62cb62545b2a89defd6dd95f7f819a6910640e9c8445e69e46d4a671d393edcb3c5c3b9b426a71e1e6a662e5712d9e264e22d843e53d122881aa215c0d7ea6ecd6b99fe83d1a374e3cf1ff6731d7ff49df0970193bcc687cfc9e607be6db01fa2b7224ae5bc76c622de0cb559e53e500d1e99e6133d2a7b818b635a53c8371ea04b108641612a14afcc6a92f19ca0ee752ef5ddff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2d4535e91f6abd977d6a0587a84f782a188bce45569548560bf09a9a749f76bd31e0420a3e26b270caa3fbf7cde86883afbed8b86d778ecf2552b4c3a8ed204e93b90ffb3035b0d5995d22626c4e7196ab0c09a5e2f516b9f3dba765eb2d71d3e909fe92abb333bfd0d72733a20412f9f57e92b2ea1ea64f3c36095a6afbcec796780080dbc61756382ebab26f8176f30207f5ff25bd858cb0a96617a99b025e1cec0eb53e5f819887e51628371cf38dd5e82b2c96ee163ba710c2bf752a36e727e55fe0594706947f6923bde880d7dbf5efd00a01916cabddde646d1c9b9605aa7166aa9055886e15525eb1defce0202e2355;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h91ec603f6e2db4e794f45c2578963bb46ff3a454c5ebc45ce71a91f0b719f3207e586c6653d9d389849d951ecabf7ef465bd76e449d481e1555bac4cbb876cffbb1f75a4fef8eacf312120d9f98ea7ce59539c01f9447f954c2173a06677ef423c07438aedebd83aa1a2428caac68a7ab47eebfeb92cfac64c478aa7697c044bc254a9089c22d4a718350dfde5c822ecc8989717e9a47f9eaa79e0402f7aa357cfbab3999dcd1ac24ab6b1e75e9d84e59a2e7d2c2e4fe6a5a023b4ade4dad2abfd4244f42240c78e932f28b1763e2a665823f9e59626a68c5d460ea3ce89a9f9b54bb9973ee1ad11245183f8a29d9f44195b6e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5fc5c2a14d630601813a1e1e0038d6eceb4d0212d1179e614609bbec997c64cb99a8e7e08e9e75303317f34c8868053e4f86ecd5e7e47204f048343db4ccf6b2c84663be3ae5fcae3c4c1af7001103145a808b547232165693b236a78ceacc91a243635e6ac969ed8a2e7aa030685a7370cc611cac4c569c269d23a79090c6a40507238d027b79856e43643e7e5fab902a0cda28d4ddb26aec9150a5007f0dc9887fe352bd1af91e2c8d09ce1f8969aaea0190c0068cdb8b63b751813c73f139e1995f6ac65ead92eeda223f08feaf1a5d7ceec748440943da479d6e4b7d0df6ffdae20c2e67247c2be67f91529357d9484257;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h206d7e5efcf0645de863ef163f0507e6fac978b0d90ecab2823c850574465513096f58544603ece1e2109f254c252fa4da08f1c7a21bf1fda69258cf1215625de846d96ec454e2dd868bd85f22a8a0a2993ece465f96d516ce2d09f65fc7efc8c0dcff907b375bd2a4b66c2109c94919e9e51c979907a5834d9ef9eeca152b6fa7df27453d142e1a8892545a01eea6d03ff0663a93d9b9325a1743f744bb361e8ec33d59316584f321aa0086c50534cd8d5800d04680b5c6956dc0d9216ddb12f8f029a85280f3bd8d2220f433f4f3d9fc9b86c8524323a0d65b5ecf331e50eab13bb4b7e7e9b6bc8b300144e208a42b63fa51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h81c7a56d0ebf2ec6fdba5302205bead6e92f6a298e3e14fdb8d202b328d4ff845f2cd910f20a832cffe691beb496b00c2e6bda82982c20790cdfcb8d4ef8aea527940ba551d7855308480e0e8b5e6c7e0f3013bf271ccb5eebe4709b00ca48fe12b8e58a46660a8dcaad780ab1027344e04462ab36f9c59d62ec7cfde2282726c42d7cc3a741db8f36ade1f4a6bfd66cad8e9a11093255498aa49da2e5b96a01fb99d08e8b03376b713c45e526fa344b9c206be01e3c073c359971b841352ea4e2b2feb869584745c32c2ff76688cd16b7f05e2156ac566cbfcf00ba2ad28ade61d15be1027d6b2ff9cb5f73d1b2101ea6c1a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he32e0ecbfe587d88d185a9b0d9f8a1b9cb0d1b430646491cab112d4db0b4db408e112f80cfe68812c6f5f492bf7af11300b4e567b7a2d92c2d0dab043062354ac4aea3b5d21d0ef032a73c9014557a02d4d911a9da97c159351f9cedbd2ad3ee67da620ba81c642de970ce647b03f9231f4a0effe4b89ad34f81fc10232c067ad89019931786174fbff2f6e350b543bd07104ca0c1ab275aeda2715fe97335bd22defc6ea8712063fdb2c8bac6e358dc9f3537e36d61dbc63c744845344efdfbf0493fa2f9472845454f4c8bdc5301c45a7186243c4691be654e92829caf793174295e3c9da8b10e5a0264e909cb844b3e4bf8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2fcb6b596c77aea881b546670dd2fe6c8d840366c713182fbf9dde993f327506a6c379450d8184ee26ddb0e524193862ff7484739f55849e18e9edc102e0251e67820469c9c79ec1d74b776c9087a41102539b2390d9d8b31897dcd94216e76c42a7eead4fcc71f947adbab1ba4660055530b6f9fb3d7e24c3635f96825e2c17e8e5312dc0865c356416d4d988d2336cfefc9f6dfd93a9bc4128e9850b23366dbe7d8f543844a351d2818b6aa28e01dcde4d591c8ddd55abaae5f91deba4230f32a9fd524f3ec6477c0bd00421cf67e3c67071a02be40ff6b93407acf04fb4d64f1223a984734a6732fa6633de4b3b37dceab4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h299bee3ee7b14b9724cfd7d1b9b61fb14e2a92e86466c69301ed27511e08ef4aa8dc668b218ccd2f89df55637efa5b20a45c20b8cd3994ed7fed5ee3e4cf62c2858f1cf4026635e9b3e648937b4179f572249e9e2733d17a7e3f84e091e6f07c995360e6ed19b50737caca2f2243f5980c0501833d56e3930f51a09a4b3fcee5dba42c2c643c661442115ff16e2ff48023478f24be3ebb8d445406dc7d137d1ec65f1427647a826c5bfe05177a1827ca7cd7071864d6817d01ce4a549cebcbe8a9dffe50647d8699e1ea33c5b4f7289052bfc6f741057c45022a50a6400b6823f9dbcb118911b4797b1db11e46aa891a7643e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h79fc2eccd19b3bd3020b3d5a2ae13c273b3f83da51623bc94f9607e686bfc5de16961055eeaed8b54f9790aa337172db47b5a87452d0a5817eb659596213bb5ec54ffdca03cb0e8cf0541a983ab5ccdab265ad4393e557d3ccd275e46f2d5933dc44d441e96d46e4eff556aa55e6cb24b3c2ec376c1e8e891c2e6541b7b5cdedec7ed26733deda6ae3e3495a272e01386013d695f1e5204afcf49c26431c8438c66be2838fed7700eefe377590febee619ff8c31799fe2a4670007ad5aca7dd0a92a0715d6e01d15d8ddac65bc9d805cf691396e41e86cb5a6d5ca7455e9cd61f5f749dc14174ecc5167cf8cd5e29970ede4a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc3b11fd578155c376d8a711fe1de8d7143096f6b1963d071a477c61287e91d6c7262b3460cc14b62fc26e7a1902017cf5f09f5d8a1f0b3c3ef4bf9dfcd7c54201f3973fd4091e97fbd4b5730b605a1fe981ab0f35cd67da95e4693b45db2d5bbeb67796e191c329835d9c768e64d02fb39d791b61414503226a4e0c3aff121a8949c25e38d593361ca9762757fd12f26845c6b1d0b8c0b8005cdfcd8f0a887030357771ab44a4a55e1dd3c0d972000301c4eb02e4c0ab0591f8f9983868b050fac3be45a77cee5141b5ee31fe74f82487f9476b0f075721c9b4f692ebcb9b6f79442bef7576cd3f24c0849b17cc2f5dfad7b3d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h38978ab8752b084239f13ada7293182b1f043bb5cb5b8bb6473ebd420d250ea4096bd1adf49ab404806c74cd66ff184ab9325f058e533027469f916bf51c81795572aaf537dc1739ba2949cfa51d0d49a0b1d782dbe337cb48d28f940496b6ed0f99da89b6c419235d7ba9244ae130815ada9986f8e211c3c04c0bca7abd3a547ab011302d2d577787d4d2bc705258e53717ad48e6b6ca45660687a563d406b0c7aefd512621886c9aeb6e9b66f5d8a1cd2c30ca149478aaa02684140d7da856ea8eb19e74552443d40274226b44de70a29d2ae189a6681309cce07db704b9942209557ad79aee70c84dfbef2c56c126d94bfa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h13780ce2fd580f70b83a3d2eb0443762c2186853e7d9fc5f41a101fe18ccfface9c00544a5f8c7a11690ee10d8c6ba91bc030781e38892f4992a6d65774c2cc8d578857e4264a22c9d0d404af690b90f482a39c40d674a79ef1b072fc08881c5f1e9ae5b16c274c9619fc61ce9ccc0df0adb7f811acdbdd092e1b2ce46f3c30aa2ffb74386942f82e52206c1dbecfb1461ab63fa091404475caaa2c5ec9e49e54c29ad6962b5b305f6c7f00a111e0d60b325b9f0854723e052d8a5790df4486529a4a22c6e8e3ab2c9a8639e4de4a0f35aedaa61dcdbb4e1ea87ac5461ed2024855db390e27b3f6d4ddf25a8f9bbd4cab6756c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha56b7adbea82636b7620ea2d15be7e67de6159f216ebc229e9221b54750e5c3985a697162196696d5972d40ec154ba95215f3ffff093ecd10a64c11780cd925f88c502e81ee3d2feb253beb6025e188d44d3acb8c701154ce1299aee992c09786995de0632cf03cbda809006438718f4731af1603845d46750ba505a5fc61cc3a836d1e77c4cf9d412b93e5cccf79d7a5a21a636e7c3561e300b092651d42bd945804f7824715440e0a49261375b9a2f57655b70ed3fccc389a9cd34f4db83692f392c5ae16a2ec2d12e4711d4776716243a7185b4a755dd05c65f1ff6de0788a499c9bbe60cbf03b2092d4773635780139939;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hb6b24dfd942507280e216b7409e88d91dc4a8605b57b05bf9095992d7ca06757e37487b3922be6c5754c4c2237e051d47bc33ef7bab51c454ca0fd20c80b226c2cdc7dafa06b87000e7551bace08c7afb72897086a3b6f8e6547e5cebb540c213a1c22f09ee5d4b57ffe39ed7f3c2bbde7df4859e78f0bcde42c49291fcf8fbf8bc37eb1998b8756afa4863098260ec5eaa9d6b4bdd9a424551551f386a2f72fdd166181f84e1ef4646bc2ee184778d58f6ccc85980e159bcb906ec9a665583a006e0ddb308509824abe0429dd51160b2cfe4acff46b4011ed2e0bb1919f13e1e9a80eb8ef5f940e9dd69b3ba61b543a3f30b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h3a223893a5f45ae036c3e299462deb1eb035aec7e2354ac704520dd15938ecbd4aa9de0391bd96d5d40e49c1cc3e55325c5a7b2d64445e0096e59c6c3665bd8650abac8df00fea036f6fcc53890502d412f5f09a25148251e27658f518a7e848b8f953a55828973be04d4adf1d811ea6d63ac4c73227de1fb7c18faaa211a63ec262cb725a31c8093b81fe33d0f371b6c68614548c3295fc1126c9f6f94f2df995b2672aadba5c43bc96a5bd31b8255dad51aa4588d75187614a89427ef9574afc719d60690d24331cc6b7d6095905da05ae97a1c748195d9e252ca1951347fbc959c0db19b4714f774f02a8d88e449b03756b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf517418cb5f15f805e7a98fc24ad828ca618b85e5df747aba2d1b8fad432df55576148f36fb64d190e461b9b9e71919e478c7653b7ea271c2a956b76558947ab85883ef4911354c7e150026053958c8056886e4f9f202f8e63c3580ecaadfa8bb477e7a42153cfbe801174ecdcda8cec22cb83d64cbc2f09c91e33e811ce415d01d40bdfd1afb63a32eab3992313fd45ad2308954b5a74b6c594a4bb10cbafd43a2b81d79d1f2e3d15ed8dad94d5a5764e2e81abdb4830462c5751b8af8b03a85e3111e8e9d1afc181f76e5083414c7f6f8d6016ba90d5799224dc6b7c7b31ded8df259de5d35b397787da030b8ee207f85172;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h15f410c6507d7e5b1386e6327cf5a6fca955350d618777cbcc60b6b34d358a7ff6c36b2a5f951b964e22d3ea5d56d974c793ba2d9d9943b7d2e847988e06549f3c88376f02da9541e5612a9980c6c05acbbba6e138539a3394e751e7dd648ff32e84b2144c762cdf0991a92b070402d7bf34fc1aa9e709c4d9257c77f7f687d4b163d4907a0777ee14c2d683e9e919740626313fedcc6e766fa2c93b6d8c0c44396fc865050d1e8156d18812591ca4ce301e5f259a30e5f8169862975490179b40dd3b65b94b87d673dd8e33596f7e545c8c77da8e1cd396271f495b36ed73f06e61c7d10de60f09f3db9132392512c55f4f4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd47d72aa515fc9839db729745de371aa23cdcf2bf8c46a024584a0e2cf7d5a5d0404a4a033fc7a19a699ab2d21ed79441949c933d709b425318f448afd5362090fb141653297ac4bd5fd4b1849a6099a5c124618d6a270e87a83192b01a208fa7ccc4231f3aa2a52183d0f975e6e49948330b87767c4eb48d918d7ecfdead053d19954ec323c84bca647866c3047cc2ed3c8aeea500156d4b6aea5f24fbfaf8c3cc25b5d4bff576a8ba551cac029949a7912cf2ace7bd1509af1562377a54266c3f3c9f75b62c5d1464e93b18b7e19a7fe2826b6624d7000786559c272593cbd9c871a552b86b2a0438305e2709a12054ab426;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc1d807c129832eea752799a911ad09ddb96ab8f6cd367bec3c41cae997b4440047f87c21bddaec9096b496a37760f50bc3324f0618619ff6be47e1bdf04ac25267f425235a5580d9a8f16de6ed4944ba475c7ff4d7c2b4bec05fa6198f16ab03f2034f7767ac44685fd19042a8dc92fac8bc9e9dcaef26505792cc925e06a7af7d52bee60ae7244aa91eee04ba987ef667dba9fa9e4b8219168916620e9672643eeac9b656821752f3ca57349ca33b867b639c02f23b3c376bc65b7846da7924ad84d41f4d0cdc71142bd23ec0be0e151125190468b4d87f3dac43743de733c461378d5acd88d84101d53d8f92e0485bf67c7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hba1fe45af6140907a9593e29599de415279040fd680234d85578fcc495ddaf42f83899a8a7354c018b98282b76c334c9cc4756d1972e2d38db4da41c4fbf3355df6a1daab0d562e2c993bc1534760b541050f879011a1b6c035383ff0022cca9a585fccba2e0526ce544bad0fdd9acaab8c22343306d1b8f44ad6b6fc74cb94f373467c0e27b2672a9adb235e72eb0979cb27c0a11e5007664f3458892461aea172c1e002b1054f56af677110501cfc1801f33486d9651291fd79710d10481e11ad6c700f9c580d676d0ce2e4157e7f9cfb5476ddddb539d26f796501e60b6633a034e3701bc43898e13a81f347cf234c14056;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hfe758861d2b7e485afc7ca24e0fdbf2d97c6947c0cfee757897a09bbf9184f80908c887fac03a0a7f14ccf4238bafe2c345b8fd6773dd78f587f2902b0320f972583ffd4c6f5803a9d3ef527559373026120a1ca9f1d30e17fcf030a34686c8c1c7a510745131940b105cd1d53de75e9e76e7cd7770c1c75a1c6a7911d6d64fb1a13fe515df4cc7c425ec917e9626fa1ae2aad25af05f11d669696ecbab96e23a45c0d7ca2d217185437a543fbd039feb99738cd621380313557b32ebcc24a0849f5276432a7bbc8984f17ae9031e551bed8fb7c3b33647c56f1620363750062a9c71990e76ddd3dcd0a1e607c6c2920af2200;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h83c3e611f0c15a554438d068d7eda391084046b4a68660540921517e4dbcc192b841a0c4ce5d7385bd4b3b3a88a1ec13a6a7456c5f05a823516e0c571de4bf206d486284b3672f7a5819bc05a7afc6def77fb8e03ffb2ec088834aa56fd9195a5483828e720edc485245fcc92abc809bda7ddfbd023f2c72d8f0fb6efcfa6942b14e2579dc8077fa0feb99aa37392fec59faf434f3069a441c4a6890147f677f2f9f80963cbf49315493f31a98150da1830014921a544f1075a04f7a4151cdf0f9f666fe813109f76703e9bc9339dbf55729bd0f75e58255c6ea1913430b5a25ec4f1164144afa920f789357471801137916ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha8cff459c7696b9c1202666851315d96a10b8a414719866e2173c27e83d05d2c74c0c31818def883de0294683f0ec2c5517e8ba36aa7e5ba785dbdefa071d7d1c5c10665574d65db242c90b19e735654b4fb941add53080e63b4618626df9d3debf098cd964021cfd1e095b3e132a8233f2a41816ae8029a72c61c1857eb3be840d6e617025ac64fa064df2052ea26db01f70b9a80a4c7145b2343eec45f17c8d9fe8f5a5bb845b13b8d8c55585076b617199b82a21732b8e117a287e1e92488c66c1ea9ca3899ec006c253490747fcffdc0e188c8703f45c020263c7756f461fa9b9c84f42f3a68b3de0eb4be8760ebe57932;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hbd849b5edaf46abce94c2387db7112214a80170608f023ddc0be8c5a0dd7a388648def8b62e6b8fdc4356292d7e80a5222d8d9b95ee67e39129e2fa51e66f479e2944a7049645a68467cdbf3cc1fbe90670526fe104253045a221856572b38e8586eb49b31232f9dba61dcb6a8904af4e7f4dbb7d00ea1c5fc6fa523f3e506906729414f26421b94cc49f22b91bddf37c060b654c688650297444aadc7e217b791389c8fd8cf006fae40c8f11c0ababd63a27e7fb192e23b5103c487db7dbf50debae1cceadf2cad83a0ef382e7a8697f496fbc2554cd962fee7592a43c9e95d31edf0243464190e1b9531431f7c4d6eacd9a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h19b5abb597c998ffb8695cbeed901431911ee04e425eacbc258979fa4673186fb15ae35640862c7a1c04cc2b6b4d4dd17f0239521cbd7d57f9cf688f1bb37312f9180baf4f0df6b47924fb8f5cb7fbf79e53f50d657599e2a824174ac45b3364ba2f51a2c1fad112e26178a39af87fad4c577e9df348e563f69587c2c786d56f50d6a457931ecdd6b12d5218e125dd09044139dd891c6d117c61b6b0046474c90ec2951eb2ce7967f1424efe312e03d8c2edb878488d36d23095c61c54ae62ca65d94d8ece7c97e67470e7355e438e0f6cb7cf17a86fed03af5b56dd46090e675ddb648155a173ee9b6e52fe57af6ee1a4b534;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha38ccf33e1dc90a48e8312b002da89177aa8b2ca3415e20ea654749e89f8e275e8dd2767aa56a05c29c3f11cb0a817027aa9fd8b9dd94744278c77d06ec44a301fe355b6f0842810350152f3b0603bed3db99b5a42525607ccefff76b8d38e5b89340f712e39ba72c7f574aa1e7c36b59734d3c920bbbb7332f16e357eb4ffc87de23438fd6a49c709ff1b860c6f0f51b1458d68cc09f69a61da9b2a066e738e7fe808722488f5e607786830de082df594b1a69a5afdb69afb6aac8599c90b10f332db0de15633cbbf40ec6a4483cbf805ded07ac827e9d8d337f875259acc76d583af349710d26b29631aa565bff8ae5e5aac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hcdcd8bcd3b93b8dfd5e16500542bdc11e8817d17c71b1684fc68ec9d37ba00fc5dc1f4c849997817eef1dd47378ee20ebe9033504e10381508b329768d2c18ecfe48064dad8501a7da9de625f844644371dd918379cb1039641795cdc6c4a3a6bed528094b175f33ed010cfa2c5754770c451f2e63d9de68961dbbffb981732326110ef7ac9e07e523776eea8f203cd3ac60a3cb544cf818b804ecbef1fe47c15914586ca6f7e6baa3c36aa4c938aaf3ce0ef4961dcb4b2e5ab89cf157895aa2fddbeb2909ec07681e2e00d03cf9cd5f390a1054c9cc1d30f2dde7189b52cd7cf4a377fff913f03996fb4fc1ed412e89c042bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h881d43d0915d84b5e03aceab6d03a84afbb7629ff25fe54f992c3fc153ad9d6411584353a5cc725922fa7b80cc5b93ca47c87be670466607d1833b1415e4cddec8464f5416f4c931dad9753973de2058c6afb8dc8134415448066544cade9e1d94e13fe8a5ae03e96dd56997d9d4a14ffdc02780147a7c71b1a6d9ebf6fbf09cd3ff4155dee9c5df4099e3207ffc6c24450f9b480003cc9fe6f58071d7400df767351650d8116f66ea0e4712f6038472693e14d09152d3f2aa92f8d61c8166e068954c6d9d2dcd37b2928a71b77c7e42c631cc74299050dded1ec23526b31b705d07b3f8fbcb4c4d905941baaaf3329f3bfe5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h188e84e0551a7290e11723176c7ceda6ca9d4ea355ca1a549fe78212a74651eabdd8a58280a1a1081100295c38a6f345446b8fc368ec6e4044f6d837fe23c1d82310bf82137dc5cb693b837500bab6a181ef02a122ebdb01e2a94fa50c6f391e20d84c09956e6262d4be49147712d36730fee2bec238c62dfe636697e94d143aa36c52b572dceb269909253591d97ccbad204bc68f606398136e2e4d651f7081582090b385a30a63d9624fc7948edca0f0833334928ab17920075debfc9870cc9c970939c77d725262240ecc6135f105e39f3ab2dba61018c3f03c2a0b5a7b4c79e4b82a7d395646a9981e9690d40f07debf3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h7d4119f6b6a7baae20f78727a7287cc2aa2ed68ed88d073972a895d5efd552d471203ee93f66be375c6ad3231cab88d1391298d3a445c014f0e08431aa3fde779150a46671615b993642e61804c10ac4c5d19a919a5c5cc6108b6c40ecb38a7d7cb789d092382ddd24c421059f7556a635b4ae72899177b59412f503d3a4a4b448dcb1d6ac88fe77956db183496a9065d137c45cf5ff8375fb28471789399650b3f9193e6e0abb2706aeee7e2797e0a8c068504eab4d9f911cc3077f8897feaeb3345525ce14eed8d2771baba788a4711e39505d6ac0b2ab886c4b373a2209f3ccb981c7db8f5792ed6477018e5283586b387b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h20d2d30612e795a56bf21c84f626195fbce88a282e981a984cd1f7a2cd563c1c312bfbbdd47a1d82454ab535ec667d9b31c8b136e2151d667963cb26541fdcad81a7e89a1479ebaae7e947f2bfcf61b2d82f7277c78f682778ed57107706087177d34e1678ec1cacf8718fbff98dd8ab0fcc0058f79457315c0327585373355d611cf61080801e54f4850af96e60f8dcb84abd270982282d66d0e77efc52a0d4a1ce765bf838dc4206fe044cd07e450a44132db18a03a497e724d6521528c1b1c2e364a4f5a4f974553e32d6a4a33d01ffa96c8c135a3a19b99896508a3a8cf163247fc965164147d9a3f8fc0676fac675d95e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h756c0e366bfd11bff5a8ae6e3be7cd4bfb1419e266ad10ea9a7695adc47db2c959e7d7d2be7b3661b1247c0448c1b41d4f80c3879d51353bf4ec9e4b69f474a1406090517e41c4ba7d006f7c9e5370fe99e920951cde096e574825a2c76fb2727e7786bb06088515a8c142b7f2d7d536b9281b77a12018c715f50bbbbd0e4a958f969d3d3f6ea74571329d68bd6c9c9f7d09f98fbb8ddc6399c72d27c1e49c09c671f775e884c6581bf4e95060bc1525ec04814fbfce4392e3d8110a4f3dcbfaace8ef7edb7b091645ae030ba90d40b8b67b325a96eddc0bfa6bc50832899f25b5709393d1afb9387862db7055055ece55bc4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h948e806bc29152bc9d2d708a7c84d66d23cbd8167ce044072c379f2096e944fe9de20df079bad6c9802cbc8c82ab2c8b6cd14542ad25b482dbe080cd553983ec2c5f172d4edfe0444b3ea22fab99c9f86b496a5ca7dbba4c084aa5359e8a9859600ddd1c40dfe2373c23053a577d2eb56b0bb37d78368e2e2b976ba36029f1cbbb96779160df7d2c3a371781e9a9f4233bf7d0350d940949fdfc56ac2827d6ffc82fa493d3bfb64d16da93d63f8f501266aff399032276e0af12b4a3f60303be5c9b75b7254e1ce5ae6a13b27beb6b7ebdbebdbac8581acb2debd0e763a21f0b856c0456b2a4bed0c78d28aaabd44ba40921b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h781318c1e32884e81456e737e9b9da7ac87f82d93812b55512b7083364f6ebdb24ceb6214c0bd3d83287cc582723193c59e38d79338a08d7a5b5d3cde29e7836b227c409296ad69348c3051a32d9f9084882a697fd740a7dfd4b970e1657a4c763e3f8596e6fd08aa9c5fe741de284e09c25cd7f7e7255cf0544b8103cce9d0e69bb68abad3083a21a35d8efb4fb38e096ad773e7dcf216e4fc88af68eb4d47c925a5570af0ba4b2925bc6cc72583659efc72d1ecced22e724b16f5d07907861aee8f909692d32c69f5b9836b6bb61007cf4e77618212d3bc6b5de16845855b9bd5479c9ae456bb751326c981404b3bd21594f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h308476d3a686b2a0971825130ab1a704d76b37d410737411ecac315ccb6bf688f0a627395194ee43f7f65b077884fb530cede5e3c5e79d74055e7f2242cc667b3a95065b50da2bd36b9cef1dd7d892f0c020218edfa5d1299a71e3a2e3109259b44d07e91d961a998112e4ef64362ad857bccfb09d1aabcb6971d42d600835e7add9cf3cc72e3b905ef442905a51718bb5b7fb1b5ded9a86939497734c90c284e65fa04b31569aa7bfbb9749d5440ebc73c9d826f285d3d5b9388b3bf6711c38e323608a9e5cb16b379c758a657a272c631d404fea0a95e9be0f524ad66776668e857c84b7766b041fea32c894496351b4748b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'heaef6c21863348eb211d3121e9446b7148cd1953e468a6a6cc91c47a1b5433723f646d816392b47c4032fc0e375868c8cda4097bfa742b62bfefc0d6abb4164296c0f9b5acbee9099085bc50cb424667b56f9c48ffe0f6b13c782c394fcd251064734009aed6eb66ad2f9a0a9463e8a9a873d93a4661de0d708b1c806e39e20598e243c4ae82691213b9955801988a0e21e470851a1b354bf7cdf101fb8353ae5b645ed288af1006fc64d50bbc6d0748295ef23a1ea2c188abe1baf267fc84c58efd1568c0165ae4443f794fdb5ef4d711db349857ece514d36c6cb29d8abb030efd9ae02fddd4ee5dddca9607e9e9db6551a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2a358ce77fea35f404db672cb7591bae65186bb4325fe32f083fcc2d7790a3d4b5d164d9ebb6ed906c5aaa2559b08d1c761cfafef2564db0238d2ce757c8072c0241bf95975d83703409dac11553e1d8cbd1b6835c3029adb0a1b95a33f2a5ba5b9cadf3ab36a6c34818fc13712a20a1af08fd16f7a6e1b66d62791943a20b9de596da13778e1451fa74b8457fc989c5a33ab35d33c76043585b1dc67e93236d7d573df0cff5fc272e78bbcf8eba5ba372f750ae39a03815515d785f5e4b830dce159d9aacdab3df194cf9d85f29e2fb1b49e3a0448fc55a6ad6eb3dda40af0e1bfc81849a0844ab58277e047b48cc2534ac54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hed2c7293ab17f28b9668523ae2fddcd6c9e3344ba174bf59f8c287072438302277518cde074d7f8fff1e0605ee2cb9bdc8a9678c3622fe7df6fce96506711e72fa6d2e0046c5b3a788631a30819b706817558e166a22810918c730bcfd85a25bd383da33bc82ca2838252faf660d2b452d5c0731aaff3af06ef5e5f73c33dfe3034ec4b9e992d1233ebb8594534ae15b1a1fb48328a34eb2fad315fbb12e3f40d6f5e06fff24d0feebe1b676fdf4eedc3d785ceea83c1eeb18b0b600ce2974cf7d33cf9dc67c2fd815866a5df5a00fe48efa6ec3f40f21100b41b9e80a4360608ff895cfc9ef0d456a3c8ebf31b3a2307cef28;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc6b32a531ef30144bb9cde6afbc7403292633461cc8a35cd562ece9b4f69434da0bbe387cbec7f9621ca101e74524f3156ad8f175f4b48b17261b47d657845acc10daa79e24527bce29f94f964f31d14fe631b4e1df2e9f9b1db539aea63d575fded40036a7ba3bfdc7b31b72f6b689ae91ca1a07e777f2b86b333eec2b855d7206b09f2a83afc0a4a1ec69083c52b6275de37e2af5a8e4e8da3552e6f2c06f1a8f8bcad920bcbf67e3f6861e979047a00fec0b4c78110afeb9805647a1649a7dc839c21d052f9ab9c29da59c0e38024b79a9358d4581db528c722d773d50037009510978ecafbb181be18e1de3ab2758f4532;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h147b50ff8e44b891dc2f611411b75939cd6fbcafa95b431ddd3926aa7dbb2d7a104f34319f6a10e1183998507669022e34849d28d05228a71f89a61af9c82a1f680406ba9aa9564c43123bdd9effcf6eca13680c8e6d50a32bb62eeffe2200e067969fd67ee8312a69bb496ccd4a1a5dc0f7855355d1b7470e778068d78c525926d90e227a8b1258d2764170fc9e64519b7667073db7b48a9d1173002ae2aee9d559f0166ca9dc2139009bc13afacbee3fe45455e094fee13a620e2db7513ae6d63afa6e713089b214e56f6127531c854fd83d345f151b1b21d05f4aa0df0d519ab70af08818824f1689d5a7490ade6b746977;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4bbf7b38d420188a39e5a7c16f60316c60ffd59be6ad1dfa2e0447cbcde5738a9b16d03d402bbfb14a1d0df5c704ec4b5bfa330a21e704da67c713f82bb9614b649316801a4c0d7c80f1721684d384ab42750a602023e8f6bc603de3429147796baefa9b8293279ead2061adad72f91584fb01ada4a2536047f1f90af462329ec92bb2d98d719e8fada86cad237a8cebad81b0c1a8352d963ef94c8b6edaf799539b21c0ddaef19fe787c20a637283a5bf8e2773b6320a28966a6ef2e16c1a52caa5e14d14943d88de12e780d7f96ad867e2f09c17285f35cf7db78607e57465cc0ea6f7e5f8de7b377bcb1a57fa61304f7459;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h90a912400c9e7834b0c3020662c8cf9bb5f85e41278be9d1be61cf2e1d4854fa9dfa5c1b7a1a778036e502ed7ce993bb338e6462661afaa169511acdb3766e926801364bfda0782d90a32f889fd49c9e9aa782a0b85419cac289d7586d1d8852aa58109507d7b6be0b81d2d27ac028b6200e078340bac692ab54788989b74074e9cbc26522c38f9270d60d358428f4020b4ad149cc214a494c24fa6e8702260caa253f62ee472553df9aed8f369b29a655117d59363868a3db7987850332bbbf677f50dc4d4869d337354e5871c1577c333c1d2c330289a5f386b18ee919fc97bdf9491c0c4f5e6e8c6508fdc638a9ca040839;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hdbe504b819640c4ef152ebab1e2e59fbc5b7b28664e212581c522304d1872b3f26def224c34825192295f5f286b29adb97ccf15990dcf07e5f74dfa107bfdce659e824c7afcf004b6df9debe4866a55fab04844efa91a95f644dc0438f907311838604773e1771b9ca7503a3275b0bba832f3811c7ebd04da0c375f1e7dc7bf9e1cdab19715c0c857cae2ec0679ad2e8ad661d2453deaf67d221ce99ab9c29473b8fc30dc93cd36dafe97ad91f47767dd2a8aee944bd620bd2624d25e82e975f53b267d3bd3177d20b643b617e82260fd3a05547ea78907b1824cbfd3983b4bb94e195d5e5626de0044a4f07ac1a137ad46353;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd4cc4a70e36deced65e4c773e9485275e6014715c1ecf797ac0980e4596815d3e2495c5b1d270cd0911c2f4ca5108b4ce1596d7433c5ff5396186321eb607a8d0cd0b2f6dd71786c284c619d9343b1eab3be5c7d22cf9daba75128cf6c41f398752cb9e3a88b6f6512d7ccb603fcf11fa05adb7b3d12bf0312e231d2b58ff31eda4da9e3319dad4ad616fcd419a6b7e6bc316c823e7a3b3cde203ab58c46bc96f859a1544161007ecbe1adb12903d461af448f655da51cd72c1113aec5a71ee9110612d3ee558f86b819ea57320ed032a1c9b7d42fce75a3b9ba4dcb048c79d90c99ee48e634723fdf576e6632f2bd2fe8f6bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf2772ef05488bb9abb74adde49b4962a240ab7f6f9c96a60b2118ef7343932c1b7777229eea6b596f3e6107ce5b894f5881d5665efb7473eca6535b4c0de1651f5a39137018e711716d52829bb9dc52b93db4998397735584fd6e5acdaeaf472a3029f1b77ad9fbcf050431252f1ec63516a2a818895225c161ef5b2358c0c098cf7bbc75e57d21be72d1419786caf4fba683acf25430783baa8d05fa882b62cb4965f25148695292ee4e20d1dfd38280ea2a4cc74bc5d4b620a6f774a19680733359945b97c25f672330dd61dd92216c4b3c3757df9f8eff92c9e229e0d7193598dc71db9368cf32612bd7eed97ab73a66bce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h1688cf10fb54d58125e6900ac8f5cb3f393e52c15435c48a23ed51d8d6643b3fb2d928ba2224ccabe1795260bfac4a94526e022cd23b1e4a2f1dc94043ab267b27ab0571e58903ec10d1ab6c66cbf7aad33fe8fc1ed5d9b058278bb3a1d8f1f21e2e0c5ef36d41a4b57dd7409a8331d6a76f99058f99480a316e29f0ffdbd22aed2577836ad3ceae1cd641850ff79e5a8f64204e967e4f90a83d3bd68379a0add2dc3ca2d4ad32097c5c1ca5e80d06764d56612e56f4ea644c46e44cf65b3046135139a3c5c5ad0e6c4db23dbdfe0cb56c852a171e0d169c08e062da14dc6537ae17248076b7781ee4cab295e35d8a54f31483;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h59f91b8a7a8124aa1d61c0b6c4fed7c03e171ac80c180c68a6dc7ba97591d5f673871b9b982b8809de718efba9a5601633168f736be5d77c3ba5a4911af65fab1dfda247dd309d7c4f420af8bcefbbb944f46fa5590f4c27b1059716387066c45ab26e4efbd0db67e5a01e186b693d4d92344b7b91575a69283b10b1f05431c40332e2ed829b1681e5d5ba9ff60b9b0ab51f7252b17303a5f57d07466293d45725a61e73ee4335af3430bfb8ed0250a97194ae067415821231d5dc9f918e240df0a81db5a21c8a118d1adc1c97c74e6102bd2176b5b0be77ded0dac2a4ea8dc696a4c759ef6c701e24a597d07492640dbf01ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4fcb4cd40bf7b0ae6bde03e2b744afd37cc68b442916e58f7cbfda4a93e209ddaa9347fe39d14de82ec0c59036064d3834804fccba68abbdc320bcdcf0e4de13699f060dfb60aa50461d1589e8d7685e0978b6f39704606afe68a3d56b0b52b855c7125a8de88ac436e46ff724a18b2d0fcb04cd94351e5bd6d56da4fa8eb8d5b2ca595cc2c25b0575ea5ca8e9472c1881aef886ab76875c7700274c2afbe3b01f13d5a29eb52f05cfac2396290792809f34e0c8245963008ec8f4f636e2466ddfb6077615862d3bb5d521f08874b9f302d22820652a3b746a07ffbd532286b9c54b9e3cafd3ca97e6f078c5653ab7bc42c4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4905bb649ef1690aa59e3f25c7243dce4be4f6980dbb46f33b6c474315768464681d965684051c7afff874865e8b17543a33a8630beab344fffc909ed8344cf5a1e21376b098045092d641efbce6a527d8a80b31b162f8488886f43a9f67e7489f04c9c016228f1072e7517776ba16fbf9d932715c51ca5b1a5ad6254b818992d520b5c263b113178f4473b511bd6cae915a6a1de68ffa5b62fadcd260b16bdeb86c2b30de3a6fbc899882df0a1fddc1a7723ed8251e9097bcbc74f2979e0464820a3ead3fe706b97249930dfa21237a3bef4460c131ec7a4a956137b5d9bdd34a3441662a0bcbdebb64f469d777bab0a6889c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h42c3eaeea20276960b2840dd407513cd03592a75b6e91ffd91f387313402f172769f00efeb2a912c7ae0f88a8192e45cb58803f332945cd468ad455e4ea13c8b17a0b5662c979e921a8eee21f46590ffbc368448757f1900b655522e634495ab6af486e75c9dea5d4d5e36de52e7b85d9d65a2c3d32591dbb52399f61fcaaa3c89ab6923f2125303c2406c80c0d7bebf566600e0d4fba15bfd9b7d0723b43f0214169b7e6c7e5e16be43595e91e26a5b106dc5376a0dae2d4341be832fae3743c6a7597a9e342f662b6cff813fb0c84b0811022412581dd17293dceaa60dfc86f5cd1d33b30bca57ddd0918d504ae72b6de1e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hb60942f755198c42efddf26fc2dabec644c0ac7a065450123fcc7f5b620d0034b5eeb5e2ecc7496c414357ba4a8009af115f5635aadf968b8cb70b8212146eb714822ca85b3b8bdea4c522dc7162dd4c185e539bf06f70b90480ce40b21c06cc43ec1085d445c0619c5c83f2900405ce6ebb0c4c5aeef852319a65c66dfdf5788d7d56bce994f76c0d42880346559a477cc25d34857849636aecea39a4d80d35c4c8ded9f865c106bd0ebcfa5d8f814954932672ebe338865dd0c58e8c218cd800e468be951d17602305daec315af8523d17deb0157b91d19aeefdd39b3f2684086b4110d941bcd3ccfff3ba62175bf98fc882;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf792da3546f2b7b738d1662a00814340c0e5072895d836b406963472e3cbdbe272440edbf69ac9f4fc00b588decbfeba55611aadd62c178a54b25a7782e3fd63e88024741f53943dce7926ba40c99d96ba63f45cb7517cac53f4856471c2ed92ceee3d40fc9abd75cb2e22d4124e0b550092330bddbdec6365168d52cd84cbe21c0f02001d6ef43da17dc4608d2ebd6adae37cb6aa651037c0957ece7a94158612ba30ea426b73711fa5f379aaee4bcbc04e94cd23846149ced16df6978643172a4e8cfc588449c25e826f41fcb9d9bb36d8f0d5e832d2deb5b6a61cfb6481c02ac9650b5268036f7b4b6d7657af1f89682d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h42648b9f73d121028869c189a15b635dd034ad35e1e32d1eb649751ec8b913a795855a91f43ebcf97207c88abc4e90b1a6eae99bb42df6296d8a63dcb8274d273684c1bc634ba411a0aea5ff55b138a6468c619686ee88de0648673d60f9d700494f1fdcef02883a78242643e879be3e63f76083bbf7de549592fb6c6f36205f8ccf39a078cbfd731652a08b5f28f9d7e4ddf0db082a2c6d265a2e5bee418bf5e67cbce376612d1fd212893c79bcfc22aef18990b4bf0eebce8852c98a1f9fceb466f9da50ec918b142c2b81fcb385890360ad1fe78a05eb71a2032848f92ba3ae970437b57ff7d694d49ffc44644e0d840498;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h516db14da032a634e802cc0725d914ad42f4d2e5e648542edd198219b6c16e393a57d615d802c74b25b5eb521e88e06149cc26e63d8acc0aa912e860309f3a27b406bcb74c3be48ad86ade51405832296772c5e0799db1ccee06fa63b7ba5544598ce10931e4c0cde390aa8f56f5c5cc705e8e47a3b07ca392174a67b99e3ad6249d78c3812c5a97b6c25a6879da16193b0c7ce201401101cd983c44f8b678f52296bc298a43f83ac1fa368dc710ac8208d8d41ea520b50880303d5f4b369d81ae932d5905a6f65980aac7dad0632c43b45ee20f5063d1480fe9a8e0e5a2ed77e9f8e36717b2ba94f2de1fba6d1204f81df426;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h55529b3ce9677fbd30de5a96a948cde2b3d5b38c8c5ba8e6df847b7fff236b6f49ddc93678a2631cd48d4b03e4d2b3c390abe15abdca39212ce88c19e722a73102e17f6b018858c1cda84c06973347ced1359dd6f2e108ab41c7ea338fa9be8032f6cddb0f7bc822617b6f48b3413a0e97bd63dffc6d2bf84c9f2f8f0d2a5f0bca2ea1904c72bf3ca0a681563c1b1019745199956b8ea08dea2e9ed32f4b9f36e21d8aa1ab655f342ec1fbde5743d5460ea5e15048e85e53d2f5964995077aa641d966a7dd4377755efd19510f1fe2d5a8995062fa0d9882fae9cf7b8eb50c9914c9c13db76c953e99c635996cbf9b4d539c5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hdc404bdaa5322fad1c8f12ba306846ab6a4becc33725f4947c22c6937023838f38abee9358b1d9e4b4df20a5e8cd4cf02b1aeb2185b3a3e5dec5ad65005214ad9eb416382180957e101d5cfb333ae510d25d2f6f9902d5da2ab5050a1e7b5c2818f30e44c822803cb6db6ef11cf418cd7525fc3f3bcacdc52680d9a25b6c3f8c11948c7c56e0568277e7234854607f48d994e9c423eb24caf5def73896f81cdaffa43fdd1a6bb0eb2aee9765ed5cb3697ad334ab166ef80ae9da13347c94e77279eca470bd988919b0c624e6b77c0618a293fad735071278d5f95870bf23424cb9c68867b82fcefb186409f01e9ce5f287853e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h86d95b0760f77aad614289841ac6cf1b8349bfc8e65d05b8419975cd4befafb2438c2dee2939d7306831859adfd32e9cbd825faa18f8cedfab7ff517f3840f8a496526e234e8d3e586dbd351c8c33394e75e49b34d455e10ab9928d55f9e982a3611d6aaa7fc1ca30a83f66f56014cfa125ab4707256a0423d426abee888b6417b06a00463f57df8207633ffcd13f7b4f1cbb8df4c7e9518a406ce057fdd031ed15b4e31adfbdde3f8fac0064e1c55f8d35c711dde789e3f1b1bdbec9dfd4d368934d6058a1c741848667edfabe08cd233bf6178ab719701e77296ae5ec5b21632a7c4623730d57e191cccff2386206fb8fbc;
        #1
        $finish();
    end
endmodule
