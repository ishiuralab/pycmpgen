module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [17:0] src19;
    reg [16:0] src20;
    reg [15:0] src21;
    reg [14:0] src22;
    reg [13:0] src23;
    reg [12:0] src24;
    reg [11:0] src25;
    reg [10:0] src26;
    reg [9:0] src27;
    reg [8:0] src28;
    reg [7:0] src29;
    reg [6:0] src30;
    reg [5:0] src31;
    reg [4:0] src32;
    reg [3:0] src33;
    reg [2:0] src34;
    reg [1:0] src35;
    reg [0:0] src36;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3])<<33) + ((src34[0] + src34[1] + src34[2])<<34) + ((src35[0] + src35[1])<<35) + ((src36[0])<<36);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c810f414fc2020dfe8e46d25439811177cdaa8a0cc8f8464788090f5211e966848e3eadc6ded25b3fa45cb392;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cabb71e055c5790312909084a1a9f7e56acea725c5a40a2d729fd06206eeeaecf0d8ed7c88fd42da225a690e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hadb3221c2b2e94ed128a315e360f2d5565475c0a7e1c0aa4fa47f0890914e765b1dc74c538d21deac66f78b9e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ece9c93f22ae9392028ac6cf365634f579c887ea6743bfdcd9745027bb502b3d61b7d30de12f44efff0546395a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34cbff662a35f5e66e0ddac86c7242474fa5a31661315a9e655e5d007207f55d464a34e112ebded275876bf1c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h723296ee05da1fa3dc17d74734b0e41f4f5d75e173df00135f50d04fc0495277bd113cb0c6d6d80da5f451c110;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1062d2e5a6a21911f7b6ca88a150dac1c7cd56187d3a3b5cf9e0e572bd5dbec4735fac04273541f9f007aa34be2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1955fe8e462bb7252eff33b9234e114e517e49bcb59fb58de03cb500a7729a8b90dd1c85fa72bcbc77cf964a7ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac1cf4b6661762c713abd3021042d81a651fef49c6cb79478ba8a0682b5655f081e657719637b524cdd42d0d1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de67e219aceb9ecfe3c10077582feb17d990318e11380148f745fb9c06636e867730478264fe026a62653839a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5c7fa5b0f543cd471f34ecb3a612784719cf01c0e662f737cbf807314dfcf65a7c72a719ab724bd5a2046c2c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b9c4930b0978d81ad1e1c101a22263bd5ef12a8f3973564de09eaa51bede27252032ba06902ad025e12148a16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8e3914054514c891467a3504d3200954c04c2b6fe9d95d947071e2f5b19db770cfbf5af964a972482b881fb3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34c50fe35ab4429b33aa9b159ce9ac7732fd4602cda4ed2eb0c5079b928795f8a981fd8f8e61b1d345a9c2f2dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc04c076ec7daad1d6f2aea276149ed23e6c0c95b77860021986603dbcf8df02c1b284a43f661713d6f934140b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ef5c33bb71c85428143409ac311db49066222a844a494c9bbd1a6412477d7e86ab97608629489fd19249b763c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d834f860cc6d4e8b97436bf8dd2c82387b531a07042a5e04799609076ff5db94435d21ccc01d984c4c20e267c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba0ace7e1883489293064397440d9e9e94ba0f1fcc06714581551497efd1c60390d3f49f71bc65952ac71478e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd43195c50a31e7c25a480e1ff12774708cf26f55d32f62444b3f33b0a1ff762dd8c8024e29216baff4ddacce16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1b91b5ef4c67378c38486276cf538adf05dc08bc56415a81a8467e044bbf592634da5a51566e0311a44d53d2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7caaca618d589fbeac161673b057aa327df934d9100964caf45bfb54208552089e3aee5a5e467b95d52fcce6b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29a90fd3ff130646aaa7d338110c61476257e7f3f01a1e257355288975e0a2b73ac3ef9b70f9db844709f3630b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc7b845eb2588af5f8320e11213a66eebf10e2af9a1f116e8ffe74b7306f214814f521478c90edbe3c4da2a2522;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82e441af12fe2f4907a7e7315ea9a4f80d0f7da1e7fa3df99e2468e53e38b511e81bbf32c033517fbb7d85f727;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf241cdf621cd560c789ff2a4f0de5c3d6621dddd08eced228da44d0e3c1bf4bbd427b1a965ff22fb72c947f9e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c347fd17be192b4af12a35a1cf0be3e87b461703089e4b9defe0293ac957f9c2ae8b46c5328040fe5a5aa3a9d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f3d745d07d6118bda24d2fe46c54e35abdd9e7f874ff386e97f5b04575e231e7708ba5bafc4c08e1c8e693219d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1081d5f6fd597b8a2384293de97aed26df564a3364466dfb3ed8be641efeb5ae8fc08bcefc775fb9666a8c68fbc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a41d6e3c05e7df3198eb66da969a91e0c07e876a82fe45cd4a87d699989b7874cd45b722ffdeab74d1f9c0b51;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181aa651d45c25022e253211893b384f8d714bcf2f0e4d08bca6598865518e14f0250178667b5e58be283fafe45;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d15de1df88de88cfc487c15bf0019ab05964a8135cc7187969a4f12976efbfb6cf39c4fcd5bb60092bbd580fe3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153f5e3fde5a667efed3c6f542c78312ece8e9fde9fb9e4cc467f7b89009babca75aee1950d1caecd19ab2bb08d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2cf25ac0da83259c468abc498e87229841419aae5d2ee189738e79daadd78cf51bc3f168fd495b920994b06d3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160ac51ca2796fbab3f701301b4f45fadf6ff0f0ec82e4198aae5477146e21ec21e1cef5adac3f8f9e0def96a2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64bb878fbd45a7018d1c94c73fb9a32a62fe81985c1047841c22a61cdf6a37ecc404d80623e482425e0449eb99;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cef0c137c0bbb410c3ed395957bba443fde0897e9ea45944250aecbc717cc8496f5bb15cc852c57f5f2cb2c7bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h179e875c50e1301fe6bb9ab37f59c5474382f39938b4541aabe2b0310558cbb9446d0954f3f51bf62624bda412d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcf6e3cb66ad23ea16c50b5d7f2da5f19337d2c551c8f5aa9047382e523922bdc39b072dfacdec3b6d5541dc8b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80822b87aa98237675dcf6d0d2fa670444a51eba9d6c3d61f93901826897da0c693cf109b43822027226a1e1cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7119d4f9fa88c55204aa1ab46460991f17746a38d44688d3636519122fe619c5bfbfaeb970a1b79ed924f41f34;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c92e96fe4473f783cec7babc097b9f0feac4c00ceb61d5f6f2ce30eb91988a3a8c9f78cb804018d27775ac9d84;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64e454c857ca968e170450f542b5ede51849a292b15f9d47a707fccd1c9617a0fb18b6d21f4953f31b27162b99;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8279f6eaed3621f483aa4c3e2029e99d8700ed8c790549b6b4154734ec33edb8ea9a76d2b3c2e9f843eccb02d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2470f1059d7a1e5b698f6b97f8d02e627840ceb309fdab0c4e56be83af6e78d3e9a84ee92539ec0a97856eeb9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h231efff511fc68ee3010603d8eb4ec7cee2e0ec29e3408c8bb835bf7f3aed4bf34db7fb862f22264c7a94017bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h635f097b92539a2c8a7a05631ed7eb41a220ca0aeb3e6e158e35188a1a98a0bf01a63e9d4d00d9b58690565566;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he563b895bed72295e1a894183067b91f2bfbfef9647069c1e4adf06963ca40ba48ebdad9599801607d8b7e91cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h674ce1cccc4dd91a29720a19634afda4ba589236495c511033be1dcb75cf75fe4cffc8eade1e59fb9dfe04ef1f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b2bfafe3887a020fad4e675296a4db9c461e5aef6ea8af13f297955da4610dae8e5da1504c11696f475f039f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c5fe92117b789738a83df7e8061bf412c237523745c75a451320b1ff09a4ce5d5d943a98ced519de93ca6091e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha78fbff66791e1b683e060461c02d6034f71b96adac523a1ff801be9a6ac9ec4face48e23245ce690fb80c757b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a25c7daed5b6133b02692844d88b7557d2bc7bcf59e839ee9a0a6656c28f26799a155f1f71ea37306801dadaa7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e724c470dcbdfcdbcedc776de0682b2c62d8c89714c8a35a5d5eccedfe76c2445f025e875f0f4cf0922e1defd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe493f5068ad001567b9aef4f7df5dc17d3660202ec3a5aae4ebaa7f1b594232e15a81b4a8b2613668c9cc72ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h130311c5485158d4eafacc11fb1d1a22752477e813cc231f14c69dfc7b7a117879124cfaeafa8d209b21581a42a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd261e88f0b7e46d13bc41ed85d395a18dc8cfb3c73a575b9e4575cdeabd8a11521b0f634e8b0cd20405024217f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b2e756cccb5482ec3ece80a64e53b1bacf6b9782d081afccdae6143a3914f35a6e892609a0263253e47cd7d23;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175bb1fe29186452d5289c9ea368558ecc3d2d5cbca2434387801ccd70b9e075040777270e93760754030cb9a50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf4071018774c4022c29c6a1322d3c232da273d62ba9b776f7b6a21dd127727dd537b2bd47ec26debed8ec93cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1048e9752c3da6b8120af392094756def50d28b4675d59ae29904c53e5dfa1613e564c63ddcc264a156717c7150;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4daef4edbbd0e8806529c64076e7f16a6f43b41cc352ce2a00d851647fb974ae55f6717a30783ce4eb2f123e05;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c098a1ef385534fea7853dd2eafe87603a91d15571768cc3300c5c69df1391a83ed82721ebfd1e77f33fe434c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143706dcdc96b5ff4df85ba1586a003b26c5c064e11045cb5d133f3558e53e13d08113cdc2e2aebc79de1dde63b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc7978a7e75dad1931eea10039110038a637da905e8f82bfac570e765d9727bbfef82f110573b68cfdfed929985;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab4a29d81701053b98ed51170ecbd115f0892b04643c9207d0736533d3c140ecfd655546a577b3cfb8b5569333;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c262d3e5e3165c896e53a2b660dd9c080356ab22f3122814afcec57c5688175355ae6167ab07cae621734b0894;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h152be95d1c0d48c4b48fff7854e312a6bf2d54c8a0e623cc7d7d9ff839244c655f0cf7ad463df510e1644ff56b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b383351bdcf678f32137bbceae2aa6c1f0b0ba99635882a51d748a87015c3cc2841ed1f5d21207df38726e90e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80331c70fc17d5038cbb389676d6a59245b72d31424df4eed10b53a33024a3f1a376eea32626584e08863092a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ba309263dcbb84fbd71b40e01c10ecc9b9131b03e80b06e0cddeb2ae1f2b74d6c7fe96b0705869661a78205ef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1034fdf1999808570d98a58e1522e04791ca7aca4e3279649b50afa74599a6598a6f7547d85c12fb2fda54b23e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he85c67900a84ebe04ce8e3d2dd6e26cd8ebc2e36918f0ec37c134488d89621d2cb2237489b8c20ef7e06e14bee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110d4ef16d7a2726430c97634ddb626c2ea913640cc73e1d14edf37873dee2ddc09289a84518dcf4878db835e81;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9fb5ff7bba75d883f29a774f6c0d4b4841cb51de81b22fa8656680f59387837234989a1441e5ee0fafc2127f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a58bf63136e19a626e33e08792cb2d985422d90c84b74617fbf04fa5de649242d265dc1f796aba9507e4be719;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15115089df14ffe991a9bafc92bb796e4c007bf4ff65f71254c2d79ed23c538eaf5cfa02c630e517caac59edc73;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c5b9fa4316b5ce46ae8dd8808f8f61e6d0beb26930de0c53e0a9b6dbe4945326bb71a620f9e59c6594bb3e90b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b52d6dc384d08faf8a35540a87c43839b5e142935469a6b775482ad33f98fa46b9ec7cc2ad6cfe7957d7cbf4f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75120e6cdef02f23031a45ac422c9ac704e3202b54a033c61f041239a22828776ad2639abe89a1e5d375c0632d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17543fcdad783c2c1cd6d4747043a2859257505ba9ee4876021f550d27b253169330af5443050c95d910f88a5af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e7e698932b4baecfa842fa15e4db8305aeec6638ddb39bc206c9d20ad51bb5e79404787266082e0c3b8f78f3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1261418d328d62b8909045510af2948df6b2b6a103bd11584f7929a8183b9d1e3d6a438879277ea64d1b0a661c0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19eed181eff538ad3d437f1615712469a18c0982c63d4cd97f9026331151b3956a8c31b9fbbaf0988d23a68e7bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1656375376f82fdd9b33a7fc100ba3886cc4d33104c0e257a7c3bb7a5842f56bc3d480aa6784396c39cd88b10;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dbdfd64692fdb95952a65f4deaf7dd82ba3866e0a1a1dcd9274fe731a671c400a13e354e36463dc3f9708966bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h180c183504b651e7fe7b34f2acdeaa896bc1bf1eb32227815ad4a83e82cb9d479ea47aa0d73493cf4756ff83ff2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9308868059b732d5908a822d5ce8545e374b99b24d71715bbf11def78e2a2b55a576b1b1cb24451760015ab97d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd9ddce68033009cc8abab8c2f2f79b5ef9a3762b9cf2ee3f29d27d9bf0fd7d36b44649ed4bdb8a8bb8943db1df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd3891424b35771971da2e651fe8792e40e6a7292a6049dcd5c4cfe14ae6e06dbf60293fc4793e86dd1ccad48d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f3da68a79bb70bd9e7bc8daf52978afc2d4de5faeb4210c10e242e41788b731507d67c0f17c7b5f2c855a89c09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca607cf1e667674b5ef5dd953c7242ccef5498b7f225b51d69b41dcf2a85713b6c2090f3ee2a248c5eba86ed50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1add2f7c086a5fd8a907b81c3d120c90aca6ac63e4e279acb4d9ccf94a76c65f79625082443325c9d11c3ee3432;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1132e653ce4be01a78c960bc33dce8386179b1260065d343709248f4d8a0f8358f6484e33194cd1e2383e4c84d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h516371be2123cc681b0b0709198e7180b4d0b13b198ca31eb2c8205b3e7675800ae7b1db59ee497a34fb049bb2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6716da30ac0af6c4d36a8b5de82fbae2f1acb3c4ade2359175c80e87d67ac33bc3f17dad831dc5b0a2fcf39fa4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2e88c63c11aefa471d99e1ac4c0b0bacc466c5b2a46c6a3c0dfc9ac6f9cc33a52aba279bf14b5e34929209f4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10320828abdff6baf24ba86c6459338c8d502e1e52d4d45e7d90b8525791ae39a471e061f2e675597219776eff3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1713070847431699f7eff165f62eada761298c82900f7e1dfb69827fb6a11cad7044b5b4baf54e889cbd4d890d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6670462315c76e6e307ce4d2934c2d7ede5eb902c9d722e429a2778213861298836cd038c0f67b5653d65e21e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1388f4e32ff3b704909600abf11e2e8a0dc41a0665ee435288ed187ade570e306c96031e61905a59fb3c97f745c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5642a3f110906d0857667db0178e47cb99a977c252f75ae32950fdc8905e85ea46d4c9791ff1ddd30f9189eca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6021379a992b915e7791cf6f4cc9359d481d3d212cb50e7034c2636994822471072c3ec8ea10d8232a0e2a4dd6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba76249299de871e64e1228182db8415c8aee941b927b0f8fc43fad8a5aeb3688c1d534a56f631231587a81926;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4af72b1a1a10e887208f2002cf816657ce05fae4a092d7a8d6fc6b8eed6df163550a0ed94609958b43b4e969af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2cda258a86565f192fa64f9de3829893333ad236ca3cde4ac252231a9acf42a0c0fcba5389fadd0d86df27f474;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4ca4717087a1a704aed5e1a0c57dd873da801473bfc825d735905024a282e5104b81df4ccd7b589dfd724793c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e54e77458b80aadf158699c2931e225356a184d45fcd3632606b226ed1477175603722fda6cd4dd09c2d9115f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f2c6012a96e607b97a60ef05837fcb09f1bea4057f303f86a3ca9829a0e9e6294634af8c642135a459f0172b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c61c1dca50c5c682bf92e6dcc0e2b430e220b18bc683c342382263e30931b04e06cd8488bd885c9031bec2bf2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6ac7b3070149238ad3f3cf932a33061eef51c4bcd1f071aacc1b205e9e78ec0ca9e15de2906aa703ead5c55ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e05a828aea6c1cf61a7c0c0d54a205b92509381b301f505189ca5516236908ce83567eaa63f691b2693b302fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16bbe76d561c171d46abc7f6d17b850eacae15df744aafcdecc9a00e24fde35771032bdd7f13aaa894a5911fb4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5c3872e64d37f90bb749534bc54c3a8dc287ea73a32f14bf1abfaa6c56c98d8e20547a71f55e9b09e46319187;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h40ca6a64919c6329ebaea2e2ea6c6e9952043a74322bfa8bfd08d3194fc8afc25566bc88c83c3c3d98287d6df2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he164b9cf9e680b4d9655428377aac9565e10df55a3cc62f23175a72901b5746994152eb18b2acdfd58833f872b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec167924e4a7b9b37c8dacfbe531c5266f7e3972f5623513367ce02b28e1098bb2cfc170fc4b0671fa79ed6e2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha038bc0d32f787b732e525bed355460748237ceeae0bc71daf25f38f93fffe8a7f40068af8397612a37bfd41df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he34106789acf5f29204de03b1a9aa75feb3ecdd60a2374b3caa45f6e94e5c2404ca71e39b05094a2031ed90d45;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1287d1740726f482adf30b511e83505e5368138c8d11b24f147a6d0661c041981a91f28e7e15540f821884c3e79;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c99d678bec656239d0074365fb3c8fdad517be9a6a91ae08e3e214831e3d49a86b87af9bf9546002ca0fafe5f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c1eb4e0c635ecadbbc8877ffdcbf698410136bea1c6539c35ab3d2bba0c9c594271956532b75f4a8415153830;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haba1a146466445ad07b832bcb1b957b7d1332457ca50f15becef6de286d4c899e7b90dc03686287c323748c6b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17105bedbb75b7a505f9fd2f4af93698f2ecb96783c635f2cca6fed494660fb404e04fa1f5178a90a010ce4aa61;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hec68880eb154d3d2e9e0b20a6e84e2006dfb2787f84877efaf92c0e9be31a0207044ee3ae99fe41074ce3bf644;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f64342a3ae33363788fc897de116ddaaa4ace0bb3f4383b2b674f35d6cea1fc5c6ebbb897715934e2952dd177;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4e0cb33ff0aea6c7bb6caf265327fbf7bfa3df9740e05672f7f72b104f9d406a228b64b5e72bac5ea20a54550;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1242be7846910637956b7bbe2a779d6ff68eb94cae081130626a62b17df0819a0677f864d637c7559a4ec740a1e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163587742688093856b013bf22cdeaa9dffd64c496cdcdadfffa323143bb9697bb5cd3d2e827b1a4e4401770b95;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6ff018923a628855c0fdae7454e7d4d884a4184514332f4d1001135c36a1db21ce34445d43671c94edf9a4be9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc222c876f4fdb1f5931e35a7e0e293be592e2f99e215961fa9a4e0c1f2dc8aab8245deb2ba8d1cdae0a169877b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ef5733630e7df1ce80d7c3acbe7cef9d9ac209c7640305b6a781a80e87fa51b94cd61b3e909cbf6c7bcd3cec7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b04ab14716212348483db2bd840c71b09f6c64d9b9be505d81bec67fb4188a5784ff0206bbc54bf5eca698fc51;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1379576d13ab1c4ab9df01319851bada63efd3179df3a11180690a0bbc35777d87a7e8a24d65d7e33b3f713e6c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67d603626724c03893f2491a1a5cfc38b8b001100b2032013161ee32e524f73736b078de4552f94c15881f2c67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1904c3bd1faef7e74929191a66350d3a6fa3f09e7bd1fc0e104223c571aaebc47482159ba3b80e2fa86a50a4432;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b63ac9592cbb8d8210fd5a3a86eadd9dfd02f5b5ab3b5c7b4d0299ed9b8e09cb82c95509a74640f2c512da2057;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc2df0dcf25e653d81175e47fa6010e2a3d77a7dd1d8824d337adfb0b97055beac0b29c59c55ce99e7fd2d206ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58ff91c04cb495b7aa2b41c051256ff81582e0df971c50496f149bd00e75a2b16268f9855a97d864b1d927cf8e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b60b9b9869e7b95a2050eec05464b7ad03d27f9262cbcc5c84db872f64d5fc882202a32f7838de2a929fa081f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc032098a0514fc6d9b12d4c91454a4f474487a93ba8e4cba0e814dfc99d94a7ce7011c40c1566251ec64c30bca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af9b58ebc0b5939fba46e7f6a70cce6daaa49f74ecdf89da714d062a082645e2f1253b9ba4c6dcd7fb53827c92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ca3e256c1d1df3f572fe31038e219af5ce242cfd102916f2ac06891faa24760dfb41151a5bfbd9bd47f4f71ef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd93b8b0b6f6519c4e070426c0694f83fee37226e034a13d328e393e11832435bf01e0a8253bbd1341f91a267ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1048306577efdbc2612cfe80d66f724668e9a16b490d3e24e4c85a962d802491c4803b8e3fe28f935a69462a7d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc3060da5c4c65f724bab96a4e47ebd116b24eb25c3efe8267827488a7dd6968a18ae549dffa188388e890182c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f93bdae2624b60a5fa4f0c52e85d594b909a81a7e82b358bb560c57613c4abc15cf2637856aae0aabae737a239;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20edb9109b807f20b0e1c30efb49779ab1de3e4cba095d4eee4284395bf9e1fb703df9aa0e0d323cbdb1fb2971;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3833d083058a830f0fbb5bf08fe088eb353f59394a6af8f29408f7f8d29e70223d91ec9a33a19b28fe68a778e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d8c1d339d6794097f3db9ef0572a3b16128324bc80f077f5f894c012687f8230fd7e90add3a55db508c6cf78f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1975d63f92f04fbc119b06a4ed82de1243cd338fc673a305013ce5ed1ab3d47ee904804bf7a3915ae7c1becb77d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f49e7daf0e585bb289f72f20b75618e3cf0058e9fe62c737fa8e811d177438a6f9bc1ce29df87cd35bb6dd5b4f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6de65044dddc8946b6b732481ef5a3f614d8ae8d7cd541e7da0161c2f8619d411fecc2ac250b87e0e1288d3d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac1bd344a158316ce84a8348db040497db4941dd7f47c6a1c3d869eb27f9732d58610cb901c1badae07dd579ba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3271319f46648ba6a7478f41172dd06b2050e2c563edac9fbd1a58c43078672647b4b503097834eb06f9e35ff9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce4607be792b94779846d4153db051f367e56089e232c62ef18a0b88a0b8038b7670d33787e2dbd13df1e4705d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h86646649aa77a83425eeecb0247fcb851efc3e6cac90391501fe29364920f11f97baf356c955cf6de0d36f6277;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2fb881ecb0f0c9b8a12cfac68265d0c7e383b3a146ab20959b60ccaa227ace0feb5e463cc2193d5dae1a6869f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a7b0f28675d5125954bc12598a674e7dca461bb80e64df7051fe4f01c2c809feb701797f3d02f80215bf29496;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17abef8fcd43effd767db9b0cd6f2a671b94d0ce5231c9321e0bc6e7b83fc79cd12f88cabe413ad2126dc7acfee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1176740cea1297abc0840a520a0c323fb97ba46a285db184681c6170c0dc5f58d438d02989edbdf693eee04cd8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a7595d30fb5dc0917661d4853b9159a20fd6e23e91f70a39403daa9db9978838ad4114f2783e0ea42c6dfaa71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffd6047a540c938ae84e2b730d1eeabb0c67a053e13eb9bb5cf42a5528f52c43711ff934264dc98a5980cc9727;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc6a4d2522721e9b21291e14681893adb9fddb745a4180d77cfda9ba47b1a3ac283c8659274b12d1b7ea6ab0bf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19390f5f44cb063cdf9b15d493ee2ad2d8e0a94ab6dbead8e3756139f363e933a99898241e862eb0e7338c7d82a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10b1ab471c083b8d7320eca5a55343ff9009b49ce760e2fac19d21a31fa0ce470bc624614314197466a39ee1171;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111018b8b4c878f90c9fb1de2ec46ceca75dd7e410aaa67907723109625262c3bdbe1862255269bf45b36887a2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5444fa728afa747f140841758e3cff715b4f30a33f504eec9a8d858e397d2bd640477d019bc9cdc8dde50f263b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f31499b5c48c407ce1d31723d9603c1d3f8fb65d6ca9aee5f7e077f261fd31cdaedf9e6671e3e7a26fadfba52;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b8a45b54392ed25ada10e2b83e2911ddade050537f9dadef9d73fd603ff821c0f31e83bdbedcf06888cbfed7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he915a402cd147145a7ca90719b189dde48a7a5bbcb92400f0baa8c2126c1cbdf879d4ddc3cc9f78c0394f2bf93;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8fccd9c1e9ae298a478886e192be136c9f246d9522f4821b455cf61d2843d0e4a0e9d9f595bf9dd70864d2621;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a477001cd507b935e02098be1362838c162cbda9f2b826d545a758a3ba090316e6ab2fa7604e2e780d73e248c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b728407c61888e8f8f3eda0809740ea65e9037e3be0f2fc1db666ec05707e2fa9f5529215d11ff0883de1bfad2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hccb54c13a8bb217f97ccae777365893973799cd6044b22f9dace5aabbca776ec00bc56d83f903a896adc07f536;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a911f02b7fa7491cb83793be8034c2c37f3dcc1f6a146f9765ede7f99264a71d7c5a2278623ddf4bbe8a2148ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae3712e2a94a26c4c98d9e9bf87ea1aa3554150ef7d5fba5a8f6fba39c206fa76c8de2f0ebc98e448c74a4e1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f5de8152763f3c0a03495e392f14032a56ae75ed6e85d015627ffba8ddde150240fab74fd547bcc98f3bfdd6f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ff7eead4287884b444ba68eba0d40160db2ce845be46ee01ec33469176ed4badfda79078472178b89066fde9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c76938b15f357f6d559baf2d7916555f411e79ab50f30215d4ea5dd190838b728fc016fc004e0e373184b0d17;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha26faf0ba603befc078ef17bbc926726d0d5a22cef36594b483879ff07050f03b86d722bb015db41a76854ad22;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d0ccc046e01755787c99a31b649891755222ab3d950bcff24c3fce25cf187987fca4ec40e8aa81746b7c237a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f6e4fd2ec0c541f4e37848a175aa27fc99b3fdf5c55eba2f9b6ec533ca3794a71ac8f985d698bbf759ca16f70;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5989506822ee6b317166ec9f792b40b76f179adcb417dd2135d8eb558d6ca9b0209e5b0d38b59eb980f140343b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11bd625fe3e64cd51310b6d1ecf1fbae80048285f775c68ed4c9c5406d296e657445dbe0e58ba1d2ac4e430d1f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1931d08947191d477fca711fd597527e400733f1ebff52a34ec976a4fe8a55920f124dd6f2a38e806133fdd2b39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68215b4e5ba504b51f19393e2d676099757dc23dcfe8c449626b7f69373e2ce7f69d1b5dee4b0b896ac74cc7f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17517eb78d02b47fd73559f23a8e1d1b2daacc7bc45e5e27cdcbd90e1e383408ef1e3d4c33adaadbfca54e850a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc250458c987168ffd97d25dc6b9138ab1bb98e71391fe909f9f5ec1d95b52dbb53cfd876b39bcd005c42aa2929;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf289398e5b6f2c029d0b18b218f081483d77d2ef2f040e006a6423ee2c5bbbb0175f650a37693dae65f97f21e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdb3f5d403aebe40681920740c2cbf484021f0783b7de12b56c5efb63274281bc2d416fd5cbd428a14207f6d8e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd5b832495fe91a5062071225dc8c99ccc15704f62c7b889415519ad13fd1e6c3c7f03e5de953201b37e5c2a57;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf72eba63383b1ea81b8f3eda08dfd3137501424669e0d2b99df5d0fcf217fe014754319dfac0e984db5a553b7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198c7084cf4d361c1fc9676adec794795dd46783a193a3b3bce7fd8adfcc01bb72405afaa080fed8f736091e60f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f883236341b13c0a9322b42c0f3b9e474354d8e4cd54370b5a7acaf9852f76f810029429818b722ecd0e9f42d3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1694cd6620a76870b1df8f65ba82823b8ad83361a1dbd5c0b18bb4031f182b76a7d9881a47c6b2220314ad415d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d144c98c40cfb55dde33fd652e7a23d7a36526e7b0bf7ccb5b61637bb7fb202a67f1658797e64f1e9e6e288e0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f43b7d282b353bda82cb0ee9fee72b2bd4f4f4593b7d16a2814b03d7a978d7604560a7d0af9b295ee65b204d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ded51df9e0528c7c69a7600646f6c2987edf17402b84c7b5d7fc97cd4b4b975feb56ddc06b4d8ce16b67bf5a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h100621658109a8f2db47a7f27d5502e33b81da04e0063b33e76fb175ebf4837d338ce776940711fc22fdab1be27;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd52bb6253678902cfc9ff34de62e0238b129de14ad2adada50af14780c84b2c19a5ac37b121dd867943c8511d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eed5c052b602e4ecdaddcede843b53fc4c46f2e5dee01aaabcd230d947f724d7aebf8e75bd2d48a975104f021d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17be99e014a0bb09082c5e2539698983cdfd8ca78bccfb37bbf6201e16ca9425bdb8307bb206775a24048cb0e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ae31281e282f20f1a37696d72e6deb1156a3de24ff775546cd67ebd2709d2798fb71d43b77194143723b4679d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd08e6519e318f24510e0201be5d596ffbbdbfd05c89cdff8ea35fc9df37b28d76e6284d35a3f36f96ec9332e3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15689a158f1b04628120f09b30756d26f1544dd10720e4e6c2eb4e2d636cb16c67624af72890ade1a74f6c2a689;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136d90b8afb113cc64ff81f552e044daca153dc2137b3dbbc8123788a230b7fba8dc71d2c4ff65e54c0a8e4206;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17617d09c12b509f9d06c7662fdb3efea0d80de64b3b558711ee28f2bd49c13f99f2d2b23b0db1beef8f3084af0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h973a62e85151cc92395fbeef01e4f94c4153a7dfacd6f5f9a283fb3a352bc4ea4f43a24b53434ed1f582e3a660;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca21cf22064fa68a5907d69b7e9396623839cef159f0aae885a3249890b2a6c6723c8c5253a88d874c846653cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114f1ad335fdcbe10faf4b9db39348bf086825ad1bd358dbc1d167d0f2c92b29d783ba150b2e3d7dea853ba318;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d6b941ab05074d87a1d6aa58dbba3066ce203541932a819cafdcfb0afa8109abb8d42b71cbfacb369f69834532;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2ae2af60f26a1c3643d860661e678482b0ea2f27351267697164f57a11367e11a999db94836572c5f0e9df066;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cd33b01308fe6cb18a6361534536c2a5b8c4df57572e34bab32576ff4107673ea2d23d570b050177ba58b6e07;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc706e0f1c314c5a77920ae43ec9ae4083f6a33a6e9071f1474d111ab0b746f28cb55dbf8a8f2f8641822855be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7b4c12469e14dce2da0818f44adcaa18ef43dc53b46738ccf7eeeb2ee8f7b9aa5e7923f4caf69b3c3402ea976;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193f3ae3a16ca1e53ebc56539598e95e0f9b210a1dcae14f03e3d31e62ef605b3cfe1d4c02a6973835d5f2f9173;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7ff87bbe5ddb28011be287ec06500fbd0744df2f6c384fe5ea613ca5d0a703d576b0c0b6b6ddcaec3affa2780;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h531b93c813d1ffe770b7bf54d8aa5b1499a68331f6b5540c264daaa237f5764407062b73e2e83f0eeeb2dc4282;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h647b11d8c0ae2a358ccc23dd0118e2af471a4c4043f086cc5ccd8bafde0c17b18639111e27219dc05d7a87e840;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf2a9203e8a0abb4fb15c983d7bfa112c3a304a0ab6965f918780dd07aa3c2d6be00a449d70e5f24d8fa27e6d27;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4217e7247cb1e7fc73d024c16cabf3e54ef2a8a4fa75187db06676ac750ed68ce8caf4282f5746853e236bd482;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae629d8f3cd62a4e802c6666e8549a9dc7ba73df7053eec87c425656b3a2684b9f3867d77bd67a691a6324c4f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ea52a7f1eb20327c3d68d14387f6129c1708926e7e6b8da9f0ed90ee308b137acd2b24ad1c473dd07ec70975c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1706aaef863e46449b548c98a4521d0867145cda14d5890d6aa430b28770a8f0b0a7da274be75c04eba304dfbb7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab991f789a38926ec928899980a6741adb4fd9fa1102a4a8050a62620e790edc33a67a9b22467c7a9d5cce305d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d5111c97bd522aad332279885977c1115c2097262119e76b7c81cd05c7a2f98103963253f8ba62f1e9577b032;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea9d42b6ca33bd2c23d39533472e1a4e4b74c6fd19d666b11b934954f112953c01f1643ab8dcc396cd56c6f513;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3bdfc174c6879a4be97b781d6a260587cfec0451bf2e9890842d142d935e47fd02a510f9f56e88fff69e84296;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a15ffe9916bb4f59801e3c1b7ff185967289c2e05e5a9f08f99c7ef14dcde4a60fda2624cc8457a23951060b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc2d977c8a5a5152596d55627bb05e2833a723b938f0f6742e1549d2eb1e266e47470c9fcbc68b6b84bb8e2d1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb93ed2f64b5270f558eb20c10ad3f8505c9c3593ef71e01e9932cfe46f5fe71e4d5aa0484f397e5ab2d9ffcd6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b188328552c28e2211b868e53f784e60d2b834ad318ab574aed752e7e88ad7d86780e7893d0290869ccd925655;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc02284c692d9c158835b224e13f83ba128f03a067909d69c316f5329992fd709d149ec817b2bf23acb2f81589;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5f63f3b9f948fdf7da8e72649a409d0603259476002979c02909da60c2c19167397f3068440189f19f05f93a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118dfcf61f65651cc7fc3637fc917ab029279691528ce1cc9e3caa5b03b765c51c90b561b299ed2a2eca5992396;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60d43fd752f41a6d76c9597bade3a804c6ba808a7947ff4c7e57bd3e30d96e9dccb977935300650c755530e805;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc613e66456d055925b82cb13b96ca51966d417635eb802a4bc148fa9c0d2b31d2e8dd0ed230b3bd739674b0a23;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc81396389f7e54f6085d66ee8ff009c4fa2f2e59b79dc15b566767b5c0217e318c2c359e177be54aaf0eb0e736;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b92a307e14cdf6ecb282186215937148d2ac12c8e6924f8a5c4157d69d0b074cb20db781f6e7dd6f3befa7020d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2187ed022bcf78be656ca773c7e59d9580ceb2bf3317e8e776f4c694f2a39df513b419c8bf2fc647a500fa5d36;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he28f0bae52fcadb561842964f512cdd6d27c84b7fa01ce8107cd2d14bec13d02d7cccd82e6d9b6e2cef33ad93d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b643b87c4ed4dc5f6f6a5b8e2307660a373a6c0ae8246707c7ce52cdd2a98de12e18b51bdb778b5b23f112f81;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43f0af7a95a6ee24c7d9ab85684a7e79153faf1f9dff3cf3b8e4334e074c0166b8f842a33267cd117320ca8aad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154a6e640fe26705ba2f1b660e34890d396da773f5cbcc0b41fc92f6b42703c9a30eec26c53dd545601d445c16f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e52fd18cfe378d86b63edd662c19456442c3dd40aec0ed837c5d90b3743ea9261857576f31089c6d2a255273c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16efa7a28ae1d30d46dc4b192d6095f201d22bd361f3d9203e0c35fe126f3da8ea8b0b60794d43a457e98c3afb0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1651ad1821ccc3ec30b70d20400bdf6d9543181a3134e77a56944cf606f4e351e8a0ebcd431aaa20141dca43d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41ab8d87a329062286561d418e40e6ab8d8c9c2bd18528192eafc3b782b0bd7a2e9407f9ee3498b7c4b5a2039c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b949c311a947987f6b8ae79c3cdf2e43a6da11483c154376f6192f813dd4f440e7201c506e35b41718e3f1aac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ce2a422aaaa579e4349afee15fbf2e281dabd8399515e11cac2f3de41661f502fc152e581fd98e8b4b23c45ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd2f04b14dc24287858559b4990b077b7cf74ddd576c7737be1f2adca7f2c3dcac7866b8484546f4968258160a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a2bf6e960131845a49f0ca9a529670d9f6edc4fd9948c22c98abc8a5e3d0c852dfcb12492b5d01ecde6e7e1fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10972be60116d9e5ae6f7b93f4aea718962c8483cb45e1bf37c9bc154757de3cff0119d573a5c42add434c15ebb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e4ac199774c83eee8aa0a3a5d585435201add57cd97f5935e19ffd509cfb3e5c6076bc45c76d0c9dc2fb79cdc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1206154cf9401c725fba3f275b5ab1d9fdee19d8393bc49afcba63fa3e7c4e7f9ed99cf785e8e09ade65253e3a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bcfd54945addb29199f3975407e659e583d2a74c778c3876f1b0ab2f1a4d1e75bfdc5618702557dc3a56af642;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170ca6b0581b057a94e8de600e4e42d455e98595fbad485c1eea4b87c143a4d97d64ecd115e5dcba2245e906d54;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e312a59b20b8097b1f5d484cf65e444e6acee87b87a9046d0d811327f25e636b349def807cc1dfe77fcc683dc6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0d13d8eedd4be01ab854d03c134b78fe7637dc1f6747ff9304a20d31b6f830754a55fcab9660757985e5049bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3512833d27460ee117ad12968a2b131c6da362c1553101cd940980ecd71fa6ed028fa690a2c91414857fc7c726;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be1343bdd1de0042c3d0a0e34bd79f8b3bb622df2a6b8690c62ad24e5171edd8cff3540d59dfb422094b43024b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42d949582806858bd8e8d43415ce36093dfb53c4ba395e37a1a8c96651dab899b14bd47b76664bb8b4c19d661;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150adfc05893dd17863f7db85f8be2835839f51ddc667f2aecc52ef42e3133b6f818c96397ab6215df5a764b4bf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1611822ca30f8da17398720dcecc363df389e12d5c18d4ee7cd16207bd84c4c0edf0f8ebdcc7c9782401fdbb10f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c932e6a1906ba685e23c1bc642603e3690c930bebc3d4465c74c6b4d807a723160e0b7420739a35e29f124812;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1119e9787e21b0d6b6e10f1bce971e30dd382c1adf5df8a8968f1b313f0efc2c8f2128b0460a23bc666baecdb05;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127025e08bd43b2d6691e54962edcb099ad6ac1d4e8dd513be842fafd2875a61f241f8c4b0f7c0319e604d7f474;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb1f4f2d72783deb41cc6e517415bd529d865774e861128fecbb1c38f7fe2a3f81834ddad9ecdfee0713471d0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33842734339df199a0da42a7511f3c039805b1729eb2bb1896fa22bf2b0eee1f0b14e4e49951ec607ad31d639a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha21812b828981a0c8e3e44cac33e7522c88e24785366e4143024f31c0d9f352a9aeb779dff905961805527ebb3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa7ce30ebb4202dcb2b9111df9d691780e1c40be82ed8ab32a9e7a4aeb4513e9dd88bec7ed3788de3a34b60c27;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd872d032e3e34d59dfa3015fab2db974ad3883b2582a2ce4886a4df5da46d9a802871f821076d937451ec91388;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h183ce517e2eb1c59ec10eb0d7dcdee8da777e765defcdeaf9323f1800a9bd21c1fe3bee6f6a778b739f7f5be5ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc3bb5300790fa5faaad16e9e32b67eebb01a409d2e008018771171a07c56161d8273764a4c76e516fea0e250b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9de15302963bcd5f5268a7dd292ead4bfd27b138004f2945c3e33640eb51cacda02951df3032c37fc7751c6c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h83d592302da7c7c35794aba287b02cc641719850ce6ba13943c09ecc9216398926a662f2f2d522e802d9682893;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a602fbc2efda331d7dbfafc3774b1ee533030cf7fc038bb8d37130861c59e7bd14df9cc9a0ff57ac59b0fac64;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1233f9326eeff9066e33e0bed540289c183fefa256b24f932718c64fbd0dea7b396a660fdb407fd9ffce29e6e30;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcbb2b3f1205056050be93d9837fcc1819d92f2901c00932436907bd3292c52df66027bd337e73a0b0c99d130d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8d048c05b92a0322300eb46ea566c4b3ca25f8024eea2090df49162a8bea6ef5a03e2347de0bf88150599e02c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h848fbb7c4e4cbac380e8fffae068559d8a603beda492a74ecd5954ea3d640a1d8ec3211120df45524459ca7209;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c60378aacc46602c10323a0d02367307ec3bd4d549e34b7f307872ebab8303a2c2afa05a18cf4b99a2a1fcbba7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2eebcb770c3cbadf8ea22953dd6ed91bfb7fa7ace7249444bb02912f23f9487856d6000ed1fff151ed381acbc2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab8c35ab86dd8547b4e1bcbdd354a5ff70cd7be7505fc77ff6fce5a88594840118c559c371bb6ff42b854d5830;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d434ee9ced8199dede56aec7c7b6c0d4ff23954c3b81e74bd31e5bc16b367f423af5b7e3e52c5cf07b30bf8456;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc0d71d6b24f73e9d885187d8d066207f29035452d3d08437543bad8e2639e824fc9b3d66f37ba9bfbb3b5abc5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ea13a4a225e003add225f7f939cd9f2102e7001153fb0230c7ad5f7a05b94e1cb4f574def39eccd1960eddb01;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba640075500d5fdf8cb6e99ab631d95b693a9deb2a92f96ff6d627d5110b20fe08bed108d1840e7d58a7783491;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10331067991b31e35555318fdd41ac1dff0bfe5ab07340d27cf8c1b61e4de0f3f226053a9afff9366f2315e4552;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca534874cabef2be26c29a50f80e049af68f0f7c14c063388b1c125dc1905c5e1522b9e05d0c6c6acc166e9b64;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ce6bf5b757c5e969ae13c9e9a482bdfc70b299913e5e90affdc6aca4f2415df496edf7eadcfeeda4fb961947c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4873bb16160d019a473e5b7601b13af2c1a8fcb95968e01604b7b90927955e17a6150fc1f107347a399c6a723a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1513cdad722504e41c86733e7b9da7cad977012041d2eb719647fb2a66efd24985afabbe9211a8f3454b2d3eac7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bc68014212eb255bb58498e4a3bd48ae885d519459f9ad406a7d18237df7814ed6e76d126817a1d17d320da12;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha45fa4e5839f688da4c1aa8ed388851329e5189309beb13434f9b5faa701d4ffa1a7f7032220dc40fcaab7d0d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4381f29899eb2c35c86c511ef893a82df8a05f981c169a729c9fcb9d2d32379f449f1c23715d4ddca8f3935d53;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1272ad30998c44eb3b39a98b739c1f7d1720fa9a765f34f00966b7840056bb64e817c8714353b485d64e8c9124b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1200f08a1af85ed850aea7828e4db698c37a08d1fa7f45327adef698126350cec4722ca088d3e254963d812ef26;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h32e21f5407e896401bdab3a31ccd7151033da3d06f7f537dcb176d97b489254a20b816bfd0fb58e6b466cd77;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cbcb14f2f5bf84fe9b2c1be6e0de8dbe35a66df4c4770b4bede0eb2fb1a844fda10623e240706dbd8e30a62ec4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1da63ccfd08a1b5c637dffd8adb991f9f25abe282c7e50b86330a1019ca681342b438327edb970d16ff8b71acbd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h158d40493d5c35fe08e721d60e5a3c0a4c446d1d09d630b1eeef10adbb1dfe67d01dd55f72e680b833b21e32a2e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b105dd858c87924ef110e821fd96e487f47ad4c9454e5b5fda80d3c3483ed725c03d422e526d84358c5e6725b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ced4ede8e55f7ef054ee719903a0eaf0771ba0c4a29e753cc2aef9fe8e49417e9353a7b674a929f3a708d393d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6158c632a7ccc2f5eec36c50f3b5e329fd8ddbc4ae8cd4bb1a3c0b9e09ef087646a529c9855492b132664257de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1482fa930209726ac3e64f29ad6bb1226370e79b4e38e3ee7b6aca51142cc82439713187dfc51e76f3ac2140631;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h518504466ee54fd9e6d7b4013a5f9fc54e237e08bc7e989f4a9bf335bf00d6fe7262c59ae02ef66664183cfb54;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h46310363adcac5d118d74c4bfd2d6cb73ac1f3ec4efd25f32834f0308318db9c8c97c34d3442d0da5bf64a791f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1adace49bb443c925613c6cdcbaf78b61a9f183c66f14c33bc4873465df173ae0c3da0d9a2ca02824157f9c3a18;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eee00e6e5fe9eb6c7b665fe94e173cb2b254bd4927652ab62d2b1621549fe6ee6664d36bae28708dbe44b9e434;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1141a9c08877ba58303693171d167be80cc933a9b85985304b6eca3a81970f70f12da94ab5056fdeee0752ff9a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25271c44e0f22640aefdc7cb83a396b2385a718fbefe56bd9a33ee79d9681a51630b4dffedda6c58b7695ee271;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3cc2bded2dc380a5bb5b62c4f55662a86988c49b9c84f3b3d73aec147917c1cbc909e1b2e0ffa6af238869340e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1034030197c9b710f80b817312a00169cdbf991df901460f6ef6063fac8e36505cdcdf4d2c3b457251259f1c1dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1977f8705f894037f7f8efde2f7a63e2c30d558e521fa86ed3b215025a1e6a8046d06f8aeaac30cc9561ef3485a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1582345892b75bf217b4f88141327f18221efb676c9ee3e68a6535926f91f105143a2b1285172dcad95867fd2a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa59c31f9fc68184ad69da9869f921b0d915e5be5def746e881b2907b68d274618c734a37157e962ff2bde97e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd283c7f19f29af925db112ab7813b3ec443156879f58de279ceee8596b01889e63f7ac8616b7f3d635e692f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193c272a8181ddd907c5ceba358df1217c1594ea94f9d221153623d79a65401dc00e064204bd45e799aea40064b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f50baee37bfb5659f7f7f5323e64b86b259e601921983f21d058fdc20bc9849802a850a36cb6616a16127a9eed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc53dc7bf52c8c51e2a2adbd23470d6a857093a119ea0efd000054798d6ed6d267d76b53a924f821e0e1920422b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a864b33130a368bb9b4e0e712f7cbe66ff91340fa32a2669ee94971979f813ebda55962c72d1cafb525d2f65d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca2ac825ffc8ba312f9ddebd1c3b2dfbff41df0285ced1db3376acb282be31297fd9c8dbb6fc1b16369a74284e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f3cb0cbd382d12590b415250151d92cdda34ef88c1a7b390b7aef0e629f4de0627fbcb31e7da665cb9c372980;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h176e9de25591a645e43266f819cf0196f9a8a4787a0741670ed24be564a0b75eb899b731dfe7c6baa494d47d23f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b037d9803f720cfb91068a2ebd3f1534d3bdcb12a33876182a921df58f3f46130bf31acf0c93933ec2707f7f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116fa5c285c6e59861f443e4ee13718767f2a49d6c1b9dea7ec042a9434af71e316deedfc1a20430fa007e923dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bb12af2d61efc1a7200d1d8dd1a387f562aaab428b680d4ffa94be79c1d4aab1dd1c9f80d4da9a39feec5c3fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5216c16d40dac0742e0777fc86d4ca818774adfa03e9a8a396be5bfe6f1083f6ae7c7849cf58e202db6964819;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h151496b1a8bcdfcc39a2014018b6d766390e507c02408f8e1395fd3263f1d62ad11c0084ab676800a13007e3e71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb10c9f6ad657dd903090df55468d075bb2060ad4175570619b3c56a39ffb5733949a46af02b7705792ccf46a1d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184069518bdb50b45c084c26b5fb5ecf3988328d0a7dfc633a7cb2462f8a77e1a911eff59ed9f7c56379544bd3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1388c98c0b1ac9c8b741b172d9723619d18527200bc09b8286d521b503e41854629c62eacd2779605495cd65ca9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5673bb20d7c1de007a334413454e02bab2bca8160804912d4bacbcf570ef84078e961c97d5f69eb00069507b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41b8437b8a8ecd7b02a032ff4fc114f847ff164e13c0466d2b1fc0f297840861f9a453afb07f5ca3293dd01339;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f906ba565ef2c86020c758a2ff953df01b6e5bca788ba7b5b5fe4bdd85b69a375ea27612a2112e5ed9f3e5778d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f68ed63bec22927eb9ffd581acf7b4bd5a49afb11229a939d6e88cbded5d477f8ca32833dceea7e17d3568f283;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5404364ea90f3e6759086a7dd1089502e7d1d3769c6aedf9a2a20a3653e0b2878ebf7cd10f6193d8fa4265b4a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b75d6ee00086aef277bb7cc9dfe1197013a88040ce1f6b260deed8c90b5e42de90459d886e86c9dbcb83935bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18432031c2a3a9ada3cf576159242db0637091f98d19696cbe3423d8344d610a8c3797e3a3f19e6f59c3ed24996;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64ea6c34f5d4c895c1c79b931d7af3d2b0c44c0db9c802125744e78da004e5621dfa7a0590e2f621ab55d22148;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33009312ab49c5faf92339195701e5a7a864a00e674911199c0eaf358388ec28f659bab9a0cab802aeb7958846;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7e1f58e84f385d6f0d49aa11214462fa98b268c9ca75f17ac1342c2821e118e98d50e94854e886fd347924df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14bebf91aa454ab77c07547f07ec79fb4ad9dde2ecfc88bf466fd437346d51d209138a4e60e8287a9403e2dd2a2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118e508661fb1b81dfa3a104def56ce808730d6c386bc1d2a675f4a570a902449ce6567f460acf3180115032178;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b99c6283977ed98205bc1cfb7ad50d340f56b0785ddb813a10359fe15f3978990e33021571ecbe25e33054f56;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134caab5d593817d3599d1c2fad1d3a51b5de9e5bd663358ed3b3c7394fd1e71c447fdb3410448345f999acdc1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fd7861f29845c04108bf3e2511f324109bf4f679007f7cad7c2123fe90d81cd9c47fcdf723b472d219b62c1916;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5e5120366fb6bf44ccd33a283e2ad67b73a1b9d18d72c1294829c7915605f7ea98dbd11cc8f87fa1047b096eb8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h710820d6d25c88303a8c46ddead39ce631c96114f0ff6b94427d338d22128fc335df72c57a7931ab6d8a10e077;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138647e24df80613d879a41a43968e493b58f93c8dee7e35bf1509a9f99c18129b0eddbb25dc0d96972226ab89;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2faef06b8307e483f3295f3f09fe97135d5c1b19048c3515ba72500f11416dbb26224c90326663c21502fc827;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185e814441f93f7ad3d2df15800743959a446622c2f8b1f3995d9022fcfbb24b5f366aae1e2c0675eec8800554c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15dd5556eeb0d58dd6d9056bca79a092349e46ce4cfe9d26059499486694feecddf3a01b383e20fe18f9dcd98db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42b6faf6ac0679531c65a614f2f29faff385607b36ed5fa5afd028154c11dd8b239f66fd5a8808d32f78695c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h123c05eaea6063419c8a9db33e7aaf6d2d7744b9ab966ed53caec35224c676bd2a12a603f01cbde98a3c3a1ba77;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h321fb799ce7fed4ddc9d51d128460706cdcec14a6084334f7a0292f064e0bf72be00e9fd9860879d783bb2cec0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ef78e3a9f3dd71618c38d51408043ac7f6bf61d024d37f9457def5b0d48b270d7388a079e96445b521791c5e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9591e70b4cb4202778b433c7ad5276ef20740536a34f8d9ce781f32f3cd7fb02ffbb5e18404cb9b5def103efa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19e4e84f53a72c2e446c720b237056e3c25519747e2f5f32765a4cf139635f89d4c7807e3ef5b37c9dcdc1f9b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128116f158b74995c1f776d52342df3d34ce5b4f8f02c5e085e64a9386488f3d2da0ac09428120328c9f586ba56;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb4a213ae18d021fbb8a1d9af842d3d7c71f80483293763d1ee94ec9217535768ca7fdcfde9e010774f465a79d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11525f1aeb1bf480bec5c9c855f2f77dc23eb06fc333ff1d29370cfc44c3239502e0628313534c8962e914751ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d70d8557b8b7d5d4cd546fa8d03591112a5690b9385289968963655b9478ed386c8b092d60fe83c77365db11a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdee4486103943b9e020b609d663e0543d510738ae0d33be10910d0470c8ab6fa8ac505776ae33be941226127df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc78f39dd37af6b6df8604d8907350cf19e54569af4d4e23007d08199d3a1fdbd6cfbdec7775c09fed19b9fe5eb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ca63b0761eceeefebffb8c82fe5547b101260c894d54c4537e4511cfc71fffa7e811f2f8f1a11843c8a0a66cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha9fb2e06191adf1ff763dd380e254567d1e1077b0a3dfbb8483fb5044a868ad6156127daba2e54415bec980cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h152757a445253c53b0be77790fce7b6843f2c533b759bdf8fd5ea76f3c700001149443a6d84f862fd467e8645e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d136757958bb05735321a1b9869b5acb49601646b9474b3d34be391f364bee42e1da44e600d9007069bfa0a5f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14db40dba51f1895d2f4e01576b94667d0cebc9bc2f694bf3c552ea2ebc4aba1aa5c7b6d25dfce1eda28b57e8d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h171cb2a70b0e673a97097013413311aadd61a39336ef14c989be64c1300a7d132bdd5954b8d127cfc5a31e2e4e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4fbfeb3df554016a0569e16b9b5bd3a5fe6ca2d3148852fc6f567434d061c31e426e6999b3beaa046b8e31a65a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187faa6c3294e144c88741ad715f57d7086186a9b1a39dec8eb4a43b0da003bdd3112d97326bae7c6066cbe48d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12be7b5b33208aea2b9baa4c9ee5c9cba2aa1deb34d8e8fd363b07b44a536793b8d33054dbf5b9686c1fa6e5ef5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142a59bf6ff5628425a24b61160d60fb8a7b4d2e69aec6698db1ce801c9ccef6a53082ed6349a763c1eb1861f39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6b248fcc44bb69ec031f1b501275a4a403e641ca14b7af39135b40506b8e37d2e63b8a55df7f6a975424617c14;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1183b69a0a019e6ca86210924abb5fab855bcec712337691abf748ec7f43a8d424ffb9fb94eb6a24603cebf82a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he9cec7cb200d81993b9087006aed063053a43ae9d87af603feebfa1f011c8a416e2431153ee808e0e63c577038;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac46a6cfdf8f862a4a4277cfac1507fdf7a03cc90cde76ba670ae0da0eabfd8f2fbfd708cf77c63bcdac50c4d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbdcb2bdaebd0671f903d88fbcf16e534edff6026c49741652ddfd28c690c32ccf4bfeaac0917aeb0b5c6438ea8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf3ea71cb3a1aaa526d215b75e9c9cef358f0cf4e8147b488eb09b25a246c7d65a4f87552d5388a2e66a96d215;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hceaafc27faf649786e813282bdf1ed5e17a9bd56be099bec905747ec5e53b256a8f445813308ab3933d0cc3236;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa90acc065fa353de73c25c3815b95601d118f090b539abffdcf97aa023f723e699f46cb7034063ba16df18395;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133ededdef98cf4c8cabdae4d127878f449e1346f549912b7fe3dc9972eb8c962757380330e32425fba3bc45983;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9dad015b2291aa84637a04f7a6b29cf4c5f491c5bcc0b99f040de1567a70973fad1303f080e00a165b306ed6fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h492a2ddc239b408086825fbcc2075b49e2b501badf748dd72a9e61f3f671ae3fb5daef334b88254772b466531e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4f30d1d7e8fc8aa6bb1f8ef03201d820a787170d5a2e4430a937aeb1ac1f7ec7db5c30ef0a5a61bcc9b8d0851;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f9ca73fb341d5467820bb933b327d7617f8f945844a3f78dd85e25d19c2695be1651170578b144e67d7a6bd57;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd9d98ef2a357057b2bb3c8c814a84616e5548411ba8cdadc7e510c0e1050ab3e2aec87963cd43dc57472f75a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2a9e7193444715bf8e890f60d7b6a65aacbe14e793a88675faddfaf31ae85c7cb77db73c23329136869917523;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe0fec8a395256693b1aa1d5ec920bf8d29e9ffc7a9baddeb74430c5b8ed7908c84f31db928210a55acdeee2a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd0aa9e3eee2dc5b4c193ce79f127e9eed2a4364f97d88c5c4d04ba5e4e1a8775b2082de0fee073235956851b14;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe5b2b04e5616b6ff90c640c61875b2a630f3871c79d6fc5bb0106aff126837765ed44bad3080bfac02714e37f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d5dd258949b7d48c105c3c44fbbf03d1af61add11c53c6484f206e0e68b9155c0cce4091e075ebd166c51fd04;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1971048825ccf0ca8a3288ad976aad0f4e23b49d5d2f8912d7e825e11aa1d2b378c991a33a822a86ebc07dfe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7e4e02c8f18877c8afda6c03195defdbbcc5b0542e74a6dac906004a9cd77b7829b4e4e51c748d6ad597e88b8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1139a51598c1944cc0f2484dfa0acc31f1205df7301d03747ad628d163208cc0bdf8789338a87734c692477c97b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b88b75b875fc27ec47b85c29c190f36f4306267e7b540083828cd5f4155caa7bd974c68126ff38c701604f3c7a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hafd88a925418f19b65e286190183d427efa2f24fae216d00dfd6dbb2c0aacc389ca9103bcd9f08cb76974a3c0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b0b00c809a526b72c5ba7af2323973a82f834e00806eccb9179dd46c46bb6598480f849c2e4f7ce85a80c54112;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118343e6247bcde52403a4e6412332fcb419e4d8d9f82c8c4f1037c0a172f94757727e9b0ac9a91084e74d0b218;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c174451c104364372c77a37cf6490911dbb0ed0c603fff02e3a00042e8e3f5ad97914b2a5c67e72554d243ecb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cbd62ed4c44fcae3e8284daaa7f0b205b8302f9e1b3f192ec1b7a1d8f27a068e5b7d7075bae6f3108de965e0a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17cabd0cde7c608fd2fd79b856cdd8f3fe5dd5ad362cd7f0bd004c96d626d6521b8a8a2b52ca48fb7ffee9b7881;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a3bbdbe11b62a9e6d469d3ef2e5a031d45ce16e940831da5f3abd2e60040141b9a13609d689a752094c854e86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138f911a266258048d559af17fad986eb0d3aec484eb8ba4bc4b7592ece0878b69c34f1e17a540260bdf86b56a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d8979858e268cf37f2b7a0a8a3836d380b9b032f9ea6c1d2c20193d777f6795b4cf75d5e01300dc81858d5137;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d9208504d3279e9ec70eb798be95f8a028c285f9e812d83b139a5c61b968660d658228cf78400e00510432f5d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b8c2923248fe823b0ee41ae7e8cf7904cedb4c34792ed43c32cbbc998ff53cfefe0e72b4ba56221ca135eb17c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11621f21630bff4ec91428f58c28449883c1d3b4234d752c3239d5765cf9da24d6484a4931a1f58f1b0e006f942;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf1d951dbffd986704ec6faffec7e2afb5af5756ce1e60383b58abac3b47d96e3b185571ce4836f407461f9a3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc65650a86726877d80df96026adb224ad9be4ddff4a2bbf71c2307602433b182609b5df68e9f25602dfc37a086;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ce3502b567664c7c26cdc1bf290d62e9065547951e3b5170a1af3467f7b2673c20133c8f887cbe4f94beaedc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b96e684a2413542248c43e0cfb744dab76b331f8644239bb646023a68665987d7c306e65889ed5fbf512c6298;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hffbe932587e46c5d670e150b0cd057936aeadcc00c5fe8e379a6e7e37b082ac1023ff59c3eeb0a9e302e2651b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2155f3f7de8ba125891b76590c6813070345956d108ffee726dcc55ada7e2615b00103aea0544c190e639be3cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34af2a209a0f8fe210485599d1b7f641acf654babb5e2a7cbabc1b9def0b7f05b8bc29beca0fc80719f89f6f0d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132c8b3df040e8fc0a2be80f7c6642356f4ceb357fa408552fc3d32c12b20e45706e86c4e188e777d5995432d7e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8de69f788d99ff6c2f3d7e3c3b0d9217914ccaae3c0aa9cda6ead1c7c838dff3967d4be4b155d1c91fa361b497;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b8f3dfcf8b860fab84e3d37436f1c3ed1aa6cf2e92b846c11be56329518a12e81f004dd6f2be57867b5ddaf78;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha859b795a15617f5984398fa92bb325e6342d043353525f7d4a7a3ff0b343af6ebc8dd7d6cb688f676799e8c7d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e5e262040ea8516c895da937aa5d39e3dc0a33559362e996bd55b6b7ec7adfaa4a2d66cf975d5c77066a4ed6d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b26bc99e939ba5d74623b91c3ddf4754582469e9bd57719e9564cce9297d1883c55be07d4fb7392f39d50c6a2b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1620113bb4c4ea646210db08fe00cb9e66e22cffa6eac905b1db384e99a08b2392e6ba268c088fafc9ad5733f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e80c68389a9d08e12db50fe1fccc5f926c01dffb7b58b98fc974deaa693ae26fd4d6fec25f7f5d2f5a4e7cf376;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51934a6bdbd305a79f798422e20da43049f6a5a6d54526a39f0d91afc2db1a9fb89f1c6d3fa8375a77e1d173cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4af72088049adb8c25e76bc1ee80bd0a30e1d302c2d31a318679e25b9b57382f0942bcf3e077de65cac9c36aaa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5256134c41d52cc7fa163be0e738b0e181ab460e353ba4a9323d443d2ce44cc8dcf4781e6b3edeb83645fb162;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b27e4ef3b05d533345187847ed4ca161acca34673bbc77c11ff10c379fc1647eb44bc9a37cf9d59d9ab4618083;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149f32e93fd965b909f6b013d06b82ea63693fc55e1fb7051414b86db4516a3f2d561e7c062263c10c51c6d1d00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199635350e9a4a3728ff5414d43f407959a1428228b52be5ab49f8faa95ae6ee582da7c47dd51cbbc0e04b9578e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2443ed3ad603a8af9bdd53b750d0fa91d758b1977179b360ecd95ada8c11ffb5c250924d950e450c37505812d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93326f479a4efa6fe70311e824f889962409e86228c9f786ed7d1b03510601d2206215e693b255775864e2d24e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b0ffb3618c09800f5f977281ac1b01996068641db74b4f7c1d8b40503850814d3efe6035643cec414bb0765b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f443a3f12adae8492b71d4c3342cc41cddb07d1725fc7ce3b649d6fc89341caf9d2e210d5d89facc017cfcbb1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a5a419542678e5c2d03fdf3dfad5d53d60824d5574d1191f6a683787e3799f065b0cdf9374247f5605d842608;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147b3c79bfc7a3e7fdf664605d9b73e30fdd951809e5d7e5ba02b7d4c2952290b2665473afe4d556a9fa9c60864;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5a21aac8b1ffad41cd7329716becb76d2648e6a7a88698497897814e7708dda920ced596a7f28c4e6b574ef74;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58242619df65b6c5f72f7b15ace8fc98a78a6262b95f868f12931913b4fa4c3a85f44728fe3a2942ca32ab8385;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc8542e04948b69a633006d3ca8d3946b6345d2de69439f258b64ba10da28b681ba7a6810425467e8038fa93546;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h173904da79e06a9ff604d2d453a22468228d770c86ea59d891a83a06c296b4b3a443c952005c74b40d7a1e3c54a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112bb5a62e872702292adb059809e5d2902ab178c925a48943bcc1d5051ef5d43823c451fe27026243b2c4cfe6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160f689e39848b5f0297731afeceb34d2184ac0b972ac81fb4ae4b3a55ecec70dcd6c70e36b805f7bbe93c38843;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16cbdfa504d6b78e43e23060cc5d0365b2d71e1022878f8cc9084475adc30d0fcbb8befb55c24e9862bb9c1b052;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20d3d3d4595729a9d387ba02820f8ec35ed4cd0b173d3233f0cd4579a149677967fd46d27669f931e05be7e90c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4b36fde23a60de7e4f3053e3b5cff9f50bfc0bba7686b9efc861016e5e968d16f6c9c4a5ab65e55ee4eb142b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h824f0c02650269b73fa48c7fe3f2d61c08fffda5bb6fdef3322dddb205c05a42915ca6f585d51f88cf05a5e8a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12e56f4ebda4065e5021338252aab59f7d8080339f0450b362ff353669b59c21168ec1418f908973be2f42ee54a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h470faf5f91a7b766c78d3c31638c2b79d869857286e05a0cd7cabf90701bd2cce9a48bb2e50f67d5720a0fe1ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h151d3ec34bb46850ffcaeec4d21cf0a209047d63807aba6e17d619532741e893ed2e49aa947c1c54b5ea8f4ea3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b690abe48d24df5473eadb9fbfc39c2deebeaf022dfc373eefc68d6acb2c76905c1abd87237f1d61bc616edcbe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae83d195a71c34da444a91c382a2d68235c3924bffcdfa0ec564d732c84d9462e23e2be5116d6b6f1e15847e40;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f41c6db59c4aab7c8978697b322703049bc83e1df003c9ceda77e897014c69a9d2b0e632ea852d72f3d26f3ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3bc7130d0079e24fcc39ac289715c50a974a901d30ece207cf09aac2ba0d79e189bac5e4b073b17f90e9b4df89;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18efb02cb5329e80594a42d4a4b4630789bd51d0f9209edbbd544bc16b7fc38c98856ddcd7a41bb6baae773679e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37e4dc55d44c29ccad5e415d71c4b9577a5d73c950ea871e657dc2758ae6dfa29f7ccbc0e646212304a61eb139;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ed3ff1730ba4e43937787e09381fbb9e75935943a7869bc35315eab4a0b73d4ea6cb257e61caf139adc0313dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd03741caed76e4f2121d660fe0e3a72a8a8ff3a79f305379c5d6cc71dc4ca1a15160b0158c58d3a6b60e4f759;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6636f3f8f760ff022277cfbbae5ad7f9045dfcd182e85512e7e93199ac8e7c93d8091517ab00e636e01460cbef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb15d4e7c0b164481153cf84670f62c98e5b2c8e03cbe3c38283479f6bcf4a86840543e0edf21e9d770ef8115e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae680370a47799de7fdd7bf2f436eb9b40f5236c905471ad78128f08b4bc9375635444bb360092d8023cc82c9d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ecde1fff44d33100f6ba6b9f90cd2edeeaf542e968422fc8e900c1d96a626ed9fbcfda6b550a19e58f40f774b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc038db36e9112b5752f9fb12eefc40ff8c6def59d3d8863fcdbe69efefb3d0bc0d7c3db55ff9f71a18b3760622;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he80d9c0e3aa3dd8b72cd545dbe156fe73e0202ecb19be6c634cc56cb0ff785887379b7362302b9d35ed1b78f91;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4ecdbedc2dd5aef93b50c71af43eaab41ba766f14d09368386df36da8d3f289068b7f81d28037835383c137341;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1866e499c3295d41555c741c51ee6cd3f5577bc00a41d15f2309a02d56d12200e0d8616d9551e2d027ce0322792;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e39c78610eded465cf19fabf4155c07a1568fd9c6c2df66edf59ea6cad47157e6eb944a51dde112b41f620b3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h445b8e14b4393640e981d2fd04d0e5717cfd272ceb18fa2ccd469df46f4f0be37ea8ccd7185928621426c2a5a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he699a2f23414f67d49b67e511df71cca516a235c13cc79549f7b2511e323b098f301ddda123a160eaa6a78bab0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c6e04f799c378eaffc58f7b276f0a505a54f7d1aa5549f6aa47524615b6ed65e47b6e7da9f6047dc4f8fcf3dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167e69a14b4416a52aea9ac42f058429de735e727847703398d77a6fc2a82817abd5e7ada8beb5c01b2f39cdb5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4fc4d5011e5833f64a312ccce95302615ae258d9d4d5d2da7f3cae19dadcdc15e7685d14b3d1a4f5b846bc42b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h32fe5e34dac471e57d0c07974be47f789b86705fa925896182c4db30f9406fa851ffa608814e8b66ad05834504;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heba11e502440ee2c7d0d375359fd84cf2608a581566c2bb2bd909835e42cb8005a41469d692e3b5f358523a6e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170e33f1133616eec13207d6f37b2245dd63ea694a2b2444b4f5ff5eafb2afdc6eded9d43d21d8e872f127fd1a8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d011e1d4bc038bb433bf43f419d564abcbd7967e2e7fc4ee674d3bd2efdce2bcf8e2b3ad6e51646511f6ca2aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cd2b97d40c151f349f00c0a1fb6936bd7bbf0f85397036b468d1891d31f2da6ba724c7b2ed927cc85656409b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc79fe857e789352232d9f8704a41cdca2f1ae97d567f56ec75e26a7f92e5e91bbd63411a24e285001d0f23c196;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4ef8794542b27b6156f512db716a0083c3eb3ca5ede7a09db0317c21459808295d85916429c411a86a7a8321f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e27c6a75b7c7dafbfd118f2de43c38af1238323259ab59cce6f7d319d257cf0baba0a22ce7ef41adb79ff781d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63cb76ac6ab31bed97be6f60f1d5a7b7277d8b61ca41818ddacb4e8173476fba7f0434de826f091c08c1d16805;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1442b5bf7804642888b9b28c91e701642a824450c527a38f2109c575770cd72085b18f2c651d5b63e523f20e2e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16f00b3c43f314826d8d3cfff66a9ece87e9951e958658ea934a8009523e53a7f92373c00462da6c1467633ad7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h970807fb8ecc1b600095271b450e7a130a920991b12b9446ec8843a1e28fbfdfb9ec8819aa88bfda471202497;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h446abe201bd9d05edd5ea092ad6dd62909d8b7411f10c98a8022ab4cf47c47255082b11ff5a34ce652380a3bd7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10dd2d59a45cdf85d4c41ce2b3bc2b0a1e9887b33d1b04c9a8302e55c36d5662e8d65d325f9bf227c609fe2388e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h126425fca7c6a97977a216dcb0b4fb998c8200088321b3f5dd460856bab09f6c00a89f011717f682687d27716c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2cff4dfec49919ab5b07141f7a989e3b2585fcf070cf13437bfdc429afae83a36cb6e69afb8cc4445a141a83ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e086dba48e6d07f25afecd57beb13fe58a0223a4b77ced8eea1f1f56de9533c7068755f70af5aa698fc123365;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha1bcedd205b3c5cd92890e0222082a759f911fbb80273023e771709685ce8d27a843f618f7878b3dc73f8b41e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e22b79480f9d638e4a95296c8f674e2820a2d08c3f59194ed27ecaa5c35e626a7ed58c476ca2d888b9d6d6b8a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c272945d64f22ec02321124381627fc3c824e626784829bd6a9a2af9ac1149bb169797178540618b343a677b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ca1dcde09e2da100dad0667c044d781b887e68521b24529c2b513acb52a1dc21a78a943e0010a4e1738adccdb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h180a9332cff00e2f6f89d916e4915a0d36e17a71bf81f4d74721319c91bfcb9e86f59d34b7838f389a02cdf9d48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161e8866dfd8dda237e8dd00acd50c80ac40d8ce44c378cc72edf032a6b568110413f9656f0a8e6a29eae383343;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e5b20d52a9b859aa69cafba82697478fa2b8fefc680e3863331eadebb88964958d220a80960b1b006c5ef79c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8dfb324f18f63ce3ecea5cf868f347986416e9148e3dd7ee0d3c2b7ac437fb2b0b1ebb5f7a16ffaab7f6b4e7bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a6113fd5a9b0f1287ef1c87fbe533c563caf32bd536ac7f60a0950beae9b319635682348cd023d24a963d0375;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc7604338964e588b540b00541d3a03ad2bfb5e22695821a6bd9f558ad062762c594fdfab61e3bd172f657c7f5a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd930b8477c7c98c4f30da912b8a1e1fab889e41e6fddd6d7f34a943ff8cdaf4a3017f4c3dc1de74f6c18e480b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f4dd59363820a2596008579a4251f685767d60f1402f2640f6aa824271e941fb435a645bd17d37ed2b5bd646d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a0ec25cd0264b543954878484865a07020e5f908a7b5416d99fb00ad87a8e4d0858b15c1579fdfbf1c642b976;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbeff7ef612cbfcc7b934d6b73f51f012785a571b3452847911e0a400dcf2f455448cf2f6d5376fc85abf5f6896;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a587109566d2b134d230f2326b02e9ea2ac2245d3bf270d133f077bcc038de967d697d1e58ddfdbbc0c0ab3b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce226e049d5152f72a737b67bcd9caa51262d8e887d47856860ef7d759c9d18c6bafbf9aac0adf330c06cbafb3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b83fd9767a508f2ab7f8c48b5ea74a28ed29e19e306497cc430920d1a735a3b16d05d8bf3ecf357251604a05e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41d463519b341cbdeb5bd9c85735e91793bed3cf772e7d11f21eced3d6158dd197a6b7c44d3270dfb60e0b8cbc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb74e06fb59b9a9db63408db30ee2bdfaca80b4c84dbfe101862044a22b2624906aae858abd1a58bd3265da7e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a5ec898eafbc3526ac06486cc3e2236245c9e4bbcd32134437ff4ef551019c7053df97c612726ed6738821076;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14403c43a2a357a235a53a437589af7abdc7405f49942e2d49ae52bd861a67ba58abf889d7d841edb8dcf168c65;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43c014925c46c50d2191c02c3ec3b3667ba93adceb66d82e62b92eb4af00eae3e5d61f9a6f866f8aaa0c64de2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13061a85946e0b91032ad3edffe796ae29b802a89763ee12d507e196f44a24e928dc2966bc97e1019808e23cf2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15776dfccd6436ea793d63c6f2bed426b2a469e8a9336e9840c4601c07270b47b6604d07c7d861a02097caf8115;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h151229a1765296ed32bd26e61b41285ccb8f01f4b309d0f8cc27295aeae824b553a0da39e6adb4156830d3aeb5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d85ee926d34e0187ddb03f4eb22a611164d88d82328d71053b03a4a7232b398d6c167a23555ace1083a7815e85;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha62e6210d0d79bb216e5b8b84f26836925457ea0af1b983f19934f7db8bd80d1621669864bd3ec8e32ddd3fda;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f847ad33df7920e2e98dd055f4a8ddb1be86a73a6392087b9d54aaa40ae9dc85669900300580b61b73eea47fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h120998fa93e5ac1e3cb6857c6de5ba4b644b553a16bcff269ae6e748469f56a03e65dcaf27f2d7ebc6f1ea4f2e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b34c150c1acac60ba1ad15ba5822db56ce48d7b2d22bf219d25585cb44ccee71bee33f58a8a9ddc7c8d7dc33;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h291a326cfb1d07ef69541110dfcc777b64e881de94dcd1ebd08dacd8e2608ef8846f25591e9f2c0206f3f4861a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee8e927101d02730e3dcd822abc6c15fa56f097a08e74edc25d1d88f1c732252645ee0360f47ca3c6b04b06f3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118b6b61fa19ed700a76e76a4c3ffb2e07455a1d8b74ba5ed0b8aa4a0e28fb987e58b303475841b50862645e9d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e73f33ae220e55132394cd22b819c4b82ebf80c0d2bf2790559f319938d3f4770174f51be7d29e4938d00d328;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf9cd274b13a79de03b79f87a719e30c6cc14487d1c212f3ccba9d4fc1318061d6a1cbe6054193b67ea70c1718;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha407f1dcb8d965f799cf466d861754dff8a7cf7af300844effd9505b6f98d4daa8b7c1a2a3780b3e19328f5af9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f244491cf449fa334628b7590449dd9a96de4f6c3d06f041a1bf3180cf8c8fcf89eb8d2fece2aea7dab8680de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd9d61eb01f93d00547c23c3215f9f67521bd122967e93188324a1731cafb01897db519ddbed15b96898ae5842;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178c2f75e856102347e05560718a198afe3de30624101c11c8d2a4a693e577c9a2398e351e460e60aa259fde52;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f3c1cc60017d9fd5c0f4c9496e3236fd3f0a00f48999a63bb470f65c5a1532855688fc2b0439d717ec8746e07;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1006189c6ce3b1ec0788d2b4033ea3577672b7aab80c12d8ef4c91669bebf5108fca846ed79e757fe76b5e23f49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a08f9fa20c2bf11b96dc1f98af65b8626707b97387baa7d02e812e2d9d0d36f918964466d4429a74d7e912ed4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6765556deb9f6562960b8073a73bf5cdfa6dbbc6c0aecddd2ba8ecbf71755edf39618cbc948837c53fe5c3c6c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c39447a6e51115aa0125ff38a9a805a16483cbf7ba0ef0e62ddde4b2b62327f77106426aaa8db51e22e5a5b65;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he821371c36f0757fc2216392eb33608c607ddb5d3e79bf3785d5849a368bb04f2f6194da4d2e3ece6c81354ebd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h144cf9ea79b66dfe545583f2532dde7ee3bea5a60edea65e5d62ee45d73e58d53da31a9386b19d5a377bbf4bb57;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10bbc7be5c89d27acf911dabecfc9b009048dfe5a5ecf2404fa7e183f3c7885d6b9bce1886bbfbef546525f441b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9bbaf9d5b96117bc5e001522f897d9a3efb30c9260ac09c86c615422ff289ab04ddeb2d6e0129fbf27bf9ed606;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d37d29647f3f560967cfa3dffdfc151b03bfb36ce5e3e3415281ab3da8649ba9085e870a0dd4955297f8495a5a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36f6c7e99a54ee8e5eb77a4d6e52e4249242ce5ac60c6a82f180008c9e86426f163e260724f18e1b0d25fa75be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9bb0bea9c77ee7ffa340e3892000bb86c39385812d70cf194c6887e17fb34510bef143aaf754310fd8b9a4a581;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h999212f4d923b003cd6936cacdbd52f46ada7c73d96a970a08986469249203910859cff18ee29a94e0d6762ef9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca497a3fe28751dd92700664884f99410040079b75c8573a4848ac5fb40da4c6960c30e66a8703036e52a91cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d7b6a35415a11904e5e5e86a4b7b58245a80aaa4a726db4a464a31896082e0044474316f74a107b2fc8b953dc1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcfb7b627b1133dd375ab78cf20cda77268c38d505a655d91dc76b77217acfea3c2c74011ff3087ab56bfc0f617;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5fd3e79828ae6fd8cd1061b1ddf1d60a790868fd35aa8bca461476ba454fe4c57f08ae97cbeeb5526b82cb02f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8869857541635ce7b6eb402c7d1674d68cd6a3fe8b2a5efb258fb0d77871a57509ab63b20ffe679765d201e393;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107727a98b06731b6c2994909cc6ee3894095479a85e6c71ef511c7da5074bee0e4eb0e83647154c5d71efa96a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116eb1fae8a43faa5b7dab518cd987aaf7e859406fbd27edc7ad555df6baada9686f072714b89f623fa8dec70a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5809ef4a9ecc864bb155e1d509c341bbbc18eb5648ad0858d6a674b7393f4531c833aa885163d52023acd10fdb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1968e4a0ab0a94e94c7141969b50758a514880a5bcc5c17c2f898c56fb6920dfec3e234a3cabd16e33057eb5bd0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e3d0ae5047233af72f634c49230fcd1cc195f5f6567884e8d800c0bd95c042202ad61830f2a2c72107b9a4b66;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h176076afbdcb433473d352813b231e9acad64e073e6e3b4f0297c9ee5dd437b55ab27a514a9e24e7813513e6cf6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89ee3911c739518fe2c7af5c4ee1be4e292a49eda45d8f21a91354b8699f213d632a5a722698075bb6cf22e2eb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h52fe17212c0569f4c986c393d1239cf9c4d80b967abcbbb4f319198746dab0d363d119cde8aa268b5d6b252316;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9168320fd4b19f88d1d2acc01dffa689c9be78f64f5e929729f83144a745c4dd8fa3f778d63d5af71099abf099;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d16bbb91227586ed31be0f34adfcb6857e49838bfe4cb13ac2978e97b9f7e91789976b7725f39be878c283c86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f21ae183e5b43e723323ef20fc801dbbe9c523cdb1d3117738ea7b6b579bf1d11abeda58a21d59d3fb54aa28c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0557422c604b94a66bfb666e2a3a534ff43ddb4f432db68e4e82a599b807b50d9e187ab35c8f129bc7a965733;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11472b86b9ae055dfa6dcd180f156d16dfde597bf1d7f4263833aae218e6aab338117a01211b67f6d97d807c1c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1878c28b113ff6b6dc3022d574dee83ad8a82741b40eb1f85239058429f11c1927206857b3e0a6e6493c6fdf9bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75555534906120c7722b75a12a9cff7b64bfda24d98cfdf41aa06284c0f0fd6df7f78cae041421ce081a328143;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170fcac75db1fda1fadd9e07efa20eb089aca747d98204baab0f074d574378636a0240e25b080beb4a2c56bac69;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h183701d34a1c467defdc836282b3257a4968eb96ea00fbddb4495d9d0099ae3e4f66340ed9f45651e6788feeaf9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf873994d1309f5b84c189e67556ec2be43d4c193c25582bf65fc6241bda5e570b0c0f83390ff9dbf69bf33ae8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0fdee4d6d67707bebc3c8a58ecf5d41a167f16c54314453e7231580b8c52186a5309de78f2c405de0dcd5f855;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191044989d90841ace7be83228a720cd6842b94c5be2eb8a0eeeeeeec4573e4d9cbb551daa28e696231398a768b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116f95a6db5cce36039ac406dd1cb374ff302178516a7dc5ec12671dc7d9253bad7ad10ef5ddf89b117ec162a26;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h563dc7b7ecc55bf903e1dda23902b25ed2cae9a162e151eadd5806a7b957b01247f387d4f764d66b2acaae2679;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11554e613aace511df1d4ed86101cf7e41ec3b8296ff74229466ee5dcce4618c66fedf2e43f51f92733117e8fd8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4c588e6ed1a24039b125190767d85f14e17ffb0ab6c0e532aa1342290fd61277674b0639a9a881079e9bae439;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b56480eb039620bc238d61cbba2ec83ab1e535095d6e64fc1a10296b1bbe6754504c80e0341cc81a90af8c3544;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147ca1949044fdb0f78d4b041ebe359c77e77a0ae4fe50f277fe334e6e3a910a5cb0197b6b82aad3a2214f7a3a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he64ce3488a093e6d16878755c2ccb374fe1f49295ed025011270871b1fcf46df8eb47f4fbce662a580c711c7dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67ae1d8d2a35d79ed73237565218d5a1e765c8dbfcbc40784c8f1cc756cd65a540c5ec2c50deeb76e81537239c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h904fd27d1b55723e9d51f300911bc5f7e02a01c1a36def72b79d2d1200a9180bb53b4494213ddc4f17bb862fe1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121de12981c7a4f42aab33d641c5207db847ec27176e5d9efd8cce001bcc0c840d009eae78f59fc7bf5f7cdff49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62ac51010149d43eeb2aff7be5f7f3a7fad9d2d47bbe3e5600e0b48dd620d100c4f9cc868f6ad7575b8a6cad60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h765fd11d8a4baaacc12d38d18a0017feeb4ffa772029d63d7fd6e2f7fa439487d6280a211e00f0698a24e780c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41a21254265726275cd32f290eaa44aacf98c2f8f71af17221518081d35a8efaa195a9652879ffe5b95d58136e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h109f9a42b097696613a673c1018f14d268cee830804d4cc35a187e66a221510628c5aae5ab77d8da407c37ef6b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f4603b92aea53ad301e65538256abd0e9accf896f92df8078665086fa703e3facd1d7cb8aa0d7263b715ae976;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1845154cb051746febb62e0c6b3d50c2695f7d436c41f6f1694e3bcd8acdc6352ad85bf79507ae8e0a3c46d9d9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15951182d918ec38c58cbec06aada156b0f6c993f7c8b0eb99b3d06cc1c5632ae206513ccbb878ce0f60267d24d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ce08dd147ffd9cfe134b348e7dd0bc1f33ac01a72bf6b39fe2ae57ea4fa7a597c0e746174a54ccb25b934dff6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a147b3fef4ea07bc4df4906795846e6ab6d7825dae4ac385b45ebd0ef5bed39571ff0ac20eae13dfc56dc9147e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc31d6b8f9a2530d48fc9643f11d250add7d058e8604549d1286f784f35441521c6e9b17ae14847c7ee4296c09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9610bc5b50e8f344bfce6e7ae7c3164bbb2d0b2a7114091d313eec6df059f21aaec21065bf603187f14aa56be6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc338366ab3afe02463ca17092805d98d7b881a8a3050115f32ae9519b6f02e0823e6060393c07af89467e29c08;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3f2dbced97368256418602ce2dcedf60c595bf74ec868177667e091475e347be756797839a255332a47c279df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4091a00ac270bae56ceec2c2762c08e62ecd670fe86a9408114b4a7db53f9aa47ed4f1871020398a6f31359fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12f91be0d7326c8f2670a29a8f66c4fdf1b36f36b61af4a4a76474f9f2df02bf1fb36b5d58cbbcbed5645960764;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f85d7b873c9ec68379ddbf98f79b5420d8b39a17a0a08762d9cd8342fc522f1a2e37ce37a3cb2c57d17287a7ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1054d5e5984d8078f09b885768dd7b0af857d18d6016a6e645c7a921fdad2ce73098dc0a34c24f5d95ab79ede68;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136db0dbefaf01f261819fffc3baee642e3e46009f11827a050bd8f0bdd75bf5424d9aff72632295bbd0caabba8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170fffc3515ef368db3e54c4df3de19bd7ee0422d4ce67308632f4d6f2e3482a148f83a3992058af158199f260b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3344012499974fa57784474eb6df998f660161e6d7932b768526ec948a8b177ddbc670733e83ff1158122cd44;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h790a219fb77e892aa491bcd10bef59df7dea6f411f756bca37f71491852f741ffaf73c0b8db63bb3a5a53a0aba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h848592fc579ebdc1becad96ccaa45b3760a7953cc87bb57bdf923f9d563682a283f47c6dd405eea4725a5a6abc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f62cb5c6fc14ec46bc62b2ee48f7b776af2f481873f9e8f61628d4019b87e34a2d3b0d3840ac678670a680811a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125ab5bc7b26202bf1d164daa87a20ddd73ca0f143c11d56e9173e9b443c40793144e91fdba0d010260d03edeb3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11115e5188acab8daf298ed7de2aa58cbbf36c902e311fdde2a5c84025829e02a13051127c3ee173b8102f82baf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15977a60f29c07cec70d5ffc87e247313f4e8c812bfb874866b53a2e517c78d77af5e09e6dc7d4133d7a0aea2a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125c5547b4731b5409974bcf6a298feb4a249d57800d470c4f11d261cb446516e85da08d4c42102e338cae64d09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e1a70e1317af9ccd23328c21723120c0a567849000b08cc6afadace3da38c8d756eefae110fdd060c637d44aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb1a3ad62da6eeaf93b9175056cab69b6b8cc18f0246ba7dd5fae147f945efd7e31a96ede6e0b7d8b0e3e6e8ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b37feba666332aa7d6c774907ff03262c9c9e25f31d76267f40432544d0881f519e5de6de58f8edd005ad5e1d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7455d7e7891756238f94c7195a93f1ce8d0e3c58add0b44747bf48b2038a8664f2644146581c2baace8546dfc7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he6ffb2c53680df8ef8a568cf0921dc81aeede818c261cf0ce02a2df6324e78f9e9bd1988b89135d6bbaae62e19;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1761f6633566f551a8861e557c2a756f2d9e53913a01967fb70a5dd32ff69ad778cbcfe0fce6e689ae77e475139;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haaaa8a8b3feac9815c7ff6d474942f2df66b0c0a6f338dae3f5c77e9ebbceb3ebfb2d40e396be4f48362f9963e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1548ae4971d445143660131c52dbcc79cb46779806b1b48e35f6c8d3d90ec652f2d182467cb52d21c5e062d72f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1640814361398ef8cc57bb25b65ec17c059b6aa1ee091940fa6c3a1db7ec8170ded040bfbe96c3c2e5df93d74d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a051296e65a53e6f2be374a8d667f95f5e6e40ca071d1f53338a24b708ae1408f46bb126918e76fa6b659a710;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1faa7462a313d9a0477af769a3209fe73255a266daedde91ec10b83c154df427ee9867e57151b17bf3731a01949;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cffd17ae24c42b7decb8c6b6f6b8dc643824a19771d15b0e36866776db4fd5e2b0a7d7c5e058e789389562db20;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8ea8aaf996320540cce783f8d7edbd36444cbe610f765cab521df408e6cc886a7965eccc4faefddc373ced230;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a3ce8b23f15b6b1deea5a6525ac1669a6674e6d5ce41a7a807358ad0774e2588f7cb3b73e079364adb81d86f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0b297e9c0d55ea36dace2ac9cf6688d2e83984fbbf31408e5102c96c24165adf9db2dfb3085f33253906c0866;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he72d40490c7e943b3be9bd23314c1dbcaca3d57463d20b9450b10e0badb73920e3f2a2e49eac7e06aa3b1ad627;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103ea05dd95361d9e587f51b48b9c6e5c0176783272233a5cf72ed9d5d37530f8075878938b3380220a03a9cb9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a68d167efff809846f56c453f77f58b86e3aa14ee99e646a0d084af47b18cf6628bc587973930963fcf3cb11b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41e8908f4e2e9e55aa757a24c4e30f4c2673f4115b20c3abe25670e4778cef47b7bbfb76bfed576ab880bfc966;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1988bf65321ed98f04f427cf04901ed3c648ab8e6907be90e8a16f8e4a056e072b2b2c112945cb43c32bdbf6e44;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63035a6aa1a988b5130af2936656a8acab4fc0b08a372b540bedf7a8880d399e3e9e79c11a28488bea5b7a8804;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9b119fd683066546c230871d567f53dee7ca7c1313f6e91266d23ea70d4adf2ab72bccbff1d1ee78426d3807e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7707e27a3427bfbe1e29672f05a265a8a5e071ab8eae01840249702647d020463d816809e5d6ff40490e9d73af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab46c0bea509ed341ff025abceb19f03c6aab8c9a037c0f35926796c04e4e8e2aaaa2b94cca880c8d263081c6f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19bc2c46a6546d9e33181f45c4da3950693bd92752600a2bdcae79d42b35eef3dbb8fa13ad30f4cc5ce118dabbd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155a9eb7878fef0bc1b665be56258643dfc9a3a8860ce64d0f89666fbb5b0db8bde46e4cea7a13a8cce10588c7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd789ab66979d35eeda4471c19d96d870de242403ce4be1bdbddf0f3652558491b58063c2ee1910d0659a79a86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec27de2871ecd6bbc035852bf4f416016125f8520c7d63a46d97f50cf263577faec17635bc5c960931ec9e6e70;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf57a9ce04698295e377f513f76184a78bc3548fb9a6444f71a22a683d3283597c1f6f4f35e6b9fd48218bce5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5520bdd6128348bed12142e6066d685cebb702f771c97c28e77a6f41bf88d26ee604e484316b6e96aa8fa10383;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76a127d6d0d041b1ef34c7989b9c0443d6be297f6a6c5cb44eb6728fc2c2f8eebb894e1a6ba74d742208d51790;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b622753a10befd34545f731ab16b701b0fa0cff9d695ca1a4934821e854710fa1fdbb7981497b2625879be2f92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df9de8d852fff5440ce267dc2c4912a1780d1377c55100425e539650b4f49cd77de3f0182352adb10ed116cd7f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd49cf44a026d15d80e197eb24a8da7fe8a54878dd7b7894bf90ecd556e3ae1a801ed022b8f083c3a0339e58195;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb9988684ab5d88166de25f2e04a4153452ca4b3979675787453dcc0236a0e50a58c8e886a59fdc9921c373da00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he727d6e74b880095321994fca05a26dd88b723f7ab9745f2b1ed8ff36b912209eba143444da29e981a37d558f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b5eec475e50fab2a65711679b41cf10d4dafc4caf923b4e09f7f7d5b3d7247d08db6720e1b91b6fd612b43bde1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4045d04a0108a30ca6711dea1e8bf721c58b28688a846d2062e622015af48f2fd027aa35ed11fc90e81790d292;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136a0eb5f558a6b1e4381bf1cd6ca7210171d4e2a066da9754c9e6f0dc25bc0fd83d62de1fdf33a901503b3806;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5dc01840db6265475a18cea599d6d3681f74bc1b478224236629e358b9ada9f7fade2f6d4e8127846fa74b75cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bb526d3b7ffa5e7efefe2768a9fa8499eba8b06e0710e23683fb9a5df55bddf2b37035c49949f8e1edb6466c0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2473255f7b1d021a6bb1dbfa4d0b9c51550c2eb87dab856eb679c074953eb3bca4eb2e417456c00c8e8e892bdf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3035c02782048922a6adc97aeda99eb4a0ba8e861ae544e349c70345cb1ad3094d4cd6d615555d6aec7f14c79e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189799c633d7e86b3730f47d0a45831e0932a742a246922c3f65e346ac5d136bbb3d4998eec6c02ff08d14832da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h101e659db102b3ac4f723f4fcb45300c630e9ef77a88ecbd71d4c774d2ee02b0fc1181bd0ef16e4234584748b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3797ad31991da58c3b7821a9e9d04b435e66337c27781cf158b698b014c5da2bd5c38aef3b58b1a40be0850e66;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff5fce7f671485026d7143df19ad7aa8254d324bde4c9bed573a2550678eaefb598efbb8a66539c53eab8a4917;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab2e17bac41f9a045c4d45370a01652043bdc74b863ded81ec78dbb735e3eb9c5e8af048ec7219a91314b3ac6f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88314fc3749d290cd7a2d4f83067f244067bff3f11eedafe3c501656088eb330725d5a5d30065aba0405140496;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ef24aaecadcbef42a22c52917c7e703afe8926894012ba2a5807b84fdf8bf50eb98d95819e024e6d57cf69728;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h657389045ee7d4d6cebeb769bab440bc8a3060661edcfc36f39f40b36606a7d931868f530e12a1fead2fc35a6a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51ee41535a896086f6ad8062e271e012c99e7f627e9da22660e1d1f4a6a970e01ec8476046ce815c27407e441;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc57d7a78c1997391fbaaceeda2de6cb7181853f6115e8d0fb2b9f4740774011234346082d2d235af8e25286a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cab0b17b96ade7b377d574aa50be9bf51755a4f00ad1b81786f94781160ce10e6a07bde745e9533be6430c6aa3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha573da03511ffa09a1b92750e21c8fd3e2c0a80a709a1fd4ecc8eea60103276cb1647998c5794aef82b0e45cec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a776b10f3dac9f6222893abe36b37de4e661124fcef88e4f105b434156729557c7ae4cfa6663d8d62937a3ffc4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa2387654018b60bfa216488ed60934416bf01f5d141d683ff7fe5cc823a96929df54d8fe643c44ae6d380cc61;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h243569e1aed6d5d4d722d3695fdc6745c96a8d60f2105460c2935517fa625dcb7c907baccb84737b666dc2525a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab0ed1609a68891444c3587b1c1cd999595adac32a1ad7966f2fb824c2edd0e97c2786aa9472d17ce65b7b5b4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ec36269a0375553564716218926e4d467a7d250e766ca2d9bd2e543b5b157ecf2e1feaf61fafdfb207a8ff51c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13adb0b68c2960d707013c03efe550279e8d10324baa10126bd5058b3ceb5a8f94e3dee2387c04d5ccb834a4144;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67a2e8b40a6138cdec42571515175ff268bab250f0bc026239ff0ed873aac12cc12309ef33e92fa0e59cf4e0a8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104e0f909fb39d318816a9591d1f2f8a60f53b32f8fc842f0251842ed90b5f5c2713422a88b92e8b6805e05f993;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d94140d04fcb0e06d382232cdfa2c062a9a7590098196bc7732eede7cbf4651bc5ac9e956f0d1ec68ea0eae4c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9116b7b6451b5f218583b1cb341d9df1b919d03252c0836b08269331c9fea80a01096433006cd45f7f2036e39b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a44586a93ade0657823c9f9b527ef7b64834258aaac84e58921acc0865b66559c780206407eb5d5b3fdab84ab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab202224e645def61078ecb0e9c82b223ebfb7958be05ab4d9000b759e11d0c0a4dbf84303a86774d1295583a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1d86c3ed9b5c91680782d78c081f6c6596168b4f8a694584b77b00c97b35b5fb9fce768d90eec8bb77253cb80;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f2498199cbcbf0f1d258394376e391acd116d57cd656a6ebf80a2d4f8957e3c76c0bd4428806ac01754cb33d7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1e75e6b045c13f3416806d9d5830d5776a7f168cde2f088e3eec3140766b171c587946218d731e3b862ef6ba8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10bc8327169c961e0096a9e5b34e8111d52955c05b7332368540889930ee41adf86681b8cc4788393099695de39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3dea8d9f2fad4271963775a509fc088afd3208ec95c688b63fd5c2dbfe0a8879fc92d6097c710579c2aedd0128;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8149039357cea90827f836ccd4fdaa2de1553cba7315aae15dd5dfa6e8dcf110a90454b2dcf1dc4eb051c90a56;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b97307c39d2a784846290cd2a982dc36f0a254a10d22441f87deb816947f9fa8f29bf1df80a8d9c843a451393c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c763354634f2d258b871c4759244605fa690e2d560ecf870052f168239b7c162c7ea8407a82c6309f39b42b203;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191a3c396ba4d0190fec197b57da02a1b9c1625f7c2af69140b4dc34ffe67c76d3dcf19d22fa0e1a3d5c1178c9e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h31fb5ce34f76f257d2b8e42c474f4fc1dd2cb380597454b0b8fe2100ada1482bd4393bbd0d487e13d0832ba357;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h144e95e1c7433fd7061815a47062dc5025745601b9a14ab653a59693b5e4b2bf8278368bcd1174c91dcbc3f4026;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43245a6526f9502a94f1a63f8ac3f091f4c4dabca37b7c830a4780b50364cfa5500c2b141626730b055918ccda;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1adf64222b2ef6bb58fe569e5fea2d2ed3a6500db6fb8a6077604b3aff444546ae62ef2e7b7dbea1a60aa3f928e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dca4a51a21fdbafa93625d85352062e75fe16e6fdb38ae8381a506d48065572131abb59fadd613a405661f0ab4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7f786222065415f3ef09f4e964624d9122e3f4392f686ebb2262ada8f30c199c6dbb9e1359718613fa72ecbeb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164979191b80624f022c771a5d01934fdb2e908e6efd18c165fbd5ff934ac2b975a2d1c100838d966b9c668311b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6a050cdc5e0a5126377fdf1b82b503a8b20094329bd34306edb586a916fb9804da8967bf26f1b3da0afdd76a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134df9c536f61494594af7c638d670ea5f21b0959f2f26ca5d090a4910b10991837d8aafbb267ac5d179eb9eb29;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66ec50ce6bdf6d945b353b561e1d654c5448fe1694d6bf1d6f3f8fb44281d1f93e5515e9ebd0f17be165cd0453;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98381ff0ce5d1635cc986df821eadfde49843e434c13226e92d7cbf6ea24bdfad67ce36981f36af7ea29aafc0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h629fbec41790b1d8f91cfc9b1f1086572ed0d4acf3c8e002a4491e2e6f856fd384d213493a30df514f7407a1ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f66177743dbe43d7eaad8b07c74971c080a29fb1ca9cf24a83726216730ab9085161d14dff6fdbc438c7aa5411;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fd1714396873431c9df90211978a10a6a77bc2c41b48608120609c62d7274bde658a881ae89c34181277b05b1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19be8d123f7e94023a9f5a927d942abff9b1de91e0bb0ae6b1b2b26983250168fa608b4d1c3ee28fa8655ca0b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6eead986129c061dceb38cfb998a5dc6ec287ad1f92d2930f5cad879bda6f6cc4f793723a9694b8843d62daf16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41a64c45eed339cf494de76d3c2591cf49bc8db222c75e323b77151749de547bbdffb5704cbd8405cefa17001b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c04126e6318c016b0f71d8faa9935976ce14ea7a9d50027d7088f7428a45bfe61612f5b72c940e7c7ba337172;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12bc397f835eaaa7f2fd3cb8259c5563d3a9007f228b80b0df28f55d9a63d9506cbc99cd3512421aea1ca6881fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10af7cfe545a555634fb6354c3e967b909dffb240001189e32c6cbe19c957b81a75f49b05596a69363010649400;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1425b04ef439c7d1d7b9734cff0165d66cf9705ddfb114744252a19d96d107b93e01b6a7dd3f8ed93d4645d6d06;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h502e1178bb5e968bbd441f318f9bd402b2223e1fcb0a319cda9cf6f5baa8c5bf42ea4e106e516a6503d6e030ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ed7f829caa7362e49c80c15fc1869ea80b66572a7363cb39268bbc9f783322f52bf0b7dc0c113abf4d0e8e46f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34b7d9e6c5c977845e28d63448010abc7407cbfd65d5dea24bdfa91e03978addb2655f995e2263f132c5ef5b4c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb0523a32449234ef7320d0f57585019ffae796c7593afbb22f65ea2bf9f0358308b355c1ad6b972dc96bfd4d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b7ec35f35615fc426d5d4a7efb78892c32012f0cff4a8d34898730634a6ef52a909b5a9706fea6cc7adf57631;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17aff4d5f386004466892e4dac08bc99fd2bd59354eb8eac3381c21a5ab26ca0c0dd511a41b127d6dc29f9949dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a97463a5a2e4f0ef7a0f8461770c1742add8c32ce172096da6eb96550c7334255f1f80da3543fdc6d4a4e095f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d3474a96eec53bc88643dec42081823aab4fbcb2751b8f6a47ceedc4cf96be922ca9c6e8b56d61da95763c126;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8c346347001d94636807c9c454c72a83ab381e6d13b8b003959bd698014ac0c649c7b1fe35b3fe0205d88ce53;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d2b5c344e1ee2d74295eaa2d2cc370042ffd7cda798d8f3c365b29285d4fa976b384602ad2e7f6b8a068fe321;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104bd1731cab7e11b8552c04a11b01dca93729915201ef2dddbc73475a699270ac1e6d7078d8e001d77b5f11ec4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb01c7a8aea83ad98c961757bd3777c346088e770acfd3d260816fbd943269a95b73f047f78cdfe381df7bd4ba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a735147679bd861af9aeb49e1ba638eab6e758703857aec19afe74d20ddc2e04cb1878d792d3f628ef6dc12641;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124dc8bed2848e2fc8d788022ece425e1c84a3571c29ae66b84422685f4eba80777074b373670b2887d9e531b87;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af6e732bbe5c42713c486b24e055c4775eb5f7b349d5c8a6defc3b0d11088ec02c208cac09f105b981759b6f35;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1623818b39095d39ba380d2852670252c81746cc22780f04aa27ae221fa3b1eabcf98b2b668bed449fbfcb01a78;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd5fcb690998366facd48d7438480a43d9657aaa21848652be6adce011a6fde7a59efe03bc2e0d9b5a9637b248e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e52a1a75b49a96564f54baed9456caa725570a43141c31136a6635c0f387aae48f2e3a3fa044ca051b841dbb50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9cb04d5161aea57945fc1fa4f6693fb24c40d3efab2cce9eaa643d45b1831a7b9e26a25836331b51a02b9c3373;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha82611c45c7a87dd47aed63f383b90562e6290080aaebe2fa32364ad21923816e7fcd22a082e212ba1bd8cc59f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14accdaad0c33fda06da556d250518f146233693c14e995a3104179d568a7679121823a33b76c274be4fd1b4d92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h102881e3329b716aae2a46d44c032b78df27aeaaac78f22802dc4510f59ff67d25e2c6e9664d2fc02b86db02ecf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ead2e98d2e0c646d534c65509d4da9eacc7217ee90a0e0759b0e5f31b6726f88e861323478a24a4422c4be0cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0cbdfa55dd3ddf7d6d38e02a238fce785bba78228d53e533d79b5595f6e561a0654ea1a7aa41cdd473e6d5862;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26224b087fa78134da809c4127828033bd1e51d9397e265ddcaab3a5ce0dfeaecdfd19f8aff858f1a7be82230c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a4c79be310b4ce631ed364f0ef41ffb974cc52ed8185973d8b9d6c3b8b10cd69996fc211e0885151bbe5e948f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182d372a5f89e268f774d0a6ee5f7325825c6b5e11cd94c9ccd9d3934fc187f022e12eacc9b2882e9f0f503cdc9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90fcb345552a87597d6000463f35d20e825ffb523e6febb2791d8168582a427aa16f260dcf36ba51e0ee908d09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5bfba9f72098f6cd7941e3953b94d6ed040bc76c3efc4eb52c4653429406efcab332b60058c6d875242d5eb1b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e682f0b3c535cdb475dc212f9e0f888dc0f794b590175e4e870e6b1029c8954e90d561808a8a7ce6b10fdc788;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h750f86dc040be6310bc26735881ffd8d86a3ee54f4fbec040f594591c8fa1105a2252b87a7d3e850ba2a1519b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb70efeeced26f58e7e3791afe686b0b019a7d24596f671f2477606c26f3918a9467b5e65541c0bf39332ecaf50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca480150036bc1955b3154e2abf0d8d61847ac892e038d5c7ef446c2cf3f53630964525e1d27d0bc509d61c759;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e43abc068a6c9e03fd98bc930669a137d2a3ad9bf5385979fd4fe12fe0105cc3d086e9358f3c11f8fb7c9fce8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6d336901f6be9aed2619bc901dc1ce0270800074ca62092b454d5469e3584fd3bbcf3f2e0f2974154386783b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60859f51c55450674c9d6f3b2920ebe449c15aac69bdbf8c80acafa2435fdbf9ae36486f8aaf2668885d972a98;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h299388a5d07dd909dd8eb8e027926acf2b06f75194a4aa531ed8b701f80e365fce3b2668abee8d52b19d4d2980;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d065975b171cbb6b180d882efa1a9f793112638d080f9dd74f892b302d33671dae5ee19f0a01650e8cbeae107d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191788821172ddd34d635a8b1e941c9e9b095713e7d93a7a333a616a0d0d6d6330bc67bd421b70061530db7388a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122db38511611d80ec3b71d7d9aeca205f97607f8a2fcfc261b449645e521deedc2e67863d0c044fbc1bf2d4fda;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f93cb599954b7438a1987a2325ddd8f1bf784dc3fc54707f0561fd394cfe5ddd8d6fa67aa64bae5094cd0b20ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be9e98e6e8498e92b6cf123f0b8882cb7641776401e71d4577335cc9ac67a54a26ec0748bbcb4b8cc86bf6f78f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd33d71bd5f70f1f2be676bcdf1c90d51aa29fb7b709cf11071ac79c17642c77ac4aa36f2b6bece05bebc5ba4c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee15b059d08ecd5b6aeecddc121c1cd8287d726324223a627bc0d0ad96cda4348ab05d199d7c7981c337fb3b55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116d389431b0c9c9b7e1756766f9e450109fb4ffad750812e02235e0a477534f21ba37a8c7cbf708b735f92ff52;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64417db96c868774fb8f4d88b54d82cab2190d42a6da528ae0b0d01b3066d964625654589b04179067a7bd7882;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a393ecf2badd8b53d8453db11e005a01fc05226960ea49cd3295d028efaa6b2d2dcaa728ffc700b9bbdfb24b9d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he30d141e8f81db6c29b3b226fec707beaf1b9c661c2c0a41d433dc56ecaadbb07910cde3ed9e25ae559dd09ee6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bba7f79c8005ac9071220255ee8ea71b8e48eab8dbf1d4e07b6b4f1d381783094cc17c1ed9f84e52567c24c989;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d142c49d01a4678b3eb38fa7592e87a1448f88bdaf9b1423326b786c56cbae95495b694d0d724364047276799;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a89b816607723679c0f8fda6d6ae86afb948efff6669d3354ff9885e6f896cdf4593b27d1bd91e48bdd16af30;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8bc5f19cadee129175a8bbc90ca250dce88297e1ea2c9c6e874d085742a0a25e52a33d0d482d795ca5ed181a58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198e77809ee4a19fabdc95816b8f66c5b3d07f9d577403ad31c1e540bfcfc3ab46051d362d004c0e981aa71f5a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d7b10044c5be8951f877db1cc0ec629d287cd15aaf2165ad9b98eaa4da3dd8e4ee8953475e6cb6d0b5ce48d98;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3bb10068f3f5680bf8de2305a031013449dd08fa6cba3294405f7fb64d29a8b06e966c6b95449cfbf4da776f5d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4dc8840de9d0cd6a2fb9236b41fe397b53097388b35e7fcad3422d356427bd08dceefe8a514ee62794ea182eaa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7930a72cae72e05697722afad1760e74aa9471d6c62eba0d2f261e91b8ae8f78f0be779da66ffe407ef9ddba8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58f3df017a3ceebb99804f937433aacd6b4ee8021fe049ab48712bcb5a2f361da5843192416e446c5ee8fb7fb7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1330371aefc4a20a16ce231fbd95681fddb9052345eb4590d54de42fe519ba4c6762cd598692dbd8803ded10349;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef9a23d173961760a380add0b6d864be8eccb4cb84b65121d4ca06021577697a7005b14c847175640d34ef20b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2631dcaafcb5ab1b646a9254b9c357d0f25d91fd725ede713d8583b0ca92dcdd34dcfc349762c2ced2e990933;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89d1815bd11a73b6c5cf653cae0d1f9e05776c2d435db906b02d33f2d3fa48ec7b438048ed5efa0a5821c4b3f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186a6b060b6b820d31ab7a96faaab1a9c0e3e9a15e8965b88033f9888b591de7eb3598a2d82d53e18890df3e5aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8354db647921a3b27ff62ba1d337e2d30be5f6ed75a8b123085758110ecc7ae7edeaee8bf1668d247fd1002e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h210b79ca46fe8033e5065f0a25d54a8c6e7834c86b3ee13c00676b72731a1727946355bc4f0b0c3c6e37aadc19;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf266957d43d3e63457032ea2a3a6c09631148675a379cb893f9d1b083214dcad42f82af24fd2838e0ed624940;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155038a1ccd381de5b6883b707ecdd0f3dd70c024e93d774de1ddb2981946b2a19528862a6f1b5e40642c6a6488;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159938fe5adc8f81d57f8d08aa28937bfdd4c36cb929a4eb31b51dc31e342f142deb465c5aff66fdc92d9b05a2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0019672a26d23b352951f827f277038cba39f55abaa56d68c842f9daa81aa9368d7f37fc4f3b73b2bd07cc138;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163bf9098d21328e785f210eacec35cc6d85114ba257f60731e1a4d7aa3eb9a2981f08e239c2fbfdbc18d6fc9b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3743a9d26ca108eda260d1a4caeafd489a5ad5cceaacb2f471f36b16bcff8cd16f4854fe4ae2ae138c1807cc5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68fb72fb77575ff228d737fd67d460ae808590610ba6d8075c3df1a0b1655ebefb17593bc101deaacd3aa1a6dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c824c58f14d06b256926049f43caea84ffcef25ed64d540fa4455b95b5b1fe977f632708374600c0d8ab64cc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha918c4e64ee0c42eaf3087139db623bdcd89b459d375f430c353d9a62b4507b899ca404f7ac42fa384e64aa84a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c9f5e46a04a9e5c0013b25b30d29f317de596131833152bff388413335f85de51ab9faf51cd151ed91070631b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbff135eaf9f3301a8630df494213d25461c751167d6205516952bd3162060e0fbc6d0eb11b1c3a4afe00299a93;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7f116d0b934b978edc49887ca694bc021144fa0c96a6ce9f7ec6bfac685f4fe4e2dc8e9a05c2946f0981fc0f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c7ae3f7f54c037a407db2ca15731b36b9920c1df45dd8c759f5e99d938c5e17ff187598b7c48ba615f9b350d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1acdda377d693356c6ba492af7ca27988191b74745dba97d0f1efcbb2afe45aeecab3670f8100feaa7c58ee9803;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f08532e11238ee3d1e79bedc8b5ae74d5c2f2176065f8a34f6d5259d83b92156046363f6adf3c2f5f9d59390c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161ebae98926957daf42a505e781ee3870be3cd92a78e7d9d55319386c6cf760425deea1ed8b54efe6d2b0a31ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ba60073da44d4a3a0ed4ac6862bc556e48cc7844691969ec43b0f6b433ddc11eb52116990d109005fb59c9d55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4101f0183ebb137c68f67a74fa8122abfe673addad434e73d2fd383b91a276ebc3fedac12dceef4ccf838e3222;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfff72a9cb9faf183e804b1eb6596294326f481deb99e43182fd066ad9fb88ed5a8b685e05160d92239f3a24bc0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a1550910eb7bae6798a2ce3ae477ed05ed444aa8dc7dd2c001c2f868ddcf6c57b7ad479f0c8c1ba81668aa196;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb02f0c86c4b9ec4971973e5fddac684cd4792052bc41eebeab7098e3246b690adf6cf86fa3150741e3a209ed4b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16aa0c048388ce0b25804e5a90e942b6674ae391ab7c9ba09922b41d6a1cb2977f3b998239fc2ea1dd9d8117da0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160c5932164acd29fbb67be60044a340048b66fe85b4cd2110166ded006bfd18c1ef7009d23a541f874918ad715;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1892bcd255e796ffaa6fb0e6f9a09aa8d2d1ccf24da51ec17c16b7da7c44ea8ac9144b43a7bebdef1c8a072a21d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he961cdca596197745b2c5c3c44fa0c21c7264da993274ef4e19c25c3950ba3bc7dbda8ad03f18a126c3f88cd95;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe8174b36c3b13b3a4bcab5cd09bb2f500642416e05693e63963879d94a0046c6469d3d117078cc5e4112d6d8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h971bb472f79938ffc405a679747e4b0f83efee744c32d86bc09cbf9ce6f219ed7312487aa77a3e3156203ac885;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fdb16078747d015b80dac2fe56b553efcb58237813dba30e2a6a503bbdfc989166158a2389b0c626d1f46a0f8b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b79c4b3ee94b9e03da614d069f8519c21bb522b4204cfbe55c4b9950dd8456e89a000aa38d18be8dd45d41c0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1504ef64d838b1a66befaced6989e0813d4b3f45aa836f8912aa69e8cceffac6dbd160b18e7370578f1fc663898;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d289d083c5417cda65e9432bf9052e7a0c23a1fde8e01f419e701b36b9d8ebd8ebfe7762125b0472381c44f34c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90be7c621bdffc3d4f35db188e27e7c1a99ea81a6012ec77b3bf7c69962b74a2a4e7e5c15c015b59e6a23d03ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54713a6f1452a3d71456eacb3763ee259f7698f618dfbbda24d25057182867dd352aef5f1204961d30a947d6f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16faa4105bbafae2a0e5ca482677da9d7034896d2a5bffc54c986c1eb32c566866c7fcf26b0b9656f49412a5911;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50dc9723c481c7c827fc0fd3cdcfaaa915e8485935a51c68f22859773543e6d1f62ed424418da8f2b47afc7c07;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha646c8501b0360586e74426f589a5dc4590062657846898f313360211626c9f3f106f65779ce1d7ad699f6c433;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ae62dbd332ca5f3ba2c58db345de724f32192b4bb3709f10118f383feda8d227eb298cd971d6cda50d959096d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he28b39684c29541f6cb19388f98eac3543b3a46e5545944dd4a48bc05a992b9c0383e9002901937982378359f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h724bb264e4313519566effc4450a542b78f741f463eb4f9f910aff2cf42b78d362793bb5b6888c8dbfab79d4d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b25527c307f62b462881c13f9c1e835a97e9cd2645b27d1b0dc572339e5aeca2fce4e373783f577af34015ffe8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16413c9ab25cbbd938f8a0ca1700a6ec9c04c958576693e89fe3c32fc5df7c47c31cc326472c965e43f9c5514a2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4a95461b6382fb763e0c0c383a53b6ca91b8be4536056c97cbed37d1654a31887dd86b602feb277546a05af4a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c7e92414dd7d3f65749b3716af82c6fd2db09fbbfb4ff9c2c1ac3ae00c63e1ac0358a464c148b0091c25157c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7effbf157aa9efa87845a93d81ba847482b67572dff0978f1613e66e46c59f1ea19557a6d0049544b70cbbfc74;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce8e447e5bece8652a94ef59a517e95de6bd831da9a71c9ea7f2334fdebda8106a22596dc612b450ee42df8cd2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142afc7dd20dcbba08e5262c09116f610a972e8404e3a8fe4c6c1783772e64770d4cc0588555f5d2b32973787d7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1305d171facf2c80fb136e4b3e2e5530a2a6f4bbadaa95217f7a6177ee9256b0ca9f2e3936ab89eeb92556fdb45;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cac4a8f985d6671efab5ab29156bcf298d863b60db28b8f4e2bae952d984e6735f5d72405279e47dd8f7662b67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e7cba06577eb2936c587fcb260e8a98163e8d49a32389893163c6ff61d5a2521fea53e71217ee2834a4c0974a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h40c0e53248511e31bb119db1eea6f41f85168dbe92a02ab7c40b7aeb5236be4bbbf32c8733dc3d297b80f247e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55975ab1d15402b33bc18b837ab810b4764da65d1c997d901e604cba43e29c09af3fa0667cff23ff1789bb95;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3254fc7c2fb8454a4bcbe45948653b3bbb0fb3e6d00dc631e025764ff594c631799c5cd367e7e477bf14c12c44;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h587958c2891902fc2547b97705310ad0bff372623af5ca36b3889043a8d7c559d6e8495dd06476229a7ec242df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he6f5bdfa77c1213f2b8a32067cc56ac08d817ed1a153c7daaa8692fdec8af98e33974a4050dc47e0f27d4b9762;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf5e6c48d47d336ffa663219179b82f82cc903a16f95c74cf2a15c43e2a8c8ec749eaa6bef4eb7f32a8c34a88f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149053cf3da1b35f57772f41a1e5b60a77febccf0c8fca2e09b8cf1e6189a48e8903385c1a944858fbe2cafb386;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa8a2e70139e700dcd7230a13f53c2a16d75e5c5c572f8df632afe331d3ca77c29e9e32c41d8fa975323bc34eb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bdc3b799abfe4ca32b9c0ccd1f9f332dfbe97b47d799e5b96e39e278fa39aa940f598d9c70d154b83336c4e50d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15318de1fbf4a0d512555bce0a39c162ff7e0b19810e205ebaaae1835f1d161848229ef551e2bd34dc24d3b891b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ef8c059ddefde4f27930529234fefd0bc18b94582bcb33cfb604935cc325a35189cce7f5521342a1801a60e67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134bb8699888450fb2fd9092f040e1eeaf60fa84b7fcda3eb526e80239e50825508ebf6580ca3e4c45182b701c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c795e9241ae9aece40cde6e1a049d7415777a502bf0885ed634340136fa0058b74deaaca65aac7f25c37c8cd6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ebc079dafbdb927068627b11627937b305a7634cd227de0111258f8a110d056b655da14b6668cd3b48ac2dcd1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc5b1e3f3500ea663af028c100e9844c6f7fb61fe7898453dc07e18475785bec7520dd4e7abf98a8c5709bdad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65cb0eab57d302b23f8d9b9c8856e49fae804d818cbeb9cafcfc47a624fb91f6a944d55c49cb23c77a19f8b69;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f3e89099095ca30bfcbca6b57836c56d0299247501d020868ad134c614fedf8593dfb5d790b51e0d2837e161;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67ed830dd2011a12826ad5fd653af51087bc077221b7d191328b01bc95b959261eee38a2957133d0d578c2b8d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1335666510de18b6ed4ec2c45fcb1b44ee64e162baad0f190a34b18f297ed9b32597b99e9a865fd7336f799620c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9862851e632193d9eacd144c86c46c03995881d83897698d14fd11757d965ab9e3a9eb05b0bb786ddd4a895ba6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66c4717eccb794d4616e2e830ec6a4b81be4055c93dcb993f4a9fc59f1494c2c5d71b970082234ad9898f90d8d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b604abf9670420444f9a462ac6934ec99bbedb5661ed0bd9f8dfbcd7dc6b6d00f0be8cc6dde7b2f67525e7befb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128633e4c6338ff35c45fca1c8bc9c6a233509dae33d0da8ff44295c791ea94d942a8981f7fddc52a2b7cdb865f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb1badc92013987b76c94e55f01c6993a554fb9dd3bda1257e174cd82c73adf03202880926e0ee77e27a90a7a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ccdc4284883785baa05b36795b69bfd9be6bd28d754c219971480389d9755564181819cc684ae5ae7b4afdb241;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b88d749276861c12666b8ca72a85d4fa9a0f9ec8357df5da5fdeced58f0c72368327454dcda992f3ddb2997485;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d767af480bfdb95e96bfa0c895b702221f36cb3a1676eb4baac2c4910ea55bed2748b8c27312e81345fc242436;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab4629ddcae28a0cddeab6875b488a2112ec2114cd3ac0a8984dfee205fa0ac983167a710af7f592fa3eecf6ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdc511cec8db3020f3595a3e10f916e3e9395a3b33aca81e90534710bdd58684e63986843cf178de2270221a99f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd423ddb25dcec6736072324f9932512f8edded8dfadb591c77d523aeb9b04c095250f997ecb8f92790e8ec657;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee1b6d2266cd28b70d5961130b5ec3c53f28282318b2ccc9f04a1b066c456a8fb2653b64e464e393ab2a20dad7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf9d925425ec7ad95adca8463b55aa0f538e25ecb0a493b2bad0763ef8879b2cf3122844f673f87e319fa5b97ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e401a733dd1effcfdd3b0f897806b936cc1a3463e703f1b6c6647fef8c3ab4485615e9088242509760c077d69;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h192747455fd7dff9df5effe4563a327b228f275bae87c8af4afd9ef3b03692b4958f93f71ef35ed7d81f791fb1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h418184785ca9819c081d724695d5aa956f14f1f0daca5ee61e1e828bcdc1918c1cc02c22d20be5bac689a10865;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf17deff441ca9875307cc5b84414d4b096b07dff08f7ea026b374dfd25595630bf97ab78e1f995820859fd44db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h770d70179f4117bdc89841f8295d0234ff9acce2823ad0df6c331b16bf1d802588a57ca30d1c2fe0f9fe8eb6e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8217973f5ea83b9157382ba1ae581b2d191e6dc7c42b362c17fd4755db5f925d351d5463104c7c06d30f60d2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c2208f89d8abb14a35f5ca4c12c5607c6757d7a812c4467fe9f55067897930886d238d474d11f2c107be7852e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154d81c56bb536e06b5e07cb94c0abba69e3e84d9e7a9a7dcfb331778513b0ac63f44ddcfa65098c5b5519cd478;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e0bafbf001a1ac08a44d256606f534721a77de55775246955430c2e355fc4fce454134ae16264584378af2944b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1afd7656aef7b60b40055d607cbbf2294c53f27911b0a558c856ef232f70f5c8d32613b0ac2d2f02b614d7f37ab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a0649f456241c970ee531300ecbdff7f41fe3e5ba7034f76b3f5702f885cfc4c51e635590806089771df34aa1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195118a9745bcc496085edd910220defadbe549cca7289e93afc8b39933572749de57ad529e010d66deead082b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a55211194767c1769e7c8c0b59b12402a39ca5b7db77f756778ba7569cf5211db290e90009389627ac3aea2ebc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12bd0af553c0189943cb443f922a6e00634a1a6b7b9e76ef6c05d5df94655f021aac01445a741cc2b27b4865bec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h85fc9b3a161fd14c309960b9e2d201309b2e984f8d61ff55cf5a6a9ae4f6a9605c628048ce072e7f167835a52f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb8e2ecddd17213b5d6016f263631de366fee4a67d1410c6a77d26fb6e30040930699c002c08b422d8b011d57a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e52fc31deeb05113556860dcebec1d376eb2030bc7ecfb6e303064a631a82a9945c3fe31a68e6d3a3e75a351;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122f2c3cae640e3e9af9b2f93956f47a2e206263561a8d5d305bde78672a67e38b68223b813484fc58b27a64782;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haca633888282e5d5f7eeb0a2f96b8d9dabec4f18a7f744859cda2cdf3bbac0f1fae230dbc5b88869241ad7ec50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1834323d30efe7189f45cb8dc3630242fbb1f90c2f991d5c422965aabc0d25af6387923ab035f898afeab04129d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc72896a476a244808ad0bba67df3704242c87579da3f1e70f46cc0f704a71778afd9629313a290dc7907ccfed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h171f83ceb8608437935a7a4dd73d0359f2f7e5cc7f06f6bc72be006cc356d99ca60928b0fb79926eddaddadaa0b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b20434e878d91d22f9e26c578b91506a8d130d476c3b7182e0f96cfaf7e4287b095704e2e25da2bc148cc0702;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163bde5c21738966d2e2849cc983cebcb89f9f6be6a93946003ea01cf5d1d777aca446d7fdb86004ad6c1b70803;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132d07f936e68d327a297ef0b2582dfef204a950878b7a4ac7250ea20e8d4eae818e06a92a6ffc969867056c049;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28680a44a6d4376b31718f2f212000e5b97404f8dfa101f068844cdbead1ca4cd58228e0524211ca93f0c94f2b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a546a530ccf23e79609c1b2fc751d3d7b521bcbaad05acfd1804ec988930dd39ed84a7e58666b1fcce85a88ce2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150e62a858fb90b265190693b37f8dd4718e90750e77a7c908e6f53459ecee1cef9a0e04e0071233b6f39ad4a90;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a377e2699165f6b49288ae53fa7ca3e3cf8924abd5d534a8608012908bb3fa01711e9aaf5437223d82dc3422e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195661c9a9d737483d6e8fc82b9f7fba4eeadf640de4f71227c4683dc2964010e1c927a3d3f90378832036b0135;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37a5591c8097b11af6f0a4b288d3fec7cb74a6fd0bcc8a41f2de8c69592feee8345ee5ec5212c237912eaf548a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e1c44fa4a457e0f33536dba4fd8b8b60adb6a3e15b1cebae563f7c2ee5e01e6a9fab1c87b1b7d62268638908c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h305cc76dda1e4d96dfb7a83119411635127764ac7f7a4eb515056dc59fd1577fd072ad9831c8f0a34dd155b472;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42c618b12017d5a20a67b4a3cd91bd933b5f04ec803d26b3ca243fe2e6a4cf03866b742d67f7ccf56368ede557;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50ee6433aff25b9575006d2afb364fcc104916c32d2f677f7400fdd3fb9bf8b393664137329460780344e94db3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1093a081ec4ef80657a7bb417593e2d0e88f80015443eddb41840415aea2a068f706dac9e4801040d947ac5438c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e94595f0b38f23380e85c66e356de29d7988fb15a147f6d923a48223eb9d217b0fc6192bfe2a848311ad0384d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf472e527173a7d99ef648800e437846e105f483d8ca5483022b55c67b021054c33b83a950cfdd33632763baef5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1227f0f1b05ceb113051a5a061e50f8f202c19eefaa2537f5ebc4339a488ec0b4355d8145af9e5b2292ddb0c9ab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d33dce34475b20f3ea1625d2e4b727f135b5e3169628777f2209ebc5208ac18e43925bc2881f394689648f7e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f21ad1e91cbc6820e2739499fc1daeaa266fda2e6f9ff0331b358ef597a7a2da30533ba7a06edfe91ab094444;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16120204c512b24d2e6ced0270826ff21d04dedeeaf4d63077f3cd9dc821544365ccc28288c0b2fb1466e324eb8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he0f4ec509ad8a9f05ebbfdcc4e759ab65eff5fc8361546975b1db38aa2f7872048dff9575a347f0ace083040bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187d07b0fd45425f6468e299488713c7b74b40bee190c00f158b1275469c28f5f0282cd55ceb8556cbd93a5aa0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19da8b255b527642b17c56cf7b6c45f692005222273e8558eae2cd2e09d725248a83839d7ce046a1fbd89d05281;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd56b74f923c89cbfab7dd83be1a7b86d8d03317cace0ed5b7b64bffc1eec90bb3faab086187f5f242892d8bbac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb9b7409675382dd3d177965db06cd8e19c63b094ceffb1dd6be458a9eebeb84fbe8c13c9371264049e35870ab8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38949a0d64ee8739d56693d842772b0234086014b86bf0541499d87f8ce8858b908a84dd081b954581c2a04c13;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h40fb958bf55bc94fbf97a17bf2b673ac9c2a5e546768ca668524fe6639dc50ddb2674459f9f36134ebb1cdc6e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11aad0bd46356cd5f800504c120a69553019f934f869e9fcff3e61631d99c22cb881d65d71186d20d4052276e5b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b7eed99d88085dad0af154d1d076c572ed543726ca3ef97f23aa312682d23e6ac170aafa56068729c5156fa17;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a9c4d8c9d2dd66370729876509a1f60ee830e3f436436ca0a18d2d6a4be73ab28e7d44b87472881193bff7d32;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e33bdf98529ea20c6030ed769f1147eeade97bc6efa5ec6bfa609fb8a58ae220d48406d31c3a3a196aa9642505;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17771a4750b0dd643a2d84376607c2d0622bdc628d1aeebff1aceb6c0a9a9326e33c7911670f20446e39a743b67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h123fe99f00f6fe9cd8380b7bb668d018f787842a4b2f5c646448dd024364aad3585a2e93db145c7d1f961d4777b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h115b6f59bd3121a81487b5e79a3eeafdbf39b74a1dce43f4706c629dd4439994e368b9aa82b9667933a0a4e0961;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf696de910e39ef2be841445adbf3a9166421f8d81722254ff29da4e6ef06e58fdb2196aa85b38d0834a0b61a47;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bde6aca84f3b3d5a16d32c37a7295404bdda382167b52cb6e4cc4566142771c0c500f29679a91c45a9d0d2fa9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e37959c16497166b7419417ce3bf08756ac9d4c4b1a79bb2f76a95b27eb87d4119263df97623ee9b66fea13e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2dd5e92b20c1df0196dd293ef32b76a2e135fa27882bfc8db41fdddd085f01028e0002af09e3bd385edfa7f26e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb74f9f8acfba11badb1a25a962e480baca52588937ed65eec2d5fcf878e27711f9ee0a91cbe0462dfb4f9f3e7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h52a41ad6f62a3c26e12746e3218903b906e004ca4c1dd04211c69a5c18c3e6425e2333f7289a88eb44f1c74100;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd26529b5bfe8661afe7ba9985911494b15b52da9b5607f6cc85fc5c8cff2fb275735ab2321db16f743b1893315;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h370eac123b4c9b49bcb1a8a1d75d9acfc9c538f803af022dc32d49e60381d9253baa0b6e97ec9525b3e9c5043a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1968d5874339005f4f6ee4b520e99b999fc19faebd0f497bdd0b9ec878ed298cb95a3c8a344f8382a06945029cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe9bf6ba156c6661e81710b82d0ba367b7a58b30aab84da2206f2bc63c6767979c54a4372a751794d3b059991f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a6d03721e05b5ad1fc0c0e668eabf31f36f7fe18b488f6bfd8349ecfdda1a727e8d3a6ca119c350f1aeba94c2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186d63735a7117e2b3c7b34610de139affcd103a7763e6c8034b77cc0924b90d3721d56c38cc7fa76cdbf450af6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12f5c0aa849395ca3fbe73767199d00c6dfee4780da4136492691986bd30e8f9d68d606d4ff77592de5ea1f7a1f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b485560a6558c142ca45094571fa7546f93735cd62909f16d1c849f5fa07c854f7c9467c2f56bcab84fb35467a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e9acace4b236fa11e974657cadc43e36af3ed6453d5cc65083b336df94ccd070288934f214ae70eac9d25a176;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13822ef2f88bed80f4ced209adf86b1f381579882fe02d5dec80cf5758699a4e2420446d81a354489517e6a3be6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5856a6cc433a1c548abae0ff30fe70b7299cb3dc78fc3efc0d5b0d608b7f95563812cc5511396dc85119508b38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff2e4fe2bd7023ebb51e567884b3e8093ac5a6694e05a089faf66b1c60c15fab059951f98fce865b2276c602de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc7d554e2002f803a36848c1c7a78fb773e1fd07a4ab87c606f3f5e795cef258f47df62cd277d227f25ac636a4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75af40f17a50d7f4a182f9844daebd2b736d51f19dd3f72bd8dcea466f245b4a23b7c27fb6123f0aa95c9778aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf8770fda1ef2db2274b249a9ccd2662ad14b4dde3cc7f45a8ae109e2739df2b76f637a388d520313decf19a6d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8ffb16b2ee32ffccee19c63776f113273ac91ec9173f61ae65dbb40b6fa83796eeae9a1a305691d7faae6fa1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14847ce106af7ed42d274d0e861707be33c832260e05569340ab0a348307920b91a4b5650a4768e5dcbf2a6de8f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12aa68bae6c04e1ddfa021b140d0219f334e2ad09f52233a4431007b0f1ca16fa5e68be51f68a38977624844cab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8097d41b646ccfd6d411d2da4721993769e9e71dc604c9d4ecf4e24578092b9469c9c969609e6e65d8f4c2cef6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165d62e93ddc663afb09f8b2b69107f51f3c0cd998669ae01bc92fc240797718bdeef49232767ccd2bb9b36f488;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c387d6cefcab6ccd80fc891ab669c27ad145b3de1e88d901cfef94365e36b3ca8a5387f633960588417b5cad5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd09d4d7495d651bf9702c27ffaac020d73771e313d920c065ec3c5b5ab0e64472905c8f170c79cf31bdd318c58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15e7ebccab24bce5c605f808088505bfbf0ef88c2224b0e12bcf3c5b14c648fca709516ad08ea8f21ebe513f6f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ba3ac5a845542386af7bf0cf2ddd407f666cd82cc731e50fca5b8606285678c51fc4f6c599cb4fffabad361cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114581c706ba0cd64420d7e6d1a757b394ff2de3b63b647aaadaa9fb340fbf06f0f77feb335cfc3ee5d539033dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h40c28de20ed1db91e700b64212b7073ec6baab7e007ef7622a5781428371d9351449ef9406edb04d9447c04088;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6cce1b88c9e057057c420d079aec60791af4644b7cb15396c460289626b9400d4f0bb67114b9d3f3943e6952aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h140a9359b547b001a2b5300a391c4c9c70bd578a9666294ff04f09ec4f95b8ab22fdc9cc6cd52304f5dd8db9efd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff6b316fd046415c255b1c403e6d5aab85317229058942241c8b517aeb0b50259159bb876a5dc74096f1492aa4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fcd7549ac12b0066288b6b276f4d97fbd87e0be9e32712666b3643482d90ac07cc3bb9aca9046f9338666204a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h21f4c9ca5422e140bdcd2af113fd5443da6615a18c7a48568b77275841ea8280989cb7e6b46442d47a4b1dc1ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1ec8c586abb235b747274b6d7a1340c33e416f3e2d5ed3486cd7b8518a7b221824776fd9f6e162f9c1e27fe90;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d6d0842129fc5dfa2f9daba9a4bec511c1c3dda830ba794bce2c9170d9930141e4b05e084806504b21fa453da2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b77f19f341bfcd6bacb43378c7baaccb45493c506c943616a706a8f70dbbbe1bb0bc79f3ba37d988ea4fba646;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha9e2b98e14c27bfdfa945eca36a62b318c44a87d990fc10453c897b0b36f8fa7216d5ae0a2b56808db394f2536;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17040bb63d44a2759b898d0aa41473cfc073b02fe334c67f55a313d79ac48c91d2fb2bba0c9142d1c766cc6517;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48609e3bc30f0c4cc713ef7c481b5897cb55b5e1211e46b65798a1509de88c1b17b3bb7a2da148a7d3cdd41e17;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h44ccaf98d5e9e8dce2112cbc5ff34422dbaf3ff0d6f08f3a0c19059d68c65d6f1cd778e52ecf8aee9562751170;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e786792fb4b1ed2150a9023cf162a434bc39f49b5dfd58811673c54811ee84f36a2b932f2bb7765f14b72eea97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h700c68615228b39724ef8e5aef334142d9557cbbaa54a9c292e522961917336f4d518c90f525d9471405eade84;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h915bc53fbf1c7be7a2f7a1470b3724b4bdfdefdb94485e4aec88356a6fc9a57d717a9b3a6f426cce59ef5fdbef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14dd11189b7eaf4d309de7418bf45a9a8549e0953f29c55532cb9230e81f7a0f2b37134c724eb20afeb68f6cf48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e413381daac508dfa06a2e17ce68974e0afa71b9f27f08cb03917ed85df0788ff2f5372e13d5f1cfd415d829f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63782b55f56b2294f05966ed20524a1aa106ba7a0a92471447ca4ce0fbc195c53388354b06d505f0f3c1e6f9cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffe8b7a1ff343594cd91484b243ed39c78033d2cd6721ac7f2b062e04dc9818d2a6749f81f087d76dca3828950;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153ac3567b2a1190577b9a584df389b3a1852609fc3dce98ba4a41de613b8340f524d09d4133a20518ee3ef063f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e745686d9342b6193dd42ec2b352602abaedd700b717da63ef3272aa9e85b62ada45956a5a6dd9c3c55865b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b748641531d2f4ac71265e7314bd156923b655c8588408c0ef750539a735d923a11f368b9a07b5e044c9d2f06b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e863744dcb96aacf5563b0df7b51c3ff0dc8a744b4cbb7f73a60aeb4eb029dd7153c5f5a79e9f83e5862feb05;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a82a8475ab6b1de1354ebe965c95c2703b82265e9e84d71caf6d18670d5e7778264e6081c3488f403f85db7789;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb83f00119db2b11795fc617c267bc04f470c09d29f806e15a1daf06caf52eeef375fc299b172270d365a16e60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122d6cfb4295a3488f26111668f065fee8abac125e64251446f25876d5969dbc0627246acb3a93c58b201ce9d9f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1384ae6c1441c028dabce966c2404fca0a0c2da42d163b74a356a2d5083e56b9de159de3a7acc18836773f536d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108c942cd36403c71c64bd5d3fc67cd31a13463b563526819d4075e6ad6df57a5c7f8866a078e87f806827f42bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25a66d86ce6f412c658b1b88bb2ccd5ec0b22c4b8f7c06316a59b2e1197ac249ba2a74c19840269478d3890398;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ffd444fd06e043ebb87f116780a8652b6d3dbd794a8f2e37b82bba7a0df9db11cc67853e7fb982c8b0499f2c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b2af9316f2109d9d1fa8c3a11e3bb4bedd64fb4152e05ce936ab36d7edb5dc2bf9dbe7a4a9d6f9103eb0ba9c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h79c7bac9bb2c23885149618578f3ae06ef9fb72b47b5c8b3eb7410d42678cd369d6fd4b5a1bcd95da1c925e5b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1379a2abdf6ef397c88691a5498d51eeadddae3b7f42a46daf591196f8c8c9bf1a92ad34bac78822f0f92d11010;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70ac104dee534bbde9951bea668a367ebacdf07a3dce8877f60cb2f0c1a8aee3e99511113302f9a0f4c061e86c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d4083e70f331349cd536f738450d5476d1b4dfee50a34d6ce919f264cc6803f207ff42570c71c3609cafcf3b11;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb11ca737ea1942b5e2cf0ae894daea54aae396864ff85d1ce438d46d0e3c51cf92439aaaf743b5e80931a1939f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha4b5aa821738a9fbc0e2dfe7777822b5563eecc0b2b3fba0844fc381b1413a94b731d8e5641ce71698ef282182;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6cf4cce7ff0fd6f3cce926342265426ded5ba60824f209b9ca86af55279af8e9cec8251a64ed1afd8f6aebe39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ce408e7e21fde79483d02fb61ed3fb647b7760081a09ac61fc1019a3a9a62840a59ed7ecb7eed96c66c56c368;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a98c722a11d0c15ad64439d6eda1a2c62565c6daacec7bf93d0fc33371bdf4798a58123f0bb595e72f788be13;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19148321b1beccce3cdc7f4438bbfd794326066478bf7e25756eaf38c65ab0b0818a9c9030c71c02a71e1ba3978;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10dfe7d3536363ed7ddecc079d159bb4fe2bc77fd67da6faf37bb6fca73c6a2d389c42fe7e06e6a08c25c3f8dcd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14534fd95583809023aa44ff1878037c6ab149b6d2fb70e6b53840fed0f653ff385c47979f9ecd827e0676fd4fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ecaef578c86837ffbba81b4b86927246f523c1fe68e5a9c249797c53c35c62f43a5c8cd38803ee333bb69955d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f7e39a10b894913c8a4a94c82c063a029be1237e596e8cac30eaed1a3858352a9ad10f1eb90a905a9ed8e6c31;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h115eecd3fbcef5807f73373e2dfbb8f4937b6c0c1f9a0537a3530baffcaf14f0a6c7adf522c23819ae09ebd2d88;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8741bd07059234723cbc741ac0e78cc827f62383435cad95716b64a1ca36d08dde31e5f647eb61108f6849c2ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b769b5ea86ca3eb71c2174b08bad85d1dcf6c891296bbbbf283a7a4e85186f06da788ed4ba567d8bfd8e31861;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h594cc39089fd3e79ac0e31c4fef57216636b92f6ad1d68c85d82192243efb441bdee882261e996d05ea539398b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d7e3b7347fd88fa66bb7582c6c4d48d411abb7664b2fd0e2944b9ad799de4271a610706c33ba394255a223f8b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10de067b7cb8acb1ac00c4bdc7c8382f854dd8dd69e3592e895c7f5feb3deb7409fc0a528dbdf73052e4ed91c76;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13de7eae6951cdcdf6bcd1cb3b617a9b00c65f35e2b57529d638122121753008c6f6af31dbb013597a32f453a2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd17557d918ca56314c320e65872dfd517ece40c82a6da7205438fd76c5665c15985e9014358890d79d7270420;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164a9703401d8bd95747d0c46c41f6f6b949afec71d3db24a3522e04d120c35bb3139ced7b41385507207129bcb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h49f371cd6a0a31f8db48c94a991c87a6c5874c008f115faab1135ec723dbed3cae8ca9e94521b7d126207eb8a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h615e90ce74d2766bba66140cfe9e5142346daac69b76a8697145f6a17d74ac88b6036f16525b6806875879e000;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3802b692062d8cbda6ab26876229dfacd4385d12c98833f7072aaa1e760cc5444a3ef77bea27a798620b230d06;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12dffe816da1f4058a2ab1583839fc7f89090cf744419b61eff1100a31c163da7ca42656884a4f3119c0e0a9738;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca42199fe3109943b0e6d5af807421c4fbdb4154a460c541f4d5d79df45ffbb2db2625f7f19326100f670b8067;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10b7d75138bfa291ccae26507b7fb5eb0dea4dd48d37f68a17acf56f347fc2156508cabfd27d02650b69b1deb04;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc279d3c5c983376e6362e9c62b2c7d4d270cde7ab180d9c439366c8a627375a6589b7a495588a256bcf5ec20e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10834c5357d2ec5b063a0ecc778cdae08a3829274a50873366cbe0e06c69deb71212bec57804740d1daa7b2ee9e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19438f6d9b338baeff587c9efa75a91eddc63510715583526d3acdd027d2d2e4c33afc8b279b4404843327b857a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33eb80a125163543f7bc13bb7f98ee02c53008d8be517354e211e44781acd7fe5b4fbe53a03cf1501c79f736ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4a36def5d3ac34c6f735dbc7cf6d80f26a825ce8742c5a21463031393952d3fc4099e00cce94ca8dc64c15752;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h942280853a4c0b6f51e1349474197408d2d6b0ae6bf596efa181434b170347f5cd6da6c670b8c0b1eedff7492e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12602ad5842795e9a638292ddb43ce564a3e0be0e05f85cc4b96300fb350cce5973f19df6245901bec2215ba765;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdbc92ddf8bae2ce6b89a833a5644864ff8104ef829f23baf1d4419be488b2aa2dd6d6bddcebc2b14d4112cbcf9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c2fa65241a05b3b35480dde13b7486f2d15b24e9cdb3fcb3027263aa019113291503fb6556de2e5720cd9d0bda;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ccbbce3c3a115d5547fb5fbd598bea6135f63788975bf505490a76dff56903a5246017c15b172cfcd1314b775;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab76d862060382033e1ec30ffed867d5f63fae05ec5604977bdeadf5846c5145286d2ce73277ff55ebf5bf1016;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17417fe138c2173bd559b6111c9726346295eb2aafb2494f9d48fe506a31925c05a25f0d8bfcf93fc7734464df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6775c7367c5fe90ed89a09a16d77d607def492c9307735e2f416f165d00ee3bbe512676ba7a4d0527c3fe9bc58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99463727abd0bd5a6bf7329f370bdd0a512b5b081898a4330c6ae534be89b66b174cbef7d9978f75afed9d9971;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1990c6450793b1290c000a55e45b5b7c8d83b18017c1a24969ffdfac59fdae789317cc5901d6a1ae6b540cd416b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba147df0563f38b90b6d0c7e2e5df928d9a7b15eb7d91bb78707b0f8ace2b70b8293c8132e4d6343ec16b85bbd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4f1a67338bf2d034a88daffd30751d44f8e0e64fe60d8b1bceede16050890304ab77c9ff1ff41dbc0541dcf1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he9323138984b3bd1977cfc00082aa5967605660ce271091ee82f11f891fa45fdd9db442f94a87038a72b58c356;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fbd966b73ac31cca6e77d3b258a0053c30b26c2505d1c2e32dfd67bcfa7a05f0304808cc43f77268e27661caac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168d750cae102fe6c501ebffc8e7e59223855319eb69b1e74cc4f0a912fde1e1d72874f58c1a67519bf871995fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec814f9de5032031e3fc77db294f9ade118035046db9df0c02ceda71eaea5b4449e2e2644814dd02b6d2005662;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1737cb5f24fa2348d30ed345421a7bf1e249e47dedec57bd2814c71a3c188626f7502bf1d19957374deda267f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d52b9b295195bd68420b4a9b4972df2d6ff19067153c4956b80d68d2dbd870e057de6478dd284bd5d5c99decd6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de8fea9e6e77e84a434c42ac8b6b136415765112df6bdaba7a58f0911bed129bbf04cb3cd288fcce5c8de8fa04;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a342277631c4c713139b5b6c7ae3b3230390436a88b8cc83dc758ef95c31d24408aa5a44f8da97c04b2072aeb5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h145e2487bbb55aeb6ce22081754d1c19f3b678766f610931a25433b6a0c24a78d6a6ca604f755ed206ec72160f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h101a2c7d261b8fa879ebaa473acd85afe665f966ceb1151305d3bca9c4780fbe6fdd316f5e2d5eb35c7210792f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153a209131c206fe013e43fdc220d8ecebdb0d185eadfa4529337d87efac5a910417c6a34492aa977737e677b7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h144b6a97c34e1c8788b2ef8818b6feae24320ee44392c2f0ea3dfbb0dd6e5b876de5fbe7ffe1d9316495a2a671c;
        #1
        $finish();
    end
endmodule
