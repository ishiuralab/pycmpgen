module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    compressor_CLA128_16 compressor_CLA128_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
        src12 <= 128'h0;
        src13 <= 128'h0;
        src14 <= 128'h0;
        src15 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA128_16(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    input [127:0]src12,
    input [127:0]src13,
    input [127:0]src14,
    input [127:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [0:0] comp_out21;
    wire [0:0] comp_out22;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      input wire [127:0] src12,
      input wire [127:0] src13,
      input wire [127:0] src14,
      input wire [127:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [0:0] dst21,
      output wire [0:0] dst22);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [127:0] stage0_12;
   wire [127:0] stage0_13;
   wire [127:0] stage0_14;
   wire [127:0] stage0_15;
   wire [45:0] stage1_0;
   wire [63:0] stage1_1;
   wire [38:0] stage1_2;
   wire [48:0] stage1_3;
   wire [59:0] stage1_4;
   wire [56:0] stage1_5;
   wire [47:0] stage1_6;
   wire [64:0] stage1_7;
   wire [55:0] stage1_8;
   wire [57:0] stage1_9;
   wire [53:0] stage1_10;
   wire [51:0] stage1_11;
   wire [56:0] stage1_12;
   wire [71:0] stage1_13;
   wire [70:0] stage1_14;
   wire [37:0] stage1_15;
   wire [35:0] stage1_16;
   wire [20:0] stage1_17;
   wire [14:0] stage2_0;
   wire [13:0] stage2_1;
   wire [19:0] stage2_2;
   wire [19:0] stage2_3;
   wire [27:0] stage2_4;
   wire [27:0] stage2_5;
   wire [16:0] stage2_6;
   wire [30:0] stage2_7;
   wire [28:0] stage2_8;
   wire [20:0] stage2_9;
   wire [17:0] stage2_10;
   wire [37:0] stage2_11;
   wire [28:0] stage2_12;
   wire [18:0] stage2_13;
   wire [34:0] stage2_14;
   wire [26:0] stage2_15;
   wire [19:0] stage2_16;
   wire [19:0] stage2_17;
   wire [6:0] stage2_18;
   wire [1:0] stage2_19;
   wire [14:0] stage3_0;
   wire [8:0] stage3_1;
   wire [12:0] stage3_2;
   wire [10:0] stage3_3;
   wire [8:0] stage3_4;
   wire [9:0] stage3_5;
   wire [10:0] stage3_6;
   wire [8:0] stage3_7;
   wire [13:0] stage3_8;
   wire [12:0] stage3_9;
   wire [7:0] stage3_10;
   wire [16:0] stage3_11;
   wire [13:0] stage3_12;
   wire [11:0] stage3_13;
   wire [15:0] stage3_14;
   wire [10:0] stage3_15;
   wire [19:0] stage3_16;
   wire [6:0] stage3_17;
   wire [5:0] stage3_18;
   wire [5:0] stage3_19;
   wire [0:0] stage3_20;
   wire [5:0] stage4_0;
   wire [9:0] stage4_1;
   wire [2:0] stage4_2;
   wire [10:0] stage4_3;
   wire [5:0] stage4_4;
   wire [4:0] stage4_5;
   wire [3:0] stage4_6;
   wire [4:0] stage4_7;
   wire [4:0] stage4_8;
   wire [6:0] stage4_9;
   wire [5:0] stage4_10;
   wire [3:0] stage4_11;
   wire [5:0] stage4_12;
   wire [5:0] stage4_13;
   wire [5:0] stage4_14;
   wire [7:0] stage4_15;
   wire [6:0] stage4_16;
   wire [5:0] stage4_17;
   wire [3:0] stage4_18;
   wire [1:0] stage4_19;
   wire [2:0] stage4_20;
   wire [0:0] stage4_21;
   wire [1:0] stage5_0;
   wire [3:0] stage5_1;
   wire [2:0] stage5_2;
   wire [6:0] stage5_3;
   wire [2:0] stage5_4;
   wire [5:0] stage5_5;
   wire [0:0] stage5_6;
   wire [4:0] stage5_7;
   wire [1:0] stage5_8;
   wire [6:0] stage5_9;
   wire [0:0] stage5_10;
   wire [4:0] stage5_11;
   wire [1:0] stage5_12;
   wire [6:0] stage5_13;
   wire [0:0] stage5_14;
   wire [4:0] stage5_15;
   wire [5:0] stage5_16;
   wire [5:0] stage5_17;
   wire [2:0] stage5_18;
   wire [0:0] stage5_19;
   wire [0:0] stage5_20;
   wire [0:0] stage5_21;
   wire [0:0] stage5_22;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [0:0] stage6_21;
   wire [0:0] stage6_22;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17]}
   );
   gpc606_5 gpc18 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18]}
   );
   gpc606_5 gpc19 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[2],stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19]}
   );
   gpc606_5 gpc20 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage1_5[3],stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20]}
   );
   gpc606_5 gpc21 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30]},
      {stage1_5[4],stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21]}
   );
   gpc606_5 gpc22 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36]},
      {stage1_5[5],stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22]}
   );
   gpc606_5 gpc23 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage1_5[6],stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48]},
      {stage1_5[7],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[8],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[9],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[10],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[11],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[12],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[13],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[14],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[15],stage1_4[32],stage1_3[32],stage1_2[32]}
   );
   gpc606_5 gpc33 (
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[16],stage1_4[33],stage1_3[33],stage1_2[33]}
   );
   gpc606_5 gpc34 (
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[17],stage1_4[34],stage1_3[34],stage1_2[34]}
   );
   gpc606_5 gpc35 (
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[18],stage1_4[35],stage1_3[35],stage1_2[35]}
   );
   gpc615_5 gpc36 (
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage0_3[91]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[19],stage1_4[36],stage1_3[36],stage1_2[36]}
   );
   gpc615_5 gpc37 (
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage0_4[30]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[5],stage1_5[20],stage1_4[37],stage1_3[37]}
   );
   gpc615_5 gpc38 (
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage0_4[31]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[6],stage1_5[21],stage1_4[38],stage1_3[38]}
   );
   gpc615_5 gpc39 (
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage0_4[32]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[7],stage1_5[22],stage1_4[39],stage1_3[39]}
   );
   gpc615_5 gpc40 (
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage0_4[33]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[8],stage1_5[23],stage1_4[40],stage1_3[40]}
   );
   gpc615_5 gpc41 (
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage0_4[34]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[9],stage1_5[24],stage1_4[41],stage1_3[41]}
   );
   gpc615_5 gpc42 (
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage0_4[35]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[10],stage1_5[25],stage1_4[42],stage1_3[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[6],stage1_6[11],stage1_5[26],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[7],stage1_6[12],stage1_5[27],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[8],stage1_6[13],stage1_5[28],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[9],stage1_6[14],stage1_5[29],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[10],stage1_6[15],stage1_5[30],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[11],stage1_6[16],stage1_5[31],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[12],stage1_6[17],stage1_5[32],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[13],stage1_6[18],stage1_5[33],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[14],stage1_6[19],stage1_5[34],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[15],stage1_6[20],stage1_5[35],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[16],stage1_6[21],stage1_5[36],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[17],stage1_6[22],stage1_5[37],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[18],stage1_6[23],stage1_5[38],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[19],stage1_6[24],stage1_5[39],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[20],stage1_6[25],stage1_5[40],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[15],stage1_7[21],stage1_6[26],stage1_5[41]}
   );
   gpc606_5 gpc59 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[16],stage1_7[22],stage1_6[27],stage1_5[42]}
   );
   gpc606_5 gpc60 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[17],stage1_7[23],stage1_6[28],stage1_5[43]}
   );
   gpc606_5 gpc61 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[18],stage1_7[24],stage1_6[29],stage1_5[44]}
   );
   gpc606_5 gpc62 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[19],stage1_7[25],stage1_6[30],stage1_5[45]}
   );
   gpc606_5 gpc63 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[20],stage1_7[26],stage1_6[31],stage1_5[46]}
   );
   gpc606_5 gpc64 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[21],stage1_7[27],stage1_6[32],stage1_5[47]}
   );
   gpc606_5 gpc65 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[22],stage1_7[28],stage1_6[33],stage1_5[48]}
   );
   gpc606_5 gpc66 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[23],stage1_7[29],stage1_6[34],stage1_5[49]}
   );
   gpc606_5 gpc67 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[24],stage1_7[30],stage1_6[35],stage1_5[50]}
   );
   gpc606_5 gpc68 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[25],stage1_7[31],stage1_6[36],stage1_5[51]}
   );
   gpc606_5 gpc69 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[26],stage1_7[32],stage1_6[37],stage1_5[52]}
   );
   gpc615_5 gpc70 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112]},
      {stage0_6[90]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[27],stage1_7[33],stage1_6[38],stage1_5[53]}
   );
   gpc615_5 gpc71 (
      {stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117]},
      {stage0_6[91]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[28],stage1_7[34],stage1_6[39],stage1_5[54]}
   );
   gpc615_5 gpc72 (
      {stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121], stage0_5[122]},
      {stage0_6[92]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[29],stage1_7[35],stage1_6[40],stage1_5[55]}
   );
   gpc615_5 gpc73 (
      {stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127]},
      {stage0_6[93]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[30],stage1_7[36],stage1_6[41],stage1_5[56]}
   );
   gpc606_5 gpc74 (
      {stage0_6[94], stage0_6[95], stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[16],stage1_8[31],stage1_7[37],stage1_6[42]}
   );
   gpc606_5 gpc75 (
      {stage0_6[100], stage0_6[101], stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[17],stage1_8[32],stage1_7[38],stage1_6[43]}
   );
   gpc606_5 gpc76 (
      {stage0_6[106], stage0_6[107], stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[18],stage1_8[33],stage1_7[39],stage1_6[44]}
   );
   gpc606_5 gpc77 (
      {stage0_6[112], stage0_6[113], stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[19],stage1_8[34],stage1_7[40],stage1_6[45]}
   );
   gpc615_5 gpc78 (
      {stage0_6[118], stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122]},
      {stage0_7[96]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[20],stage1_8[35],stage1_7[41],stage1_6[46]}
   );
   gpc615_5 gpc79 (
      {stage0_6[123], stage0_6[124], stage0_6[125], stage0_6[126], stage0_6[127]},
      {stage0_7[97]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[21],stage1_8[36],stage1_7[42],stage1_6[47]}
   );
   gpc615_5 gpc80 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[36]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[6],stage1_9[22],stage1_8[37],stage1_7[43]}
   );
   gpc615_5 gpc81 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[37]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[7],stage1_9[23],stage1_8[38],stage1_7[44]}
   );
   gpc606_5 gpc82 (
      {stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[2],stage1_10[8],stage1_9[24],stage1_8[39]}
   );
   gpc606_5 gpc83 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[3],stage1_10[9],stage1_9[25],stage1_8[40]}
   );
   gpc606_5 gpc84 (
      {stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[4],stage1_10[10],stage1_9[26],stage1_8[41]}
   );
   gpc606_5 gpc85 (
      {stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[5],stage1_10[11],stage1_9[27],stage1_8[42]}
   );
   gpc606_5 gpc86 (
      {stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66], stage0_8[67]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[6],stage1_10[12],stage1_9[28],stage1_8[43]}
   );
   gpc606_5 gpc87 (
      {stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[7],stage1_10[13],stage1_9[29],stage1_8[44]}
   );
   gpc606_5 gpc88 (
      {stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[8],stage1_10[14],stage1_9[30],stage1_8[45]}
   );
   gpc606_5 gpc89 (
      {stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[9],stage1_10[15],stage1_9[31],stage1_8[46]}
   );
   gpc606_5 gpc90 (
      {stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[10],stage1_10[16],stage1_9[32],stage1_8[47]}
   );
   gpc606_5 gpc91 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[11],stage1_10[17],stage1_9[33],stage1_8[48]}
   );
   gpc606_5 gpc92 (
      {stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[12],stage1_10[18],stage1_9[34],stage1_8[49]}
   );
   gpc606_5 gpc93 (
      {stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[13],stage1_10[19],stage1_9[35],stage1_8[50]}
   );
   gpc606_5 gpc94 (
      {stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[14],stage1_10[20],stage1_9[36],stage1_8[51]}
   );
   gpc615_5 gpc95 (
      {stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_9[12]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[15],stage1_10[21],stage1_9[37],stage1_8[52]}
   );
   gpc615_5 gpc96 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_9[13]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[16],stage1_10[22],stage1_9[38],stage1_8[53]}
   );
   gpc606_5 gpc97 (
      {stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[15],stage1_11[17],stage1_10[23],stage1_9[39]}
   );
   gpc606_5 gpc98 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[16],stage1_11[18],stage1_10[24],stage1_9[40]}
   );
   gpc606_5 gpc99 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[17],stage1_11[19],stage1_10[25],stage1_9[41]}
   );
   gpc606_5 gpc100 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[18],stage1_11[20],stage1_10[26],stage1_9[42]}
   );
   gpc606_5 gpc101 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[19],stage1_11[21],stage1_10[27],stage1_9[43]}
   );
   gpc606_5 gpc102 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[20],stage1_11[22],stage1_10[28],stage1_9[44]}
   );
   gpc606_5 gpc103 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[21],stage1_11[23],stage1_10[29],stage1_9[45]}
   );
   gpc606_5 gpc104 (
      {stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[22],stage1_11[24],stage1_10[30],stage1_9[46]}
   );
   gpc606_5 gpc105 (
      {stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[23],stage1_11[25],stage1_10[31],stage1_9[47]}
   );
   gpc606_5 gpc106 (
      {stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[24],stage1_11[26],stage1_10[32],stage1_9[48]}
   );
   gpc606_5 gpc107 (
      {stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[25],stage1_11[27],stage1_10[33],stage1_9[49]}
   );
   gpc606_5 gpc108 (
      {stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[26],stage1_11[28],stage1_10[34],stage1_9[50]}
   );
   gpc606_5 gpc109 (
      {stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[27],stage1_11[29],stage1_10[35],stage1_9[51]}
   );
   gpc606_5 gpc110 (
      {stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[28],stage1_11[30],stage1_10[36],stage1_9[52]}
   );
   gpc606_5 gpc111 (
      {stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[29],stage1_11[31],stage1_10[37],stage1_9[53]}
   );
   gpc606_5 gpc112 (
      {stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[30],stage1_11[32],stage1_10[38],stage1_9[54]}
   );
   gpc606_5 gpc113 (
      {stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[31],stage1_11[33],stage1_10[39],stage1_9[55]}
   );
   gpc606_5 gpc114 (
      {stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[32],stage1_11[34],stage1_10[40],stage1_9[56]}
   );
   gpc606_5 gpc115 (
      {stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[33],stage1_11[35],stage1_10[41],stage1_9[57]}
   );
   gpc606_5 gpc116 (
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[19],stage1_12[34],stage1_11[36],stage1_10[42]}
   );
   gpc606_5 gpc117 (
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[20],stage1_12[35],stage1_11[37],stage1_10[43]}
   );
   gpc615_5 gpc118 (
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106]},
      {stage0_11[114]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[21],stage1_12[36],stage1_11[38],stage1_10[44]}
   );
   gpc615_5 gpc119 (
      {stage0_10[107], stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111]},
      {stage0_11[115]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[22],stage1_12[37],stage1_11[39],stage1_10[45]}
   );
   gpc615_5 gpc120 (
      {stage0_10[112], stage0_10[113], stage0_10[114], stage0_10[115], stage0_10[116]},
      {stage0_11[116]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[23],stage1_12[38],stage1_11[40],stage1_10[46]}
   );
   gpc615_5 gpc121 (
      {stage0_10[117], stage0_10[118], stage0_10[119], stage0_10[120], stage0_10[121]},
      {stage0_11[117]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[24],stage1_12[39],stage1_11[41],stage1_10[47]}
   );
   gpc606_5 gpc122 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[6],stage1_13[25],stage1_12[40]}
   );
   gpc606_5 gpc123 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[1],stage1_14[7],stage1_13[26],stage1_12[41]}
   );
   gpc606_5 gpc124 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[2],stage1_14[8],stage1_13[27],stage1_12[42]}
   );
   gpc606_5 gpc125 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[3],stage1_14[9],stage1_13[28],stage1_12[43]}
   );
   gpc606_5 gpc126 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[4],stage1_14[10],stage1_13[29],stage1_12[44]}
   );
   gpc606_5 gpc127 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[5],stage1_14[11],stage1_13[30],stage1_12[45]}
   );
   gpc606_5 gpc128 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[6],stage1_14[12],stage1_13[31],stage1_12[46]}
   );
   gpc606_5 gpc129 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[7],stage1_14[13],stage1_13[32],stage1_12[47]}
   );
   gpc606_5 gpc130 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[8],stage1_14[14],stage1_13[33],stage1_12[48]}
   );
   gpc606_5 gpc131 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[9],stage1_14[15],stage1_13[34],stage1_12[49]}
   );
   gpc606_5 gpc132 (
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[10],stage1_14[16],stage1_13[35],stage1_12[50]}
   );
   gpc606_5 gpc133 (
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[11],stage1_14[17],stage1_13[36],stage1_12[51]}
   );
   gpc606_5 gpc134 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[12],stage1_14[18],stage1_13[37],stage1_12[52]}
   );
   gpc606_5 gpc135 (
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[13],stage1_14[19],stage1_13[38],stage1_12[53]}
   );
   gpc606_5 gpc136 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[14],stage1_14[20],stage1_13[39],stage1_12[54]}
   );
   gpc606_5 gpc137 (
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[15],stage1_15[15],stage1_14[21],stage1_13[40]}
   );
   gpc606_5 gpc138 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[16],stage1_15[16],stage1_14[22],stage1_13[41]}
   );
   gpc606_5 gpc139 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[17],stage1_15[17],stage1_14[23],stage1_13[42]}
   );
   gpc606_5 gpc140 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[18],stage1_15[18],stage1_14[24],stage1_13[43]}
   );
   gpc606_5 gpc141 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[19],stage1_15[19],stage1_14[25],stage1_13[44]}
   );
   gpc606_5 gpc142 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[20],stage1_15[20],stage1_14[26],stage1_13[45]}
   );
   gpc606_5 gpc143 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[21],stage1_15[21],stage1_14[27],stage1_13[46]}
   );
   gpc606_5 gpc144 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[22],stage1_15[22],stage1_14[28],stage1_13[47]}
   );
   gpc606_5 gpc145 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[23],stage1_15[23],stage1_14[29],stage1_13[48]}
   );
   gpc606_5 gpc146 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[24],stage1_15[24],stage1_14[30],stage1_13[49]}
   );
   gpc606_5 gpc147 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[25],stage1_15[25],stage1_14[31],stage1_13[50]}
   );
   gpc606_5 gpc148 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[26],stage1_15[26],stage1_14[32],stage1_13[51]}
   );
   gpc615_5 gpc149 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76]},
      {stage0_14[90]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[27],stage1_15[27],stage1_14[33],stage1_13[52]}
   );
   gpc615_5 gpc150 (
      {stage0_13[77], stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81]},
      {stage0_14[91]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[28],stage1_15[28],stage1_14[34],stage1_13[53]}
   );
   gpc615_5 gpc151 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86]},
      {stage0_14[92]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[29],stage1_15[29],stage1_14[35],stage1_13[54]}
   );
   gpc615_5 gpc152 (
      {stage0_13[87], stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91]},
      {stage0_14[93]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[30],stage1_15[30],stage1_14[36],stage1_13[55]}
   );
   gpc615_5 gpc153 (
      {stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95], stage0_13[96]},
      {stage0_14[94]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[31],stage1_15[31],stage1_14[37],stage1_13[56]}
   );
   gpc615_5 gpc154 (
      {stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_14[95]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[32],stage1_15[32],stage1_14[38],stage1_13[57]}
   );
   gpc615_5 gpc155 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106]},
      {stage0_14[96]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[33],stage1_15[33],stage1_14[39],stage1_13[58]}
   );
   gpc615_5 gpc156 (
      {stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111]},
      {stage0_14[97]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[34],stage1_15[34],stage1_14[40],stage1_13[59]}
   );
   gpc615_5 gpc157 (
      {stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115], stage0_13[116]},
      {stage0_14[98]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[35],stage1_15[35],stage1_14[41],stage1_13[60]}
   );
   gpc1_1 gpc158 (
      {stage0_0[99]},
      {stage1_0[17]}
   );
   gpc1_1 gpc159 (
      {stage0_0[100]},
      {stage1_0[18]}
   );
   gpc1_1 gpc160 (
      {stage0_0[101]},
      {stage1_0[19]}
   );
   gpc1_1 gpc161 (
      {stage0_0[102]},
      {stage1_0[20]}
   );
   gpc1_1 gpc162 (
      {stage0_0[103]},
      {stage1_0[21]}
   );
   gpc1_1 gpc163 (
      {stage0_0[104]},
      {stage1_0[22]}
   );
   gpc1_1 gpc164 (
      {stage0_0[105]},
      {stage1_0[23]}
   );
   gpc1_1 gpc165 (
      {stage0_0[106]},
      {stage1_0[24]}
   );
   gpc1_1 gpc166 (
      {stage0_0[107]},
      {stage1_0[25]}
   );
   gpc1_1 gpc167 (
      {stage0_0[108]},
      {stage1_0[26]}
   );
   gpc1_1 gpc168 (
      {stage0_0[109]},
      {stage1_0[27]}
   );
   gpc1_1 gpc169 (
      {stage0_0[110]},
      {stage1_0[28]}
   );
   gpc1_1 gpc170 (
      {stage0_0[111]},
      {stage1_0[29]}
   );
   gpc1_1 gpc171 (
      {stage0_0[112]},
      {stage1_0[30]}
   );
   gpc1_1 gpc172 (
      {stage0_0[113]},
      {stage1_0[31]}
   );
   gpc1_1 gpc173 (
      {stage0_0[114]},
      {stage1_0[32]}
   );
   gpc1_1 gpc174 (
      {stage0_0[115]},
      {stage1_0[33]}
   );
   gpc1_1 gpc175 (
      {stage0_0[116]},
      {stage1_0[34]}
   );
   gpc1_1 gpc176 (
      {stage0_0[117]},
      {stage1_0[35]}
   );
   gpc1_1 gpc177 (
      {stage0_0[118]},
      {stage1_0[36]}
   );
   gpc1_1 gpc178 (
      {stage0_0[119]},
      {stage1_0[37]}
   );
   gpc1_1 gpc179 (
      {stage0_0[120]},
      {stage1_0[38]}
   );
   gpc1_1 gpc180 (
      {stage0_0[121]},
      {stage1_0[39]}
   );
   gpc1_1 gpc181 (
      {stage0_0[122]},
      {stage1_0[40]}
   );
   gpc1_1 gpc182 (
      {stage0_0[123]},
      {stage1_0[41]}
   );
   gpc1_1 gpc183 (
      {stage0_0[124]},
      {stage1_0[42]}
   );
   gpc1_1 gpc184 (
      {stage0_0[125]},
      {stage1_0[43]}
   );
   gpc1_1 gpc185 (
      {stage0_0[126]},
      {stage1_0[44]}
   );
   gpc1_1 gpc186 (
      {stage0_0[127]},
      {stage1_0[45]}
   );
   gpc1_1 gpc187 (
      {stage0_1[96]},
      {stage1_1[32]}
   );
   gpc1_1 gpc188 (
      {stage0_1[97]},
      {stage1_1[33]}
   );
   gpc1_1 gpc189 (
      {stage0_1[98]},
      {stage1_1[34]}
   );
   gpc1_1 gpc190 (
      {stage0_1[99]},
      {stage1_1[35]}
   );
   gpc1_1 gpc191 (
      {stage0_1[100]},
      {stage1_1[36]}
   );
   gpc1_1 gpc192 (
      {stage0_1[101]},
      {stage1_1[37]}
   );
   gpc1_1 gpc193 (
      {stage0_1[102]},
      {stage1_1[38]}
   );
   gpc1_1 gpc194 (
      {stage0_1[103]},
      {stage1_1[39]}
   );
   gpc1_1 gpc195 (
      {stage0_1[104]},
      {stage1_1[40]}
   );
   gpc1_1 gpc196 (
      {stage0_1[105]},
      {stage1_1[41]}
   );
   gpc1_1 gpc197 (
      {stage0_1[106]},
      {stage1_1[42]}
   );
   gpc1_1 gpc198 (
      {stage0_1[107]},
      {stage1_1[43]}
   );
   gpc1_1 gpc199 (
      {stage0_1[108]},
      {stage1_1[44]}
   );
   gpc1_1 gpc200 (
      {stage0_1[109]},
      {stage1_1[45]}
   );
   gpc1_1 gpc201 (
      {stage0_1[110]},
      {stage1_1[46]}
   );
   gpc1_1 gpc202 (
      {stage0_1[111]},
      {stage1_1[47]}
   );
   gpc1_1 gpc203 (
      {stage0_1[112]},
      {stage1_1[48]}
   );
   gpc1_1 gpc204 (
      {stage0_1[113]},
      {stage1_1[49]}
   );
   gpc1_1 gpc205 (
      {stage0_1[114]},
      {stage1_1[50]}
   );
   gpc1_1 gpc206 (
      {stage0_1[115]},
      {stage1_1[51]}
   );
   gpc1_1 gpc207 (
      {stage0_1[116]},
      {stage1_1[52]}
   );
   gpc1_1 gpc208 (
      {stage0_1[117]},
      {stage1_1[53]}
   );
   gpc1_1 gpc209 (
      {stage0_1[118]},
      {stage1_1[54]}
   );
   gpc1_1 gpc210 (
      {stage0_1[119]},
      {stage1_1[55]}
   );
   gpc1_1 gpc211 (
      {stage0_1[120]},
      {stage1_1[56]}
   );
   gpc1_1 gpc212 (
      {stage0_1[121]},
      {stage1_1[57]}
   );
   gpc1_1 gpc213 (
      {stage0_1[122]},
      {stage1_1[58]}
   );
   gpc1_1 gpc214 (
      {stage0_1[123]},
      {stage1_1[59]}
   );
   gpc1_1 gpc215 (
      {stage0_1[124]},
      {stage1_1[60]}
   );
   gpc1_1 gpc216 (
      {stage0_1[125]},
      {stage1_1[61]}
   );
   gpc1_1 gpc217 (
      {stage0_1[126]},
      {stage1_1[62]}
   );
   gpc1_1 gpc218 (
      {stage0_1[127]},
      {stage1_1[63]}
   );
   gpc1_1 gpc219 (
      {stage0_2[126]},
      {stage1_2[37]}
   );
   gpc1_1 gpc220 (
      {stage0_2[127]},
      {stage1_2[38]}
   );
   gpc1_1 gpc221 (
      {stage0_3[122]},
      {stage1_3[43]}
   );
   gpc1_1 gpc222 (
      {stage0_3[123]},
      {stage1_3[44]}
   );
   gpc1_1 gpc223 (
      {stage0_3[124]},
      {stage1_3[45]}
   );
   gpc1_1 gpc224 (
      {stage0_3[125]},
      {stage1_3[46]}
   );
   gpc1_1 gpc225 (
      {stage0_3[126]},
      {stage1_3[47]}
   );
   gpc1_1 gpc226 (
      {stage0_3[127]},
      {stage1_3[48]}
   );
   gpc1_1 gpc227 (
      {stage0_4[126]},
      {stage1_4[58]}
   );
   gpc1_1 gpc228 (
      {stage0_4[127]},
      {stage1_4[59]}
   );
   gpc1_1 gpc229 (
      {stage0_7[108]},
      {stage1_7[45]}
   );
   gpc1_1 gpc230 (
      {stage0_7[109]},
      {stage1_7[46]}
   );
   gpc1_1 gpc231 (
      {stage0_7[110]},
      {stage1_7[47]}
   );
   gpc1_1 gpc232 (
      {stage0_7[111]},
      {stage1_7[48]}
   );
   gpc1_1 gpc233 (
      {stage0_7[112]},
      {stage1_7[49]}
   );
   gpc1_1 gpc234 (
      {stage0_7[113]},
      {stage1_7[50]}
   );
   gpc1_1 gpc235 (
      {stage0_7[114]},
      {stage1_7[51]}
   );
   gpc1_1 gpc236 (
      {stage0_7[115]},
      {stage1_7[52]}
   );
   gpc1_1 gpc237 (
      {stage0_7[116]},
      {stage1_7[53]}
   );
   gpc1_1 gpc238 (
      {stage0_7[117]},
      {stage1_7[54]}
   );
   gpc1_1 gpc239 (
      {stage0_7[118]},
      {stage1_7[55]}
   );
   gpc1_1 gpc240 (
      {stage0_7[119]},
      {stage1_7[56]}
   );
   gpc1_1 gpc241 (
      {stage0_7[120]},
      {stage1_7[57]}
   );
   gpc1_1 gpc242 (
      {stage0_7[121]},
      {stage1_7[58]}
   );
   gpc1_1 gpc243 (
      {stage0_7[122]},
      {stage1_7[59]}
   );
   gpc1_1 gpc244 (
      {stage0_7[123]},
      {stage1_7[60]}
   );
   gpc1_1 gpc245 (
      {stage0_7[124]},
      {stage1_7[61]}
   );
   gpc1_1 gpc246 (
      {stage0_7[125]},
      {stage1_7[62]}
   );
   gpc1_1 gpc247 (
      {stage0_7[126]},
      {stage1_7[63]}
   );
   gpc1_1 gpc248 (
      {stage0_7[127]},
      {stage1_7[64]}
   );
   gpc1_1 gpc249 (
      {stage0_8[126]},
      {stage1_8[54]}
   );
   gpc1_1 gpc250 (
      {stage0_8[127]},
      {stage1_8[55]}
   );
   gpc1_1 gpc251 (
      {stage0_10[122]},
      {stage1_10[48]}
   );
   gpc1_1 gpc252 (
      {stage0_10[123]},
      {stage1_10[49]}
   );
   gpc1_1 gpc253 (
      {stage0_10[124]},
      {stage1_10[50]}
   );
   gpc1_1 gpc254 (
      {stage0_10[125]},
      {stage1_10[51]}
   );
   gpc1_1 gpc255 (
      {stage0_10[126]},
      {stage1_10[52]}
   );
   gpc1_1 gpc256 (
      {stage0_10[127]},
      {stage1_10[53]}
   );
   gpc1_1 gpc257 (
      {stage0_11[118]},
      {stage1_11[42]}
   );
   gpc1_1 gpc258 (
      {stage0_11[119]},
      {stage1_11[43]}
   );
   gpc1_1 gpc259 (
      {stage0_11[120]},
      {stage1_11[44]}
   );
   gpc1_1 gpc260 (
      {stage0_11[121]},
      {stage1_11[45]}
   );
   gpc1_1 gpc261 (
      {stage0_11[122]},
      {stage1_11[46]}
   );
   gpc1_1 gpc262 (
      {stage0_11[123]},
      {stage1_11[47]}
   );
   gpc1_1 gpc263 (
      {stage0_11[124]},
      {stage1_11[48]}
   );
   gpc1_1 gpc264 (
      {stage0_11[125]},
      {stage1_11[49]}
   );
   gpc1_1 gpc265 (
      {stage0_11[126]},
      {stage1_11[50]}
   );
   gpc1_1 gpc266 (
      {stage0_11[127]},
      {stage1_11[51]}
   );
   gpc1_1 gpc267 (
      {stage0_12[126]},
      {stage1_12[55]}
   );
   gpc1_1 gpc268 (
      {stage0_12[127]},
      {stage1_12[56]}
   );
   gpc1_1 gpc269 (
      {stage0_13[117]},
      {stage1_13[61]}
   );
   gpc1_1 gpc270 (
      {stage0_13[118]},
      {stage1_13[62]}
   );
   gpc1_1 gpc271 (
      {stage0_13[119]},
      {stage1_13[63]}
   );
   gpc1_1 gpc272 (
      {stage0_13[120]},
      {stage1_13[64]}
   );
   gpc1_1 gpc273 (
      {stage0_13[121]},
      {stage1_13[65]}
   );
   gpc1_1 gpc274 (
      {stage0_13[122]},
      {stage1_13[66]}
   );
   gpc1_1 gpc275 (
      {stage0_13[123]},
      {stage1_13[67]}
   );
   gpc1_1 gpc276 (
      {stage0_13[124]},
      {stage1_13[68]}
   );
   gpc1_1 gpc277 (
      {stage0_13[125]},
      {stage1_13[69]}
   );
   gpc1_1 gpc278 (
      {stage0_13[126]},
      {stage1_13[70]}
   );
   gpc1_1 gpc279 (
      {stage0_13[127]},
      {stage1_13[71]}
   );
   gpc1_1 gpc280 (
      {stage0_14[99]},
      {stage1_14[42]}
   );
   gpc1_1 gpc281 (
      {stage0_14[100]},
      {stage1_14[43]}
   );
   gpc1_1 gpc282 (
      {stage0_14[101]},
      {stage1_14[44]}
   );
   gpc1_1 gpc283 (
      {stage0_14[102]},
      {stage1_14[45]}
   );
   gpc1_1 gpc284 (
      {stage0_14[103]},
      {stage1_14[46]}
   );
   gpc1_1 gpc285 (
      {stage0_14[104]},
      {stage1_14[47]}
   );
   gpc1_1 gpc286 (
      {stage0_14[105]},
      {stage1_14[48]}
   );
   gpc1_1 gpc287 (
      {stage0_14[106]},
      {stage1_14[49]}
   );
   gpc1_1 gpc288 (
      {stage0_14[107]},
      {stage1_14[50]}
   );
   gpc1_1 gpc289 (
      {stage0_14[108]},
      {stage1_14[51]}
   );
   gpc1_1 gpc290 (
      {stage0_14[109]},
      {stage1_14[52]}
   );
   gpc1_1 gpc291 (
      {stage0_14[110]},
      {stage1_14[53]}
   );
   gpc1_1 gpc292 (
      {stage0_14[111]},
      {stage1_14[54]}
   );
   gpc1_1 gpc293 (
      {stage0_14[112]},
      {stage1_14[55]}
   );
   gpc1_1 gpc294 (
      {stage0_14[113]},
      {stage1_14[56]}
   );
   gpc1_1 gpc295 (
      {stage0_14[114]},
      {stage1_14[57]}
   );
   gpc1_1 gpc296 (
      {stage0_14[115]},
      {stage1_14[58]}
   );
   gpc1_1 gpc297 (
      {stage0_14[116]},
      {stage1_14[59]}
   );
   gpc1_1 gpc298 (
      {stage0_14[117]},
      {stage1_14[60]}
   );
   gpc1_1 gpc299 (
      {stage0_14[118]},
      {stage1_14[61]}
   );
   gpc1_1 gpc300 (
      {stage0_14[119]},
      {stage1_14[62]}
   );
   gpc1_1 gpc301 (
      {stage0_14[120]},
      {stage1_14[63]}
   );
   gpc1_1 gpc302 (
      {stage0_14[121]},
      {stage1_14[64]}
   );
   gpc1_1 gpc303 (
      {stage0_14[122]},
      {stage1_14[65]}
   );
   gpc1_1 gpc304 (
      {stage0_14[123]},
      {stage1_14[66]}
   );
   gpc1_1 gpc305 (
      {stage0_14[124]},
      {stage1_14[67]}
   );
   gpc1_1 gpc306 (
      {stage0_14[125]},
      {stage1_14[68]}
   );
   gpc1_1 gpc307 (
      {stage0_14[126]},
      {stage1_14[69]}
   );
   gpc1_1 gpc308 (
      {stage0_14[127]},
      {stage1_14[70]}
   );
   gpc1_1 gpc309 (
      {stage0_15[126]},
      {stage1_15[36]}
   );
   gpc1_1 gpc310 (
      {stage0_15[127]},
      {stage1_15[37]}
   );
   gpc1163_5 gpc311 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc312 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc313 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc314 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc315 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc316 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc317 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc318 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc319 (
      {stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc320 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc321 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1406_5 gpc322 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage1_4[0]},
      {stage2_5[0],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc615_5 gpc323 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58]},
      {stage1_2[26]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[1],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc615_5 gpc324 (
      {stage1_1[59], stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63]},
      {stage1_2[27]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[2],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc325 (
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage2_6[0],stage2_5[3],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc326 (
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28]},
      {stage1_4[7]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[1],stage2_5[4],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc327 (
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_4[8]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[2],stage2_5[5],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc328 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[9]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[3],stage2_5[6],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc329 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[10]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[4],stage2_5[7],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc330 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[11]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[5],stage2_5[8],stage2_4[19],stage2_3[19]}
   );
   gpc606_5 gpc331 (
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[5],stage2_6[6],stage2_5[9],stage2_4[20]}
   );
   gpc606_5 gpc332 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[6],stage2_6[7],stage2_5[10],stage2_4[21]}
   );
   gpc606_5 gpc333 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[7],stage2_6[8],stage2_5[11],stage2_4[22]}
   );
   gpc606_5 gpc334 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[8],stage2_6[9],stage2_5[12],stage2_4[23]}
   );
   gpc606_5 gpc335 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[9],stage2_6[10],stage2_5[13],stage2_4[24]}
   );
   gpc606_5 gpc336 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[10],stage2_6[11],stage2_5[14],stage2_4[25]}
   );
   gpc606_5 gpc337 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[11],stage2_6[12],stage2_5[15],stage2_4[26]}
   );
   gpc606_5 gpc338 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[12],stage2_6[13],stage2_5[16],stage2_4[27]}
   );
   gpc207_4 gpc339 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[8],stage2_7[13],stage2_6[14],stage2_5[17]}
   );
   gpc606_5 gpc340 (
      {stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42]},
      {stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage2_9[0],stage2_8[9],stage2_7[14],stage2_6[15],stage2_5[18]}
   );
   gpc606_5 gpc341 (
      {stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48]},
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[10],stage2_7[15],stage2_6[16],stage2_5[19]}
   );
   gpc615_5 gpc342 (
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[2],stage2_8[11],stage2_7[16]}
   );
   gpc615_5 gpc343 (
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[3],stage2_8[12],stage2_7[17]}
   );
   gpc615_5 gpc344 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28]},
      {stage1_8[2]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[2],stage2_9[4],stage2_8[13],stage2_7[18]}
   );
   gpc615_5 gpc345 (
      {stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[3]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[3],stage2_9[5],stage2_8[14],stage2_7[19]}
   );
   gpc615_5 gpc346 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38]},
      {stage1_8[4]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[4],stage2_9[6],stage2_8[15],stage2_7[20]}
   );
   gpc615_5 gpc347 (
      {stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_8[5]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[5],stage2_9[7],stage2_8[16],stage2_7[21]}
   );
   gpc615_5 gpc348 (
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage1_8[6]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[6],stage2_9[8],stage2_8[17],stage2_7[22]}
   );
   gpc615_5 gpc349 (
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_8[7]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[7],stage2_9[9],stage2_8[18],stage2_7[23]}
   );
   gpc615_5 gpc350 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58]},
      {stage1_8[8]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[8],stage2_9[10],stage2_8[19],stage2_7[24]}
   );
   gpc606_5 gpc351 (
      {stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13], stage1_8[14]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[9],stage2_10[9],stage2_9[11],stage2_8[20]}
   );
   gpc606_5 gpc352 (
      {stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[10],stage2_10[10],stage2_9[12],stage2_8[21]}
   );
   gpc606_5 gpc353 (
      {stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[11],stage2_10[11],stage2_9[13],stage2_8[22]}
   );
   gpc606_5 gpc354 (
      {stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[12],stage2_10[12],stage2_9[14],stage2_8[23]}
   );
   gpc606_5 gpc355 (
      {stage1_8[33], stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37], stage1_8[38]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[13],stage2_10[13],stage2_9[15],stage2_8[24]}
   );
   gpc606_5 gpc356 (
      {stage1_8[39], stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43], stage1_8[44]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[14],stage2_10[14],stage2_9[16],stage2_8[25]}
   );
   gpc615_5 gpc357 (
      {stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49]},
      {stage1_9[54]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[15],stage2_10[15],stage2_9[17],stage2_8[26]}
   );
   gpc615_5 gpc358 (
      {stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54]},
      {stage1_9[55]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[16],stage2_10[16],stage2_9[18],stage2_8[27]}
   );
   gpc606_5 gpc359 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[8],stage2_11[17],stage2_10[17]}
   );
   gpc615_5 gpc360 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[1],stage2_12[9],stage2_11[18]}
   );
   gpc615_5 gpc361 (
      {stage1_11[5], stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9]},
      {stage1_12[7]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[2],stage2_13[2],stage2_12[10],stage2_11[19]}
   );
   gpc615_5 gpc362 (
      {stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13], stage1_11[14]},
      {stage1_12[8]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[3],stage2_13[3],stage2_12[11],stage2_11[20]}
   );
   gpc615_5 gpc363 (
      {stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19]},
      {stage1_12[9]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[4],stage2_13[4],stage2_12[12],stage2_11[21]}
   );
   gpc615_5 gpc364 (
      {stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_12[10]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[5],stage2_13[5],stage2_12[13],stage2_11[22]}
   );
   gpc615_5 gpc365 (
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage1_12[11]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[6],stage2_13[6],stage2_12[14],stage2_11[23]}
   );
   gpc615_5 gpc366 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[12]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[7],stage2_13[7],stage2_12[15],stage2_11[24]}
   );
   gpc615_5 gpc367 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[13]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[8],stage2_13[8],stage2_12[16],stage2_11[25]}
   );
   gpc207_4 gpc368 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19], stage1_12[20]},
      {stage1_14[0], stage1_14[1]},
      {stage2_15[8],stage2_14[9],stage2_13[9],stage2_12[17]}
   );
   gpc606_5 gpc369 (
      {stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25], stage1_12[26]},
      {stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage2_16[0],stage2_15[9],stage2_14[10],stage2_13[10],stage2_12[18]}
   );
   gpc606_5 gpc370 (
      {stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31], stage1_12[32]},
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage2_16[1],stage2_15[10],stage2_14[11],stage2_13[11],stage2_12[19]}
   );
   gpc606_5 gpc371 (
      {stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38]},
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18], stage1_14[19]},
      {stage2_16[2],stage2_15[11],stage2_14[12],stage2_13[12],stage2_12[20]}
   );
   gpc606_5 gpc372 (
      {stage1_12[39], stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43], stage1_12[44]},
      {stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage2_16[3],stage2_15[12],stage2_14[13],stage2_13[13],stage2_12[21]}
   );
   gpc606_5 gpc373 (
      {stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49], stage1_12[50]},
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31]},
      {stage2_16[4],stage2_15[13],stage2_14[14],stage2_13[14],stage2_12[22]}
   );
   gpc606_5 gpc374 (
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[5],stage2_15[14],stage2_14[15],stage2_13[15]}
   );
   gpc606_5 gpc375 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[6],stage2_15[15],stage2_14[16],stage2_13[16]}
   );
   gpc606_5 gpc376 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[7],stage2_15[16],stage2_14[17],stage2_13[17]}
   );
   gpc606_5 gpc377 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[8],stage2_15[17],stage2_14[18],stage2_13[18]}
   );
   gpc606_5 gpc378 (
      {stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[4],stage2_16[9],stage2_15[18],stage2_14[19]}
   );
   gpc606_5 gpc379 (
      {stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42], stage1_14[43]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[5],stage2_16[10],stage2_15[19],stage2_14[20]}
   );
   gpc606_5 gpc380 (
      {stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48], stage1_14[49]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[6],stage2_16[11],stage2_15[20],stage2_14[21]}
   );
   gpc615_5 gpc381 (
      {stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_15[24]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[7],stage2_16[12],stage2_15[21],stage2_14[22]}
   );
   gpc615_5 gpc382 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_15[25]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[8],stage2_16[13],stage2_15[22],stage2_14[23]}
   );
   gpc615_5 gpc383 (
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30]},
      {stage1_16[30]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[5],stage2_17[9],stage2_16[14],stage2_15[23]}
   );
   gpc615_5 gpc384 (
      {stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage1_16[31]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[6],stage2_17[10],stage2_16[15],stage2_15[24]}
   );
   gpc1_1 gpc385 (
      {stage1_0[42]},
      {stage2_0[11]}
   );
   gpc1_1 gpc386 (
      {stage1_0[43]},
      {stage2_0[12]}
   );
   gpc1_1 gpc387 (
      {stage1_0[44]},
      {stage2_0[13]}
   );
   gpc1_1 gpc388 (
      {stage1_0[45]},
      {stage2_0[14]}
   );
   gpc1_1 gpc389 (
      {stage1_2[34]},
      {stage2_2[15]}
   );
   gpc1_1 gpc390 (
      {stage1_2[35]},
      {stage2_2[16]}
   );
   gpc1_1 gpc391 (
      {stage1_2[36]},
      {stage2_2[17]}
   );
   gpc1_1 gpc392 (
      {stage1_2[37]},
      {stage2_2[18]}
   );
   gpc1_1 gpc393 (
      {stage1_2[38]},
      {stage2_2[19]}
   );
   gpc1_1 gpc394 (
      {stage1_5[49]},
      {stage2_5[20]}
   );
   gpc1_1 gpc395 (
      {stage1_5[50]},
      {stage2_5[21]}
   );
   gpc1_1 gpc396 (
      {stage1_5[51]},
      {stage2_5[22]}
   );
   gpc1_1 gpc397 (
      {stage1_5[52]},
      {stage2_5[23]}
   );
   gpc1_1 gpc398 (
      {stage1_5[53]},
      {stage2_5[24]}
   );
   gpc1_1 gpc399 (
      {stage1_5[54]},
      {stage2_5[25]}
   );
   gpc1_1 gpc400 (
      {stage1_5[55]},
      {stage2_5[26]}
   );
   gpc1_1 gpc401 (
      {stage1_5[56]},
      {stage2_5[27]}
   );
   gpc1_1 gpc402 (
      {stage1_7[59]},
      {stage2_7[25]}
   );
   gpc1_1 gpc403 (
      {stage1_7[60]},
      {stage2_7[26]}
   );
   gpc1_1 gpc404 (
      {stage1_7[61]},
      {stage2_7[27]}
   );
   gpc1_1 gpc405 (
      {stage1_7[62]},
      {stage2_7[28]}
   );
   gpc1_1 gpc406 (
      {stage1_7[63]},
      {stage2_7[29]}
   );
   gpc1_1 gpc407 (
      {stage1_7[64]},
      {stage2_7[30]}
   );
   gpc1_1 gpc408 (
      {stage1_8[55]},
      {stage2_8[28]}
   );
   gpc1_1 gpc409 (
      {stage1_9[56]},
      {stage2_9[19]}
   );
   gpc1_1 gpc410 (
      {stage1_9[57]},
      {stage2_9[20]}
   );
   gpc1_1 gpc411 (
      {stage1_11[40]},
      {stage2_11[26]}
   );
   gpc1_1 gpc412 (
      {stage1_11[41]},
      {stage2_11[27]}
   );
   gpc1_1 gpc413 (
      {stage1_11[42]},
      {stage2_11[28]}
   );
   gpc1_1 gpc414 (
      {stage1_11[43]},
      {stage2_11[29]}
   );
   gpc1_1 gpc415 (
      {stage1_11[44]},
      {stage2_11[30]}
   );
   gpc1_1 gpc416 (
      {stage1_11[45]},
      {stage2_11[31]}
   );
   gpc1_1 gpc417 (
      {stage1_11[46]},
      {stage2_11[32]}
   );
   gpc1_1 gpc418 (
      {stage1_11[47]},
      {stage2_11[33]}
   );
   gpc1_1 gpc419 (
      {stage1_11[48]},
      {stage2_11[34]}
   );
   gpc1_1 gpc420 (
      {stage1_11[49]},
      {stage2_11[35]}
   );
   gpc1_1 gpc421 (
      {stage1_11[50]},
      {stage2_11[36]}
   );
   gpc1_1 gpc422 (
      {stage1_11[51]},
      {stage2_11[37]}
   );
   gpc1_1 gpc423 (
      {stage1_12[51]},
      {stage2_12[23]}
   );
   gpc1_1 gpc424 (
      {stage1_12[52]},
      {stage2_12[24]}
   );
   gpc1_1 gpc425 (
      {stage1_12[53]},
      {stage2_12[25]}
   );
   gpc1_1 gpc426 (
      {stage1_12[54]},
      {stage2_12[26]}
   );
   gpc1_1 gpc427 (
      {stage1_12[55]},
      {stage2_12[27]}
   );
   gpc1_1 gpc428 (
      {stage1_12[56]},
      {stage2_12[28]}
   );
   gpc1_1 gpc429 (
      {stage1_14[60]},
      {stage2_14[24]}
   );
   gpc1_1 gpc430 (
      {stage1_14[61]},
      {stage2_14[25]}
   );
   gpc1_1 gpc431 (
      {stage1_14[62]},
      {stage2_14[26]}
   );
   gpc1_1 gpc432 (
      {stage1_14[63]},
      {stage2_14[27]}
   );
   gpc1_1 gpc433 (
      {stage1_14[64]},
      {stage2_14[28]}
   );
   gpc1_1 gpc434 (
      {stage1_14[65]},
      {stage2_14[29]}
   );
   gpc1_1 gpc435 (
      {stage1_14[66]},
      {stage2_14[30]}
   );
   gpc1_1 gpc436 (
      {stage1_14[67]},
      {stage2_14[31]}
   );
   gpc1_1 gpc437 (
      {stage1_14[68]},
      {stage2_14[32]}
   );
   gpc1_1 gpc438 (
      {stage1_14[69]},
      {stage2_14[33]}
   );
   gpc1_1 gpc439 (
      {stage1_14[70]},
      {stage2_14[34]}
   );
   gpc1_1 gpc440 (
      {stage1_15[36]},
      {stage2_15[25]}
   );
   gpc1_1 gpc441 (
      {stage1_15[37]},
      {stage2_15[26]}
   );
   gpc1_1 gpc442 (
      {stage1_16[32]},
      {stage2_16[16]}
   );
   gpc1_1 gpc443 (
      {stage1_16[33]},
      {stage2_16[17]}
   );
   gpc1_1 gpc444 (
      {stage1_16[34]},
      {stage2_16[18]}
   );
   gpc1_1 gpc445 (
      {stage1_16[35]},
      {stage2_16[19]}
   );
   gpc1_1 gpc446 (
      {stage1_17[12]},
      {stage2_17[11]}
   );
   gpc1_1 gpc447 (
      {stage1_17[13]},
      {stage2_17[12]}
   );
   gpc1_1 gpc448 (
      {stage1_17[14]},
      {stage2_17[13]}
   );
   gpc1_1 gpc449 (
      {stage1_17[15]},
      {stage2_17[14]}
   );
   gpc1_1 gpc450 (
      {stage1_17[16]},
      {stage2_17[15]}
   );
   gpc1_1 gpc451 (
      {stage1_17[17]},
      {stage2_17[16]}
   );
   gpc1_1 gpc452 (
      {stage1_17[18]},
      {stage2_17[17]}
   );
   gpc1_1 gpc453 (
      {stage1_17[19]},
      {stage2_17[18]}
   );
   gpc1_1 gpc454 (
      {stage1_17[20]},
      {stage2_17[19]}
   );
   gpc606_5 gpc455 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc615_5 gpc456 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc615_5 gpc457 (
      {stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9]},
      {stage2_3[7]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc1163_5 gpc458 (
      {stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[3]}
   );
   gpc1163_5 gpc459 (
      {stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage2_5[1]},
      {stage2_6[1]},
      {stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4],stage3_3[4]}
   );
   gpc606_5 gpc460 (
      {stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[2],stage3_6[4],stage3_5[5]}
   );
   gpc615_5 gpc461 (
      {stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12]},
      {stage2_6[2]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[1],stage3_7[3],stage3_6[5],stage3_5[6]}
   );
   gpc615_5 gpc462 (
      {stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_6[3]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[2],stage3_7[4],stage3_6[6],stage3_5[7]}
   );
   gpc615_5 gpc463 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22]},
      {stage2_6[4]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[3],stage3_7[5],stage3_6[7],stage3_5[8]}
   );
   gpc615_5 gpc464 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27]},
      {stage2_6[5]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[4],stage3_7[6],stage3_6[8],stage3_5[9]}
   );
   gpc606_5 gpc465 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[5],stage3_8[5],stage3_7[7],stage3_6[9]}
   );
   gpc615_5 gpc466 (
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16]},
      {stage2_7[30]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[6],stage3_8[6],stage3_7[8],stage3_6[10]}
   );
   gpc606_5 gpc467 (
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[2],stage3_9[7],stage3_8[7]}
   );
   gpc606_5 gpc468 (
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[1],stage3_10[3],stage3_9[8],stage3_8[8]}
   );
   gpc1163_5 gpc469 (
      {stage2_9[0], stage2_9[1], stage2_9[2]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage2_11[0]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[2],stage3_11[2],stage3_10[4],stage3_9[9]}
   );
   gpc606_5 gpc470 (
      {stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6], stage2_9[7], stage2_9[8]},
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage3_13[1],stage3_12[3],stage3_11[3],stage3_10[5],stage3_9[10]}
   );
   gpc606_5 gpc471 (
      {stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12]},
      {stage3_13[2],stage3_12[4],stage3_11[4],stage3_10[6],stage3_9[11]}
   );
   gpc606_5 gpc472 (
      {stage2_9[15], stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18]},
      {stage3_13[3],stage3_12[5],stage3_11[5],stage3_10[7],stage3_9[12]}
   );
   gpc615_5 gpc473 (
      {stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage2_12[1]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[4],stage3_12[6],stage3_11[6]}
   );
   gpc615_5 gpc474 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28]},
      {stage2_12[2]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[5],stage3_12[7],stage3_11[7]}
   );
   gpc606_5 gpc475 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[2],stage3_13[6],stage3_12[8]}
   );
   gpc606_5 gpc476 (
      {stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[3],stage3_14[3],stage3_13[7],stage3_12[9]}
   );
   gpc606_5 gpc477 (
      {stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[4],stage3_14[4],stage3_13[8],stage3_12[10]}
   );
   gpc606_5 gpc478 (
      {stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[5],stage3_14[5],stage3_13[9],stage3_12[11]}
   );
   gpc606_5 gpc479 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[6],stage3_14[6],stage3_13[10]}
   );
   gpc1163_5 gpc480 (
      {stage2_14[24], stage2_14[25], stage2_14[26]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage2_16[0]},
      {stage2_17[0]},
      {stage3_18[0],stage3_17[1],stage3_16[5],stage3_15[7],stage3_14[7]}
   );
   gpc615_5 gpc481 (
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16]},
      {stage2_16[1]},
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage3_19[0],stage3_18[1],stage3_17[2],stage3_16[6],stage3_15[8]}
   );
   gpc615_5 gpc482 (
      {stage2_15[17], stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21]},
      {stage2_16[2]},
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage3_19[1],stage3_18[2],stage3_17[3],stage3_16[7],stage3_15[9]}
   );
   gpc615_5 gpc483 (
      {stage2_15[22], stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26]},
      {stage2_16[3]},
      {stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18]},
      {stage3_19[2],stage3_18[3],stage3_17[4],stage3_16[8],stage3_15[10]}
   );
   gpc606_5 gpc484 (
      {stage2_16[4], stage2_16[5], stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[3],stage3_18[4],stage3_17[5],stage3_16[9]}
   );
   gpc1_1 gpc485 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc486 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc487 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc488 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc489 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc490 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc491 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc492 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc493 (
      {stage2_0[8]},
      {stage3_0[8]}
   );
   gpc1_1 gpc494 (
      {stage2_0[9]},
      {stage3_0[9]}
   );
   gpc1_1 gpc495 (
      {stage2_0[10]},
      {stage3_0[10]}
   );
   gpc1_1 gpc496 (
      {stage2_0[11]},
      {stage3_0[11]}
   );
   gpc1_1 gpc497 (
      {stage2_0[12]},
      {stage3_0[12]}
   );
   gpc1_1 gpc498 (
      {stage2_0[13]},
      {stage3_0[13]}
   );
   gpc1_1 gpc499 (
      {stage2_0[14]},
      {stage3_0[14]}
   );
   gpc1_1 gpc500 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc501 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc502 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc503 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc504 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc505 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc506 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc507 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc508 (
      {stage2_2[10]},
      {stage3_2[3]}
   );
   gpc1_1 gpc509 (
      {stage2_2[11]},
      {stage3_2[4]}
   );
   gpc1_1 gpc510 (
      {stage2_2[12]},
      {stage3_2[5]}
   );
   gpc1_1 gpc511 (
      {stage2_2[13]},
      {stage3_2[6]}
   );
   gpc1_1 gpc512 (
      {stage2_2[14]},
      {stage3_2[7]}
   );
   gpc1_1 gpc513 (
      {stage2_2[15]},
      {stage3_2[8]}
   );
   gpc1_1 gpc514 (
      {stage2_2[16]},
      {stage3_2[9]}
   );
   gpc1_1 gpc515 (
      {stage2_2[17]},
      {stage3_2[10]}
   );
   gpc1_1 gpc516 (
      {stage2_2[18]},
      {stage3_2[11]}
   );
   gpc1_1 gpc517 (
      {stage2_2[19]},
      {stage3_2[12]}
   );
   gpc1_1 gpc518 (
      {stage2_3[14]},
      {stage3_3[5]}
   );
   gpc1_1 gpc519 (
      {stage2_3[15]},
      {stage3_3[6]}
   );
   gpc1_1 gpc520 (
      {stage2_3[16]},
      {stage3_3[7]}
   );
   gpc1_1 gpc521 (
      {stage2_3[17]},
      {stage3_3[8]}
   );
   gpc1_1 gpc522 (
      {stage2_3[18]},
      {stage3_3[9]}
   );
   gpc1_1 gpc523 (
      {stage2_3[19]},
      {stage3_3[10]}
   );
   gpc1_1 gpc524 (
      {stage2_4[24]},
      {stage3_4[5]}
   );
   gpc1_1 gpc525 (
      {stage2_4[25]},
      {stage3_4[6]}
   );
   gpc1_1 gpc526 (
      {stage2_4[26]},
      {stage3_4[7]}
   );
   gpc1_1 gpc527 (
      {stage2_4[27]},
      {stage3_4[8]}
   );
   gpc1_1 gpc528 (
      {stage2_8[24]},
      {stage3_8[9]}
   );
   gpc1_1 gpc529 (
      {stage2_8[25]},
      {stage3_8[10]}
   );
   gpc1_1 gpc530 (
      {stage2_8[26]},
      {stage3_8[11]}
   );
   gpc1_1 gpc531 (
      {stage2_8[27]},
      {stage3_8[12]}
   );
   gpc1_1 gpc532 (
      {stage2_8[28]},
      {stage3_8[13]}
   );
   gpc1_1 gpc533 (
      {stage2_11[29]},
      {stage3_11[8]}
   );
   gpc1_1 gpc534 (
      {stage2_11[30]},
      {stage3_11[9]}
   );
   gpc1_1 gpc535 (
      {stage2_11[31]},
      {stage3_11[10]}
   );
   gpc1_1 gpc536 (
      {stage2_11[32]},
      {stage3_11[11]}
   );
   gpc1_1 gpc537 (
      {stage2_11[33]},
      {stage3_11[12]}
   );
   gpc1_1 gpc538 (
      {stage2_11[34]},
      {stage3_11[13]}
   );
   gpc1_1 gpc539 (
      {stage2_11[35]},
      {stage3_11[14]}
   );
   gpc1_1 gpc540 (
      {stage2_11[36]},
      {stage3_11[15]}
   );
   gpc1_1 gpc541 (
      {stage2_11[37]},
      {stage3_11[16]}
   );
   gpc1_1 gpc542 (
      {stage2_12[27]},
      {stage3_12[12]}
   );
   gpc1_1 gpc543 (
      {stage2_12[28]},
      {stage3_12[13]}
   );
   gpc1_1 gpc544 (
      {stage2_13[18]},
      {stage3_13[11]}
   );
   gpc1_1 gpc545 (
      {stage2_14[27]},
      {stage3_14[8]}
   );
   gpc1_1 gpc546 (
      {stage2_14[28]},
      {stage3_14[9]}
   );
   gpc1_1 gpc547 (
      {stage2_14[29]},
      {stage3_14[10]}
   );
   gpc1_1 gpc548 (
      {stage2_14[30]},
      {stage3_14[11]}
   );
   gpc1_1 gpc549 (
      {stage2_14[31]},
      {stage3_14[12]}
   );
   gpc1_1 gpc550 (
      {stage2_14[32]},
      {stage3_14[13]}
   );
   gpc1_1 gpc551 (
      {stage2_14[33]},
      {stage3_14[14]}
   );
   gpc1_1 gpc552 (
      {stage2_14[34]},
      {stage3_14[15]}
   );
   gpc1_1 gpc553 (
      {stage2_16[10]},
      {stage3_16[10]}
   );
   gpc1_1 gpc554 (
      {stage2_16[11]},
      {stage3_16[11]}
   );
   gpc1_1 gpc555 (
      {stage2_16[12]},
      {stage3_16[12]}
   );
   gpc1_1 gpc556 (
      {stage2_16[13]},
      {stage3_16[13]}
   );
   gpc1_1 gpc557 (
      {stage2_16[14]},
      {stage3_16[14]}
   );
   gpc1_1 gpc558 (
      {stage2_16[15]},
      {stage3_16[15]}
   );
   gpc1_1 gpc559 (
      {stage2_16[16]},
      {stage3_16[16]}
   );
   gpc1_1 gpc560 (
      {stage2_16[17]},
      {stage3_16[17]}
   );
   gpc1_1 gpc561 (
      {stage2_16[18]},
      {stage3_16[18]}
   );
   gpc1_1 gpc562 (
      {stage2_16[19]},
      {stage3_16[19]}
   );
   gpc1_1 gpc563 (
      {stage2_17[19]},
      {stage3_17[6]}
   );
   gpc1_1 gpc564 (
      {stage2_18[6]},
      {stage3_18[5]}
   );
   gpc1_1 gpc565 (
      {stage2_19[0]},
      {stage3_19[4]}
   );
   gpc1_1 gpc566 (
      {stage2_19[1]},
      {stage3_19[5]}
   );
   gpc606_5 gpc567 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc568 (
      {stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9], stage3_0[10]},
      {stage3_1[0]},
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc1163_5 gpc569 (
      {stage3_3[0], stage3_3[1], stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_5[0]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2]}
   );
   gpc606_5 gpc570 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc615_5 gpc571 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[2],stage4_6[2]}
   );
   gpc615_5 gpc572 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[7]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[2],stage4_7[3],stage4_6[3]}
   );
   gpc606_5 gpc573 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[2],stage4_9[3]}
   );
   gpc615_5 gpc574 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10]},
      {stage3_10[0]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[1],stage4_10[3],stage4_9[4]}
   );
   gpc606_5 gpc575 (
      {stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[2],stage4_11[2],stage4_10[4]}
   );
   gpc615_5 gpc576 (
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16]},
      {stage3_12[6]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[1],stage4_13[3],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc577 (
      {stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11], stage3_12[12]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[2],stage4_13[4],stage4_12[4]}
   );
   gpc606_5 gpc578 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[3],stage4_13[5]}
   );
   gpc615_5 gpc579 (
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage3_15[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[1],stage4_16[2],stage4_15[3],stage4_14[4]}
   );
   gpc615_5 gpc580 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[7]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[2],stage4_16[3],stage4_15[4],stage4_14[5]}
   );
   gpc606_5 gpc581 (
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[2],stage4_17[3],stage4_16[4]}
   );
   gpc606_5 gpc582 (
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[1],stage4_19[1],stage4_18[3],stage4_17[4]}
   );
   gpc1_1 gpc583 (
      {stage3_0[11]},
      {stage4_0[2]}
   );
   gpc1_1 gpc584 (
      {stage3_0[12]},
      {stage4_0[3]}
   );
   gpc1_1 gpc585 (
      {stage3_0[13]},
      {stage4_0[4]}
   );
   gpc1_1 gpc586 (
      {stage3_0[14]},
      {stage4_0[5]}
   );
   gpc1_1 gpc587 (
      {stage3_1[1]},
      {stage4_1[2]}
   );
   gpc1_1 gpc588 (
      {stage3_1[2]},
      {stage4_1[3]}
   );
   gpc1_1 gpc589 (
      {stage3_1[3]},
      {stage4_1[4]}
   );
   gpc1_1 gpc590 (
      {stage3_1[4]},
      {stage4_1[5]}
   );
   gpc1_1 gpc591 (
      {stage3_1[5]},
      {stage4_1[6]}
   );
   gpc1_1 gpc592 (
      {stage3_1[6]},
      {stage4_1[7]}
   );
   gpc1_1 gpc593 (
      {stage3_1[7]},
      {stage4_1[8]}
   );
   gpc1_1 gpc594 (
      {stage3_1[8]},
      {stage4_1[9]}
   );
   gpc1_1 gpc595 (
      {stage3_2[12]},
      {stage4_2[2]}
   );
   gpc1_1 gpc596 (
      {stage3_3[3]},
      {stage4_3[3]}
   );
   gpc1_1 gpc597 (
      {stage3_3[4]},
      {stage4_3[4]}
   );
   gpc1_1 gpc598 (
      {stage3_3[5]},
      {stage4_3[5]}
   );
   gpc1_1 gpc599 (
      {stage3_3[6]},
      {stage4_3[6]}
   );
   gpc1_1 gpc600 (
      {stage3_3[7]},
      {stage4_3[7]}
   );
   gpc1_1 gpc601 (
      {stage3_3[8]},
      {stage4_3[8]}
   );
   gpc1_1 gpc602 (
      {stage3_3[9]},
      {stage4_3[9]}
   );
   gpc1_1 gpc603 (
      {stage3_3[10]},
      {stage4_3[10]}
   );
   gpc1_1 gpc604 (
      {stage3_4[6]},
      {stage4_4[3]}
   );
   gpc1_1 gpc605 (
      {stage3_4[7]},
      {stage4_4[4]}
   );
   gpc1_1 gpc606 (
      {stage3_4[8]},
      {stage4_4[5]}
   );
   gpc1_1 gpc607 (
      {stage3_5[7]},
      {stage4_5[2]}
   );
   gpc1_1 gpc608 (
      {stage3_5[8]},
      {stage4_5[3]}
   );
   gpc1_1 gpc609 (
      {stage3_5[9]},
      {stage4_5[4]}
   );
   gpc1_1 gpc610 (
      {stage3_7[8]},
      {stage4_7[4]}
   );
   gpc1_1 gpc611 (
      {stage3_8[12]},
      {stage4_8[3]}
   );
   gpc1_1 gpc612 (
      {stage3_8[13]},
      {stage4_8[4]}
   );
   gpc1_1 gpc613 (
      {stage3_9[11]},
      {stage4_9[5]}
   );
   gpc1_1 gpc614 (
      {stage3_9[12]},
      {stage4_9[6]}
   );
   gpc1_1 gpc615 (
      {stage3_10[7]},
      {stage4_10[5]}
   );
   gpc1_1 gpc616 (
      {stage3_12[13]},
      {stage4_12[5]}
   );
   gpc1_1 gpc617 (
      {stage3_15[8]},
      {stage4_15[5]}
   );
   gpc1_1 gpc618 (
      {stage3_15[9]},
      {stage4_15[6]}
   );
   gpc1_1 gpc619 (
      {stage3_15[10]},
      {stage4_15[7]}
   );
   gpc1_1 gpc620 (
      {stage3_16[18]},
      {stage4_16[5]}
   );
   gpc1_1 gpc621 (
      {stage3_16[19]},
      {stage4_16[6]}
   );
   gpc1_1 gpc622 (
      {stage3_17[6]},
      {stage4_17[5]}
   );
   gpc1_1 gpc623 (
      {stage3_20[0]},
      {stage4_20[2]}
   );
   gpc2135_5 gpc624 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc1415_5 gpc625 (
      {stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6], stage4_1[7]},
      {stage4_2[1]},
      {stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage4_4[0]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1415_5 gpc626 (
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[0]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[1],stage5_4[2]}
   );
   gpc615_5 gpc627 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[0],stage5_8[1]}
   );
   gpc606_5 gpc628 (
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[1]}
   );
   gpc135_4 gpc629 (
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1]}
   );
   gpc1343_5 gpc630 (
      {stage4_18[0], stage4_18[1], stage4_18[2]},
      {stage4_19[0], stage4_19[1], 1'b0, 1'b0},
      {stage4_20[0], stage4_20[1], stage4_20[2]},
      {stage4_21[0]},
      {stage5_22[0],stage5_21[0],stage5_20[0],stage5_19[0],stage5_18[1]}
   );
   gpc1_1 gpc631 (
      {stage4_0[5]},
      {stage5_0[1]}
   );
   gpc1_1 gpc632 (
      {stage4_1[8]},
      {stage5_1[2]}
   );
   gpc1_1 gpc633 (
      {stage4_1[9]},
      {stage5_1[3]}
   );
   gpc1_1 gpc634 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc635 (
      {stage4_3[6]},
      {stage5_3[2]}
   );
   gpc1_1 gpc636 (
      {stage4_3[7]},
      {stage5_3[3]}
   );
   gpc1_1 gpc637 (
      {stage4_3[8]},
      {stage5_3[4]}
   );
   gpc1_1 gpc638 (
      {stage4_3[9]},
      {stage5_3[5]}
   );
   gpc1_1 gpc639 (
      {stage4_3[10]},
      {stage5_3[6]}
   );
   gpc1_1 gpc640 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc641 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc642 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc643 (
      {stage4_5[4]},
      {stage5_5[5]}
   );
   gpc1_1 gpc644 (
      {stage4_7[1]},
      {stage5_7[1]}
   );
   gpc1_1 gpc645 (
      {stage4_7[2]},
      {stage5_7[2]}
   );
   gpc1_1 gpc646 (
      {stage4_7[3]},
      {stage5_7[3]}
   );
   gpc1_1 gpc647 (
      {stage4_7[4]},
      {stage5_7[4]}
   );
   gpc1_1 gpc648 (
      {stage4_9[1]},
      {stage5_9[1]}
   );
   gpc1_1 gpc649 (
      {stage4_9[2]},
      {stage5_9[2]}
   );
   gpc1_1 gpc650 (
      {stage4_9[3]},
      {stage5_9[3]}
   );
   gpc1_1 gpc651 (
      {stage4_9[4]},
      {stage5_9[4]}
   );
   gpc1_1 gpc652 (
      {stage4_9[5]},
      {stage5_9[5]}
   );
   gpc1_1 gpc653 (
      {stage4_9[6]},
      {stage5_9[6]}
   );
   gpc1_1 gpc654 (
      {stage4_11[0]},
      {stage5_11[1]}
   );
   gpc1_1 gpc655 (
      {stage4_11[1]},
      {stage5_11[2]}
   );
   gpc1_1 gpc656 (
      {stage4_11[2]},
      {stage5_11[3]}
   );
   gpc1_1 gpc657 (
      {stage4_11[3]},
      {stage5_11[4]}
   );
   gpc1_1 gpc658 (
      {stage4_13[0]},
      {stage5_13[1]}
   );
   gpc1_1 gpc659 (
      {stage4_13[1]},
      {stage5_13[2]}
   );
   gpc1_1 gpc660 (
      {stage4_13[2]},
      {stage5_13[3]}
   );
   gpc1_1 gpc661 (
      {stage4_13[3]},
      {stage5_13[4]}
   );
   gpc1_1 gpc662 (
      {stage4_13[4]},
      {stage5_13[5]}
   );
   gpc1_1 gpc663 (
      {stage4_13[5]},
      {stage5_13[6]}
   );
   gpc1_1 gpc664 (
      {stage4_15[5]},
      {stage5_15[2]}
   );
   gpc1_1 gpc665 (
      {stage4_15[6]},
      {stage5_15[3]}
   );
   gpc1_1 gpc666 (
      {stage4_15[7]},
      {stage5_15[4]}
   );
   gpc1_1 gpc667 (
      {stage4_16[3]},
      {stage5_16[2]}
   );
   gpc1_1 gpc668 (
      {stage4_16[4]},
      {stage5_16[3]}
   );
   gpc1_1 gpc669 (
      {stage4_16[5]},
      {stage5_16[4]}
   );
   gpc1_1 gpc670 (
      {stage4_16[6]},
      {stage5_16[5]}
   );
   gpc1_1 gpc671 (
      {stage4_17[1]},
      {stage5_17[1]}
   );
   gpc1_1 gpc672 (
      {stage4_17[2]},
      {stage5_17[2]}
   );
   gpc1_1 gpc673 (
      {stage4_17[3]},
      {stage5_17[3]}
   );
   gpc1_1 gpc674 (
      {stage4_17[4]},
      {stage5_17[4]}
   );
   gpc1_1 gpc675 (
      {stage4_17[5]},
      {stage5_17[5]}
   );
   gpc1_1 gpc676 (
      {stage4_18[3]},
      {stage5_18[2]}
   );
   gpc2223_5 gpc677 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1]},
      {stage5_3[0], stage5_3[1]},
      {stage5_4[0], stage5_4[1]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc615_5 gpc678 (
      {stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5], stage5_3[6]},
      {stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc615_5 gpc679 (
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4]},
      {stage5_8[0]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1]}
   );
   gpc615_5 gpc680 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4]},
      {stage5_12[0]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1]}
   );
   gpc615_5 gpc681 (
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4]},
      {stage5_16[0]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage6_19[0],stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1]}
   );
   gpc1415_5 gpc682 (
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {1'b0},
      {stage5_18[0], stage5_18[1], stage5_18[2], 1'b0},
      {stage5_19[0]},
      {stage6_20[0],stage6_19[1],stage6_18[1],stage6_17[1],stage6_16[1]}
   );
   gpc1_1 gpc683 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc684 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc685 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc686 (
      {stage5_2[2]},
      {stage6_2[1]}
   );
   gpc1_1 gpc687 (
      {stage5_6[0]},
      {stage6_6[1]}
   );
   gpc1_1 gpc688 (
      {stage5_8[1]},
      {stage6_8[1]}
   );
   gpc1_1 gpc689 (
      {stage5_9[6]},
      {stage6_9[1]}
   );
   gpc1_1 gpc690 (
      {stage5_10[0]},
      {stage6_10[1]}
   );
   gpc1_1 gpc691 (
      {stage5_12[1]},
      {stage6_12[1]}
   );
   gpc1_1 gpc692 (
      {stage5_13[6]},
      {stage6_13[1]}
   );
   gpc1_1 gpc693 (
      {stage5_14[0]},
      {stage6_14[1]}
   );
   gpc1_1 gpc694 (
      {stage5_20[0]},
      {stage6_20[1]}
   );
   gpc1_1 gpc695 (
      {stage5_21[0]},
      {stage6_21[0]}
   );
   gpc1_1 gpc696 (
      {stage5_22[0]},
      {stage6_22[0]}
   );
endmodule

module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [22:0] srcsum;
    wire [22:0] dstsum;
    wire test;
    compressor_CLA128_16 compressor_CLA128_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h32f659af754e888f9268cedb7f8f04754edcd6d05ba1ddc9050037b1341c80f1e8b5d3cf60cd79eeffeeeda276ad2678a1edd859f20547d43e954a6fd3051ee634a14f7e6c7ba1f6108b539c5f5321106c4c3f74b111084207d9695fbbf2bedf095854b6ee5b18386b82527492e66d2b3b5d58e98cb9a7da7dc15077e90fd712e0f9682dba0ed318cca693ebcd22db884ab285e9fd9b7cc8f6a99a43e1d4025a47503c5ddf9e6e2a5e1d38eff558d208920823e53b09cbdc5204d952a29f24b176f1037a719cab038b6c2c50619e9ea190d70767198b3316b39a9d0109618dc834a283310fc1f1db4f839a795adfcd076a8b95bd0c8ca7134fa71750609e7323;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h11e62edc525b53c8c91db0934b67b65b052347648861f6137520a22f7c31f788b298e4c6fd564643eb8285a222e1eeeeec5a420e71d8125f6e98aacfb111c39256df0999870f06b3fabaea52ccd99419879ae0a6dd739c18d02b88d25541d61da6acc12074e541f346dc15e9d9d59b20cc1a19eca448ec826ba33f32a9eafa4aeecc97bc04ca81612b8ffa4aa8aeae3060ab378acb4cc376f359739a2428f75bd78f98ee7f5d350442050d538afc8e9d4888ece586c56493e6ee64266c210808bb68670bf0c5497be15ec01d8ec21069b5c0787e1ad97fe33a653b74bc77578eb450661a86edf156e2d0cbb18fb6ec9676a99927b380c9e08c0e22fbf2db8c4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4431e54224cc740dabb82fb382feb0c1a66f8a51e85317352e1b1f6894d2c631569439ee4d915d75a347717cd7bef6e2a2e377750c7a911e33dd1dd76c228751e5a2c0969f7eebe7eaff6a47af34bbca43f88d8024ea1b8608001201e82c69a60df307681d094d1578f163ec5c5825e3b00080daef707666f3e7b7bfc8a2eaba8e4b343c930681cd5fee3bc3f03da5c0d900208027b2bbdaedc598ed2e59e827df6da169902a1683c495b54cc6b7591118db91ece6288c2fc5655dc9ae52aa7ff4ee7453b6f76777d54451aa1f7dd11a046504b326f0db7d587ff71d04df0aa22edd81d8547a0fed7899d761a10c2572ef98cdcfac9cf171dc3d23783024fc2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha20f5ce8273e3285913216b3da21436eb8bb4a7704214d717c090f4e94f4bb3e79398b30ee98d01f10448ef425f522372191382f9b045b41f201127b0f047ca058a5cb0aad0fa21b161602f5a714fa66a7e56d7a1a4060d08b941858741e0e9c8ff65c7c9cab64331e9debdf150ef805b96159548bf34d8a72a79596c880e9b91d92061406e0a71c4a1a0463eebdeddfeac6bc32e28a454056b1ed256b9c4a7e336b27872360614d0927cad3166008d50eba0ef2d06fc8033a6dc95bc0dbb0052d4e80904bace3ce808c3b26140a9fe72d151c05ea750add2c16f7ac34978c1f3b47ef722c2faee35968e7e6cf920797ffcb65aab0f7f32feaf8c3f0489d76ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3f1e7b59b3c6067ec9941e214cac7292b121c1ec6c3e1c9097309029c03c4fbfe936d50c5414315cacab999e7384d27a493c4d5d1b682de26d7472770d4cef11efeee806975ab90f6b8164a3815959a0ffbe58c26abaabf0ca72b3c7ef1ed2545fd0f4472bad390e6bf09b342dd6d23ac1922a54660267c46f34a2dfb8d1e2ed59f479a0b39fb3414651d1731c5f304cf34d722354a839b8af5d791478a9997d1d607c84b3e268bc0b8134175983b030a291f7a4ac3793658c50770ff2ded28f4c591abd8fd5e95fba2a9494719eaae27b0a47ea143ffa2447904ec4b5ff54c930a6c9d51bc68f3865c5b273b50fa9464bc2abf94962bedfdf78c7850ed5b305;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h57c69f3511ce43494590510596565b0a5e558bebbc5170d94d7344ef8365d74fcea8ff97c8770d4a47bbb2de49871d9e0c6609c085e67acb3f5dd87728934dadc642bb6056959201dc634f519e826c90c6c573344903769179a4408ff9f5e15f88304db3dc64333ab4725f7fa06794b3514dbb8d5da07e6e708d436f36b589137c9a5a387a97abaa8fb00551c8f32447a9195b2afe8f27604646a07e9132150e4ca5cd91e2054f5e09f573b707fc0e897a4e57184bd03a4affbc343a0b69a98d253e1cf64496dd465864fa81d6cb4e0ab68ea957d858ef218065ced3104b056a90e55e8682a980e00ffb02df5e974c018c2c65248f860830591d71471aef5e42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h242c4d3218bf0006f901116be950ebeefa63a2de20a7834fd0fd9fc36c4534cecaaf0c396055760b69eececbd006b52f9c3a417f1a9bd911ee4889f96c9dacf5d0c05bf1e3b7fb7ff56a79314cf1fa3c009b0c56b99873945ce2d745cac5853af7ea883942cc0b8432e58c971dc8589d556978af1695661ea2acf16ad7b08d6591689bcd72ab6ff9076f01eac3228e46e4ed7c3a8de81a4f77864df8d91803d299f17095b084be73c941653a90411a5e2fcd108476ae3ef6b614fa67d57630555fc5fb13c37b51e9a00ec18ac89226243dc02484158b40abdf42c490e8f07357d6c80c1a2ec2673bd882f7d16ca57b985d400552b475efb96ce8302c87d04760;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hca4babe972a5c867462d66aaa39f9e15ea398e1749b4606e74d5f41ca604918e19a81638e7f2b438af036d9f3926977553c4a754346d2d964f7ef98a622aea110fdd1ca3091070674051ce0d926eb661644358faae02cfd6afc5b7d794076e37328a60ebd9f0ae4196f3daeb3e676d942969eb75756ae4e9e6267700950b2eaf7dc5b514b12e9f4f0139c1629f45fbdf9ecd3e639288e7c5a93865a1543c9e44024f37e61109fa1ad8c87c4eab91a964ead211a49eb5efa2e20b716d6aa35f83ef3c3bbb1683c33287f9684e88340a2cb5984dbbc42e1731d02ab4ad30bff244dacaea0a69571f0a3c6d1d113d3e78f828c155aeb6afa5f18da4f15b1e00bea2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc14908002c0d7761d4eaa6d9e2f93be9c67f4510d8f9cad56b5c0c5bbc342dbe369b15640b9c95b2c67b46e72f48ab3ef689e21bce101458e41ff2b9eb9ccfb380db2ae7ec3e14f367d717cfe03a7f4a8737fe60c11329cddefb00f4b98a9c47ce2ec59ea10441aeb711d7d0b2ab560b51d0cb72f1d6052da8b00d47bb6e2c2ca38e7a5d107f1ff2b0934df2eccf6a171a4a7b4355e6029fa1fe7c89fe743df4b5be1ea7839046eff6cea07c533653a19cc0b1f0be125394603823bbea87eef182cdb1a69ed8618209cc0bb6bed9ecc87e5310fcf4b151140c3112298c909e86f8634afc5ee05b68416b40931a8ccdace9d91c196e199e7c2eefdd6019a2d59f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc7ae7593d3074a201368ceb0d9f2c2cbdd8def1cd429a069d0e986a06c022c65b06b3a577544eb74d7be86fc3067fda137da6017286a5644fdf775b20cac07c8f758f66b2bcabf7e8837436ad10294720b6f255fa1887e19ff8b4133400817a51839c472b79abb7e258850ba45b3761cf53ad94270c0de063d7b44a75fd1cdda6d04de2750d3cff9f1aa50bc83cd5e383f7fc6eff57aa49a549eee9863dff56f60b0d54ba15a94da848c299d4a8f549760f9d0ee78edabfd400d44b8e4c0e5687ed254d35213c35afb76f02f8a5435de912e5a3ef616c7774fdda704375127fa9df883062204941c7436f9867664b251a7f75e9a6bb2dbb05126144ddb386a56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hdb230a007bfcf56e27ae85330a358a8089d0332e3ee154f1f8bb1dc78f7a427c6ca81c3caf7c4d21e782f1d0dead6d4dff52aec21948d4f2efd65ad0a16346e6587cb4c9f9273a2610beaf421a54c4739492d911d932c5b6f8f00653f323c8c35195f95f4fb490452274b9dda9f6edf50d8f3423fa488fef55842233cfe4d1b93597473c53687c2c4fa774bff4ab6b713a83ed0a79dd1c1433cb484a88f051123b8772f1d957f11853fbe9ad42289ba5ba4424aed880dbe7d13a128aa7ebbfb28f39d299f81c8ba1eabd7b4b55a7afcf345e779397460b332e2b420f9b2061d006cb471395959437bd03025c88340b8491ae198f0de77402e6e0c472bb4a2ddb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd7cf0ba5fac9467df493c1550338b781c9e7c9137f83cf2e7d13317b935237c072d221b175410047b0887df87d0940b2f5ad266d1f5421c7d1b0be049b7a65db2e88286e025742b3438dd391deb0e07674db875fd7186ff5a9f5d2d525e2e35910bb3c27929e9c2f0af9c897ebab41e0d9f7f411eecf1de99ca28ff0c0d12accca6f4a652d96df42553b8779a1ef4699cf07dbfa958c9fc0038ae4fbc4a030c9246ad24fa979e2ac3bb7265332df956d33d9db19c2676325df51b54b401b64e41b2ea0fbc97aceba688932700b89688f6f39eb7c522599341679aa99be9cc88d053df3d78b5cfd2b7bd4d6ae9951d2101a9148ffa2f799ba3cc199fec59d69f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h481fc18728f2eb7e65896dafc5c261f7697cca5acacbfc984d6da6ca9e91e382070bf2e9d177e3b3432c254f45cd9a297994d41b88674df504a0a6992cc0604f67faf65d82c71ba02ffdb4b8c5f7ac7fdfd89b88a54fd2f5cce9833b52baf6601093932593a93a4e486284afa7dc06a6a8c11a76702d52593f2d9d58a34fafe5ac10b339aedd6ac82ab923109c0f1012754827d0ecab6c2870034e5e1ab5ff75197710adccf455de94f939e03ad0a1243225066f8827a9ea520272a05e8a39f610c938f53fa0f040089a4805711c6842f1f24b88611ef8aca9a5afa4a173fb89501d1d11124e004000f10ad94587ba2a5cf8c89619ac9d73c50afef8c0fac5ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb09f69fc1b39578f1814d05469de093a1ead2d8e96c48dfe8724d2b9f82ddb7f1c5d6296519b1d46c5633d8d1167a43c842b646a8ca81244670fa96f5137b403dde1cfbdd0ff6287e81d671350353e8a6e94216ef3041efa96391e582723f956d1244ea00c8a886364402d30f90fe6ad033e65070b7e948b7a1c96d5fb7a0bb8d49dfe4781069cfa6b82ca6f60bdd5ae7c56c153f3cb703fa203a918367cb3dbdda782d2b55a2f34f8873784d6198289b5ebdbfaf3c2ecc1ebf5440587944039a8e020da901ce1fc2144ff18842e706dae85577e4d2fc7f44aadb5f542074f7e681e3985885dc651a2fb7fc58bfe53d9a95452d285261ee221ec15ac36db5a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h17aca8e551fd2a5afb02b692aebcb35eda9bea227c479b8d6a5c58da33e9822aafdb65605e026235772311fb45b00c14802a33a6e67ef99d4d06c96c131bd134398d535dc5501d762412796d258e269d4e8f465b86c4d747f7bf4af51bce2b0b33e16df678c04cb1970be498f2291f7f6412f81ad443db82286d25c318d680d71c8df73b8e74da9bfb2cc21bebc55f08b4d67a6503d9b2c514b51893f22a1c4f795bf08cba16aacf18cbbd2c3a38fbb8ca725d8404fa19cf033981f72fd2f3c19aadb5e665eb4bebf9ed648cefce094ac8a15299b7366a1a274d8e63bb0a76541109772a5c2b1617d7806016e898b0baf492be30282cde65a63aa714bc99bfa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h210a87840ff77bf63a419b833a18ff1b63e43d5cfba1135cf473142262b50e342edb9895600380cba6aa98be4936468e9ce0787c42a1f23d97a19c7c465b5097485f1a4b80bae9d7e002f151ffd58cd1f26826031b33e26088100d3e57bcad0e67213a3a74422df89a4f0d0f5abdea68bf5d763158cc958a4a660766713d05aef4a84314d53a6586d502202c4c98b5c661a8a773c56343e43fdb56cd7849a90a1351bc1af78a25d0ebb11d215074154dd85417a12ec31aaa3139ed7c177260534d365ed5f9e6ecf291dd2332cdffeec181cf6b01b1fd76ca70a98edbd065749aa951e09692834ab3bcd737950228a953c8e0856e0abe07aaaec256f9b830172b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hff8972bfaf51ed1a8070ac903ebee716bbc134a51152a720a3a190a588a67e4ff326490ffb6b68f37aeac1297a6b47d36a4f10d9764758cd08286f12453bd875539bf91918dacc93d6dcb241e55a6654e61301485cdcd6871c18908f1f876915bab572b78bf7db283c8d69b393ca8a67b8ef5c738744912216d01b8fb86876ed103c9fd228210398edbc29c07025d70a751ebe215f5e05750fd3e5ac4625080e0160c1a096cd7b4cfe2f8da825e5092ae9624f98010f982f4ca7e4a6687e03d7c604b5313b3a63238d62a820a9a01f8707c5e55c9a0315c0b975bbc60847caaac0f096e78d1985546b5356f73fb73b9c5d6a56726909cbf5642343c8caa07eb5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4164f8b028921684b38c846fbee19576c00b8edc7c44b766425aafe37931612412ec134d5fa066cc7c7ca7a6fe5fa965ea0546326624e696ced89083e8e5bcfa666f4a3aa13699863aabb0ce72f2155bb6e215e58e57173c2922434e907b6bab30f3b54d4c960f7cdf9c20671affcb35ed5f6d170115e2598536a4ea40bf4d216ad2e35f935c11ce4c44f2d9822c1f13cf78fc41ee5397156803e44cd479056acccce76ab6b636f3cb37eac47c401bab3553244d465af3ebfe221739cde9aad3b8916efcbf38268fe77e783f20c57d24ef00f4a089a920eeaca3e7c814cd07764e80f9a5bfe66c67e0836cfdd0084b286700739d6fa2739ce64ee0927403d022;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hea42c907adca1eb9405afb0aa2d5b971e260596e64c499cba3742154b6671f787ca8af5571e3bc453a2f7d0daa6e95efcff59f7a745d9b6a17d5afcb3fb3ed170c1531cfb727991f8beda335878fa405b2b84acd80f7cc9f58620ff5755e2c654ba98b5dab0e3d7fe2f7ccfd9c140ab12329ac5db43b1eb56b74e426334fb524352d3bc007266e3d98df02370958c82626e24e386bee1c1856c5cb0c82d35326087f3bb8e215434e8d5c30b1decaf77e8fc22473ea957c42ab3746dc099444ab01c50485223af326d8e7551f3cc4bcccc590f4254a08951e5bf4c23c38c7cfc771e72c73868c359cb89a5f0b3a93bd144d90d8664b3ef9e26ee55efaebe4b6bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h17a970e364db92be294d2298b23c94f911aca5bdb9a0f0700598592fa33848d04a0bd82fe6ca2bea7e26f8e78dc3748c690154f8faf66d7ab258c69ff1695e17d820f8c583977c6bb26d019777368e7f7656abc50f5cba04fef68d8bc953ce405de6cf05660972f272ed82530e2863149d6815ada36bb4b53afaab8a9727a4431d73ada1369390bcdb93112ec37be946f4ef5dc2d96892f3e5787959545f716a9b480dde5c7787e9621e9091d142009c8845c19502d146821f2f2c46e1f4fb7b90e84db5198cd07a67a291211754a1f6c6cdac74266d93582b7cf2f7949e483f07a2f7f443118b759726cc8ec4b6fea1b1f364b43457278814e03851b69c465f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hae49217c9af34a1e3d65b1fc89edc070df4739cab1cd194a5a0efd7b1e2080f4696a3e34198f917320163e92813236511cd199de5e1907b91af09be29268af56c56329fa7055786bbc9f5a926a234ef6b97d910d1e0ab80fb35ee4ba4a9d8cd64c871dc3e46cc4795bfed943ab1009676d1684701857c54728c92ff9c19cb4077eb96902a17b9ea4547bf6f5d0fda8ec2987334683bc88a252cd9a067cd38c87a2d040cd3f77b94d2340da6ce7ad7e2fdeb788474ed31cca6b1d09aa89f58960e30342827daac9b88adb5e86f7be4c26512ea810d1bf696b9c9cf5581b115b322430962c30b2f18050305d0eff850a358020faca262376091bf35b1427a2796f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7ab4bbe60916841d24da115d3e0373e9eeedbaf78c5e700ccdf2241bdf7f5c5ddf6e8085ab916fc33a1ac9e36f83a04a565030b2f4a1ec3d2e54d746cb30b40f40c42f05a9f9b32df7d28c7554271d1e1b7a51e763d88e220deff537a17ea9d2f2a89e8eab8b8793233fca2f10db078172868fef0b77d31529ea6a1c47eeefa7fd619fc0515fb84141ad14ef4cd89aace2608902ac5c974bd2c3d00960fb3ed5cc7da70b38c47d56e36fea43078677a1dd9f8d6ea6ae77fb42aa06b6094ae1574dee7f29caf9722780d4edc2cb1627f988af91ed685189c31cce840a25a4bb6539ae2aaaa8a770239a2a4c03ea7143a2578ab8515e6076d9eba018bea010b6fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8945ecc761aa6f9dbb3b74093c5f98717c46aa9ccc9b7b51f9c20a951c75a8efd12028bce98c72cbeae0b0611f51069262f2de9215a0a61ff3d18b648b6601ca4a46b1ede4d9d57e287fc40e4688578a0f18a1f315c928d2d0e26097edb0af96806e21ca879568b3fd793111a5879bdbb819f8356bc176614f63d0ed6ea5ae38882d73f9475f0e449072d69dcabecaae7b0d1882512277dd9fb52a46d323f216d7a1f67eceb43e56e4b95fcdd3d4206e314a5c70431763d021fc3c20a8e8a29694b74dbf40cc8dd3b45087e65ba5db19f984a24c07bec0eac56f56cc9bb767556faedec57849f9c1a905e2476e75b59d13d6fea447d22cfc4882ce2199ef7360;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3c5dee5ce48dadb1e2fbfa35a8748bfc9a4ffc899f977e72fcde0c7f2ea3962907579bac7b0db480069e0659bc3389f684b9df308c3f0d6d097e009f17fb6a23d4995063a70183826296300486288f6fe1e7f6babe4d2662ed9ee73e4488bb0765fc02a5caef5e076d32606e19bc6db3e0b8dbbccd00b20c736ef438bff67809e33812d2e6e405e9139c3e5e4085681dd9649800bdab839b84fee9cb11f0404c3777578ceb39389bdfa9af9769b4a96ca38754361b00ddbde1bc531bc8f4d52f8ff2e2165d36848618b197751f8df83d6529eba1b56e68f42246ea8bde4a9d5261cfadbc413de7fcc7722b20bff6258e3a887709d38c28548e7948250420ee7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h77661229904178aa40906bf01be6655081670db1d9b6678bde350f0854313d92dec3ca9853e1e2a9e8cff4f50f4b7c312a8d384633ac3f268eb655381be099fb16267d29fdf6a2971ca4ecaee8dde7feb0c24bf2acbc5bdf9dfc3830e2e8ceb47e7b2a88ab0d1d9ec009a709c74cbeb80b65343a3615483d3bc97533b8eb1ad75db7c9edabcdb8f8f7c4df2ab204a8972bb8819a5dbf743ad614a90ab0cecfb310b51e2ea1426a3aa5823f3c5340f6f575e0652e60720d7ff5050b645e576059ac2976cb3ea635b432f60f3ec20616c5f24c4bd1d1bce710eb785244a9758bd0243d2710d92fdc6fb62d56e9fae133f2c34e6904a8d3e3c7a417ba03996070f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8c1e075d6428ed533666cc85ddeef340edcb601a0e088b000f0e016206d20a6131141dd6aa7bd9c456dfd25bf2d6a3d360ba197026dd9da5c74a225043953030c731e78dce71282779143ed055752384c03252e4abb0a460583990a7673fb62faea77364813a375d1cf6b8a1b67a85e074dec8b2d9b4adb79ee35b3d05f6a12346ff2d8a39658346a1578cc997b0cc44eab61b4f9aa517c70d9e746ba4198c3bcd76d3a313afbecf3e6a0008e37ae002cfaaafbd92c19d045d9db044d3b1f7e1cae5c700ad4ed589b09d0dfad41fa10b594574f2821b7eacc2fb849993b04139c13eea873289ce96d4bc799337205410d53300668ae9e5862c59cf18da0af0e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8812ad047a3f19ea767c2b2a6ac58355edbaf4c6f67a0e975d1da0502e59338a0701a5458e94bfb26d7b2154ba053090e20cf85e774bd001f4e34da08342772f287381dcdd144cd6135dd0613b619a00fd154c1f804ca286428ddf59a348dc3ef2d79b253f8c93cf2ed363955d5ced318d612da3def31ff32b941f976aa008eab7367cb4e675aaa50f4f9749053e18a2f16283a3417c05fe9084c8e3d72888d81e49c2904c23f3d842dde9555cfb425a6d2ed0912b4f3904a4fba697e1477d4dec022ab7e84860382fa0756553e3644b74531909436fd2216a5a0a353e3ccbf17bb32c2d8f4fc4f3aeaf2d391c96884badf4932a69c08fe971a56821ef0aef6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h32f13f70baa93084ff6a3492e072daf3151e0abee3920b60fd3814ba9f1f50f26c59fceb3e70ed70fe456d0e2682803eb55e4885f4a4372e65c1f33e620da1d549bf73b3c132ab636e2f6b391f8874345754f060a035a2b5487daa2fcf0982a140551be187f71e5d70e2cd21b5e78c51825bd835cdc49a0d4fdbc2a4b12d3bc0d91f079553020e2cea79d99a9c12b334aabac658991a6c99a5631c52726151cd734703b607bb874d6c3b093c8d4b9cbb3ec3113fcc5f1870a0e60aefae7b3a1c8967e38bf6f64fac3151f55e40a3760df08c410237ff3f71f99a6f1406d143d93203e0b6f4ad0ea6f4a051e31d05aa37467710aeda82d44586cadb2f1eb94f05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7b70a33d2571e8e103dbafd31b04f3d2c9592fde3c67a94f4ac8595a45ce4cd80b11a0503222686b14020f475910b088a1305f6664deb83fd122f72bfeaa907628276b1f20d6ca0d5be0b19ccd61e264a71db1d1ca45ecaff03bcc2005e795c6cf4926f93d15c33be2149d78b17f96abd25f539ff07bb71199939b8374849b45cba60bcd3a211f15675edda11fe77242944ee69e30e723d1c63b39ebbd4161aa1fce8be68c92648b2a039634ee390b169ecf28842fcba92248f515a17c71c24e1c24f6e7f58a810d43e5a7a486714196ec93239fe115a9c8b850d41f920a535a52979dfe654ab2a221f6c57d328fb66897d2aa27c7a2c7f74f7074727988f143;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'heec45059ec03632455cbc21336d3e160ee9d814852ad0497cbafc5a883c07d9b7b976d710224c7c38c100c33019084984378311231eee868d696355ccb1bf9fa82cff6e436e508b5446d96d58b2b800753171f7948185267ee0ff525cef1cc48e83e37c7045f9412106d35a4e68229e1f8a9e70b881d22af5e6dd5006d3ae89acf9b7f6780842eeb72cda0d3d3307f529eac34b1436ff0a48132346b94090c7e0cdd5a0baa76cd171ea1334b99ce439eaba71fd1607b7094434eab0050f535d59c85199143a4425a9483cb4f92a2f666fcc6c81ccfb4fcdb868cd3e57bb71c365575b006f86ec6ffc367e65f34825f1e536115b9a3a31cc154b2a8d5ae278bfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h96dcf7016303debfa88b7db0732e1613d18d65f3b4e1c971b25d35dfb40e0d0b971221be3456f75fadb142cda618c13476d1246a8752f248ff89ce5a390d9d957e22843a1396c9b0682c519c0fd6da273fe958760e6a06313fec6f58cacdc67249811055507026a6d75f786fb428aed8f006cefee832a8111d1e655d8ab957c5f1ffbda01e22b8e4a2367de806e80bae0c5874a1f37f844e0702fcebc16dca0deb7342ae8151e867c488ad10299860f51b3798c308951e62dc2a56fcf6384fc0c9fbe151b17b7a57126d224a52c6bec8c2ecae0d9ff78c39b58c23aade5bd9192bbf22e23845488c03b39fe4bcbbbe48817ea84f69ef6b46881e62c775f17ff4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2075eac51d527e6c0cd5478e50ab4ac2ef63bd3127677c9d1a076452d3fd688c765064e47a89f3d5c7e148f2cf589874e632e1d9ab92de77bfd7818e465a24acbb6538c7add03211d5d9c9fe38d5079502b0b1c6bcc99d3f528f73712486f434e7c2fbee53227eec29852eafe5bc0664871b6c99cecfb78520ab3af5b58f25f8d3ce9dec5529fdc832d961d898c8ec8e2a1e3d8f8e3c8372e7c5c94f60080c7a9eaffb8bbef67319fe4c552108accb01f2308f4a6027e433c10c4aa2af499f7591922e4c7f8e709ee7be7cf0eb43b7d5b7b7f64fa3c2982de3110238ffc0ba03233af769464ddf11830e08218a5c3d742e06b9a6e9985f686341952bd75583c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb64caca8b3eced95ff6dd94b30ded7684860aedb24598282f6c4ee3e4c762a16bbb6ba4a26378544f201900ab32bb8f087a0d059cb6756bf69098d46f33bdbee1d2c315c40360fdff2b2f2d2868b749847bbfaeb9139e214c50d337a065a47a94fcc461f14d11dff724b26354aa2def92fc837d1580ed764710376883904b744ca6256e34faf89ed698828a80ba5529985d6de07ffe9bc8d9da3e473a18167c0a2030dbb2dce941467ca3f553c36968bc1087e92982068fe3dd5a4d33f63b6fb535235a450c5e8f1e0194b8841a0360ddaa639e80e407d7316b1ebb3a41a4d8d94f682a4986468e18ee0e84bbc0cb14c7584f5906a981e5a93248075ee974599;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4193d1a085ea39ff9c4d7232019787cde758e8604a5794c5587c4a28d6361824a8cf9ebed81f587f3473f5656450e3d15d43d0e99bdfd914e0ca345ff33e52653a0d6cea76aa9efd8a818608be677dfd602d4451f4cd09fe67f5d1adab6d6c65468d11855f84222e0314d09ea5f0926ff4c4e0d66018d8b911bda740abe5d4e797876e0a87c6fe8892c0c8c2409d8280072e54edd2fa78b964321b2f0763c678a5ca93b6285d078c26ed118f7bfaad2c35d8dad39e0dad368611ab06c3f5bf63b40e0b27140a059e917b8602c531eb050adab9e471b2ef30f72b044ceac0d3f5cf6bf4ecd9dff6843a93aacc4e9e4ca440422290e6716e0995e4caf54ee3df82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hddd23104ab51afd9f3571bcd86e8b79c3a4149d1febc0c9125cd299a645280bc88e8c7127ccdfd9600cf2f17733649d3de1620291d8e9c0772f90dcacc76d97416d7ffe9ee575aa29a3d4a2cf94f0a014d06b2fcbc878382cea4776aa68ec18a77b28d90481d5569fa28b042a2ec0c68dd0b94061c964551991b7932bffa1b661f76931256d5b38af1d1e0c5a1182345ae19e5ea31f0dde5adebaccb114a87666b7b985952b3271fd86977d7db42f02c18772bb28d3c93458b82a649beeb3d063eb3a222e547bbc985d5e7297cc9e9f708b791e3ceb0225b800ef53d686eb4e1b2a3b5051187302a90b8cd7bf520580a1e6af140cf4ddafd9083d44c9d6966e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb6154057298b726f6d2914f20ed58ee6ad5428a1e2f79a6c0e44788551b3224ab44f75b90f53c2c50c2fe630b5e04ec825f4ba3818183018c407957ca8653f417de59c3633af7653e777cf14b434ef9397b9773eefa935b839f2f439f914d978d04b41b552597d45d33c602bcab0284d1df517fed371a385cf7ff8fc48ef9f9821e985e74922d8a7832adcec01f0a8b49a9cefaabc5f5f92d6cb24a99bba7ce31953189684ddf5ea0f318d957840c4fa7bec6f7078eb3a6f0c037e651d303514a6c7c6c77902d4fbe37ddf811771efb4bdac4d3c50722995287101eb5e780232720e8a03dfafc3927cd84660510b94cc97f807aabdba9fcbe69653a35cac88c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h47aff2c219b9b45b4095499bfea66ca5884a887e38479282a060e046bef0e16753431e2cbcd9fa3acd27f23859af84f2b08ebec6bb42df86d898f27cb2d5642f4b26fbddfc9e9109744ab5124e69ab0e9de07f8f5723bd8e6ecd57f6524dd92f534adfa64d86bdf830505ecf924e13b397ae4ffbaef7da347fc34c6f8c86fb071cb7d1905b65be9611c031887fe8cd112b612fb52604b33a5edfc54c0f635a53b10750d7af8f943d08b244f216a101e89aebb6166a95ff31cb1eafa9cca5f5a1f8e724db46f82ee02fcb836b1e9500e451dd7bb1e320c0c646224c9605dd05f7d45a11a0e6f8cbd91b29fcc2dddfdfdf378dd1e6294e769e2ed56221fabd4db5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd27adebb08e90b516802433817b7ce16630875aaa16c02ceba6063fcec7149aeb5bbbede3bd66a5b54e2d0679f01babd2daf983e80d3e9023e0fefbbd47ab3bddec2f1e085e57c1b07872760e155e7b3df56ae62d66f25757b79117483fc566ff00e20433ae8066c40e73c34433869a0ddccdf9b48fd5eb34307e3cc3168f4673b9b5272429ff94e833752a484b7075220592835644ed0dbc7127516f4b4dee310d0d15bf10dbb5f95272a37af66ef881b6b5a2700ac913e80573423fc9c8834c251a624b937b934ed583587f96c736ab37ee2157ce236b3ee765b1af185856bdd8e9fad6c6e89f745e7a015f8d87620bb1fa97216df30691d0396effe57c100;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9d0f505ce565195bfb3f7010d5dc410f765b3f6f39986c63d4ad311a2203b53b3c0da8a983e258228c0fd4da59e7ed9f02a199b71a4653c4a28646d522a839125d160f260068fcd245bab5480fc2f1b7b915e17b28b702f41a0a00b029c1a23fc6e099618cd2314a461f42ee4ca1898c0886c1bf683f5e052ec2b0074bf64a835b86095358d196059ff49d077900b3b7c38567cedc76a0b7f21add909d1493c2c20182ebb43b1b2ed4664ce12a5cb853571d7327f4e0509474bd7c3f52c152776cf05e8bca8a988eac7e5b0db099b6a43e1d4e69821c06d9192a778947407288d6fa05b52c5657630c6e6dafdcd94d923789e05c03bd3e56398aaf6d6369e5f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h46e9b950d76879c0c252501e4ae5a81467f4ff5ddec3cf37e89f38e4021276171ff2b6b375038fc18262ed865f391a4123c72af57f42870bfb35f6e7945dcb4abf6a8164261dd4984837af148dd9882a85bfb0962d8e426c790d85e8f9794f16e835f642b452f7116a9e79d4944730efe1e24c77b18471204095abfef0c65f65cce3e4b0a3e59f0aa5a312a8d7f9718f639d74a398ff1d45ef3b28bb7dd974a604186ed9abdf0e77fdc04f223bdf4755b47c81f6ad156c8752273e6c0e7d7de1a43ae76c39f1e36ac84da75b582288855d47a54d87e6d23baca9e36444acc226f81882c405e76756e4f0bb4451ea72f28a19fb9b1c4666e2ac9dadc584fb7a10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h56349cc6bb97d130e445782175f0e9187f86f352eff50b6936ccb44b21c6cc6bccf3162ad677b45be5fbee5da72ea764a2eee640fa29dd14fb46afb6d66f1aefa1ee1eb5540449082d89e6e93297531ca20bcab913a67a53ca1bf79bfa18f48b806812e95af07b18254556264deea585f3354f76448b99cece46cb3bc6c066182c51688a3e57c0953fa43d44f0d75222f2c15df4f519554090db1c2eea841cb942481dece7a42075c5d8b3dcc604a5f557355d7a34fb50d0313990af2dd8f660a62d039db7ca32c6eeda4fc219adcde3a9ef55f6a66faafdd3da8f3ded049e6cbc113e8fcb0dca65e7a8f0a63def87b3a7b24edb3c9f124611e9affb4d3da106;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5c2c58bdeb3b752f99b6b7832f83452d021e9872b4b697c41bb8f490986b8866882ff97a2cef5c0373dcfcfe2aaba34734e766d76cbe89b8b17c3aaf009b6150b9cfb90b9777bd747616af52df1a6371c03348dbd5696de39961eaea53ae9d84fde2a564be1d14a61fe222159eef9873d3b6a9cf6f345ea01f7d31a461c7eb25f31ee899dc8578ad97ce6b28f434048d999466e5eaa2abc5950de7ce50de003931640062c1399d4a1ba0e112278297798a6d1f5d61de802f0014f0aa9a3fc682572f6b2eecf6ef4d6b015c684d0c8404edc00dcd257ae6470deb6cd1043bddcb0de96f38b3b6bc020f5e5ec52e68c39122e6a51664f31ee32801db9bfe809729;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h86bd0abf12dc3894084a80f926b98fd260e4f567c7de27e43959eaf89e4751129642af8e93ed777d6a4e70d3def88e1b13fbb970d5afafcd64a43ae543114214625c2bb6d32d0976779af3fc558ea21e87a659c1106bb8990630f0827936f68335767210e660b52a85ba8a20bcb865fb450124233ef4b906658a52a667890c6d67a7d2fa2aab80fb821ba988f3253185e1d24f611701d1fce5e99de23d693ff3baf6edfc2ca0260006c7c2fb735b008d410a90cd9d90118dacd7987d7ef8e508f340fac5831b40b00088f2359875d1cd4bc07c120bd35959d6406f21e82bdfa0c6b055d93ecb220f3a6b2126a2ea752e510a972cd3ad0bd9b2f9dc8c4edf8b39;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha6bf10e0bac83861764f3af4e76282d69b53637f853d17377703facfa07a5683900963687d64a29be25a0d7b76336cb4a17d438fa0194a83b124dd8670edb41616d708bc7ab4bf2db9970acea9299e6e109c7a402ca7ea6e4f23e7eea7d931cca5e1d9c50c1ac27503db530a8b30eeafa4e4430cd5b9eadfdd2de2570ad4b5a74a30812d940f5b7bbd4ee894e02b56cfcfe3f72045f4e2e87ff08b5909357a5bb927ffeb499b4916c176bd09f1f3ad5f3606e12cc3003dd91377f97daee28c76148db51102ae5e3de1c66bb12e303f06547af565a2c630ecfc979a2a3b34a2554a280e5db60d8cd228df2abdf4307603829df3ecadfc35c9068b9c7034d3d5fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haa8bc1451fe861ae567f075ad33593eed0f9808d5059520a2f0d4e0d1db975440a0503be306d373e08d1a1c6a6607fec1261441b055d11174ccdb351af8c799b1e117fd706cdc385e458f4daed608c7b64f15f934229423a5da5829a693fd0c3116a64acfdc1efc072bf81afdb8ea91e594c087b530fc02d357a9a4cf540d924c617c5e137193afa4f2bceb8eae4facb4e86d9a4c07ae3ffd26ad3abbe73f5009f2a97399006c5473e4e534eb55f7d393ada36076b534f570e7e008e8e137d55809e07b1580a18516947496f1a5592184748a54c9c1399e89384bc212a6c9be1472a27494420d30cbaa09b986b19bca54a3a04b8774722299549d11221103bf9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5dca4773b08b8774d847e2a1bc80c76b9228ef24ddeb92876afa3d2550c994a7905ea7676636a8fde64a539e3d4bfcc48d84dce4a727bb412b9575e97879edd504d855ceab993d3c98d21013129e405bfcb78ba91ffd3e29d2951f3056ae565c7560809891b97f35378e4dcd55d812e4bcebdd626ad1c55d8b49d786245d9de97c0264571cfa5d8153fa5b7053cbfb2ea37bd06d4544b5be398dd57c3e9fbb3b9984a8802772f56fe37e3edd0ffd8d7cd7c3078bb67cc411031bb663f12b2e3d57fc57c561ae6961f39b5fccb580fbc0d65404ad386d9ed75c5b2d4cafe63eb6aa42af9345f557760e4f3ffb097c4f0f7ee665c2eed5682a24cf1b74c72391fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha780fc378244030c93cf4ee734b37f1ecaa5014c17e0cf014956bb50bf0ef377da0ddf0b126747608f36d5e8c6d0d2d15c43604c6b56d41982ef2aedfa206938b6262af170e2cfe484111cdbd2673ac3d28b0849ef4e967ba4af38252f2423c332a31493608e3e307033527425cca416db5f6529fdb867708124277ce3065309e0946231f87a7d1c548b11bc32cb46ddf958f015b4a9316ad6f07557cf33f542d890daaa3dad3bd1d85a37ab8e655aa90be3bb984f0506f2695427daa67277c7e9c6c19d21b9a1291aff81b798779e90afdb6e729feb6cd113fa3b3b349462eb26a826f8e448a481cd96a5440d5bbbcfdaced891f04c86ceaa13f1ec2c9f5a78;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haae9c9e167bc545c8c993797112e825980cfb155ad6bd88fe8f79df0209ebe85a08da5bb1ae1c10002b8436e619fd47e5aa4d6a1dda05b22aa5f62b4e56266551ad349ab838abf779ef38c939a4525e26124c99e539fa50689d0933c9b33c57389bc32ecd9cc4c5509d4d3b414cd71df55044db7921c67dd48bed47eebd1c196a1e844a245246b0fd2156d58ee77003f7f3c71ecb33fbb733331589e1df807fb6ed631321a723e7fc1f31c7ee32434ad4609ccb91bccfcbcf796ad0bf69e0979ca88259deb4212dfe5fec6a48d2939610a7d2cb798e5f8a6a6ff8c70e69db793cbffa693bef9132c18a86779274e1f1717afc866f827cdc176f7572b2c30ee75;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5bd5f0e52a58c9ae5e745e793b131d1726b66772717c5443f50b0781fbfd16f4dbfb57ef893815d7abd4ece7a482a6f50accd3fca762567953dc7a7f8c40860ef24dd06c09f2d59a1c03019b69793d0a6c4133e782a93eefb4f70fde95b542b5f4ff1ebd9810a1f0ed3fc91dfd9db25f6b9f7d3e6c13e696dfe09039cd3e5294321db3d1d25a2fd5c0b0f90fa64e86b3a6257b08635697265282769e0536432fa07ff125404a7027b8e6529724c5c78844bdcc0cb85ae28a3458c8cdfe34060fa4cde85eaef3cc480be73b32615ef527a52d0f37ec5ac07bdd7705c417bced62c70b59db11e301bc3f128739acbb2d3ea419a82ff10dd8a26e291d328afcb94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1f74ab851379028164580c68300ecdb12c5ca138e94549b5a5b4280150dbd18cc2c480d2e109896a27d74e025d3dc3c42b553a37b63bb755e141df675320ae0511d8de8282fbc6e5173558f6edb5587e66ce73a047a6c441169e22558f9b4a7849371ccfbc638a05a50c6c204122e28af87efac47ad940550ffebbf80b88d7ceb405e540ae319b24313449c631e5a7756b7f15f7fcdc23f98c1c21bba18d30ff08bfca5c29fdcc6e4a03bdb4ef37da9172676edff47acb817b7371a53d54c7f71a812ceae37d6bc231cb858f42126012b41553dbde00c3e2deaf99423b0eeb9e135c89823b8fbb27852d0e35041e0013cfc0adb4ea51682420eb508c18ba52fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h739ccb7edf189a696a6d1ba90c17892a2be73eff16357dbddcdf25939c4b00c63e14a23e19d5ae050d260f7f8eecf10eda8e75b3c5c6d9a197823556e3ce16278951747ef0b0ae458ebeb1d3b43b3d9ac769599c1163ce82fb7f96ad5d8cc48b6757abe99022c552c62ae1f27b17a71850c15b11a31781c5f971e390dba997854b889794cc1adf8e0d1f9bc6fb0e77f958cbdb1b30d0d530262fe56cc8ee02c7d11b543900b902b0f75008e0cad0043aa6e8af14fda1c725acf1b736a634dc67b15067474a781b356a6f94ce74bef6cb260854f10be6f0df40af80729f7903cd6ca166111c95a7344c576a9e84c13ed2bb09f0c38b71aacc741281a2e9992945;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4807ea7737ac38a2f57a91b43207874c12166c6075fa5a4d02ac08ccb272c62666da0b1a36bb5c755e5d353363b5d96ecd68e39cdad63c8d813624a5525530a921dd2c185ff4f80f05e456fa7b03d1b98851941cc217602c9fdce2eece98a1bf2ed531518e0ffc17e492ac8d3d035cec734bc07c9ed097865d3766e27fc29b43ffe2eb47d06ca61e828b89521076da1fe1ae8584527f9599dc53479d2c02e224818e2ef777cae320283a6bac350d4de45da3145e3f64d44d1c68e89edc5baf4ac59b9cbce6beeeb0321f9cfbddd938c87b930c80b56d8c2b8c5326ae075b599d03a5e534c578309d02201794b331490355942f7b2f3af357f79711d0c17283d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h31995ec98dc023afdf5ecb519a72c9aae9c386f4c4c5d0474749a75b61a37fbd92278a85ae6c5e57b6e4b2b94f1a088a3f53b52a4587282d04396e17136fef8a02d121e1a83cfd93d2680be31ae5048443e915264c10957bff1373da908fc620ea2f31c767ab2ca84356a4b42931a4d8055764b6953031e7347a98b46a2a9a7fdb485ddc58ed094547fd6ea6659ecb217e0ecf51acbda50a6f49dc68086b93341c00302b9f3d1422c5149644429c2634ccc2d408e3125f25f0833efda03548a555331e4621db98f5631a9e0b091cc52eb9dbc62978fd9603f87c48acccb361f6408f9ef218098bbd44b5e8f1cc453e924f170dbf0f38f5bf5e0b40e798e505cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7e7670af8a6e6178a07a71eb02c72ec8c9ad29b21fc250390b6d426db2896cc3202c4af7dc2af2fdf8606ca5a3c111888b13d85f3ec971c010bd69d013a95e65f2d7f28697a4f24c76a5abca46cf8db5a28bee391179d40c42eff9a06be0d2d19981200934bacba5721088872dc083ab7bd59fb9b32d3a6807d5f16845cf20f902d9523fa346f67a022a8bc17591b6bcbb9c1f844b7854571c335bf1bf9ad23e40e57cbb34246e67255577171fdbc6e58c180ae786ca329442e8791642039523e19a28714c0eea5dc9de3829576989e9b5055be00ddedb2bd0dd8c3e26672978791253726c1c2f9f9f8239a8bc1ee3d961fdab66791ae51251976ced562d888c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h29c23846a4588b78da4f1361f7ee004167c8b18bed75329770cc5dc6487d12dfa5df4773e4f64c2a8319b5fdb843788ef988de2ca2e2a2e6fac4b89fc2be12c387b9a76a63d95bcd1cc8e621a5374c584023901cb849f861e75b087a88c37709d206f04436baf782dd01f14b119b271fc8bc580cc6cd4b34135e01a5dd3f3c408ae7b8a099f3c4dcf45a3a1b476ae34c4f345e6b0b2adb055488c41733c7384a2b86db8c18de47dff7009977252dc2a607615bf8624054c9d0e921020e8e307233304dcd7450fc05a39a668588ce55d252baee3316476c823368ecf01889516268ad8d444c5bdc092765fe349737e59f7aae4f958b8e9c4b0dbd9b4a545e7712;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h334bdc77148d4ccd0f0f0eafb865348e7ee88d779582ee40444c8c0b5b44759595d397b14a71277810c663908df927587209d8292962b8fa28b383a58acfff3a33adc9c1fa77c6f51400fa06b50af8c16b6fd526605fdd8703d1d761e5607182abf0d6c4c0103b116a6bb7d2cbb2fc33f20d50bf623320a71a478bab4f7fb7038835e908d56dfb5fb70f919e99c13544a4d267a80919c5a7598f6b7291ef432558a9e2017366e2f5f5f19dc29c355679e1108b85a2ea8d6dedc463845a61fd3911de31df682133fbebae7c51537f4b5445c0e2912227488da06a662de003d66a2712736cfb9e6f881ab4f01357269003b3917a9a45f6663d42f43e45df052217;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h143997f661c44bf909ff9e86e62d44dc95a16dfe6b85df226f6a990270235b88a69438360c5b33dbdc968176f7e6858b82344f7650fcc97650cbfd00b466b111ab231ef0de4d49c4f082f91df10e86b517f9d5f538fec838bef90c1ede9537f6fee02041d5cf5997772e9ea51e525303fabfd3925fec4a3994d301c63cd53a4f2b9832dcad9890f6f717539917951facd459f1f2e32ad196b5673f6f7a4edb9d104a735fcdd0ae6c25a3c7e4c54f2d767bd5242291622ad006ad8326ae396b44cf01f4da86cce8647318057493546d546ef4fe6077a8327bdfffa8544d728e2e260ac2b363eceffaaf309e34d6c8f04a7d70eeda3ca245708042f71145c52142;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8bde214da2c213678614c26d9dc271f31e4b99b07ed9d3ca0bf3107adc897dffbc815d1a68597f8c04614515948cd5e5e310b27e7244b117bc33a3cb479739000af6ea4eb0dd09e684452638d760efc201836b7c5d0d0146df22eb1fd41c50daf0bd39f68da6b39e482b96910fe103b954b520dfe22c89705e4ef3138367d2771c87a826e7e76763721608eea37c7712dadf4dd34a3db4be4aeabdf19db118a3ffd725b07f41cf1bcb49b23f3a1ce9650661ce00a453c3ebe214fd7b0ff7a626ffdd7447285f4d923688407c8b89a3690156ca7209e11c29be2dbc8c4b82b5419c09e6e2dc04720124e770aebc1dd53833def0875338c19edeacfa57dc9602f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h82a07fdc8f34b63c429a12ee83f20767025137d5a4c5ed2def3436ac5976e07ff11cb08ab5fb3dbfa5d93f50ae7079f06c0633e61d2960b3d2d2cdedbdeea47e7130635b7d6e14f1a4db5d132a689959932d863be9939806c5ca1045fddb3024d238a46308306b72f5c99deea740165f3bfc4741379240cd1fa1326cb0acb1382090577da4f26970030a46e15f1c081d14432d0a355d654d42afabe4fb2eb21336b049db7a95411a5e7aca5d0110097f5f670c68b322cdd7fa39907fa47d6d493c773e8718db1e72dd1d175a1fb9b4f1e5c3da8935bf73aeca65be870320efcc2f0a4e1853a1bc72d0dc54d392ea82e3ad5c7f4ff5ef5241fd74c7afcd1a8c5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6c69fa40d503dc5390dd4a2083b94bf8970c2e68e1c579f09c84e41a735dc9fcf8b50ea94b939489d88648d88fd9ea815acf4be9ce8f430c744c4f0b470f737bf1073054153b49dc2c604bc99dfa48f7df58cd09c4cc953d01f66f7ef1a6680d137ad30a53024e224d85066082e369d30de1c4e76c83fd1d13d5720c1de56a9fe9bac75242723a1c522ccfd07d1ba865f6062daa4a6e7f60403ad443cd1700588d87c145499f6b343f6340ceb4948d6b00da5649db8d97214446f9ede0c98091b4b403c8758aa6dce30186f8ec129c7db1eec6062ccca13a865cf3ff9ccfeb1ce60ab5fc4d366d4dda76a67b43b7581207b3bcd117aa22bfaa7060d22eac7ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h666ab57e9a826e09a34713005ecc1229d7d39351a27e0b514e2b8ac3d7db94f2393f46a726efad40d2171e80e4720012e2a8b7ea46229aa73cf6a8cdaaf9fe81d696c40dc8f3f74475795d71eefed4a5b0e11e0a1d6602fe395bfd143875cc282d170b2e3d45d33994fe094b0dcaa094e3deac951eef54f50607bf41a7a02619cd9477a986679320918397f969be724d1b8d584854948db43b176465c0d55a8a166aaba85d8371c0a0db479c8a607846a8334c18d313d5f4b1526c34d0ac849724e5a64874d11f238b2341ffde4e0784e8a0dfbd86e99955972d8690a7139cdc1db8660a359cdba1235af8e737bc97a102b38e9df4b73c58df9d10c1e016430e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd80ae1522de539518e52931457b2368c67915fbf7848bc38906cf8bb9d04a1311608a19653d15946925db1b5c1129f4ac4463cf41ae717146ee26d083040ab6f88f72b3879a223205866cc5c0abe1b58b473823f6de93a9133ceae91480d48ceb5364f036881f1a33e5a7bd3b7588b1eb962739fc96822338253d9004ad3ffda46fa5a93dc97519c6a42541276a2eed11925ce7a14e1b355ae74aa3303b86048130842fdb02715c7b62ad418425a9a3e286e8beca24d66fc35fb4a56619d8b77368608e97ae634830f821b8c442ea603721512bdf211caae9a2ec0acf79d7b2760d3dda213de5c6f252bb568bcdcf3a497df26b240e2acdba4eab5930b7637e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h61f606ced816e0f881ff7eb31f72a1b84e4507be1d1b673a78472a7fa6ce243ad83aa56c256bc7449861eb8c39a7ac51739c8aa56b70122451e40d65e3713d36c48b11047f7d94cddc7579713cf7090d1823d0e77d8e00914e17abd471b1bf51a9ce8936c6ca5bfaea5c25479720101a90f55fc54aef68735c29d166fe25370c9fee5b7d41a0e7dfd3d8c4604386a7344abae3784160a45f95557de30aea66063290188cc851bc33fa04763bb0745282edad7ae6d834f53ef6ef33cf5213c81a2ceeff35a9e1fb8d775d71d364a1bba1337ecaa7e6fc5dc2727b0e9ca67b3b993881054f629fda0ad54a8cfb57790301fbc25ffb74b8b32cdb17054ad05de521;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h70a1d3ee3f29a7e55b30168a6e8dd4440b8d076829afb75f9e431ac627ebd281862a1407e43937b42e42f6433c5093d1b54f883227eef82be08192891c475370acd9499647d02d5fac24f1e06b34ca82f761194ff91f07748cf190c89a5681b07c25f183ab9b4392417c9a8875115a7ff6a368c117294f33d41360bfc923f4c8858026be0fa63c9a624081041c02d7fd7c49c30608b7e6589ebe315104f09ae080b693a2081030e96b46e461e29c200c6c221f6183d80037bd17f4f14a57d45ac37537cb69bf358f576b3d8f1b7ce9df7898a7c516ccf73b0e8ec6287962a717c69eec62cb141d20909441ad693d51e259a828b5d83f9f1d122b3a1199262c6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfbb652ca6486751f5bc935ff098e0f7071c8c7a41f43cc229789e4330f312dea40361717cad2e33ad0bb11f1d51a152be1fbf86e3c1fb1c53f1f2c4f56b28a00da9acd9bc454832adf3743c59bb2e24b28774587d084fda31adecb349071951ea9e45ec95c1b18e7ce07210037160f27c2a36d01aba22e1cf1b1529d764f616c27f5480e18d6d013885e9692f08d801945989e15f1ed95b8f3e61595c9fa9fadd1cfb48aa9ad69c1b862b89a021b04f8a34d082b988364ee8cc149eefc16dcb5340e07f7a62a95cb814bd89124a7fde86196603a8ad65a1c70531b3fa1be41f3e778c990dd46431201e837164aaaba5450bdfac6710d74451e2784d205cbe5a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h690e60901cc952c57fb476d3b4d62c8b3cec033a5daeca8b31093c62cea445cd28732a9918156ce86f4c5ddd83c7d2d62f85e4812a31f4dd48e33c78befc2209a8bdef0a8c2d5d4217a8cb5a6b29435d8f398f3764c8c10bdd6c8a54407b36f6bcbbd3be5e3611c632d63d6aabc6bf452fb429a8c6ee9f0f84b83653229b5d6b594da5d40065525d6c09f620934a9ea89df254c3c486e50e383179b0db2d5a9afdeac7b0f628e1927e2deee20ff21af116db9ff1c73229c710fbda449db90131589481c4657e3428447128e894be3578455939e03b935a37fc8e8b498423c86f86a515a5bb9188938b886b1625bab769b01f2464454b80f6548e1d0dfb3cbffd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h47ba84d530f222d67f14934f35c92de5293dcbbb781970917a0b19218630af0a70b9f5319f5236e044a6b038d8995fd74184adaab3f00144875e9990c7cbb6ee3ea74521f41d93db44905d0fb2e4bbb9824e614a427bc399f5088bfbb4ac1ce2ab8b2378523047b8867dfc2372e808dd1e2e8bdae6f9c12b442845b1d8176f21f720f190aec068fbf49a4240678bb6d6481994fee729682c1be252da1a65f6b5ad95f2cbce12fd020284ff7c5186e9b588aeb29427e62bded21023a62d14939caa08de642514886121631ece1c465205244a10c6be8802ae77ce2c95c703f89e2d288452505b86b76a7047b8e4c2eca76368c29f569f600be2bc8e333fae6b16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haf0ec98f8cdc5776b28b4c521f4480cca24fbbda9c4168777f133982c727a338322cbf876e205269d1930db7ca092c46f329e149194608262def2c38416ef7709eb7e8c773904a465801b6b6f51b194ea21be54e34898b1ee588214f9a9efb09eec270b9ab5e8f2d67e820417a0a6a259c5fd5b138e399d1e65ab4d391fd0c1a482d25b30cf7610c7399937a3d321f820b92a31127dc1f16ebf336530cccad979de189a7bb9e80e31fe4e5e8de7c56244dcee705e5e38ced30892968412a1afaa5ed3b2546d95abf6606898a85f850c8f60f64e4ab133b4c985fd43cafa80eb94de0c14208acbeab661335684f2a9789354600660009a26677a6752f4ff248ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3f9bcf86b36b6ab480102acf1bf850f311505a46ef9026efff6976ea80e6b64ed4a1d8e64e8d30c2723e68242fdf63de99827cddb4c22266f78cb40a4efa9bc19754a3f1653036236a2b5c44d5c2509f2624377c9730ce061e5f7c9754d936fa58346f3015ce96cdbedace5a3d940481bd820ad85c141ab667f36ff9ff0d5451080aaf66ad8dea0bec38d620216ab546c85003b477c06febbbb658a082230e1c6f761cf73307cbcc559b9c3c2343b2eb4d94ec28bb041e8b2f0640e8132bc6b64c81c22b601f4169369dde32d00831cff704c195b658d7a56574ca86c47350ec47429d650f318d5081ac82aaeaf96c6622b5364b88b9a826254f31ff6d56badf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h81e8a9326664745bc988ce5d3b5a8979db1a7d71780565273978d5baf0a5c8e1a04db1c29797d2ae77fa1e4660a543d2c31dbeeb3151e2d5f056f66a9afd5da24fe94461994912da5929f5512083e5e63922b4e8447de5d77c07cd099a4975a74589b0a747cbd93b80f2c370c53666bba4a8a717dee09e689ae8ec7cf8b05799bdbb41226eb20e71a9f142572b8ed111cf710f3d13f46876dac69fd1604f8ab0c763e795fef1c5d86ff3b998b6a9e4da118d4ec4723c29ecd83e3deeaebbc1cc4ba5e46793f86395de6097f3d324fb7ae1e6b15eab5a1f2d3ac8124222962cff6f5191949a27ffc0d519675b8d9b0e8c42a14c8ab566b099e16ffbfe3d59f85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he39d1e10a877a088b938fb32866752cd4208006ca5627aa0b01b82ee5600af12feac2f519518c8a24686ffe5e6812f6ca3f4fe8ce4707bee69e511df6df5e000c3c122ad20e587e6bbb3fb2175feb8f5be4f62c0dc491a9947774a51f3e21121361b666b7b529d1baf70f87b0b5a82eba7fc5b8f0bba17a8e269ad634b8994bcc99c9aceca86f19f5d86cbe3d284861ced603b416ed7a786d3838012aa95738ce6d97ce628f58cb5905e04707104a1d5c8be23f4dfcee5dc1db2554658c3788ea7e9585f17b3b62ea23625c71977aed0616735976c467349edbac4d24a74094521a03b4018ca38ad8ca47e3669cfef54b507c5f139de21d40f869dcaaf77ee64;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he6111f7dbdf5a5d199a0fd99027e73691058a5e0834f8e75ac041e80f0ae1326f1460ae0749771623ca7a1e13fce5029a1f0c01cf6d92a50eb67f8db6c876dabfd81575e1db351e1bb1074f6c42cc78c57a1f8b6538ac4dbe3c4c4e9d466dad11c6bf9176c8531d47da3058b0920a5e1059809dc92a57abc256fc0f5381066e132de26cdffd0963bc91e4e685e270e0fd2339103f117484404866db99fd6d54ac99761d1cc9315853168e81da7a49e5b1da93fb635a34ba05afc3e1a4362f6e4448fa7e5e4085e6bbb146529db344a9dbec82abca673b9f511fd334fc37369dc41bf206411646a1718412f9b460f5f8fef206797049d230a1d34e96a451c792f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7487400a58f141fdb37b7d65ab89ac736e7827610916bf70c02fc8c338f079bdebc2a2d9c16761aa0f840415b78c93fded2be19c932897fb67f170f6b075774562af8e9cecc1868058bed01299e85b8a3b57f91d6038221323854d9af787ef69f5adc98a784baa1ca47c4224e34c44456fb8d08795fd18080b1cc9f84876db13fd05633aca594dfd29001abf1298093f589ae6a6d3818bc79e57c1ec26d38c6ede097f78e9a543e0e1c818c414b6c8aae6244d3f8ec1bc21fb5ed2213430054a30725ffaedbe5cf9861485ef3e9ccff557b23db6d17dd8ee2fb2426fe40abcedb3234c80179ae1a0c22fe347c2f0b32b0c11e73b448dcb5850dca6a9c5b3a861;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hea97a9be0f4648cb3c48d930d13f7135753b18061f9a5fa4902e7093ae9e8b468bdcfe33eca3ddc71954d945a785b13fd06b4d581ab08f4245878e929dc4af3598a52724015fae62a7fb57aed1beac3c4e55d6d5067d6203ed8ec3f59e7c52b39f83ad15732210db8fa7b97183310ee628465c2ee5e34264a4abe1c32c8bdaae047c396a21e6dc13dc4511d0aea944af33859969d60888d2aeecc9c0c3d7b6615d86a1105cd0699139bc0804a618ccf4dc5bf72b5ead86fe43500b3ac697f8ae3e54de5f41617ee880d0d919662378ed9155884d457be01ab62f50f5c848601c92cef0063af899367238c90ffffb73dde5d9046d9e1ac22f6bf77f9ac7e5093f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4358e121e9090d742afd6bccdb3a60d1e2312997d872d0c77422a9a658b32c93821586626d748f2bd5e489ef28f7ebbd606bd6a4cdc09e98ab2ce0a5deb246c8e7cbe31f437efa0d34934f5bed5509fa63cd163bedd7e5975855dc4367461e3174a47c48c4a1fc516aa86cc4b88e9a304f2a412f3cef2a7ee30257e14e1b00c9e7e335e222112b56b8f4b34d7ad75b4209f9f8211dfb115992aefe02433605116a852c54695fed79cdfda15f52899cf6d946d57f57357967dbc8f10522ad589ce5cc76b5fe6cda5e3a4d17810674ca6a4c97958a1dbabbfb2ab4f122f303dabcc22e1ff9a6a82b131092cb5051d6c41e006d6eedd38a29241c8b5a16fd99395c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9bff738667ab4c8acc308a4d8bbd23c7e5987234b9faece8b61709035287ce09484c587d7b7e622b4ea5c3e4eda780ce0005c9ceb4b382d6d60b41e60589c095b0e8bb907c0ea8e0d067db186f5995625698b11cac75b3054463b76df5d48be63a82dc0442ad48ceb2be222a2ef7ee6bb9320dde573fdb8901380a36ae5034618dc88549ea7a91e97ac55f41a76d8af971bacd92edf8cd0186ec494463e0c066c9a6faa548c1801feb40e02a8de4f339a59f62e154222f66a68ffec8881c9e0f1c44e7609b1f8626a25810e948925b54f5a752b57e6951aa1247c1e748e7f0b2be13a22ea94f132ca50d1c41200177d3a32599fdb066692be507f147b3d2d0d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3a683477bafb1fdf6f6b59c4df31b891d98d5fd54a8da0d573e88fe003192c860943ff5f06ae3fb4be15c183d4465a2431c14fb746e2fb31d5564d60e1d533006b145e0590dc9eb3206bc108e7b6ddea20c2e15c4096315f37c690c318b44c88eb94293f7f55a8b433daaaf1bef59b97e1d6537081c3a0b2b4c120320d023e5e97eaec819e07207ee29ffee318793617d6a92b1a0a1128bfc176a201b73df6a5452389868f3123fd5fd1e8ef15dead874a1e590c71443d37e67473e3b083aa3a48b045b3afb41c691fd8f46c9a2cf28bc8df9eb211f45b30ff6b7c7d93660fec4c5433fa3b62040076ecee24b6354039250fd65675fbd5ec83f5b5c0aac7ff4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h486cecfbede4a1b7b05e84c83e6b33643e71361dab92cb0042ef4ce6ded30560f0085f3b1d033796dcaba5b65253b41228ce5aa83f5ae808d221507c6d1d5e7c642d4f333176bb23e1de4bccb51059e914a0362015836a2d365cced0e4a3c919aa873fb509f2b7ade11f48f03d18a4a38da03883439d32a6a629514fb7e094e25c2faf6e905add882475bb85af393585b500be5ac3d1b5e605ede243995d0f6cdd2fbe62785f7ca7e333b8d4b846384a58db1f9cc30cb30dc5e8e7a96481566101e832674e7c149be8f60ee4e9bcd117feb064d33cf36e49725e71b6ef51ec2f9b5663e0a344a915609811cfc93de090919f94c20883b3a28ab2e1f90a6eb0de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h125e927a9ad9d63c10b4c43efb56b6db0e722f1a3a855cce81bb65c265881fedf915354a582e6ae2f25b1e3c54c93a143db2ad0d324a5e60dfec4d13bcc2e94d0a2a6dffcb1d996549d1521b6220063dff198959128ce7f908f18b3cf855c0311e0da6e6d37d018d94f0d9ae214c7e482e689132fae43aaa1b296d490e9b3a63fca6080e633784be36da7901b928a6e74c711eb301bfc75ba77e0b696b8d966f7d74c8a0bb397a3f996679f4176b1fea1fa8fc7fccd2394502b6affa11151e5d356b0497cd49873908c7c345d3a6604239c0708b82cfeb68a9baa094daea9bbaf1529513659f556d4f1e8988d2ed1031e71ebdcd038a795f3bc2a440c8cd2297;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbf6fb253c697c62919ab01b6cd62075d7072af66ac89a7c71e86f0a95cfbd2a28396876681ecf4ccbcf4198b729ed4a470a52fd8486dcfa253aad56e00d38f3426457e00e7f66a2f18cef4812889199958507a377519dd5b2f71a00b45c2d56c5235d8d86c51ca964d07e9a5f458930242dea20bb4f2125781201be5ab29688bdf64c549f4121c69d50cab9f4b6086a201066128476c13c3cd3e266de3f59dfd3701fe5dda1bbb94be1624bc0b94e4f013b9def529520c183917ede5c446321d70f8481632e7c1ad531b7fef0571df891feef36869fa52b9237126c9a53cb323e36e67c9962c8392bf0da0fb8c30da06c694f3fdd8489bf5246ff7c395f0a843;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he8af24b3bc172ff05f82363108396a741d088e59f2ea56e7935ac223bfc872802a4c9b52cc82ec9c9268374f4f6cc1dba0442732af928c64dbca5b4b2d3fba4fef2a58758f75b37aa11c47660c49638fc606957b8d26d6f2d7052aa15d92013469bd83e2358536f8e491c98175b2f60445ebd57267d16bb1cc953a6fde4416ebd83afe18897866122a790737467f1dd290cbb4506e57f27018c43b5d514d15f4231e545d4397d28c9840c31b6bdca58d9b4d5863cd752f10e74e576f10fc05039ed0bc80d6b0b6044704a043aade6284880677ff24ac67f00a82897fd06912875af1e049de1f1a54640439d597c84de66d71dfd6a35a74da39767b5a3c964b1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbbd80ed4ab46322cfed3244325e6f03e2c7169511edcdc1a67bbdb09902981b531ad527579e842ca757873592d550e9e647509a9a8cf5d42cc6a472aea79563aec417bb8a22c8da2a944fbc90cd658bbfc6352c9c756fb968eb7cab4efe5d19aafefdac3c2d5cff798d687c6294325a64bd1221c9d6aa65d85b1172020fd21605c30d02bea33caebf210095afdc9c3d628d9540b8d9603cc8e0a30b7967d005d0b0faf31c081981db0b7edff4d7f12a05d063b5683bcc0073c6662f8156bd426fbde3086b8aeaf24c62c10e92a8edfd71d758c9a4e7a764a723278bd140b2c0273a6c127aa0847922b726d340960811719118d6dea267cd9aea563e2f4ee960f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha528eb479d0b062a37234844ad8637262cc7aaea6d14eb58f2bcf47f256d3d01c538668b23bbc6af4651c3bd4c1e06885bb095cfd9a043edfe7e9343f00842b6ea4c1f717f0cb71d328833963a772e3176237db76376f0cb8c91a3f860ecc4bfcc93de170710c320a6402ce71db489be9d36d78b9e65ab4ec2c72350399e7d94ed29e41f341c0d5cfaab4754fb4e4066b755f6d3aeb6c9da7ab8e33b098ab5f8c421e99e8f9d80937325d5e886d5af0cb2adf63ffd72f70820575539348feae5cf30a9dbd9f49f907726e4b2f4ec0104b92f28f58954971f7b897cb4639bfaf3af2c64d3c615827d819fb8f51b69b7173f5ff7739c7e509e5f589b9a30c55695;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4377502f27f2a541cbbb358ee4c0a7562e06fc5c986f496737465ac4e42dd21f37f11a061f58282a586f9eaa854b6800af84375c5a43637e19235b6958c48834e98d40dfbd93c316897e014847fd261d9384a362a4f9109a016f6fcbd2e64399e5a2c15c677088f39c19bc826a8807b6c2d2b58394b3c13e328f25a79ad2caa2eac239763cbce76af807253f379349fff22c805dcd37d58705fa2fe743d7f9642c66c6ad5c54cdadab1d01a3a853665cad903eb68f15ee9395bd79640274d07a13d244d5418d9ecb2c6a49261509bc6805bf1221de10f6d816c7816c095cdf0bc1c342204c52903837b58b173bdd4d473a93b8bd9310a40651a64e472afb7ef9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h85cbb083f500850f2abe743a4d6cd022e892b8b680daa222c818bd42a8457952e6ed1356c6b68bf48f92ea1514ad5039361314591bdaa46b0e2af14a8d53c69d91843fc565ceffa00a84e7ef52224e0b8fedf1932db493d2eda56dd57ae64ab6d33568848c5b73501f05b36fe261295c8af0d231234eb541501290a2c697d44d1a2d26555047e53df0d74c8d9c318d683813823ffdc2e6aa535b0ee2ec865a098ee1d4d7dc3fd3f027bfcf998bfc3608b8f64631305a8d55ac7f50fe69f089c3a5d92914b702e43e05328a69794733debc5be52b85a7d872cc78ec35c582757211de7896b4c682ce50fde46e002040ae33ba9235fb9bf84e99a593fcfc8237de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h93ab609a0be4f6e66a6e0b68f26774bf536cba48cdb7d69aaae5423184e1a286bef92d1d5cb85541975a0e288e849374cfd5cb2f2623194e81ccfe4e2fcb2df156cb90f59a0beb6d69986b29747fb3551a17e5e8d8e3c66ef13f7a575c6ae54036b124bff84a66aa16e8fb89f2007b2f531851e996da005ce0f256d011e17f682e393f997df236b6cd3d43352aa9d557073db4d4e320682a7e9c2d028e5800f3129895a524723538fb5a96532405e100f607a2b935f7fa07e1b842e83d379476c977fa6e2cc7c90b56a356c30e0116f89db7bab8b7d3854b043ca40d4c9d8100d0a9b641752e2c1fc5894a5a709e413488f8b109513074fadc8de6264335c818;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h472a80877c090c4f438eca22304e5f293113c15f0f07d26df30f153cd3cfc8e6a260b14745a895623e5927d10bcde20a3aa02e9518a8b0d34a86fd633a68dacffad3f5c7ec12f3335722818aebcab0bc5e4a965b7866d765e6c24b4f6f0d68f9dfcedff7f4168a608839740b67c1f21a70141fe4a2feaabf7570d53dd6781d2d0e38e553a6d8d2371540dbd4890ae8cb200e94bbf78843dcc07ee32a6fa1f6e5f1e331e5e4aa544ca06f9f67c40fc5ad7d2f42c3070842af7bcd0b5a1463e38d7483b53814927d61dbdec5adf23447559a861d862dd57de4960de4da9ab57e70a307d7831035fd55428918f91f64289fdbb2cd97f3cc77505288929f5a9d3a5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8255e54c261b64581c7ea2e8e7b4012f539aeb41db3497bf1b4b42eadde47befaba19ebc816f68c1445144b23d5ca12f97395bec980cb8ad99a378df6b2ccd2eb25a714687d26c66d44a7e7e83b7981d7145efbedbaed2ae6c65de646700d394398af9f02f0f7ce38045c2fa8e73e28ad8ced997cce5a202abd497a2984c4e617e3915f94d2e88ba9ea252352428321858fc921d72cf692fda1019d4fe3823156ec3b79ed3e0098a871880ce182556c80fd2607a462cd9828a06fae0b93fcfff54d0bf8dc6acba6267edf100539f3afa5773e34bd81f9efdb45e63d092316c295ac6028e4b5e5539b764369804786979e5fa52a5e70c8b677c213b4d7f129c04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha1fb1ef11fce9be0196d84e376a962e6244d02e0b436b911f858dd70d67bfff0ebd0b5bc99f5941be756d97f2c69721a29003b9a872dea1a2f359ce083c01974171a057b1fb3c176c6e6453e0e9ee21ce27a4f5b68cfe6624ff16cc00d9aaf35538e465ee54bd7940246a97726141c011a51c4da5d7904b904baf3599b39416e654b3a0c95b18975d30d2bb1815abd9e2514b0d1a1a02bf4b1d6ee8ac5cbeafd20aa8a380c3cb4d6469c3a6c9e33353faccb46b6a50312216260ace3df08d59d204e6c3b1515fc67320866b10bccf48e5d41c327973530a4a73fc56b1c3b60fa464a8953b4e740b375879a1c79e48cc506b3a14c1172173904d53020311bb549;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h78c2e576deb6b25d90a1417df93108f072ae0fc312356112c979150b405007b76731b97e8741cf0e05fc5c81fdb5ae7d5b56adf0073af2c684903fa255b42219f480af9ce214e99a0705ab7165c580fe7fcbeb07d0c786b90288edcd0f512c3cf26d5c509ce8d677ccdc082b21ce10ac0a5ed02664ead69f18e58e17ca2ce40f56c72597811913f22390ffbbd7c38b039cfe5b9c525081bdd624d9a5f346c61adb76699d1367c6611b194c657382afe96703116305dbea54e082eed2ada89009ae6692d88894339724b655c0739f7b8d52771e00a734ad848a6d507d51de6b1f7e383efcd396fc9466a9a1f43e270ee9ef772e236667407dab4bfe7169d295e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6ce6dd8b1a411f5a7f4f8bc82e10aea687f8c31f547fc2dd6cbcb34d2ee92abcc4ca273e6c8dc0e9a4b036060a6adbe3cb75f351296dc2ed1d58e6dae55eb84ed4c2228db1311f6df3c28e360973bdaeb11cc6695c7d952fa7a84c69825a979c365abc480e837295cc097d9dc676ffdac6f7857272286ae1d74d19a018708603993c61618091f7df11ead8767b07c2b1f18e42be459d0c56bfbc12612df574fcde4e6f9e7c28901a412d1124c914c31b8418d3f43349ab74faf2b0c713ed81ed667d193ee2d02d185b0c7d8cbb12a6e45263aea80e0de4c74622960dac7c82a43a07f8e1ec609205d11a807f00c0308614ab324675f3c29ac9166f432e53b549;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'heeca38888f460f52b5af5b7b02e6d112f29b731150a5e28d9387ca5578462598e2eed81396a1f2ded86712870ea9828f2ec1f60beaa3d393f77955b1ba38bfc1ceaf7d648f4191a6d08e093d838d543dcf189c8fa895384b3541a99c691c6fa1264921e67da270f19ed05451274376a8332584257f512d6ef8c658d8161b62623d51f810f81d54337ff0a0bf68a8ffac7e5a7f3a17dd642d4d889426370f7252e1b02fd38a2341cf6f390b0c933c091f82b49ee9a970cab2d3eac6262da115fd1bc0a297dc6dc179efbb9ca425de009a78348a58dcc26469bf6849b3ec2f5c7df0bda8bb75c3635b7292abe4cb4add9e97eca955e2a3b6be3b6b36e657b81430;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hca761149406a0b079998ce2faf79e4252c9b7c566ea18a8dd89da0727e04b80bef6b1feffc1edbf432322c22b0353ac8699715eddf4022e3f9a4eebda484b2fb80e9175adc691f06a8d99c4ddebceaff091ed1c138924072b5a9da7b1404dd6566e3ba8709b2cef150b37af679c14814794860204ee0c4c5ed419167f9ef2676a20037fad7357908e7aa141c6e266c852feb5fa09c3fdd5bc17c16fa24528eb9579bc98b2a160fae8960a4caf6b101101eba8c931652b200c74da3e8cfa8474a0de54711f87d04996b24edabd3798b76b53947d73211fe92fd5c5b8e3cd4e05ab7bc164f83956737c809542b2fc8969f5a36a6aadda9af4c354173c5c5023e5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h900c2d3dfc49cf01933ad9b46cad03853468a7296b9978844db748be6620afc6a8bb4ee61eca726a5b3fa0b2d490c009e4973419af594d6740dc2b5abbdc0e6ed83cdaf0e1f03025047b110efb8849f88dbde65f590142db54231bbb2bef8aae0cfd72cea5ff525ecc0750210a7893199b160e511a07aafec110ea7390346da570316afc8c1785aadb286b59199c59d1fe89058eb4338da8f037cfec76d94202238cf58c0b438161fe37e92b1765ab92f6910600cdbbbc6474966e0d93de21324c74baec21223e01443180695fb1c2ff6e22c25973e3c535b93bcc99ff21775cef3ba407f1db2fa042e57e36f82b4871582f0657a3ee865ddb49abf38c5f95b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfc683ef686879010d083af83b8930db9184deb585b28e1ea5498318f85795369a5d38523124ab3006b62c9de9b43c3c2ad9a367f2506bba0d64a4991c361b7f23bf2f450b049741dac249d35944136fe07af5ad406b2e1e1d0ad120ab0510b5b7a14ec8c43867b414559a1e3ef6480eb3846a50b3aa52b7b80309c344c71b4fba4f2a337b990763bd7698561acd05744a4e4f5d5b304add6439486f6959719f199070e2c0cdadfb23a7dd9b20e53ac07c6c1f3a261bfdc8f189bd9c8e424383a4030e375a573bb91509eb9059d6c617e4c8ba5ce4aef9a6f8de157a8a2008991d438ae41a186f0d45f2de7fb4395b3f58ffe2960ee3986e7546475db8522209c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7a631997287eaca7242661f6b9b7dc04475dbebc2804a7a86dc181d5d529b0c42b05943eec97ad660f1204e204e293e923cae10f25f1b6bd9a587b24167ea37c5766f3ebc30aa6afec4ca128c23d242c75aed82791fd3744234d38bd852b5d552dc405351b3d1e1caa0f2d30d4ff88d572ab016510c98502a9ac2503b4b17b102947930559d6c5a5d63e4a68716687979049e6dfd9430b848a50f4bfa3a4a21b1d8c1d206a07f6c443e5fcec9cfd6775f9ad0a3a318cc1718ca9510c29cb91141f85e6d549f25a8b4692c826eb300b328326e575af4edee65201bd04efa4f61209a42a2c37edc73c08d223ad73056acffd5165429d1589647192dd55b7efa982;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h78dc7a6583b9a880989d3dab16db4f2aeff26c78c99bf02acdd15bfeb5283b099dfc967eb223f07a21a6b53c40bc889c62a4a028b2f7fe01ff2ee6c0543b4d2716c8a737a0e8f048d5e59e1fd70da24cb1cbfe0334fdf25489097a0b770842942e0105571de5b489716250f7031ba22b52c91ce049f7a4254302851532a42825ded44a8ab4a627d19b7bc30378ef768803af9d767a9c9f91d27da325013069ffc4e89409c926a0b5788874b78ea5f2171abd611be8fa696a87b42399f05907f0daa4ec894e2090fa0c5c15945313a15dd54fe99828d81d26a452c4c5268147a2e5cdd223e284c821c47912d87ed4160617eaad91b784a5ec7958c69cd2d9f527;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbe5c9ec5a9e20f8aeee649535318a0845fc06a1bf70bc0e461042a65740e5f418729d27e209c01815849f1b420d7126f5040da5bf528fb68b74263780ad5b6eb86598391e94732db8d4c336d1a493990cfa171ce084d8726de50415b9e2851173f13d66828c7154ee651f161b18b3e86156ce2ca83f3cab95c706d10d136578ce3674efe218c22ac3f4a586fbda30b9181406d74603a19db18136b0611e1c715d885224fea9b1ed27d5691aa2389cd1d2d787f422c8af1c6caf16fbc499bb36fbe604f506195a848dce7cf4d26a003cbac988e8f6910c29688d4a50369571fcd7c0c2eb22f5cd44cd47d26b0848817e3f25ae5cf7864de78772f429fe286ef7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8bf62cf00d0f758b8ba689fc56282e7a44b586da4b7032f727b77bf095065410dd4be43155d4430f6ea116e708c55a295cb1bae51734019ba15006227259f431018e999369c6952538ceb52e1fad26cc3e039f89a1516f63dc124cb8642d3fc83ca741f59ac7c172e5068dee1249b14a8c84cc848eb098068cd2fc8c2d9be42b3f04171e203fb33d28f7d0a58adc8f1a45ebaf1f2cee86d46db37fec686c84502ddd691215d4f942925090bb5d446b6291100189d9ab3e87046eb558d342839b4c906c30a186dd92bb6f0c901aa01f0c62e34d41b1162e3ef3c9208110df8c89f888db24923dd9c1c446471de1ad26f124aebd860fcf31127718f56959b034b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5867a7a8857b94bfc1ae7c185563dc138e948fe5c955e25541ab8ac916ffdcf388d6f7417ef01612e2882292fb2a17b7757dbd1ad457ebfa8048bac9d40e118e40190772554356ddc7d78f7af860fe66fb73027755420dcb5c4da35790d8f34d60d692e6ab7a47df67288349e5f1e9260763457854f869f475125e71d7bdd4f2819df086ea353d2302a9e23db96b26f02900cd8138623329bff8326131ce569fcfb397a2ea205362a8e299238205fe5cf4c04c7990fc3938721368588536c9503befcf90ac72de1a291014146bdbd83814aa63c8f94b345eca44a69540291bd6cec6f83267e029c5ae475ad9680c4c9cdc6fa49402d6e04292c91421cbf5fe2c;
        #1
        $finish();
    end
endmodule
