module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    reg [53:0] src32;
    reg [53:0] src33;
    reg [53:0] src34;
    reg [53:0] src35;
    reg [53:0] src36;
    reg [53:0] src37;
    reg [53:0] src38;
    reg [53:0] src39;
    reg [53:0] src40;
    reg [53:0] src41;
    reg [53:0] src42;
    reg [53:0] src43;
    reg [53:0] src44;
    reg [53:0] src45;
    reg [53:0] src46;
    reg [53:0] src47;
    reg [53:0] src48;
    reg [53:0] src49;
    reg [53:0] src50;
    reg [53:0] src51;
    reg [53:0] src52;
    reg [53:0] src53;
    reg [53:0] src54;
    reg [53:0] src55;
    reg [53:0] src56;
    reg [53:0] src57;
    reg [53:0] src58;
    reg [53:0] src59;
    reg [53:0] src60;
    reg [53:0] src61;
    reg [53:0] src62;
    reg [53:0] src63;
    compressor2_1_54_64 compressor2_1_54_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
        src12 <= 54'h0;
        src13 <= 54'h0;
        src14 <= 54'h0;
        src15 <= 54'h0;
        src16 <= 54'h0;
        src17 <= 54'h0;
        src18 <= 54'h0;
        src19 <= 54'h0;
        src20 <= 54'h0;
        src21 <= 54'h0;
        src22 <= 54'h0;
        src23 <= 54'h0;
        src24 <= 54'h0;
        src25 <= 54'h0;
        src26 <= 54'h0;
        src27 <= 54'h0;
        src28 <= 54'h0;
        src29 <= 54'h0;
        src30 <= 54'h0;
        src31 <= 54'h0;
        src32 <= 54'h0;
        src33 <= 54'h0;
        src34 <= 54'h0;
        src35 <= 54'h0;
        src36 <= 54'h0;
        src37 <= 54'h0;
        src38 <= 54'h0;
        src39 <= 54'h0;
        src40 <= 54'h0;
        src41 <= 54'h0;
        src42 <= 54'h0;
        src43 <= 54'h0;
        src44 <= 54'h0;
        src45 <= 54'h0;
        src46 <= 54'h0;
        src47 <= 54'h0;
        src48 <= 54'h0;
        src49 <= 54'h0;
        src50 <= 54'h0;
        src51 <= 54'h0;
        src52 <= 54'h0;
        src53 <= 54'h0;
        src54 <= 54'h0;
        src55 <= 54'h0;
        src56 <= 54'h0;
        src57 <= 54'h0;
        src58 <= 54'h0;
        src59 <= 54'h0;
        src60 <= 54'h0;
        src61 <= 54'h0;
        src62 <= 54'h0;
        src63 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor2_1_54_64(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    input [53:0]src12,
    input [53:0]src13,
    input [53:0]src14,
    input [53:0]src15,
    input [53:0]src16,
    input [53:0]src17,
    input [53:0]src18,
    input [53:0]src19,
    input [53:0]src20,
    input [53:0]src21,
    input [53:0]src22,
    input [53:0]src23,
    input [53:0]src24,
    input [53:0]src25,
    input [53:0]src26,
    input [53:0]src27,
    input [53:0]src28,
    input [53:0]src29,
    input [53:0]src30,
    input [53:0]src31,
    input [53:0]src32,
    input [53:0]src33,
    input [53:0]src34,
    input [53:0]src35,
    input [53:0]src36,
    input [53:0]src37,
    input [53:0]src38,
    input [53:0]src39,
    input [53:0]src40,
    input [53:0]src41,
    input [53:0]src42,
    input [53:0]src43,
    input [53:0]src44,
    input [53:0]src45,
    input [53:0]src46,
    input [53:0]src47,
    input [53:0]src48,
    input [53:0]src49,
    input [53:0]src50,
    input [53:0]src51,
    input [53:0]src52,
    input [53:0]src53,
    input [53:0]src54,
    input [53:0]src55,
    input [53:0]src56,
    input [53:0]src57,
    input [53:0]src58,
    input [53:0]src59,
    input [53:0]src60,
    input [53:0]src61,
    input [53:0]src62,
    input [53:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [0:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [0:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [0:0] comp_out68;
    wire [0:0] comp_out69;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69)
    );
    rowadder2_1_70 rowadder2_1inst(
        .src0({comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], 1'h0, comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], 1'h0, comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst0({dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      input wire [53:0] src16,
      input wire [53:0] src17,
      input wire [53:0] src18,
      input wire [53:0] src19,
      input wire [53:0] src20,
      input wire [53:0] src21,
      input wire [53:0] src22,
      input wire [53:0] src23,
      input wire [53:0] src24,
      input wire [53:0] src25,
      input wire [53:0] src26,
      input wire [53:0] src27,
      input wire [53:0] src28,
      input wire [53:0] src29,
      input wire [53:0] src30,
      input wire [53:0] src31,
      input wire [53:0] src32,
      input wire [53:0] src33,
      input wire [53:0] src34,
      input wire [53:0] src35,
      input wire [53:0] src36,
      input wire [53:0] src37,
      input wire [53:0] src38,
      input wire [53:0] src39,
      input wire [53:0] src40,
      input wire [53:0] src41,
      input wire [53:0] src42,
      input wire [53:0] src43,
      input wire [53:0] src44,
      input wire [53:0] src45,
      input wire [53:0] src46,
      input wire [53:0] src47,
      input wire [53:0] src48,
      input wire [53:0] src49,
      input wire [53:0] src50,
      input wire [53:0] src51,
      input wire [53:0] src52,
      input wire [53:0] src53,
      input wire [53:0] src54,
      input wire [53:0] src55,
      input wire [53:0] src56,
      input wire [53:0] src57,
      input wire [53:0] src58,
      input wire [53:0] src59,
      input wire [53:0] src60,
      input wire [53:0] src61,
      input wire [53:0] src62,
      input wire [53:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [0:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [0:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [0:0] dst68,
      output wire [0:0] dst69);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [53:0] stage0_16;
   wire [53:0] stage0_17;
   wire [53:0] stage0_18;
   wire [53:0] stage0_19;
   wire [53:0] stage0_20;
   wire [53:0] stage0_21;
   wire [53:0] stage0_22;
   wire [53:0] stage0_23;
   wire [53:0] stage0_24;
   wire [53:0] stage0_25;
   wire [53:0] stage0_26;
   wire [53:0] stage0_27;
   wire [53:0] stage0_28;
   wire [53:0] stage0_29;
   wire [53:0] stage0_30;
   wire [53:0] stage0_31;
   wire [53:0] stage0_32;
   wire [53:0] stage0_33;
   wire [53:0] stage0_34;
   wire [53:0] stage0_35;
   wire [53:0] stage0_36;
   wire [53:0] stage0_37;
   wire [53:0] stage0_38;
   wire [53:0] stage0_39;
   wire [53:0] stage0_40;
   wire [53:0] stage0_41;
   wire [53:0] stage0_42;
   wire [53:0] stage0_43;
   wire [53:0] stage0_44;
   wire [53:0] stage0_45;
   wire [53:0] stage0_46;
   wire [53:0] stage0_47;
   wire [53:0] stage0_48;
   wire [53:0] stage0_49;
   wire [53:0] stage0_50;
   wire [53:0] stage0_51;
   wire [53:0] stage0_52;
   wire [53:0] stage0_53;
   wire [53:0] stage0_54;
   wire [53:0] stage0_55;
   wire [53:0] stage0_56;
   wire [53:0] stage0_57;
   wire [53:0] stage0_58;
   wire [53:0] stage0_59;
   wire [53:0] stage0_60;
   wire [53:0] stage0_61;
   wire [53:0] stage0_62;
   wire [53:0] stage0_63;
   wire [16:0] stage1_0;
   wire [19:0] stage1_1;
   wire [24:0] stage1_2;
   wire [23:0] stage1_3;
   wire [32:0] stage1_4;
   wire [35:0] stage1_5;
   wire [18:0] stage1_6;
   wire [24:0] stage1_7;
   wire [30:0] stage1_8;
   wire [17:0] stage1_9;
   wire [25:0] stage1_10;
   wire [28:0] stage1_11;
   wire [20:0] stage1_12;
   wire [29:0] stage1_13;
   wire [23:0] stage1_14;
   wire [42:0] stage1_15;
   wire [23:0] stage1_16;
   wire [17:0] stage1_17;
   wire [33:0] stage1_18;
   wire [20:0] stage1_19;
   wire [19:0] stage1_20;
   wire [25:0] stage1_21;
   wire [22:0] stage1_22;
   wire [21:0] stage1_23;
   wire [31:0] stage1_24;
   wire [24:0] stage1_25;
   wire [31:0] stage1_26;
   wire [23:0] stage1_27;
   wire [17:0] stage1_28;
   wire [25:0] stage1_29;
   wire [34:0] stage1_30;
   wire [33:0] stage1_31;
   wire [18:0] stage1_32;
   wire [45:0] stage1_33;
   wire [18:0] stage1_34;
   wire [27:0] stage1_35;
   wire [33:0] stage1_36;
   wire [24:0] stage1_37;
   wire [23:0] stage1_38;
   wire [30:0] stage1_39;
   wire [38:0] stage1_40;
   wire [19:0] stage1_41;
   wire [20:0] stage1_42;
   wire [22:0] stage1_43;
   wire [21:0] stage1_44;
   wire [31:0] stage1_45;
   wire [29:0] stage1_46;
   wire [33:0] stage1_47;
   wire [17:0] stage1_48;
   wire [23:0] stage1_49;
   wire [42:0] stage1_50;
   wire [47:0] stage1_51;
   wire [21:0] stage1_52;
   wire [40:0] stage1_53;
   wire [16:0] stage1_54;
   wire [37:0] stage1_55;
   wire [20:0] stage1_56;
   wire [40:0] stage1_57;
   wire [14:0] stage1_58;
   wire [34:0] stage1_59;
   wire [22:0] stage1_60;
   wire [20:0] stage1_61;
   wire [23:0] stage1_62;
   wire [34:0] stage1_63;
   wire [13:0] stage1_64;
   wire [5:0] stage1_65;
   wire [5:0] stage2_0;
   wire [6:0] stage2_1;
   wire [13:0] stage2_2;
   wire [8:0] stage2_3;
   wire [22:0] stage2_4;
   wire [9:0] stage2_5;
   wire [10:0] stage2_6;
   wire [12:0] stage2_7;
   wire [10:0] stage2_8;
   wire [19:0] stage2_9;
   wire [9:0] stage2_10;
   wire [12:0] stage2_11;
   wire [9:0] stage2_12;
   wire [9:0] stage2_13;
   wire [14:0] stage2_14;
   wire [13:0] stage2_15;
   wire [10:0] stage2_16;
   wire [11:0] stage2_17;
   wire [19:0] stage2_18;
   wire [8:0] stage2_19;
   wire [8:0] stage2_20;
   wire [21:0] stage2_21;
   wire [10:0] stage2_22;
   wire [20:0] stage2_23;
   wire [9:0] stage2_24;
   wire [12:0] stage2_25;
   wire [18:0] stage2_26;
   wire [6:0] stage2_27;
   wire [13:0] stage2_28;
   wire [17:0] stage2_29;
   wire [9:0] stage2_30;
   wire [16:0] stage2_31;
   wire [11:0] stage2_32;
   wire [15:0] stage2_33;
   wire [15:0] stage2_34;
   wire [10:0] stage2_35;
   wire [18:0] stage2_36;
   wire [16:0] stage2_37;
   wire [12:0] stage2_38;
   wire [16:0] stage2_39;
   wire [11:0] stage2_40;
   wire [12:0] stage2_41;
   wire [13:0] stage2_42;
   wire [9:0] stage2_43;
   wire [14:0] stage2_44;
   wire [11:0] stage2_45;
   wire [17:0] stage2_46;
   wire [21:0] stage2_47;
   wire [12:0] stage2_48;
   wire [17:0] stage2_49;
   wire [10:0] stage2_50;
   wire [16:0] stage2_51;
   wire [18:0] stage2_52;
   wire [12:0] stage2_53;
   wire [14:0] stage2_54;
   wire [18:0] stage2_55;
   wire [12:0] stage2_56;
   wire [12:0] stage2_57;
   wire [17:0] stage2_58;
   wire [12:0] stage2_59;
   wire [12:0] stage2_60;
   wire [11:0] stage2_61;
   wire [17:0] stage2_62;
   wire [16:0] stage2_63;
   wire [5:0] stage2_64;
   wire [9:0] stage2_65;
   wire [3:0] stage2_66;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [4:0] stage3_2;
   wire [5:0] stage3_3;
   wire [14:0] stage3_4;
   wire [8:0] stage3_5;
   wire [4:0] stage3_6;
   wire [13:0] stage3_7;
   wire [6:0] stage3_8;
   wire [10:0] stage3_9;
   wire [6:0] stage3_10;
   wire [3:0] stage3_11;
   wire [4:0] stage3_12;
   wire [7:0] stage3_13;
   wire [3:0] stage3_14;
   wire [5:0] stage3_15;
   wire [5:0] stage3_16;
   wire [7:0] stage3_17;
   wire [5:0] stage3_18;
   wire [7:0] stage3_19;
   wire [4:0] stage3_20;
   wire [6:0] stage3_21;
   wire [6:0] stage3_22;
   wire [4:0] stage3_23;
   wire [5:0] stage3_24;
   wire [7:0] stage3_25;
   wire [5:0] stage3_26;
   wire [4:0] stage3_27;
   wire [4:0] stage3_28;
   wire [11:0] stage3_29;
   wire [5:0] stage3_30;
   wire [6:0] stage3_31;
   wire [3:0] stage3_32;
   wire [14:0] stage3_33;
   wire [8:0] stage3_34;
   wire [3:0] stage3_35;
   wire [5:0] stage3_36;
   wire [6:0] stage3_37;
   wire [6:0] stage3_38;
   wire [5:0] stage3_39;
   wire [6:0] stage3_40;
   wire [6:0] stage3_41;
   wire [5:0] stage3_42;
   wire [7:0] stage3_43;
   wire [7:0] stage3_44;
   wire [4:0] stage3_45;
   wire [5:0] stage3_46;
   wire [8:0] stage3_47;
   wire [12:0] stage3_48;
   wire [5:0] stage3_49;
   wire [10:0] stage3_50;
   wire [7:0] stage3_51;
   wire [10:0] stage3_52;
   wire [6:0] stage3_53;
   wire [5:0] stage3_54;
   wire [5:0] stage3_55;
   wire [10:0] stage3_56;
   wire [7:0] stage3_57;
   wire [3:0] stage3_58;
   wire [13:0] stage3_59;
   wire [5:0] stage3_60;
   wire [9:0] stage3_61;
   wire [3:0] stage3_62;
   wire [9:0] stage3_63;
   wire [4:0] stage3_64;
   wire [6:0] stage3_65;
   wire [5:0] stage3_66;
   wire [0:0] stage3_67;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [0:0] stage4_2;
   wire [1:0] stage4_3;
   wire [5:0] stage4_4;
   wire [2:0] stage4_5;
   wire [3:0] stage4_6;
   wire [5:0] stage4_7;
   wire [3:0] stage4_8;
   wire [2:0] stage4_9;
   wire [3:0] stage4_10;
   wire [3:0] stage4_11;
   wire [3:0] stage4_12;
   wire [1:0] stage4_13;
   wire [2:0] stage4_14;
   wire [4:0] stage4_15;
   wire [3:0] stage4_16;
   wire [1:0] stage4_17;
   wire [6:0] stage4_18;
   wire [2:0] stage4_19;
   wire [2:0] stage4_20;
   wire [3:0] stage4_21;
   wire [1:0] stage4_22;
   wire [2:0] stage4_23;
   wire [2:0] stage4_24;
   wire [2:0] stage4_25;
   wire [3:0] stage4_26;
   wire [5:0] stage4_27;
   wire [0:0] stage4_28;
   wire [5:0] stage4_29;
   wire [2:0] stage4_30;
   wire [1:0] stage4_31;
   wire [2:0] stage4_32;
   wire [5:0] stage4_33;
   wire [2:0] stage4_34;
   wire [3:0] stage4_35;
   wire [2:0] stage4_36;
   wire [5:0] stage4_37;
   wire [6:0] stage4_38;
   wire [0:0] stage4_39;
   wire [2:0] stage4_40;
   wire [2:0] stage4_41;
   wire [2:0] stage4_42;
   wire [3:0] stage4_43;
   wire [5:0] stage4_44;
   wire [1:0] stage4_45;
   wire [2:0] stage4_46;
   wire [3:0] stage4_47;
   wire [3:0] stage4_48;
   wire [2:0] stage4_49;
   wire [3:0] stage4_50;
   wire [4:0] stage4_51;
   wire [3:0] stage4_52;
   wire [2:0] stage4_53;
   wire [2:0] stage4_54;
   wire [3:0] stage4_55;
   wire [5:0] stage4_56;
   wire [2:0] stage4_57;
   wire [2:0] stage4_58;
   wire [5:0] stage4_59;
   wire [2:0] stage4_60;
   wire [5:0] stage4_61;
   wire [2:0] stage4_62;
   wire [5:0] stage4_63;
   wire [2:0] stage4_64;
   wire [2:0] stage4_65;
   wire [2:0] stage4_66;
   wire [2:0] stage4_67;
   wire [0:0] stage4_68;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [0:0] stage5_2;
   wire [1:0] stage5_3;
   wire [0:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [1:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [0:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [1:0] stage5_36;
   wire [1:0] stage5_37;
   wire [1:0] stage5_38;
   wire [1:0] stage5_39;
   wire [1:0] stage5_40;
   wire [1:0] stage5_41;
   wire [1:0] stage5_42;
   wire [1:0] stage5_43;
   wire [1:0] stage5_44;
   wire [1:0] stage5_45;
   wire [1:0] stage5_46;
   wire [1:0] stage5_47;
   wire [1:0] stage5_48;
   wire [1:0] stage5_49;
   wire [1:0] stage5_50;
   wire [1:0] stage5_51;
   wire [1:0] stage5_52;
   wire [1:0] stage5_53;
   wire [1:0] stage5_54;
   wire [1:0] stage5_55;
   wire [1:0] stage5_56;
   wire [1:0] stage5_57;
   wire [1:0] stage5_58;
   wire [1:0] stage5_59;
   wire [1:0] stage5_60;
   wire [1:0] stage5_61;
   wire [1:0] stage5_62;
   wire [1:0] stage5_63;
   wire [1:0] stage5_64;
   wire [1:0] stage5_65;
   wire [1:0] stage5_66;
   wire [1:0] stage5_67;
   wire [0:0] stage5_68;
   wire [0:0] stage5_69;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;
   assign dst38 = stage5_38;
   assign dst39 = stage5_39;
   assign dst40 = stage5_40;
   assign dst41 = stage5_41;
   assign dst42 = stage5_42;
   assign dst43 = stage5_43;
   assign dst44 = stage5_44;
   assign dst45 = stage5_45;
   assign dst46 = stage5_46;
   assign dst47 = stage5_47;
   assign dst48 = stage5_48;
   assign dst49 = stage5_49;
   assign dst50 = stage5_50;
   assign dst51 = stage5_51;
   assign dst52 = stage5_52;
   assign dst53 = stage5_53;
   assign dst54 = stage5_54;
   assign dst55 = stage5_55;
   assign dst56 = stage5_56;
   assign dst57 = stage5_57;
   assign dst58 = stage5_58;
   assign dst59 = stage5_59;
   assign dst60 = stage5_60;
   assign dst61 = stage5_61;
   assign dst62 = stage5_62;
   assign dst63 = stage5_63;
   assign dst64 = stage5_64;
   assign dst65 = stage5_65;
   assign dst66 = stage5_66;
   assign dst67 = stage5_67;
   assign dst68 = stage5_68;
   assign dst69 = stage5_69;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc7_3 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15]},
      {stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage1_4[3],stage1_3[3],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[4],stage1_3[4],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[5],stage1_3[5],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[6],stage1_3[6],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[7],stage1_3[7],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[14]}
   );
   gpc606_5 gpc15 (
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[15]}
   );
   gpc615_5 gpc16 (
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[7],stage1_4[15],stage1_3[15]}
   );
   gpc615_5 gpc17 (
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage0_4[13]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[3],stage1_5[8],stage1_4[16],stage1_3[16]}
   );
   gpc615_5 gpc18 (
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage0_4[14]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[4],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc615_5 gpc19 (
      {stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_5[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[3],stage1_6[5],stage1_5[10],stage1_4[18]}
   );
   gpc615_5 gpc20 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_5[19]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[4],stage1_6[6],stage1_5[11],stage1_4[19]}
   );
   gpc615_5 gpc21 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage0_5[20]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[5],stage1_6[7],stage1_5[12],stage1_4[20]}
   );
   gpc615_5 gpc22 (
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_5[21]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[6],stage1_6[8],stage1_5[13],stage1_4[21]}
   );
   gpc615_5 gpc23 (
      {stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39]},
      {stage0_5[22]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[7],stage1_6[9],stage1_5[14],stage1_4[22]}
   );
   gpc615_5 gpc24 (
      {stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44]},
      {stage0_5[23]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[8],stage1_6[10],stage1_5[15],stage1_4[23]}
   );
   gpc606_5 gpc25 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[6],stage1_7[9],stage1_6[11],stage1_5[16]}
   );
   gpc606_5 gpc26 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[7],stage1_7[10],stage1_6[12],stage1_5[17]}
   );
   gpc615_5 gpc27 (
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40]},
      {stage0_7[12]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[2],stage1_8[8],stage1_7[11],stage1_6[13]}
   );
   gpc615_5 gpc28 (
      {stage0_6[41], stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45]},
      {stage0_7[13]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[3],stage1_8[9],stage1_7[12],stage1_6[14]}
   );
   gpc615_5 gpc29 (
      {stage0_6[46], stage0_6[47], stage0_6[48], stage0_6[49], stage0_6[50]},
      {stage0_7[14]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[4],stage1_8[10],stage1_7[13],stage1_6[15]}
   );
   gpc606_5 gpc30 (
      {stage0_7[15], stage0_7[16], stage0_7[17], stage0_7[18], stage0_7[19], stage0_7[20]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[5],stage1_8[11],stage1_7[14]}
   );
   gpc606_5 gpc31 (
      {stage0_7[21], stage0_7[22], stage0_7[23], stage0_7[24], stage0_7[25], stage0_7[26]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[6],stage1_8[12],stage1_7[15]}
   );
   gpc606_5 gpc32 (
      {stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30], stage0_7[31], stage0_7[32]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[5],stage1_9[7],stage1_8[13],stage1_7[16]}
   );
   gpc606_5 gpc33 (
      {stage0_7[33], stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37], stage0_7[38]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[6],stage1_9[8],stage1_8[14],stage1_7[17]}
   );
   gpc615_5 gpc34 (
      {stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43]},
      {stage0_8[18]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[7],stage1_9[9],stage1_8[15],stage1_7[18]}
   );
   gpc615_5 gpc35 (
      {stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47], stage0_7[48]},
      {stage0_8[19]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[8],stage1_9[10],stage1_8[16],stage1_7[19]}
   );
   gpc606_5 gpc36 (
      {stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[6],stage1_10[9],stage1_9[11],stage1_8[17]}
   );
   gpc606_5 gpc37 (
      {stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[7],stage1_10[10],stage1_9[12],stage1_8[18]}
   );
   gpc606_5 gpc38 (
      {stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[8],stage1_10[11],stage1_9[13],stage1_8[19]}
   );
   gpc606_5 gpc39 (
      {stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[9],stage1_10[12],stage1_9[14],stage1_8[20]}
   );
   gpc606_5 gpc40 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[4],stage1_11[10],stage1_10[13],stage1_9[15]}
   );
   gpc606_5 gpc41 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[5],stage1_11[11],stage1_10[14],stage1_9[16]}
   );
   gpc606_5 gpc42 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[6],stage1_11[12],stage1_10[15],stage1_9[17]}
   );
   gpc615_5 gpc43 (
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28]},
      {stage0_11[18]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[3],stage1_12[7],stage1_11[13],stage1_10[16]}
   );
   gpc615_5 gpc44 (
      {stage0_10[29], stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33]},
      {stage0_11[19]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[4],stage1_12[8],stage1_11[14],stage1_10[17]}
   );
   gpc615_5 gpc45 (
      {stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37], stage0_10[38]},
      {stage0_11[20]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[5],stage1_12[9],stage1_11[15],stage1_10[18]}
   );
   gpc615_5 gpc46 (
      {stage0_10[39], stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43]},
      {stage0_11[21]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[6],stage1_12[10],stage1_11[16],stage1_10[19]}
   );
   gpc615_5 gpc47 (
      {stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48]},
      {stage0_11[22]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[7],stage1_12[11],stage1_11[17],stage1_10[20]}
   );
   gpc615_5 gpc48 (
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27]},
      {stage0_12[30]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[5],stage1_13[8],stage1_12[12],stage1_11[18]}
   );
   gpc615_5 gpc49 (
      {stage0_11[28], stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32]},
      {stage0_12[31]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[6],stage1_13[9],stage1_12[13],stage1_11[19]}
   );
   gpc615_5 gpc50 (
      {stage0_11[33], stage0_11[34], stage0_11[35], stage0_11[36], stage0_11[37]},
      {stage0_12[32]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[7],stage1_13[10],stage1_12[14],stage1_11[20]}
   );
   gpc615_5 gpc51 (
      {stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41], stage0_11[42]},
      {stage0_12[33]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[8],stage1_13[11],stage1_12[15],stage1_11[21]}
   );
   gpc615_5 gpc52 (
      {stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage0_12[34]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[9],stage1_13[12],stage1_12[16],stage1_11[22]}
   );
   gpc606_5 gpc53 (
      {stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[5],stage1_14[10],stage1_13[13],stage1_12[17]}
   );
   gpc606_5 gpc54 (
      {stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[6],stage1_14[11],stage1_13[14],stage1_12[18]}
   );
   gpc606_5 gpc55 (
      {stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[7],stage1_14[12],stage1_13[15],stage1_12[19]}
   );
   gpc606_5 gpc56 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[3],stage1_15[8],stage1_14[13],stage1_13[16]}
   );
   gpc606_5 gpc57 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[4],stage1_15[9],stage1_14[14],stage1_13[17]}
   );
   gpc606_5 gpc58 (
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[2],stage1_16[5],stage1_15[10],stage1_14[15]}
   );
   gpc606_5 gpc59 (
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[3],stage1_16[6],stage1_15[11],stage1_14[16]}
   );
   gpc606_5 gpc60 (
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[4],stage1_16[7],stage1_15[12],stage1_14[17]}
   );
   gpc615_5 gpc61 (
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40]},
      {stage0_15[12]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[5],stage1_16[8],stage1_15[13],stage1_14[18]}
   );
   gpc615_5 gpc62 (
      {stage0_14[41], stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45]},
      {stage0_15[13]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[6],stage1_16[9],stage1_15[14],stage1_14[19]}
   );
   gpc615_5 gpc63 (
      {stage0_14[46], stage0_14[47], stage0_14[48], stage0_14[49], stage0_14[50]},
      {stage0_15[14]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[7],stage1_16[10],stage1_15[15],stage1_14[20]}
   );
   gpc615_5 gpc64 (
      {stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18], stage0_15[19]},
      {stage0_16[36]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[6],stage1_17[8],stage1_16[11],stage1_15[16]}
   );
   gpc615_5 gpc65 (
      {stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24]},
      {stage0_16[37]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[7],stage1_17[9],stage1_16[12],stage1_15[17]}
   );
   gpc615_5 gpc66 (
      {stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage0_16[38]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[8],stage1_17[10],stage1_16[13],stage1_15[18]}
   );
   gpc606_5 gpc67 (
      {stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43], stage0_16[44]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[3],stage1_18[9],stage1_17[11],stage1_16[14]}
   );
   gpc606_5 gpc68 (
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[1],stage1_19[4],stage1_18[10],stage1_17[12]}
   );
   gpc606_5 gpc69 (
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[2],stage1_19[5],stage1_18[11],stage1_17[13]}
   );
   gpc606_5 gpc70 (
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[3],stage1_19[6],stage1_18[12],stage1_17[14]}
   );
   gpc606_5 gpc71 (
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[4],stage1_19[7],stage1_18[13],stage1_17[15]}
   );
   gpc606_5 gpc72 (
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[5],stage1_19[8],stage1_18[14],stage1_17[16]}
   );
   gpc606_5 gpc73 (
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[6],stage1_19[9],stage1_18[15],stage1_17[17]}
   );
   gpc606_5 gpc74 (
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[6],stage1_20[7],stage1_19[10],stage1_18[16]}
   );
   gpc606_5 gpc75 (
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[7],stage1_20[8],stage1_19[11],stage1_18[17]}
   );
   gpc606_5 gpc76 (
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[8],stage1_20[9],stage1_19[12],stage1_18[18]}
   );
   gpc606_5 gpc77 (
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[9],stage1_20[10],stage1_19[13],stage1_18[19]}
   );
   gpc606_5 gpc78 (
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[10],stage1_20[11],stage1_19[14],stage1_18[20]}
   );
   gpc606_5 gpc79 (
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[11],stage1_20[12],stage1_19[15],stage1_18[21]}
   );
   gpc606_5 gpc80 (
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[6],stage1_21[12],stage1_20[13],stage1_19[16]}
   );
   gpc615_5 gpc81 (
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46]},
      {stage0_20[36]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[7],stage1_21[13],stage1_20[14],stage1_19[17]}
   );
   gpc615_5 gpc82 (
      {stage0_19[47], stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51]},
      {stage0_20[37]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[8],stage1_21[14],stage1_20[15],stage1_19[18]}
   );
   gpc615_5 gpc83 (
      {stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42]},
      {stage0_21[18]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[3],stage1_22[9],stage1_21[15],stage1_20[16]}
   );
   gpc615_5 gpc84 (
      {stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage0_21[19]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[4],stage1_22[10],stage1_21[16],stage1_20[17]}
   );
   gpc615_5 gpc85 (
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[20]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[5],stage1_22[11],stage1_21[17],stage1_20[18]}
   );
   gpc606_5 gpc86 (
      {stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25], stage0_21[26]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[3],stage1_23[6],stage1_22[12],stage1_21[18]}
   );
   gpc606_5 gpc87 (
      {stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31], stage0_21[32]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[4],stage1_23[7],stage1_22[13],stage1_21[19]}
   );
   gpc606_5 gpc88 (
      {stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36], stage0_21[37], stage0_21[38]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[5],stage1_23[8],stage1_22[14],stage1_21[20]}
   );
   gpc606_5 gpc89 (
      {stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43], stage0_21[44]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[6],stage1_23[9],stage1_22[15],stage1_21[21]}
   );
   gpc606_5 gpc90 (
      {stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48], stage0_21[49], stage0_21[50]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[7],stage1_23[10],stage1_22[16],stage1_21[22]}
   );
   gpc606_5 gpc91 (
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[5],stage1_24[8],stage1_23[11],stage1_22[17]}
   );
   gpc606_5 gpc92 (
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[6],stage1_24[9],stage1_23[12],stage1_22[18]}
   );
   gpc606_5 gpc93 (
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[7],stage1_24[10],stage1_23[13],stage1_22[19]}
   );
   gpc606_5 gpc94 (
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[8],stage1_24[11],stage1_23[14],stage1_22[20]}
   );
   gpc606_5 gpc95 (
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[9],stage1_24[12],stage1_23[15],stage1_22[21]}
   );
   gpc606_5 gpc96 (
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[10],stage1_24[13],stage1_23[16],stage1_22[22]}
   );
   gpc615_5 gpc97 (
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34]},
      {stage0_24[36]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[6],stage1_25[11],stage1_24[14],stage1_23[17]}
   );
   gpc615_5 gpc98 (
      {stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39]},
      {stage0_24[37]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[7],stage1_25[12],stage1_24[15],stage1_23[18]}
   );
   gpc615_5 gpc99 (
      {stage0_23[40], stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44]},
      {stage0_24[38]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[8],stage1_25[13],stage1_24[16],stage1_23[19]}
   );
   gpc615_5 gpc100 (
      {stage0_23[45], stage0_23[46], stage0_23[47], stage0_23[48], stage0_23[49]},
      {stage0_24[39]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[9],stage1_25[14],stage1_24[17],stage1_23[20]}
   );
   gpc615_5 gpc101 (
      {stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53], 1'b0},
      {stage0_24[40]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[10],stage1_25[15],stage1_24[18],stage1_23[21]}
   );
   gpc606_5 gpc102 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[0],stage1_27[5],stage1_26[11],stage1_25[16]}
   );
   gpc606_5 gpc103 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[1],stage1_27[6],stage1_26[12],stage1_25[17]}
   );
   gpc606_5 gpc104 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[2],stage1_27[7],stage1_26[13],stage1_25[18]}
   );
   gpc2135_5 gpc105 (
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4]},
      {stage0_27[18], stage0_27[19], stage0_27[20]},
      {stage0_28[0]},
      {stage0_29[0], stage0_29[1]},
      {stage1_30[0],stage1_29[3],stage1_28[3],stage1_27[8],stage1_26[14]}
   );
   gpc2135_5 gpc106 (
      {stage0_26[5], stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9]},
      {stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage0_28[1]},
      {stage0_29[2], stage0_29[3]},
      {stage1_30[1],stage1_29[4],stage1_28[4],stage1_27[9],stage1_26[15]}
   );
   gpc2135_5 gpc107 (
      {stage0_26[10], stage0_26[11], stage0_26[12], stage0_26[13], stage0_26[14]},
      {stage0_27[24], stage0_27[25], stage0_27[26]},
      {stage0_28[2]},
      {stage0_29[4], stage0_29[5]},
      {stage1_30[2],stage1_29[5],stage1_28[5],stage1_27[10],stage1_26[16]}
   );
   gpc2135_5 gpc108 (
      {stage0_26[15], stage0_26[16], stage0_26[17], stage0_26[18], stage0_26[19]},
      {stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage0_28[3]},
      {stage0_29[6], stage0_29[7]},
      {stage1_30[3],stage1_29[6],stage1_28[6],stage1_27[11],stage1_26[17]}
   );
   gpc615_5 gpc109 (
      {stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23], stage0_26[24]},
      {stage0_27[30]},
      {stage0_28[4], stage0_28[5], stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9]},
      {stage1_30[4],stage1_29[7],stage1_28[7],stage1_27[12],stage1_26[18]}
   );
   gpc615_5 gpc110 (
      {stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage0_27[31]},
      {stage0_28[10], stage0_28[11], stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15]},
      {stage1_30[5],stage1_29[8],stage1_28[8],stage1_27[13],stage1_26[19]}
   );
   gpc615_5 gpc111 (
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34]},
      {stage0_27[32]},
      {stage0_28[16], stage0_28[17], stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21]},
      {stage1_30[6],stage1_29[9],stage1_28[9],stage1_27[14],stage1_26[20]}
   );
   gpc615_5 gpc112 (
      {stage0_26[35], stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39]},
      {stage0_27[33]},
      {stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27]},
      {stage1_30[7],stage1_29[10],stage1_28[10],stage1_27[15],stage1_26[21]}
   );
   gpc615_5 gpc113 (
      {stage0_26[40], stage0_26[41], stage0_26[42], stage0_26[43], stage0_26[44]},
      {stage0_27[34]},
      {stage0_28[28], stage0_28[29], stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33]},
      {stage1_30[8],stage1_29[11],stage1_28[11],stage1_27[16],stage1_26[22]}
   );
   gpc615_5 gpc114 (
      {stage0_27[35], stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39]},
      {stage0_28[34]},
      {stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12], stage0_29[13]},
      {stage1_31[0],stage1_30[9],stage1_29[12],stage1_28[12],stage1_27[17]}
   );
   gpc615_5 gpc115 (
      {stage0_27[40], stage0_27[41], stage0_27[42], stage0_27[43], stage0_27[44]},
      {stage0_28[35]},
      {stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17], stage0_29[18], stage0_29[19]},
      {stage1_31[1],stage1_30[10],stage1_29[13],stage1_28[13],stage1_27[18]}
   );
   gpc615_5 gpc116 (
      {stage0_27[45], stage0_27[46], stage0_27[47], stage0_27[48], stage0_27[49]},
      {stage0_28[36]},
      {stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23], stage0_29[24], stage0_29[25]},
      {stage1_31[2],stage1_30[11],stage1_29[14],stage1_28[14],stage1_27[19]}
   );
   gpc606_5 gpc117 (
      {stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[3],stage1_30[12],stage1_29[15],stage1_28[15]}
   );
   gpc606_5 gpc118 (
      {stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47], stage0_28[48]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[4],stage1_30[13],stage1_29[16],stage1_28[16]}
   );
   gpc606_5 gpc119 (
      {stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53], 1'b0},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[5],stage1_30[14],stage1_29[17],stage1_28[17]}
   );
   gpc606_5 gpc120 (
      {stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29], stage0_29[30], stage0_29[31]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[3],stage1_31[6],stage1_30[15],stage1_29[18]}
   );
   gpc606_5 gpc121 (
      {stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35], stage0_29[36], stage0_29[37]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[4],stage1_31[7],stage1_30[16],stage1_29[19]}
   );
   gpc606_5 gpc122 (
      {stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41], stage0_29[42], stage0_29[43]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[5],stage1_31[8],stage1_30[17],stage1_29[20]}
   );
   gpc606_5 gpc123 (
      {stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[6],stage1_31[9],stage1_30[18],stage1_29[21]}
   );
   gpc606_5 gpc124 (
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[4],stage1_32[7],stage1_31[10],stage1_30[19]}
   );
   gpc606_5 gpc125 (
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[5],stage1_32[8],stage1_31[11],stage1_30[20]}
   );
   gpc606_5 gpc126 (
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage1_34[2],stage1_33[6],stage1_32[9],stage1_31[12],stage1_30[21]}
   );
   gpc606_5 gpc127 (
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21], stage0_32[22], stage0_32[23]},
      {stage1_34[3],stage1_33[7],stage1_32[10],stage1_31[13],stage1_30[22]}
   );
   gpc606_5 gpc128 (
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[4],stage1_33[8],stage1_32[11],stage1_31[14]}
   );
   gpc606_5 gpc129 (
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[5],stage1_33[9],stage1_32[12],stage1_31[15]}
   );
   gpc606_5 gpc130 (
      {stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27], stage0_32[28], stage0_32[29]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[2],stage1_34[6],stage1_33[10],stage1_32[13]}
   );
   gpc606_5 gpc131 (
      {stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33], stage0_32[34], stage0_32[35]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[3],stage1_34[7],stage1_33[11],stage1_32[14]}
   );
   gpc606_5 gpc132 (
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[4],stage1_34[8],stage1_33[12],stage1_32[15]}
   );
   gpc606_5 gpc133 (
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[5],stage1_34[9],stage1_33[13],stage1_32[16]}
   );
   gpc615_5 gpc134 (
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52]},
      {stage0_33[12]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[6],stage1_34[10],stage1_33[14],stage1_32[17]}
   );
   gpc606_5 gpc135 (
      {stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17], stage0_33[18]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[5],stage1_35[7],stage1_34[11],stage1_33[15]}
   );
   gpc606_5 gpc136 (
      {stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23], stage0_33[24]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[6],stage1_35[8],stage1_34[12],stage1_33[16]}
   );
   gpc117_4 gpc137 (
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35], stage0_34[36]},
      {stage0_35[12]},
      {stage0_36[0]},
      {stage1_37[2],stage1_36[7],stage1_35[9],stage1_34[13]}
   );
   gpc117_4 gpc138 (
      {stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41], stage0_34[42], stage0_34[43]},
      {stage0_35[13]},
      {stage0_36[1]},
      {stage1_37[3],stage1_36[8],stage1_35[10],stage1_34[14]}
   );
   gpc117_4 gpc139 (
      {stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47], stage0_34[48], stage0_34[49], stage0_34[50]},
      {stage0_35[14]},
      {stage0_36[2]},
      {stage1_37[4],stage1_36[9],stage1_35[11],stage1_34[15]}
   );
   gpc606_5 gpc140 (
      {stage0_35[15], stage0_35[16], stage0_35[17], stage0_35[18], stage0_35[19], stage0_35[20]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[0],stage1_37[5],stage1_36[10],stage1_35[12]}
   );
   gpc606_5 gpc141 (
      {stage0_35[21], stage0_35[22], stage0_35[23], stage0_35[24], stage0_35[25], stage0_35[26]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[1],stage1_37[6],stage1_36[11],stage1_35[13]}
   );
   gpc606_5 gpc142 (
      {stage0_35[27], stage0_35[28], stage0_35[29], stage0_35[30], stage0_35[31], stage0_35[32]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[2],stage1_37[7],stage1_36[12],stage1_35[14]}
   );
   gpc615_5 gpc143 (
      {stage0_35[33], stage0_35[34], stage0_35[35], stage0_35[36], stage0_35[37]},
      {stage0_36[3]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[3],stage1_37[8],stage1_36[13],stage1_35[15]}
   );
   gpc615_5 gpc144 (
      {stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41], stage0_35[42]},
      {stage0_36[4]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[4],stage1_37[9],stage1_36[14],stage1_35[16]}
   );
   gpc606_5 gpc145 (
      {stage0_36[5], stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[5],stage1_38[5],stage1_37[10],stage1_36[15]}
   );
   gpc606_5 gpc146 (
      {stage0_36[11], stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[6],stage1_38[6],stage1_37[11],stage1_36[16]}
   );
   gpc606_5 gpc147 (
      {stage0_36[17], stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[7],stage1_38[7],stage1_37[12],stage1_36[17]}
   );
   gpc606_5 gpc148 (
      {stage0_36[23], stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[8],stage1_38[8],stage1_37[13],stage1_36[18]}
   );
   gpc606_5 gpc149 (
      {stage0_36[29], stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[9],stage1_38[9],stage1_37[14],stage1_36[19]}
   );
   gpc606_5 gpc150 (
      {stage0_36[35], stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[10],stage1_38[10],stage1_37[15],stage1_36[20]}
   );
   gpc606_5 gpc151 (
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[6],stage1_39[11],stage1_38[11],stage1_37[16]}
   );
   gpc606_5 gpc152 (
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[7],stage1_39[12],stage1_38[12],stage1_37[17]}
   );
   gpc606_5 gpc153 (
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[8],stage1_39[13],stage1_38[13],stage1_37[18]}
   );
   gpc615_5 gpc154 (
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40]},
      {stage0_39[18]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[3],stage1_40[9],stage1_39[14],stage1_38[14]}
   );
   gpc615_5 gpc155 (
      {stage0_38[41], stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45]},
      {stage0_39[19]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[4],stage1_40[10],stage1_39[15],stage1_38[15]}
   );
   gpc606_5 gpc156 (
      {stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23], stage0_39[24], stage0_39[25]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[2],stage1_41[5],stage1_40[11],stage1_39[16]}
   );
   gpc606_5 gpc157 (
      {stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29], stage0_39[30], stage0_39[31]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[3],stage1_41[6],stage1_40[12],stage1_39[17]}
   );
   gpc606_5 gpc158 (
      {stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35], stage0_39[36], stage0_39[37]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[4],stage1_41[7],stage1_40[13],stage1_39[18]}
   );
   gpc615_5 gpc159 (
      {stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41], stage0_39[42]},
      {stage0_40[12]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[5],stage1_41[8],stage1_40[14],stage1_39[19]}
   );
   gpc1406_5 gpc160 (
      {stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17], stage0_40[18]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3]},
      {stage0_43[0]},
      {stage1_44[0],stage1_43[4],stage1_42[6],stage1_41[9],stage1_40[15]}
   );
   gpc615_5 gpc161 (
      {stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage0_41[24]},
      {stage0_42[4], stage0_42[5], stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9]},
      {stage1_44[1],stage1_43[5],stage1_42[7],stage1_41[10],stage1_40[16]}
   );
   gpc615_5 gpc162 (
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28]},
      {stage0_41[25]},
      {stage0_42[10], stage0_42[11], stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15]},
      {stage1_44[2],stage1_43[6],stage1_42[8],stage1_41[11],stage1_40[17]}
   );
   gpc615_5 gpc163 (
      {stage0_40[29], stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33]},
      {stage0_41[26]},
      {stage0_42[16], stage0_42[17], stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21]},
      {stage1_44[3],stage1_43[7],stage1_42[9],stage1_41[12],stage1_40[18]}
   );
   gpc606_5 gpc164 (
      {stage0_41[27], stage0_41[28], stage0_41[29], stage0_41[30], stage0_41[31], stage0_41[32]},
      {stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5], stage0_43[6]},
      {stage1_45[0],stage1_44[4],stage1_43[8],stage1_42[10],stage1_41[13]}
   );
   gpc606_5 gpc165 (
      {stage0_41[33], stage0_41[34], stage0_41[35], stage0_41[36], stage0_41[37], stage0_41[38]},
      {stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11], stage0_43[12]},
      {stage1_45[1],stage1_44[5],stage1_43[9],stage1_42[11],stage1_41[14]}
   );
   gpc606_5 gpc166 (
      {stage0_41[39], stage0_41[40], stage0_41[41], stage0_41[42], stage0_41[43], stage0_41[44]},
      {stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17], stage0_43[18]},
      {stage1_45[2],stage1_44[6],stage1_43[10],stage1_42[12],stage1_41[15]}
   );
   gpc606_5 gpc167 (
      {stage0_41[45], stage0_41[46], stage0_41[47], stage0_41[48], stage0_41[49], stage0_41[50]},
      {stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23], stage0_43[24]},
      {stage1_45[3],stage1_44[7],stage1_43[11],stage1_42[13],stage1_41[16]}
   );
   gpc606_5 gpc168 (
      {stage0_42[22], stage0_42[23], stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[4],stage1_44[8],stage1_43[12],stage1_42[14]}
   );
   gpc606_5 gpc169 (
      {stage0_42[28], stage0_42[29], stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[5],stage1_44[9],stage1_43[13],stage1_42[15]}
   );
   gpc606_5 gpc170 (
      {stage0_42[34], stage0_42[35], stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[6],stage1_44[10],stage1_43[14],stage1_42[16]}
   );
   gpc606_5 gpc171 (
      {stage0_42[40], stage0_42[41], stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[7],stage1_44[11],stage1_43[15],stage1_42[17]}
   );
   gpc606_5 gpc172 (
      {stage0_42[46], stage0_42[47], stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[8],stage1_44[12],stage1_43[16],stage1_42[18]}
   );
   gpc615_5 gpc173 (
      {stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage0_44[30]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[5],stage1_45[9],stage1_44[13],stage1_43[17]}
   );
   gpc615_5 gpc174 (
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34]},
      {stage0_44[31]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[6],stage1_45[10],stage1_44[14],stage1_43[18]}
   );
   gpc615_5 gpc175 (
      {stage0_43[35], stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39]},
      {stage0_44[32]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[7],stage1_45[11],stage1_44[15],stage1_43[19]}
   );
   gpc615_5 gpc176 (
      {stage0_43[40], stage0_43[41], stage0_43[42], stage0_43[43], stage0_43[44]},
      {stage0_44[33]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[8],stage1_45[12],stage1_44[16],stage1_43[20]}
   );
   gpc615_5 gpc177 (
      {stage0_43[45], stage0_43[46], stage0_43[47], stage0_43[48], stage0_43[49]},
      {stage0_44[34]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[9],stage1_45[13],stage1_44[17],stage1_43[21]}
   );
   gpc615_5 gpc178 (
      {stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53], 1'b0},
      {stage0_44[35]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[10],stage1_45[14],stage1_44[18],stage1_43[22]}
   );
   gpc606_5 gpc179 (
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[6],stage1_46[11],stage1_45[15],stage1_44[19]}
   );
   gpc606_5 gpc180 (
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[7],stage1_46[12],stage1_45[16],stage1_44[20]}
   );
   gpc606_5 gpc181 (
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[8],stage1_46[13],stage1_45[17],stage1_44[21]}
   );
   gpc615_5 gpc182 (
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40]},
      {stage0_46[18]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[3],stage1_47[9],stage1_46[14],stage1_45[18]}
   );
   gpc615_5 gpc183 (
      {stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage0_47[6]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[1],stage1_48[4],stage1_47[10],stage1_46[15]}
   );
   gpc615_5 gpc184 (
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28]},
      {stage0_47[7]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[2],stage1_48[5],stage1_47[11],stage1_46[16]}
   );
   gpc615_5 gpc185 (
      {stage0_46[29], stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33]},
      {stage0_47[8]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[3],stage1_48[6],stage1_47[12],stage1_46[17]}
   );
   gpc615_5 gpc186 (
      {stage0_46[34], stage0_46[35], stage0_46[36], stage0_46[37], stage0_46[38]},
      {stage0_47[9]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[4],stage1_48[7],stage1_47[13],stage1_46[18]}
   );
   gpc615_5 gpc187 (
      {stage0_46[39], stage0_46[40], stage0_46[41], stage0_46[42], stage0_46[43]},
      {stage0_47[10]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[5],stage1_48[8],stage1_47[14],stage1_46[19]}
   );
   gpc615_5 gpc188 (
      {stage0_47[11], stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15]},
      {stage0_48[30]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[5],stage1_49[6],stage1_48[9],stage1_47[15]}
   );
   gpc615_5 gpc189 (
      {stage0_47[16], stage0_47[17], stage0_47[18], stage0_47[19], stage0_47[20]},
      {stage0_48[31]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[6],stage1_49[7],stage1_48[10],stage1_47[16]}
   );
   gpc615_5 gpc190 (
      {stage0_47[21], stage0_47[22], stage0_47[23], stage0_47[24], stage0_47[25]},
      {stage0_48[32]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[7],stage1_49[8],stage1_48[11],stage1_47[17]}
   );
   gpc615_5 gpc191 (
      {stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29], stage0_47[30]},
      {stage0_48[33]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[8],stage1_49[9],stage1_48[12],stage1_47[18]}
   );
   gpc615_5 gpc192 (
      {stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage0_48[34]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[9],stage1_49[10],stage1_48[13],stage1_47[19]}
   );
   gpc615_5 gpc193 (
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40]},
      {stage0_48[35]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[10],stage1_49[11],stage1_48[14],stage1_47[20]}
   );
   gpc606_5 gpc194 (
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[6],stage1_50[11],stage1_49[12],stage1_48[15]}
   );
   gpc606_5 gpc195 (
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[7],stage1_50[12],stage1_49[13],stage1_48[16]}
   );
   gpc606_5 gpc196 (
      {stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[8],stage1_50[13],stage1_49[14],stage1_48[17]}
   );
   gpc606_5 gpc197 (
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[3],stage1_51[9],stage1_50[14],stage1_49[15]}
   );
   gpc615_5 gpc198 (
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46]},
      {stage0_50[18]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[4],stage1_51[10],stage1_50[15],stage1_49[16]}
   );
   gpc615_5 gpc199 (
      {stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage0_51[12]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[2],stage1_52[5],stage1_51[11],stage1_50[16]}
   );
   gpc615_5 gpc200 (
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28]},
      {stage0_51[13]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[3],stage1_52[6],stage1_51[12],stage1_50[17]}
   );
   gpc606_5 gpc201 (
      {stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17], stage0_51[18], stage0_51[19]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[2],stage1_53[4],stage1_52[7],stage1_51[13]}
   );
   gpc615_5 gpc202 (
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16]},
      {stage0_53[6]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[1],stage1_54[3],stage1_53[5],stage1_52[8]}
   );
   gpc615_5 gpc203 (
      {stage0_52[17], stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21]},
      {stage0_53[7]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[2],stage1_54[4],stage1_53[6],stage1_52[9]}
   );
   gpc615_5 gpc204 (
      {stage0_52[22], stage0_52[23], stage0_52[24], stage0_52[25], stage0_52[26]},
      {stage0_53[8]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[3],stage1_54[5],stage1_53[7],stage1_52[10]}
   );
   gpc615_5 gpc205 (
      {stage0_52[27], stage0_52[28], stage0_52[29], stage0_52[30], stage0_52[31]},
      {stage0_53[9]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[4],stage1_54[6],stage1_53[8],stage1_52[11]}
   );
   gpc615_5 gpc206 (
      {stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35], stage0_52[36]},
      {stage0_53[10]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[5],stage1_54[7],stage1_53[9],stage1_52[12]}
   );
   gpc615_5 gpc207 (
      {stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage0_53[11]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[6],stage1_54[8],stage1_53[10],stage1_52[13]}
   );
   gpc615_5 gpc208 (
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46]},
      {stage0_53[12]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[7],stage1_54[9],stage1_53[11],stage1_52[14]}
   );
   gpc615_5 gpc209 (
      {stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage0_54[42]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[7],stage1_55[8],stage1_54[10],stage1_53[12]}
   );
   gpc615_5 gpc210 (
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22]},
      {stage0_54[43]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[8],stage1_55[9],stage1_54[11],stage1_53[13]}
   );
   gpc615_5 gpc211 (
      {stage0_53[23], stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27]},
      {stage0_54[44]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[9],stage1_55[10],stage1_54[12],stage1_53[14]}
   );
   gpc606_5 gpc212 (
      {stage0_54[45], stage0_54[46], stage0_54[47], stage0_54[48], stage0_54[49], stage0_54[50]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[3],stage1_56[10],stage1_55[11],stage1_54[13]}
   );
   gpc606_5 gpc213 (
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[1],stage1_57[4],stage1_56[11],stage1_55[12]}
   );
   gpc606_5 gpc214 (
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[2],stage1_57[5],stage1_56[12],stage1_55[13]}
   );
   gpc606_5 gpc215 (
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[2],stage1_58[3],stage1_57[6],stage1_56[13]}
   );
   gpc606_5 gpc216 (
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[3],stage1_58[4],stage1_57[7],stage1_56[14]}
   );
   gpc606_5 gpc217 (
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[4],stage1_58[5],stage1_57[8],stage1_56[15]}
   );
   gpc606_5 gpc218 (
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[5],stage1_58[6],stage1_57[9],stage1_56[16]}
   );
   gpc606_5 gpc219 (
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[6],stage1_58[7],stage1_57[10],stage1_56[17]}
   );
   gpc606_5 gpc220 (
      {stage0_56[36], stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[7],stage1_58[8],stage1_57[11],stage1_56[18]}
   );
   gpc606_5 gpc221 (
      {stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[8],stage1_58[9],stage1_57[12],stage1_56[19]}
   );
   gpc606_5 gpc222 (
      {stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[9],stage1_58[10],stage1_57[13],stage1_56[20]}
   );
   gpc606_5 gpc223 (
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[8],stage1_59[10],stage1_58[11],stage1_57[14]}
   );
   gpc606_5 gpc224 (
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[9],stage1_59[11],stage1_58[12],stage1_57[15]}
   );
   gpc606_5 gpc225 (
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[10],stage1_59[12],stage1_58[13],stage1_57[16]}
   );
   gpc606_5 gpc226 (
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[3],stage1_60[11],stage1_59[13],stage1_58[14]}
   );
   gpc606_5 gpc227 (
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage1_63[0],stage1_62[1],stage1_61[4],stage1_60[12],stage1_59[14]}
   );
   gpc606_5 gpc228 (
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage1_63[1],stage1_62[2],stage1_61[5],stage1_60[13],stage1_59[15]}
   );
   gpc606_5 gpc229 (
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage1_63[2],stage1_62[3],stage1_61[6],stage1_60[14],stage1_59[16]}
   );
   gpc606_5 gpc230 (
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[3],stage1_62[4],stage1_61[7],stage1_60[15]}
   );
   gpc606_5 gpc231 (
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[4],stage1_62[5],stage1_61[8],stage1_60[16]}
   );
   gpc606_5 gpc232 (
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[5],stage1_62[6],stage1_61[9],stage1_60[17]}
   );
   gpc606_5 gpc233 (
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[6],stage1_62[7],stage1_61[10],stage1_60[18]}
   );
   gpc606_5 gpc234 (
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[7],stage1_62[8],stage1_61[11],stage1_60[19]}
   );
   gpc606_5 gpc235 (
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[8],stage1_62[9],stage1_61[12],stage1_60[20]}
   );
   gpc606_5 gpc236 (
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[9],stage1_62[10],stage1_61[13],stage1_60[21]}
   );
   gpc606_5 gpc237 (
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[10],stage1_62[11],stage1_61[14],stage1_60[22]}
   );
   gpc606_5 gpc238 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22], stage0_61[23]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[8],stage1_63[11],stage1_62[12],stage1_61[15]}
   );
   gpc606_5 gpc239 (
      {stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27], stage0_61[28], stage0_61[29]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[9],stage1_63[12],stage1_62[13],stage1_61[16]}
   );
   gpc606_5 gpc240 (
      {stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33], stage0_61[34], stage0_61[35]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[10],stage1_63[13],stage1_62[14],stage1_61[17]}
   );
   gpc606_5 gpc241 (
      {stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[11],stage1_63[14],stage1_62[15],stage1_61[18]}
   );
   gpc606_5 gpc242 (
      {stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[12],stage1_63[15],stage1_62[16],stage1_61[19]}
   );
   gpc606_5 gpc243 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52], stage0_61[53]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[13],stage1_63[16],stage1_62[17],stage1_61[20]}
   );
   gpc1_1 gpc244 (
      {stage0_0[46]},
      {stage1_0[9]}
   );
   gpc1_1 gpc245 (
      {stage0_0[47]},
      {stage1_0[10]}
   );
   gpc1_1 gpc246 (
      {stage0_0[48]},
      {stage1_0[11]}
   );
   gpc1_1 gpc247 (
      {stage0_0[49]},
      {stage1_0[12]}
   );
   gpc1_1 gpc248 (
      {stage0_0[50]},
      {stage1_0[13]}
   );
   gpc1_1 gpc249 (
      {stage0_0[51]},
      {stage1_0[14]}
   );
   gpc1_1 gpc250 (
      {stage0_0[52]},
      {stage1_0[15]}
   );
   gpc1_1 gpc251 (
      {stage0_0[53]},
      {stage1_0[16]}
   );
   gpc1_1 gpc252 (
      {stage0_1[48]},
      {stage1_1[14]}
   );
   gpc1_1 gpc253 (
      {stage0_1[49]},
      {stage1_1[15]}
   );
   gpc1_1 gpc254 (
      {stage0_1[50]},
      {stage1_1[16]}
   );
   gpc1_1 gpc255 (
      {stage0_1[51]},
      {stage1_1[17]}
   );
   gpc1_1 gpc256 (
      {stage0_1[52]},
      {stage1_1[18]}
   );
   gpc1_1 gpc257 (
      {stage0_1[53]},
      {stage1_1[19]}
   );
   gpc1_1 gpc258 (
      {stage0_2[45]},
      {stage1_2[16]}
   );
   gpc1_1 gpc259 (
      {stage0_2[46]},
      {stage1_2[17]}
   );
   gpc1_1 gpc260 (
      {stage0_2[47]},
      {stage1_2[18]}
   );
   gpc1_1 gpc261 (
      {stage0_2[48]},
      {stage1_2[19]}
   );
   gpc1_1 gpc262 (
      {stage0_2[49]},
      {stage1_2[20]}
   );
   gpc1_1 gpc263 (
      {stage0_2[50]},
      {stage1_2[21]}
   );
   gpc1_1 gpc264 (
      {stage0_2[51]},
      {stage1_2[22]}
   );
   gpc1_1 gpc265 (
      {stage0_2[52]},
      {stage1_2[23]}
   );
   gpc1_1 gpc266 (
      {stage0_2[53]},
      {stage1_2[24]}
   );
   gpc1_1 gpc267 (
      {stage0_3[48]},
      {stage1_3[18]}
   );
   gpc1_1 gpc268 (
      {stage0_3[49]},
      {stage1_3[19]}
   );
   gpc1_1 gpc269 (
      {stage0_3[50]},
      {stage1_3[20]}
   );
   gpc1_1 gpc270 (
      {stage0_3[51]},
      {stage1_3[21]}
   );
   gpc1_1 gpc271 (
      {stage0_3[52]},
      {stage1_3[22]}
   );
   gpc1_1 gpc272 (
      {stage0_3[53]},
      {stage1_3[23]}
   );
   gpc1_1 gpc273 (
      {stage0_4[45]},
      {stage1_4[24]}
   );
   gpc1_1 gpc274 (
      {stage0_4[46]},
      {stage1_4[25]}
   );
   gpc1_1 gpc275 (
      {stage0_4[47]},
      {stage1_4[26]}
   );
   gpc1_1 gpc276 (
      {stage0_4[48]},
      {stage1_4[27]}
   );
   gpc1_1 gpc277 (
      {stage0_4[49]},
      {stage1_4[28]}
   );
   gpc1_1 gpc278 (
      {stage0_4[50]},
      {stage1_4[29]}
   );
   gpc1_1 gpc279 (
      {stage0_4[51]},
      {stage1_4[30]}
   );
   gpc1_1 gpc280 (
      {stage0_4[52]},
      {stage1_4[31]}
   );
   gpc1_1 gpc281 (
      {stage0_4[53]},
      {stage1_4[32]}
   );
   gpc1_1 gpc282 (
      {stage0_5[36]},
      {stage1_5[18]}
   );
   gpc1_1 gpc283 (
      {stage0_5[37]},
      {stage1_5[19]}
   );
   gpc1_1 gpc284 (
      {stage0_5[38]},
      {stage1_5[20]}
   );
   gpc1_1 gpc285 (
      {stage0_5[39]},
      {stage1_5[21]}
   );
   gpc1_1 gpc286 (
      {stage0_5[40]},
      {stage1_5[22]}
   );
   gpc1_1 gpc287 (
      {stage0_5[41]},
      {stage1_5[23]}
   );
   gpc1_1 gpc288 (
      {stage0_5[42]},
      {stage1_5[24]}
   );
   gpc1_1 gpc289 (
      {stage0_5[43]},
      {stage1_5[25]}
   );
   gpc1_1 gpc290 (
      {stage0_5[44]},
      {stage1_5[26]}
   );
   gpc1_1 gpc291 (
      {stage0_5[45]},
      {stage1_5[27]}
   );
   gpc1_1 gpc292 (
      {stage0_5[46]},
      {stage1_5[28]}
   );
   gpc1_1 gpc293 (
      {stage0_5[47]},
      {stage1_5[29]}
   );
   gpc1_1 gpc294 (
      {stage0_5[48]},
      {stage1_5[30]}
   );
   gpc1_1 gpc295 (
      {stage0_5[49]},
      {stage1_5[31]}
   );
   gpc1_1 gpc296 (
      {stage0_5[50]},
      {stage1_5[32]}
   );
   gpc1_1 gpc297 (
      {stage0_5[51]},
      {stage1_5[33]}
   );
   gpc1_1 gpc298 (
      {stage0_5[52]},
      {stage1_5[34]}
   );
   gpc1_1 gpc299 (
      {stage0_5[53]},
      {stage1_5[35]}
   );
   gpc1_1 gpc300 (
      {stage0_6[51]},
      {stage1_6[16]}
   );
   gpc1_1 gpc301 (
      {stage0_6[52]},
      {stage1_6[17]}
   );
   gpc1_1 gpc302 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc303 (
      {stage0_7[49]},
      {stage1_7[20]}
   );
   gpc1_1 gpc304 (
      {stage0_7[50]},
      {stage1_7[21]}
   );
   gpc1_1 gpc305 (
      {stage0_7[51]},
      {stage1_7[22]}
   );
   gpc1_1 gpc306 (
      {stage0_7[52]},
      {stage1_7[23]}
   );
   gpc1_1 gpc307 (
      {stage0_7[53]},
      {stage1_7[24]}
   );
   gpc1_1 gpc308 (
      {stage0_8[44]},
      {stage1_8[21]}
   );
   gpc1_1 gpc309 (
      {stage0_8[45]},
      {stage1_8[22]}
   );
   gpc1_1 gpc310 (
      {stage0_8[46]},
      {stage1_8[23]}
   );
   gpc1_1 gpc311 (
      {stage0_8[47]},
      {stage1_8[24]}
   );
   gpc1_1 gpc312 (
      {stage0_8[48]},
      {stage1_8[25]}
   );
   gpc1_1 gpc313 (
      {stage0_8[49]},
      {stage1_8[26]}
   );
   gpc1_1 gpc314 (
      {stage0_8[50]},
      {stage1_8[27]}
   );
   gpc1_1 gpc315 (
      {stage0_8[51]},
      {stage1_8[28]}
   );
   gpc1_1 gpc316 (
      {stage0_8[52]},
      {stage1_8[29]}
   );
   gpc1_1 gpc317 (
      {stage0_8[53]},
      {stage1_8[30]}
   );
   gpc1_1 gpc318 (
      {stage0_10[49]},
      {stage1_10[21]}
   );
   gpc1_1 gpc319 (
      {stage0_10[50]},
      {stage1_10[22]}
   );
   gpc1_1 gpc320 (
      {stage0_10[51]},
      {stage1_10[23]}
   );
   gpc1_1 gpc321 (
      {stage0_10[52]},
      {stage1_10[24]}
   );
   gpc1_1 gpc322 (
      {stage0_10[53]},
      {stage1_10[25]}
   );
   gpc1_1 gpc323 (
      {stage0_11[48]},
      {stage1_11[23]}
   );
   gpc1_1 gpc324 (
      {stage0_11[49]},
      {stage1_11[24]}
   );
   gpc1_1 gpc325 (
      {stage0_11[50]},
      {stage1_11[25]}
   );
   gpc1_1 gpc326 (
      {stage0_11[51]},
      {stage1_11[26]}
   );
   gpc1_1 gpc327 (
      {stage0_11[52]},
      {stage1_11[27]}
   );
   gpc1_1 gpc328 (
      {stage0_11[53]},
      {stage1_11[28]}
   );
   gpc1_1 gpc329 (
      {stage0_12[53]},
      {stage1_12[20]}
   );
   gpc1_1 gpc330 (
      {stage0_13[42]},
      {stage1_13[18]}
   );
   gpc1_1 gpc331 (
      {stage0_13[43]},
      {stage1_13[19]}
   );
   gpc1_1 gpc332 (
      {stage0_13[44]},
      {stage1_13[20]}
   );
   gpc1_1 gpc333 (
      {stage0_13[45]},
      {stage1_13[21]}
   );
   gpc1_1 gpc334 (
      {stage0_13[46]},
      {stage1_13[22]}
   );
   gpc1_1 gpc335 (
      {stage0_13[47]},
      {stage1_13[23]}
   );
   gpc1_1 gpc336 (
      {stage0_13[48]},
      {stage1_13[24]}
   );
   gpc1_1 gpc337 (
      {stage0_13[49]},
      {stage1_13[25]}
   );
   gpc1_1 gpc338 (
      {stage0_13[50]},
      {stage1_13[26]}
   );
   gpc1_1 gpc339 (
      {stage0_13[51]},
      {stage1_13[27]}
   );
   gpc1_1 gpc340 (
      {stage0_13[52]},
      {stage1_13[28]}
   );
   gpc1_1 gpc341 (
      {stage0_13[53]},
      {stage1_13[29]}
   );
   gpc1_1 gpc342 (
      {stage0_14[51]},
      {stage1_14[21]}
   );
   gpc1_1 gpc343 (
      {stage0_14[52]},
      {stage1_14[22]}
   );
   gpc1_1 gpc344 (
      {stage0_14[53]},
      {stage1_14[23]}
   );
   gpc1_1 gpc345 (
      {stage0_15[30]},
      {stage1_15[19]}
   );
   gpc1_1 gpc346 (
      {stage0_15[31]},
      {stage1_15[20]}
   );
   gpc1_1 gpc347 (
      {stage0_15[32]},
      {stage1_15[21]}
   );
   gpc1_1 gpc348 (
      {stage0_15[33]},
      {stage1_15[22]}
   );
   gpc1_1 gpc349 (
      {stage0_15[34]},
      {stage1_15[23]}
   );
   gpc1_1 gpc350 (
      {stage0_15[35]},
      {stage1_15[24]}
   );
   gpc1_1 gpc351 (
      {stage0_15[36]},
      {stage1_15[25]}
   );
   gpc1_1 gpc352 (
      {stage0_15[37]},
      {stage1_15[26]}
   );
   gpc1_1 gpc353 (
      {stage0_15[38]},
      {stage1_15[27]}
   );
   gpc1_1 gpc354 (
      {stage0_15[39]},
      {stage1_15[28]}
   );
   gpc1_1 gpc355 (
      {stage0_15[40]},
      {stage1_15[29]}
   );
   gpc1_1 gpc356 (
      {stage0_15[41]},
      {stage1_15[30]}
   );
   gpc1_1 gpc357 (
      {stage0_15[42]},
      {stage1_15[31]}
   );
   gpc1_1 gpc358 (
      {stage0_15[43]},
      {stage1_15[32]}
   );
   gpc1_1 gpc359 (
      {stage0_15[44]},
      {stage1_15[33]}
   );
   gpc1_1 gpc360 (
      {stage0_15[45]},
      {stage1_15[34]}
   );
   gpc1_1 gpc361 (
      {stage0_15[46]},
      {stage1_15[35]}
   );
   gpc1_1 gpc362 (
      {stage0_15[47]},
      {stage1_15[36]}
   );
   gpc1_1 gpc363 (
      {stage0_15[48]},
      {stage1_15[37]}
   );
   gpc1_1 gpc364 (
      {stage0_15[49]},
      {stage1_15[38]}
   );
   gpc1_1 gpc365 (
      {stage0_15[50]},
      {stage1_15[39]}
   );
   gpc1_1 gpc366 (
      {stage0_15[51]},
      {stage1_15[40]}
   );
   gpc1_1 gpc367 (
      {stage0_15[52]},
      {stage1_15[41]}
   );
   gpc1_1 gpc368 (
      {stage0_15[53]},
      {stage1_15[42]}
   );
   gpc1_1 gpc369 (
      {stage0_16[45]},
      {stage1_16[15]}
   );
   gpc1_1 gpc370 (
      {stage0_16[46]},
      {stage1_16[16]}
   );
   gpc1_1 gpc371 (
      {stage0_16[47]},
      {stage1_16[17]}
   );
   gpc1_1 gpc372 (
      {stage0_16[48]},
      {stage1_16[18]}
   );
   gpc1_1 gpc373 (
      {stage0_16[49]},
      {stage1_16[19]}
   );
   gpc1_1 gpc374 (
      {stage0_16[50]},
      {stage1_16[20]}
   );
   gpc1_1 gpc375 (
      {stage0_16[51]},
      {stage1_16[21]}
   );
   gpc1_1 gpc376 (
      {stage0_16[52]},
      {stage1_16[22]}
   );
   gpc1_1 gpc377 (
      {stage0_16[53]},
      {stage1_16[23]}
   );
   gpc1_1 gpc378 (
      {stage0_18[42]},
      {stage1_18[22]}
   );
   gpc1_1 gpc379 (
      {stage0_18[43]},
      {stage1_18[23]}
   );
   gpc1_1 gpc380 (
      {stage0_18[44]},
      {stage1_18[24]}
   );
   gpc1_1 gpc381 (
      {stage0_18[45]},
      {stage1_18[25]}
   );
   gpc1_1 gpc382 (
      {stage0_18[46]},
      {stage1_18[26]}
   );
   gpc1_1 gpc383 (
      {stage0_18[47]},
      {stage1_18[27]}
   );
   gpc1_1 gpc384 (
      {stage0_18[48]},
      {stage1_18[28]}
   );
   gpc1_1 gpc385 (
      {stage0_18[49]},
      {stage1_18[29]}
   );
   gpc1_1 gpc386 (
      {stage0_18[50]},
      {stage1_18[30]}
   );
   gpc1_1 gpc387 (
      {stage0_18[51]},
      {stage1_18[31]}
   );
   gpc1_1 gpc388 (
      {stage0_18[52]},
      {stage1_18[32]}
   );
   gpc1_1 gpc389 (
      {stage0_18[53]},
      {stage1_18[33]}
   );
   gpc1_1 gpc390 (
      {stage0_19[52]},
      {stage1_19[19]}
   );
   gpc1_1 gpc391 (
      {stage0_19[53]},
      {stage1_19[20]}
   );
   gpc1_1 gpc392 (
      {stage0_20[53]},
      {stage1_20[19]}
   );
   gpc1_1 gpc393 (
      {stage0_21[51]},
      {stage1_21[23]}
   );
   gpc1_1 gpc394 (
      {stage0_21[52]},
      {stage1_21[24]}
   );
   gpc1_1 gpc395 (
      {stage0_21[53]},
      {stage1_21[25]}
   );
   gpc1_1 gpc396 (
      {stage0_24[41]},
      {stage1_24[19]}
   );
   gpc1_1 gpc397 (
      {stage0_24[42]},
      {stage1_24[20]}
   );
   gpc1_1 gpc398 (
      {stage0_24[43]},
      {stage1_24[21]}
   );
   gpc1_1 gpc399 (
      {stage0_24[44]},
      {stage1_24[22]}
   );
   gpc1_1 gpc400 (
      {stage0_24[45]},
      {stage1_24[23]}
   );
   gpc1_1 gpc401 (
      {stage0_24[46]},
      {stage1_24[24]}
   );
   gpc1_1 gpc402 (
      {stage0_24[47]},
      {stage1_24[25]}
   );
   gpc1_1 gpc403 (
      {stage0_24[48]},
      {stage1_24[26]}
   );
   gpc1_1 gpc404 (
      {stage0_24[49]},
      {stage1_24[27]}
   );
   gpc1_1 gpc405 (
      {stage0_24[50]},
      {stage1_24[28]}
   );
   gpc1_1 gpc406 (
      {stage0_24[51]},
      {stage1_24[29]}
   );
   gpc1_1 gpc407 (
      {stage0_24[52]},
      {stage1_24[30]}
   );
   gpc1_1 gpc408 (
      {stage0_24[53]},
      {stage1_24[31]}
   );
   gpc1_1 gpc409 (
      {stage0_25[48]},
      {stage1_25[19]}
   );
   gpc1_1 gpc410 (
      {stage0_25[49]},
      {stage1_25[20]}
   );
   gpc1_1 gpc411 (
      {stage0_25[50]},
      {stage1_25[21]}
   );
   gpc1_1 gpc412 (
      {stage0_25[51]},
      {stage1_25[22]}
   );
   gpc1_1 gpc413 (
      {stage0_25[52]},
      {stage1_25[23]}
   );
   gpc1_1 gpc414 (
      {stage0_25[53]},
      {stage1_25[24]}
   );
   gpc1_1 gpc415 (
      {stage0_26[45]},
      {stage1_26[23]}
   );
   gpc1_1 gpc416 (
      {stage0_26[46]},
      {stage1_26[24]}
   );
   gpc1_1 gpc417 (
      {stage0_26[47]},
      {stage1_26[25]}
   );
   gpc1_1 gpc418 (
      {stage0_26[48]},
      {stage1_26[26]}
   );
   gpc1_1 gpc419 (
      {stage0_26[49]},
      {stage1_26[27]}
   );
   gpc1_1 gpc420 (
      {stage0_26[50]},
      {stage1_26[28]}
   );
   gpc1_1 gpc421 (
      {stage0_26[51]},
      {stage1_26[29]}
   );
   gpc1_1 gpc422 (
      {stage0_26[52]},
      {stage1_26[30]}
   );
   gpc1_1 gpc423 (
      {stage0_26[53]},
      {stage1_26[31]}
   );
   gpc1_1 gpc424 (
      {stage0_27[50]},
      {stage1_27[20]}
   );
   gpc1_1 gpc425 (
      {stage0_27[51]},
      {stage1_27[21]}
   );
   gpc1_1 gpc426 (
      {stage0_27[52]},
      {stage1_27[22]}
   );
   gpc1_1 gpc427 (
      {stage0_27[53]},
      {stage1_27[23]}
   );
   gpc1_1 gpc428 (
      {stage0_29[50]},
      {stage1_29[22]}
   );
   gpc1_1 gpc429 (
      {stage0_29[51]},
      {stage1_29[23]}
   );
   gpc1_1 gpc430 (
      {stage0_29[52]},
      {stage1_29[24]}
   );
   gpc1_1 gpc431 (
      {stage0_29[53]},
      {stage1_29[25]}
   );
   gpc1_1 gpc432 (
      {stage0_30[42]},
      {stage1_30[23]}
   );
   gpc1_1 gpc433 (
      {stage0_30[43]},
      {stage1_30[24]}
   );
   gpc1_1 gpc434 (
      {stage0_30[44]},
      {stage1_30[25]}
   );
   gpc1_1 gpc435 (
      {stage0_30[45]},
      {stage1_30[26]}
   );
   gpc1_1 gpc436 (
      {stage0_30[46]},
      {stage1_30[27]}
   );
   gpc1_1 gpc437 (
      {stage0_30[47]},
      {stage1_30[28]}
   );
   gpc1_1 gpc438 (
      {stage0_30[48]},
      {stage1_30[29]}
   );
   gpc1_1 gpc439 (
      {stage0_30[49]},
      {stage1_30[30]}
   );
   gpc1_1 gpc440 (
      {stage0_30[50]},
      {stage1_30[31]}
   );
   gpc1_1 gpc441 (
      {stage0_30[51]},
      {stage1_30[32]}
   );
   gpc1_1 gpc442 (
      {stage0_30[52]},
      {stage1_30[33]}
   );
   gpc1_1 gpc443 (
      {stage0_30[53]},
      {stage1_30[34]}
   );
   gpc1_1 gpc444 (
      {stage0_31[36]},
      {stage1_31[16]}
   );
   gpc1_1 gpc445 (
      {stage0_31[37]},
      {stage1_31[17]}
   );
   gpc1_1 gpc446 (
      {stage0_31[38]},
      {stage1_31[18]}
   );
   gpc1_1 gpc447 (
      {stage0_31[39]},
      {stage1_31[19]}
   );
   gpc1_1 gpc448 (
      {stage0_31[40]},
      {stage1_31[20]}
   );
   gpc1_1 gpc449 (
      {stage0_31[41]},
      {stage1_31[21]}
   );
   gpc1_1 gpc450 (
      {stage0_31[42]},
      {stage1_31[22]}
   );
   gpc1_1 gpc451 (
      {stage0_31[43]},
      {stage1_31[23]}
   );
   gpc1_1 gpc452 (
      {stage0_31[44]},
      {stage1_31[24]}
   );
   gpc1_1 gpc453 (
      {stage0_31[45]},
      {stage1_31[25]}
   );
   gpc1_1 gpc454 (
      {stage0_31[46]},
      {stage1_31[26]}
   );
   gpc1_1 gpc455 (
      {stage0_31[47]},
      {stage1_31[27]}
   );
   gpc1_1 gpc456 (
      {stage0_31[48]},
      {stage1_31[28]}
   );
   gpc1_1 gpc457 (
      {stage0_31[49]},
      {stage1_31[29]}
   );
   gpc1_1 gpc458 (
      {stage0_31[50]},
      {stage1_31[30]}
   );
   gpc1_1 gpc459 (
      {stage0_31[51]},
      {stage1_31[31]}
   );
   gpc1_1 gpc460 (
      {stage0_31[52]},
      {stage1_31[32]}
   );
   gpc1_1 gpc461 (
      {stage0_31[53]},
      {stage1_31[33]}
   );
   gpc1_1 gpc462 (
      {stage0_32[53]},
      {stage1_32[18]}
   );
   gpc1_1 gpc463 (
      {stage0_33[25]},
      {stage1_33[17]}
   );
   gpc1_1 gpc464 (
      {stage0_33[26]},
      {stage1_33[18]}
   );
   gpc1_1 gpc465 (
      {stage0_33[27]},
      {stage1_33[19]}
   );
   gpc1_1 gpc466 (
      {stage0_33[28]},
      {stage1_33[20]}
   );
   gpc1_1 gpc467 (
      {stage0_33[29]},
      {stage1_33[21]}
   );
   gpc1_1 gpc468 (
      {stage0_33[30]},
      {stage1_33[22]}
   );
   gpc1_1 gpc469 (
      {stage0_33[31]},
      {stage1_33[23]}
   );
   gpc1_1 gpc470 (
      {stage0_33[32]},
      {stage1_33[24]}
   );
   gpc1_1 gpc471 (
      {stage0_33[33]},
      {stage1_33[25]}
   );
   gpc1_1 gpc472 (
      {stage0_33[34]},
      {stage1_33[26]}
   );
   gpc1_1 gpc473 (
      {stage0_33[35]},
      {stage1_33[27]}
   );
   gpc1_1 gpc474 (
      {stage0_33[36]},
      {stage1_33[28]}
   );
   gpc1_1 gpc475 (
      {stage0_33[37]},
      {stage1_33[29]}
   );
   gpc1_1 gpc476 (
      {stage0_33[38]},
      {stage1_33[30]}
   );
   gpc1_1 gpc477 (
      {stage0_33[39]},
      {stage1_33[31]}
   );
   gpc1_1 gpc478 (
      {stage0_33[40]},
      {stage1_33[32]}
   );
   gpc1_1 gpc479 (
      {stage0_33[41]},
      {stage1_33[33]}
   );
   gpc1_1 gpc480 (
      {stage0_33[42]},
      {stage1_33[34]}
   );
   gpc1_1 gpc481 (
      {stage0_33[43]},
      {stage1_33[35]}
   );
   gpc1_1 gpc482 (
      {stage0_33[44]},
      {stage1_33[36]}
   );
   gpc1_1 gpc483 (
      {stage0_33[45]},
      {stage1_33[37]}
   );
   gpc1_1 gpc484 (
      {stage0_33[46]},
      {stage1_33[38]}
   );
   gpc1_1 gpc485 (
      {stage0_33[47]},
      {stage1_33[39]}
   );
   gpc1_1 gpc486 (
      {stage0_33[48]},
      {stage1_33[40]}
   );
   gpc1_1 gpc487 (
      {stage0_33[49]},
      {stage1_33[41]}
   );
   gpc1_1 gpc488 (
      {stage0_33[50]},
      {stage1_33[42]}
   );
   gpc1_1 gpc489 (
      {stage0_33[51]},
      {stage1_33[43]}
   );
   gpc1_1 gpc490 (
      {stage0_33[52]},
      {stage1_33[44]}
   );
   gpc1_1 gpc491 (
      {stage0_33[53]},
      {stage1_33[45]}
   );
   gpc1_1 gpc492 (
      {stage0_34[51]},
      {stage1_34[16]}
   );
   gpc1_1 gpc493 (
      {stage0_34[52]},
      {stage1_34[17]}
   );
   gpc1_1 gpc494 (
      {stage0_34[53]},
      {stage1_34[18]}
   );
   gpc1_1 gpc495 (
      {stage0_35[43]},
      {stage1_35[17]}
   );
   gpc1_1 gpc496 (
      {stage0_35[44]},
      {stage1_35[18]}
   );
   gpc1_1 gpc497 (
      {stage0_35[45]},
      {stage1_35[19]}
   );
   gpc1_1 gpc498 (
      {stage0_35[46]},
      {stage1_35[20]}
   );
   gpc1_1 gpc499 (
      {stage0_35[47]},
      {stage1_35[21]}
   );
   gpc1_1 gpc500 (
      {stage0_35[48]},
      {stage1_35[22]}
   );
   gpc1_1 gpc501 (
      {stage0_35[49]},
      {stage1_35[23]}
   );
   gpc1_1 gpc502 (
      {stage0_35[50]},
      {stage1_35[24]}
   );
   gpc1_1 gpc503 (
      {stage0_35[51]},
      {stage1_35[25]}
   );
   gpc1_1 gpc504 (
      {stage0_35[52]},
      {stage1_35[26]}
   );
   gpc1_1 gpc505 (
      {stage0_35[53]},
      {stage1_35[27]}
   );
   gpc1_1 gpc506 (
      {stage0_36[41]},
      {stage1_36[21]}
   );
   gpc1_1 gpc507 (
      {stage0_36[42]},
      {stage1_36[22]}
   );
   gpc1_1 gpc508 (
      {stage0_36[43]},
      {stage1_36[23]}
   );
   gpc1_1 gpc509 (
      {stage0_36[44]},
      {stage1_36[24]}
   );
   gpc1_1 gpc510 (
      {stage0_36[45]},
      {stage1_36[25]}
   );
   gpc1_1 gpc511 (
      {stage0_36[46]},
      {stage1_36[26]}
   );
   gpc1_1 gpc512 (
      {stage0_36[47]},
      {stage1_36[27]}
   );
   gpc1_1 gpc513 (
      {stage0_36[48]},
      {stage1_36[28]}
   );
   gpc1_1 gpc514 (
      {stage0_36[49]},
      {stage1_36[29]}
   );
   gpc1_1 gpc515 (
      {stage0_36[50]},
      {stage1_36[30]}
   );
   gpc1_1 gpc516 (
      {stage0_36[51]},
      {stage1_36[31]}
   );
   gpc1_1 gpc517 (
      {stage0_36[52]},
      {stage1_36[32]}
   );
   gpc1_1 gpc518 (
      {stage0_36[53]},
      {stage1_36[33]}
   );
   gpc1_1 gpc519 (
      {stage0_37[48]},
      {stage1_37[19]}
   );
   gpc1_1 gpc520 (
      {stage0_37[49]},
      {stage1_37[20]}
   );
   gpc1_1 gpc521 (
      {stage0_37[50]},
      {stage1_37[21]}
   );
   gpc1_1 gpc522 (
      {stage0_37[51]},
      {stage1_37[22]}
   );
   gpc1_1 gpc523 (
      {stage0_37[52]},
      {stage1_37[23]}
   );
   gpc1_1 gpc524 (
      {stage0_37[53]},
      {stage1_37[24]}
   );
   gpc1_1 gpc525 (
      {stage0_38[46]},
      {stage1_38[16]}
   );
   gpc1_1 gpc526 (
      {stage0_38[47]},
      {stage1_38[17]}
   );
   gpc1_1 gpc527 (
      {stage0_38[48]},
      {stage1_38[18]}
   );
   gpc1_1 gpc528 (
      {stage0_38[49]},
      {stage1_38[19]}
   );
   gpc1_1 gpc529 (
      {stage0_38[50]},
      {stage1_38[20]}
   );
   gpc1_1 gpc530 (
      {stage0_38[51]},
      {stage1_38[21]}
   );
   gpc1_1 gpc531 (
      {stage0_38[52]},
      {stage1_38[22]}
   );
   gpc1_1 gpc532 (
      {stage0_38[53]},
      {stage1_38[23]}
   );
   gpc1_1 gpc533 (
      {stage0_39[43]},
      {stage1_39[20]}
   );
   gpc1_1 gpc534 (
      {stage0_39[44]},
      {stage1_39[21]}
   );
   gpc1_1 gpc535 (
      {stage0_39[45]},
      {stage1_39[22]}
   );
   gpc1_1 gpc536 (
      {stage0_39[46]},
      {stage1_39[23]}
   );
   gpc1_1 gpc537 (
      {stage0_39[47]},
      {stage1_39[24]}
   );
   gpc1_1 gpc538 (
      {stage0_39[48]},
      {stage1_39[25]}
   );
   gpc1_1 gpc539 (
      {stage0_39[49]},
      {stage1_39[26]}
   );
   gpc1_1 gpc540 (
      {stage0_39[50]},
      {stage1_39[27]}
   );
   gpc1_1 gpc541 (
      {stage0_39[51]},
      {stage1_39[28]}
   );
   gpc1_1 gpc542 (
      {stage0_39[52]},
      {stage1_39[29]}
   );
   gpc1_1 gpc543 (
      {stage0_39[53]},
      {stage1_39[30]}
   );
   gpc1_1 gpc544 (
      {stage0_40[34]},
      {stage1_40[19]}
   );
   gpc1_1 gpc545 (
      {stage0_40[35]},
      {stage1_40[20]}
   );
   gpc1_1 gpc546 (
      {stage0_40[36]},
      {stage1_40[21]}
   );
   gpc1_1 gpc547 (
      {stage0_40[37]},
      {stage1_40[22]}
   );
   gpc1_1 gpc548 (
      {stage0_40[38]},
      {stage1_40[23]}
   );
   gpc1_1 gpc549 (
      {stage0_40[39]},
      {stage1_40[24]}
   );
   gpc1_1 gpc550 (
      {stage0_40[40]},
      {stage1_40[25]}
   );
   gpc1_1 gpc551 (
      {stage0_40[41]},
      {stage1_40[26]}
   );
   gpc1_1 gpc552 (
      {stage0_40[42]},
      {stage1_40[27]}
   );
   gpc1_1 gpc553 (
      {stage0_40[43]},
      {stage1_40[28]}
   );
   gpc1_1 gpc554 (
      {stage0_40[44]},
      {stage1_40[29]}
   );
   gpc1_1 gpc555 (
      {stage0_40[45]},
      {stage1_40[30]}
   );
   gpc1_1 gpc556 (
      {stage0_40[46]},
      {stage1_40[31]}
   );
   gpc1_1 gpc557 (
      {stage0_40[47]},
      {stage1_40[32]}
   );
   gpc1_1 gpc558 (
      {stage0_40[48]},
      {stage1_40[33]}
   );
   gpc1_1 gpc559 (
      {stage0_40[49]},
      {stage1_40[34]}
   );
   gpc1_1 gpc560 (
      {stage0_40[50]},
      {stage1_40[35]}
   );
   gpc1_1 gpc561 (
      {stage0_40[51]},
      {stage1_40[36]}
   );
   gpc1_1 gpc562 (
      {stage0_40[52]},
      {stage1_40[37]}
   );
   gpc1_1 gpc563 (
      {stage0_40[53]},
      {stage1_40[38]}
   );
   gpc1_1 gpc564 (
      {stage0_41[51]},
      {stage1_41[17]}
   );
   gpc1_1 gpc565 (
      {stage0_41[52]},
      {stage1_41[18]}
   );
   gpc1_1 gpc566 (
      {stage0_41[53]},
      {stage1_41[19]}
   );
   gpc1_1 gpc567 (
      {stage0_42[52]},
      {stage1_42[19]}
   );
   gpc1_1 gpc568 (
      {stage0_42[53]},
      {stage1_42[20]}
   );
   gpc1_1 gpc569 (
      {stage0_45[41]},
      {stage1_45[19]}
   );
   gpc1_1 gpc570 (
      {stage0_45[42]},
      {stage1_45[20]}
   );
   gpc1_1 gpc571 (
      {stage0_45[43]},
      {stage1_45[21]}
   );
   gpc1_1 gpc572 (
      {stage0_45[44]},
      {stage1_45[22]}
   );
   gpc1_1 gpc573 (
      {stage0_45[45]},
      {stage1_45[23]}
   );
   gpc1_1 gpc574 (
      {stage0_45[46]},
      {stage1_45[24]}
   );
   gpc1_1 gpc575 (
      {stage0_45[47]},
      {stage1_45[25]}
   );
   gpc1_1 gpc576 (
      {stage0_45[48]},
      {stage1_45[26]}
   );
   gpc1_1 gpc577 (
      {stage0_45[49]},
      {stage1_45[27]}
   );
   gpc1_1 gpc578 (
      {stage0_45[50]},
      {stage1_45[28]}
   );
   gpc1_1 gpc579 (
      {stage0_45[51]},
      {stage1_45[29]}
   );
   gpc1_1 gpc580 (
      {stage0_45[52]},
      {stage1_45[30]}
   );
   gpc1_1 gpc581 (
      {stage0_45[53]},
      {stage1_45[31]}
   );
   gpc1_1 gpc582 (
      {stage0_46[44]},
      {stage1_46[20]}
   );
   gpc1_1 gpc583 (
      {stage0_46[45]},
      {stage1_46[21]}
   );
   gpc1_1 gpc584 (
      {stage0_46[46]},
      {stage1_46[22]}
   );
   gpc1_1 gpc585 (
      {stage0_46[47]},
      {stage1_46[23]}
   );
   gpc1_1 gpc586 (
      {stage0_46[48]},
      {stage1_46[24]}
   );
   gpc1_1 gpc587 (
      {stage0_46[49]},
      {stage1_46[25]}
   );
   gpc1_1 gpc588 (
      {stage0_46[50]},
      {stage1_46[26]}
   );
   gpc1_1 gpc589 (
      {stage0_46[51]},
      {stage1_46[27]}
   );
   gpc1_1 gpc590 (
      {stage0_46[52]},
      {stage1_46[28]}
   );
   gpc1_1 gpc591 (
      {stage0_46[53]},
      {stage1_46[29]}
   );
   gpc1_1 gpc592 (
      {stage0_47[41]},
      {stage1_47[21]}
   );
   gpc1_1 gpc593 (
      {stage0_47[42]},
      {stage1_47[22]}
   );
   gpc1_1 gpc594 (
      {stage0_47[43]},
      {stage1_47[23]}
   );
   gpc1_1 gpc595 (
      {stage0_47[44]},
      {stage1_47[24]}
   );
   gpc1_1 gpc596 (
      {stage0_47[45]},
      {stage1_47[25]}
   );
   gpc1_1 gpc597 (
      {stage0_47[46]},
      {stage1_47[26]}
   );
   gpc1_1 gpc598 (
      {stage0_47[47]},
      {stage1_47[27]}
   );
   gpc1_1 gpc599 (
      {stage0_47[48]},
      {stage1_47[28]}
   );
   gpc1_1 gpc600 (
      {stage0_47[49]},
      {stage1_47[29]}
   );
   gpc1_1 gpc601 (
      {stage0_47[50]},
      {stage1_47[30]}
   );
   gpc1_1 gpc602 (
      {stage0_47[51]},
      {stage1_47[31]}
   );
   gpc1_1 gpc603 (
      {stage0_47[52]},
      {stage1_47[32]}
   );
   gpc1_1 gpc604 (
      {stage0_47[53]},
      {stage1_47[33]}
   );
   gpc1_1 gpc605 (
      {stage0_49[47]},
      {stage1_49[17]}
   );
   gpc1_1 gpc606 (
      {stage0_49[48]},
      {stage1_49[18]}
   );
   gpc1_1 gpc607 (
      {stage0_49[49]},
      {stage1_49[19]}
   );
   gpc1_1 gpc608 (
      {stage0_49[50]},
      {stage1_49[20]}
   );
   gpc1_1 gpc609 (
      {stage0_49[51]},
      {stage1_49[21]}
   );
   gpc1_1 gpc610 (
      {stage0_49[52]},
      {stage1_49[22]}
   );
   gpc1_1 gpc611 (
      {stage0_49[53]},
      {stage1_49[23]}
   );
   gpc1_1 gpc612 (
      {stage0_50[29]},
      {stage1_50[18]}
   );
   gpc1_1 gpc613 (
      {stage0_50[30]},
      {stage1_50[19]}
   );
   gpc1_1 gpc614 (
      {stage0_50[31]},
      {stage1_50[20]}
   );
   gpc1_1 gpc615 (
      {stage0_50[32]},
      {stage1_50[21]}
   );
   gpc1_1 gpc616 (
      {stage0_50[33]},
      {stage1_50[22]}
   );
   gpc1_1 gpc617 (
      {stage0_50[34]},
      {stage1_50[23]}
   );
   gpc1_1 gpc618 (
      {stage0_50[35]},
      {stage1_50[24]}
   );
   gpc1_1 gpc619 (
      {stage0_50[36]},
      {stage1_50[25]}
   );
   gpc1_1 gpc620 (
      {stage0_50[37]},
      {stage1_50[26]}
   );
   gpc1_1 gpc621 (
      {stage0_50[38]},
      {stage1_50[27]}
   );
   gpc1_1 gpc622 (
      {stage0_50[39]},
      {stage1_50[28]}
   );
   gpc1_1 gpc623 (
      {stage0_50[40]},
      {stage1_50[29]}
   );
   gpc1_1 gpc624 (
      {stage0_50[41]},
      {stage1_50[30]}
   );
   gpc1_1 gpc625 (
      {stage0_50[42]},
      {stage1_50[31]}
   );
   gpc1_1 gpc626 (
      {stage0_50[43]},
      {stage1_50[32]}
   );
   gpc1_1 gpc627 (
      {stage0_50[44]},
      {stage1_50[33]}
   );
   gpc1_1 gpc628 (
      {stage0_50[45]},
      {stage1_50[34]}
   );
   gpc1_1 gpc629 (
      {stage0_50[46]},
      {stage1_50[35]}
   );
   gpc1_1 gpc630 (
      {stage0_50[47]},
      {stage1_50[36]}
   );
   gpc1_1 gpc631 (
      {stage0_50[48]},
      {stage1_50[37]}
   );
   gpc1_1 gpc632 (
      {stage0_50[49]},
      {stage1_50[38]}
   );
   gpc1_1 gpc633 (
      {stage0_50[50]},
      {stage1_50[39]}
   );
   gpc1_1 gpc634 (
      {stage0_50[51]},
      {stage1_50[40]}
   );
   gpc1_1 gpc635 (
      {stage0_50[52]},
      {stage1_50[41]}
   );
   gpc1_1 gpc636 (
      {stage0_50[53]},
      {stage1_50[42]}
   );
   gpc1_1 gpc637 (
      {stage0_51[20]},
      {stage1_51[14]}
   );
   gpc1_1 gpc638 (
      {stage0_51[21]},
      {stage1_51[15]}
   );
   gpc1_1 gpc639 (
      {stage0_51[22]},
      {stage1_51[16]}
   );
   gpc1_1 gpc640 (
      {stage0_51[23]},
      {stage1_51[17]}
   );
   gpc1_1 gpc641 (
      {stage0_51[24]},
      {stage1_51[18]}
   );
   gpc1_1 gpc642 (
      {stage0_51[25]},
      {stage1_51[19]}
   );
   gpc1_1 gpc643 (
      {stage0_51[26]},
      {stage1_51[20]}
   );
   gpc1_1 gpc644 (
      {stage0_51[27]},
      {stage1_51[21]}
   );
   gpc1_1 gpc645 (
      {stage0_51[28]},
      {stage1_51[22]}
   );
   gpc1_1 gpc646 (
      {stage0_51[29]},
      {stage1_51[23]}
   );
   gpc1_1 gpc647 (
      {stage0_51[30]},
      {stage1_51[24]}
   );
   gpc1_1 gpc648 (
      {stage0_51[31]},
      {stage1_51[25]}
   );
   gpc1_1 gpc649 (
      {stage0_51[32]},
      {stage1_51[26]}
   );
   gpc1_1 gpc650 (
      {stage0_51[33]},
      {stage1_51[27]}
   );
   gpc1_1 gpc651 (
      {stage0_51[34]},
      {stage1_51[28]}
   );
   gpc1_1 gpc652 (
      {stage0_51[35]},
      {stage1_51[29]}
   );
   gpc1_1 gpc653 (
      {stage0_51[36]},
      {stage1_51[30]}
   );
   gpc1_1 gpc654 (
      {stage0_51[37]},
      {stage1_51[31]}
   );
   gpc1_1 gpc655 (
      {stage0_51[38]},
      {stage1_51[32]}
   );
   gpc1_1 gpc656 (
      {stage0_51[39]},
      {stage1_51[33]}
   );
   gpc1_1 gpc657 (
      {stage0_51[40]},
      {stage1_51[34]}
   );
   gpc1_1 gpc658 (
      {stage0_51[41]},
      {stage1_51[35]}
   );
   gpc1_1 gpc659 (
      {stage0_51[42]},
      {stage1_51[36]}
   );
   gpc1_1 gpc660 (
      {stage0_51[43]},
      {stage1_51[37]}
   );
   gpc1_1 gpc661 (
      {stage0_51[44]},
      {stage1_51[38]}
   );
   gpc1_1 gpc662 (
      {stage0_51[45]},
      {stage1_51[39]}
   );
   gpc1_1 gpc663 (
      {stage0_51[46]},
      {stage1_51[40]}
   );
   gpc1_1 gpc664 (
      {stage0_51[47]},
      {stage1_51[41]}
   );
   gpc1_1 gpc665 (
      {stage0_51[48]},
      {stage1_51[42]}
   );
   gpc1_1 gpc666 (
      {stage0_51[49]},
      {stage1_51[43]}
   );
   gpc1_1 gpc667 (
      {stage0_51[50]},
      {stage1_51[44]}
   );
   gpc1_1 gpc668 (
      {stage0_51[51]},
      {stage1_51[45]}
   );
   gpc1_1 gpc669 (
      {stage0_51[52]},
      {stage1_51[46]}
   );
   gpc1_1 gpc670 (
      {stage0_51[53]},
      {stage1_51[47]}
   );
   gpc1_1 gpc671 (
      {stage0_52[47]},
      {stage1_52[15]}
   );
   gpc1_1 gpc672 (
      {stage0_52[48]},
      {stage1_52[16]}
   );
   gpc1_1 gpc673 (
      {stage0_52[49]},
      {stage1_52[17]}
   );
   gpc1_1 gpc674 (
      {stage0_52[50]},
      {stage1_52[18]}
   );
   gpc1_1 gpc675 (
      {stage0_52[51]},
      {stage1_52[19]}
   );
   gpc1_1 gpc676 (
      {stage0_52[52]},
      {stage1_52[20]}
   );
   gpc1_1 gpc677 (
      {stage0_52[53]},
      {stage1_52[21]}
   );
   gpc1_1 gpc678 (
      {stage0_53[28]},
      {stage1_53[15]}
   );
   gpc1_1 gpc679 (
      {stage0_53[29]},
      {stage1_53[16]}
   );
   gpc1_1 gpc680 (
      {stage0_53[30]},
      {stage1_53[17]}
   );
   gpc1_1 gpc681 (
      {stage0_53[31]},
      {stage1_53[18]}
   );
   gpc1_1 gpc682 (
      {stage0_53[32]},
      {stage1_53[19]}
   );
   gpc1_1 gpc683 (
      {stage0_53[33]},
      {stage1_53[20]}
   );
   gpc1_1 gpc684 (
      {stage0_53[34]},
      {stage1_53[21]}
   );
   gpc1_1 gpc685 (
      {stage0_53[35]},
      {stage1_53[22]}
   );
   gpc1_1 gpc686 (
      {stage0_53[36]},
      {stage1_53[23]}
   );
   gpc1_1 gpc687 (
      {stage0_53[37]},
      {stage1_53[24]}
   );
   gpc1_1 gpc688 (
      {stage0_53[38]},
      {stage1_53[25]}
   );
   gpc1_1 gpc689 (
      {stage0_53[39]},
      {stage1_53[26]}
   );
   gpc1_1 gpc690 (
      {stage0_53[40]},
      {stage1_53[27]}
   );
   gpc1_1 gpc691 (
      {stage0_53[41]},
      {stage1_53[28]}
   );
   gpc1_1 gpc692 (
      {stage0_53[42]},
      {stage1_53[29]}
   );
   gpc1_1 gpc693 (
      {stage0_53[43]},
      {stage1_53[30]}
   );
   gpc1_1 gpc694 (
      {stage0_53[44]},
      {stage1_53[31]}
   );
   gpc1_1 gpc695 (
      {stage0_53[45]},
      {stage1_53[32]}
   );
   gpc1_1 gpc696 (
      {stage0_53[46]},
      {stage1_53[33]}
   );
   gpc1_1 gpc697 (
      {stage0_53[47]},
      {stage1_53[34]}
   );
   gpc1_1 gpc698 (
      {stage0_53[48]},
      {stage1_53[35]}
   );
   gpc1_1 gpc699 (
      {stage0_53[49]},
      {stage1_53[36]}
   );
   gpc1_1 gpc700 (
      {stage0_53[50]},
      {stage1_53[37]}
   );
   gpc1_1 gpc701 (
      {stage0_53[51]},
      {stage1_53[38]}
   );
   gpc1_1 gpc702 (
      {stage0_53[52]},
      {stage1_53[39]}
   );
   gpc1_1 gpc703 (
      {stage0_53[53]},
      {stage1_53[40]}
   );
   gpc1_1 gpc704 (
      {stage0_54[51]},
      {stage1_54[14]}
   );
   gpc1_1 gpc705 (
      {stage0_54[52]},
      {stage1_54[15]}
   );
   gpc1_1 gpc706 (
      {stage0_54[53]},
      {stage1_54[16]}
   );
   gpc1_1 gpc707 (
      {stage0_55[30]},
      {stage1_55[14]}
   );
   gpc1_1 gpc708 (
      {stage0_55[31]},
      {stage1_55[15]}
   );
   gpc1_1 gpc709 (
      {stage0_55[32]},
      {stage1_55[16]}
   );
   gpc1_1 gpc710 (
      {stage0_55[33]},
      {stage1_55[17]}
   );
   gpc1_1 gpc711 (
      {stage0_55[34]},
      {stage1_55[18]}
   );
   gpc1_1 gpc712 (
      {stage0_55[35]},
      {stage1_55[19]}
   );
   gpc1_1 gpc713 (
      {stage0_55[36]},
      {stage1_55[20]}
   );
   gpc1_1 gpc714 (
      {stage0_55[37]},
      {stage1_55[21]}
   );
   gpc1_1 gpc715 (
      {stage0_55[38]},
      {stage1_55[22]}
   );
   gpc1_1 gpc716 (
      {stage0_55[39]},
      {stage1_55[23]}
   );
   gpc1_1 gpc717 (
      {stage0_55[40]},
      {stage1_55[24]}
   );
   gpc1_1 gpc718 (
      {stage0_55[41]},
      {stage1_55[25]}
   );
   gpc1_1 gpc719 (
      {stage0_55[42]},
      {stage1_55[26]}
   );
   gpc1_1 gpc720 (
      {stage0_55[43]},
      {stage1_55[27]}
   );
   gpc1_1 gpc721 (
      {stage0_55[44]},
      {stage1_55[28]}
   );
   gpc1_1 gpc722 (
      {stage0_55[45]},
      {stage1_55[29]}
   );
   gpc1_1 gpc723 (
      {stage0_55[46]},
      {stage1_55[30]}
   );
   gpc1_1 gpc724 (
      {stage0_55[47]},
      {stage1_55[31]}
   );
   gpc1_1 gpc725 (
      {stage0_55[48]},
      {stage1_55[32]}
   );
   gpc1_1 gpc726 (
      {stage0_55[49]},
      {stage1_55[33]}
   );
   gpc1_1 gpc727 (
      {stage0_55[50]},
      {stage1_55[34]}
   );
   gpc1_1 gpc728 (
      {stage0_55[51]},
      {stage1_55[35]}
   );
   gpc1_1 gpc729 (
      {stage0_55[52]},
      {stage1_55[36]}
   );
   gpc1_1 gpc730 (
      {stage0_55[53]},
      {stage1_55[37]}
   );
   gpc1_1 gpc731 (
      {stage0_57[30]},
      {stage1_57[17]}
   );
   gpc1_1 gpc732 (
      {stage0_57[31]},
      {stage1_57[18]}
   );
   gpc1_1 gpc733 (
      {stage0_57[32]},
      {stage1_57[19]}
   );
   gpc1_1 gpc734 (
      {stage0_57[33]},
      {stage1_57[20]}
   );
   gpc1_1 gpc735 (
      {stage0_57[34]},
      {stage1_57[21]}
   );
   gpc1_1 gpc736 (
      {stage0_57[35]},
      {stage1_57[22]}
   );
   gpc1_1 gpc737 (
      {stage0_57[36]},
      {stage1_57[23]}
   );
   gpc1_1 gpc738 (
      {stage0_57[37]},
      {stage1_57[24]}
   );
   gpc1_1 gpc739 (
      {stage0_57[38]},
      {stage1_57[25]}
   );
   gpc1_1 gpc740 (
      {stage0_57[39]},
      {stage1_57[26]}
   );
   gpc1_1 gpc741 (
      {stage0_57[40]},
      {stage1_57[27]}
   );
   gpc1_1 gpc742 (
      {stage0_57[41]},
      {stage1_57[28]}
   );
   gpc1_1 gpc743 (
      {stage0_57[42]},
      {stage1_57[29]}
   );
   gpc1_1 gpc744 (
      {stage0_57[43]},
      {stage1_57[30]}
   );
   gpc1_1 gpc745 (
      {stage0_57[44]},
      {stage1_57[31]}
   );
   gpc1_1 gpc746 (
      {stage0_57[45]},
      {stage1_57[32]}
   );
   gpc1_1 gpc747 (
      {stage0_57[46]},
      {stage1_57[33]}
   );
   gpc1_1 gpc748 (
      {stage0_57[47]},
      {stage1_57[34]}
   );
   gpc1_1 gpc749 (
      {stage0_57[48]},
      {stage1_57[35]}
   );
   gpc1_1 gpc750 (
      {stage0_57[49]},
      {stage1_57[36]}
   );
   gpc1_1 gpc751 (
      {stage0_57[50]},
      {stage1_57[37]}
   );
   gpc1_1 gpc752 (
      {stage0_57[51]},
      {stage1_57[38]}
   );
   gpc1_1 gpc753 (
      {stage0_57[52]},
      {stage1_57[39]}
   );
   gpc1_1 gpc754 (
      {stage0_57[53]},
      {stage1_57[40]}
   );
   gpc1_1 gpc755 (
      {stage0_59[36]},
      {stage1_59[17]}
   );
   gpc1_1 gpc756 (
      {stage0_59[37]},
      {stage1_59[18]}
   );
   gpc1_1 gpc757 (
      {stage0_59[38]},
      {stage1_59[19]}
   );
   gpc1_1 gpc758 (
      {stage0_59[39]},
      {stage1_59[20]}
   );
   gpc1_1 gpc759 (
      {stage0_59[40]},
      {stage1_59[21]}
   );
   gpc1_1 gpc760 (
      {stage0_59[41]},
      {stage1_59[22]}
   );
   gpc1_1 gpc761 (
      {stage0_59[42]},
      {stage1_59[23]}
   );
   gpc1_1 gpc762 (
      {stage0_59[43]},
      {stage1_59[24]}
   );
   gpc1_1 gpc763 (
      {stage0_59[44]},
      {stage1_59[25]}
   );
   gpc1_1 gpc764 (
      {stage0_59[45]},
      {stage1_59[26]}
   );
   gpc1_1 gpc765 (
      {stage0_59[46]},
      {stage1_59[27]}
   );
   gpc1_1 gpc766 (
      {stage0_59[47]},
      {stage1_59[28]}
   );
   gpc1_1 gpc767 (
      {stage0_59[48]},
      {stage1_59[29]}
   );
   gpc1_1 gpc768 (
      {stage0_59[49]},
      {stage1_59[30]}
   );
   gpc1_1 gpc769 (
      {stage0_59[50]},
      {stage1_59[31]}
   );
   gpc1_1 gpc770 (
      {stage0_59[51]},
      {stage1_59[32]}
   );
   gpc1_1 gpc771 (
      {stage0_59[52]},
      {stage1_59[33]}
   );
   gpc1_1 gpc772 (
      {stage0_59[53]},
      {stage1_59[34]}
   );
   gpc1_1 gpc773 (
      {stage0_62[48]},
      {stage1_62[18]}
   );
   gpc1_1 gpc774 (
      {stage0_62[49]},
      {stage1_62[19]}
   );
   gpc1_1 gpc775 (
      {stage0_62[50]},
      {stage1_62[20]}
   );
   gpc1_1 gpc776 (
      {stage0_62[51]},
      {stage1_62[21]}
   );
   gpc1_1 gpc777 (
      {stage0_62[52]},
      {stage1_62[22]}
   );
   gpc1_1 gpc778 (
      {stage0_62[53]},
      {stage1_62[23]}
   );
   gpc1_1 gpc779 (
      {stage0_63[36]},
      {stage1_63[17]}
   );
   gpc1_1 gpc780 (
      {stage0_63[37]},
      {stage1_63[18]}
   );
   gpc1_1 gpc781 (
      {stage0_63[38]},
      {stage1_63[19]}
   );
   gpc1_1 gpc782 (
      {stage0_63[39]},
      {stage1_63[20]}
   );
   gpc1_1 gpc783 (
      {stage0_63[40]},
      {stage1_63[21]}
   );
   gpc1_1 gpc784 (
      {stage0_63[41]},
      {stage1_63[22]}
   );
   gpc1_1 gpc785 (
      {stage0_63[42]},
      {stage1_63[23]}
   );
   gpc1_1 gpc786 (
      {stage0_63[43]},
      {stage1_63[24]}
   );
   gpc1_1 gpc787 (
      {stage0_63[44]},
      {stage1_63[25]}
   );
   gpc1_1 gpc788 (
      {stage0_63[45]},
      {stage1_63[26]}
   );
   gpc1_1 gpc789 (
      {stage0_63[46]},
      {stage1_63[27]}
   );
   gpc1_1 gpc790 (
      {stage0_63[47]},
      {stage1_63[28]}
   );
   gpc1_1 gpc791 (
      {stage0_63[48]},
      {stage1_63[29]}
   );
   gpc1_1 gpc792 (
      {stage0_63[49]},
      {stage1_63[30]}
   );
   gpc1_1 gpc793 (
      {stage0_63[50]},
      {stage1_63[31]}
   );
   gpc1_1 gpc794 (
      {stage0_63[51]},
      {stage1_63[32]}
   );
   gpc1_1 gpc795 (
      {stage0_63[52]},
      {stage1_63[33]}
   );
   gpc1_1 gpc796 (
      {stage0_63[53]},
      {stage1_63[34]}
   );
   gpc1163_5 gpc797 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc798 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc799 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13]},
      {stage1_1[6]},
      {stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc800 (
      {stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage1_3[1]},
      {stage1_4[0], stage1_4[1]},
      {stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc801 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4]}
   );
   gpc615_5 gpc802 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[2]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[2],stage2_4[5],stage2_3[5]}
   );
   gpc615_5 gpc803 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[3]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc804 (
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22]},
      {stage1_4[4]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[2],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc2135_5 gpc805 (
      {stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9]},
      {stage1_5[18], stage1_5[19], stage1_5[20]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[0],stage2_7[3],stage2_6[3],stage2_5[5],stage2_4[8]}
   );
   gpc2135_5 gpc806 (
      {stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_6[1]},
      {stage1_7[2], stage1_7[3]},
      {stage2_8[1],stage2_7[4],stage2_6[4],stage2_5[6],stage2_4[9]}
   );
   gpc606_5 gpc807 (
      {stage1_4[15], stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[2],stage2_7[5],stage2_6[5],stage2_5[7],stage2_4[10]}
   );
   gpc606_5 gpc808 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9]},
      {stage2_9[0],stage2_8[3],stage2_7[6],stage2_6[6],stage2_5[8]}
   );
   gpc606_5 gpc809 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15]},
      {stage2_9[1],stage2_8[4],stage2_7[7],stage2_6[7],stage2_5[9]}
   );
   gpc615_5 gpc810 (
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage1_7[16]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[5],stage2_7[8],stage2_6[8]}
   );
   gpc615_5 gpc811 (
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_7[17]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[6],stage2_7[9],stage2_6[9]}
   );
   gpc615_5 gpc812 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[12]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[4],stage2_8[7],stage2_7[10]}
   );
   gpc606_5 gpc813 (
      {stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[3],stage2_9[5],stage2_8[8]}
   );
   gpc606_5 gpc814 (
      {stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[2],stage2_10[4],stage2_9[6],stage2_8[9]}
   );
   gpc606_5 gpc815 (
      {stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[3],stage2_10[5],stage2_9[7],stage2_8[10]}
   );
   gpc615_5 gpc816 (
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22]},
      {stage1_11[0]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[3],stage2_11[4],stage2_10[6]}
   );
   gpc1415_5 gpc817 (
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[1],stage2_12[4],stage2_11[5]}
   );
   gpc1415_5 gpc818 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10]},
      {stage1_12[7]},
      {stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7]},
      {stage1_14[1]},
      {stage2_15[1],stage2_14[2],stage2_13[2],stage2_12[5],stage2_11[6]}
   );
   gpc1163_5 gpc819 (
      {stage1_11[11], stage1_11[12], stage1_11[13]},
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage1_13[8]},
      {stage1_14[2]},
      {stage2_15[2],stage2_14[3],stage2_13[3],stage2_12[6],stage2_11[7]}
   );
   gpc1163_5 gpc820 (
      {stage1_11[14], stage1_11[15], stage1_11[16]},
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage1_13[9]},
      {stage1_14[3]},
      {stage2_15[3],stage2_14[4],stage2_13[4],stage2_12[7],stage2_11[8]}
   );
   gpc615_5 gpc821 (
      {stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_12[20]},
      {stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15]},
      {stage2_15[4],stage2_14[5],stage2_13[5],stage2_12[8],stage2_11[9]}
   );
   gpc615_5 gpc822 (
      {stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25], stage1_11[26]},
      {1'b0},
      {stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21]},
      {stage2_15[5],stage2_14[6],stage2_13[6],stage2_12[9],stage2_11[10]}
   );
   gpc606_5 gpc823 (
      {stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[6],stage2_14[7],stage2_13[7]}
   );
   gpc1343_5 gpc824 (
      {stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9]},
      {stage1_16[0], stage1_16[1], stage1_16[2]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[1],stage2_16[1],stage2_15[7],stage2_14[8]}
   );
   gpc1343_5 gpc825 (
      {stage1_14[7], stage1_14[8], stage1_14[9]},
      {stage1_15[10], stage1_15[11], stage1_15[12], stage1_15[13]},
      {stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage1_17[1]},
      {stage2_18[1],stage2_17[2],stage2_16[2],stage2_15[8],stage2_14[9]}
   );
   gpc1163_5 gpc826 (
      {stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19]},
      {stage1_16[6]},
      {stage1_17[2]},
      {stage2_18[2],stage2_17[3],stage2_16[3],stage2_15[9],stage2_14[10]}
   );
   gpc1163_5 gpc827 (
      {stage1_14[13], stage1_14[14], stage1_14[15]},
      {stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25]},
      {stage1_16[7]},
      {stage1_17[3]},
      {stage2_18[3],stage2_17[4],stage2_16[4],stage2_15[10],stage2_14[11]}
   );
   gpc1163_5 gpc828 (
      {stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31]},
      {stage1_16[8]},
      {stage1_17[4]},
      {stage2_18[4],stage2_17[5],stage2_16[5],stage2_15[11],stage2_14[12]}
   );
   gpc1163_5 gpc829 (
      {stage1_14[19], stage1_14[20], stage1_14[21]},
      {stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage1_16[9]},
      {stage1_17[5]},
      {stage2_18[5],stage2_17[6],stage2_16[6],stage2_15[12],stage2_14[13]}
   );
   gpc1163_5 gpc830 (
      {stage1_14[22], stage1_14[23], 1'b0},
      {stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], 1'b0},
      {stage1_16[10]},
      {stage1_17[6]},
      {stage2_18[6],stage2_17[7],stage2_16[7],stage2_15[13],stage2_14[14]}
   );
   gpc606_5 gpc831 (
      {stage1_16[11], stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[7],stage2_17[8],stage2_16[8]}
   );
   gpc606_5 gpc832 (
      {stage1_16[17], stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[1],stage2_18[8],stage2_17[9],stage2_16[9]}
   );
   gpc606_5 gpc833 (
      {stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[9],stage2_17[10]}
   );
   gpc615_5 gpc834 (
      {stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage1_18[12]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[10],stage2_17[11]}
   );
   gpc615_5 gpc835 (
      {stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage1_19[12]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[11]}
   );
   gpc615_5 gpc836 (
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22]},
      {stage1_19[13]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[3],stage2_20[5],stage2_19[5],stage2_18[12]}
   );
   gpc615_5 gpc837 (
      {stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27]},
      {stage1_19[14]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[4],stage2_20[6],stage2_19[6],stage2_18[13]}
   );
   gpc615_5 gpc838 (
      {stage1_19[15], stage1_19[16], stage1_19[17], stage1_19[18], stage1_19[19]},
      {stage1_20[18]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[5],stage2_20[7],stage2_19[7]}
   );
   gpc1343_5 gpc839 (
      {stage1_21[6], stage1_21[7], stage1_21[8]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3]},
      {stage1_23[0], stage1_23[1], stage1_23[2]},
      {stage1_24[0]},
      {stage2_25[0],stage2_24[0],stage2_23[1],stage2_22[4],stage2_21[6]}
   );
   gpc1343_5 gpc840 (
      {stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage1_22[4], stage1_22[5], stage1_22[6], stage1_22[7]},
      {stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage1_24[1]},
      {stage2_25[1],stage2_24[1],stage2_23[2],stage2_22[5],stage2_21[7]}
   );
   gpc606_5 gpc841 (
      {stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11], stage1_22[12], stage1_22[13]},
      {stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6], stage1_24[7]},
      {stage2_26[0],stage2_25[2],stage2_24[2],stage2_23[3],stage2_22[6]}
   );
   gpc606_5 gpc842 (
      {stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17], stage1_22[18], stage1_22[19]},
      {stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13]},
      {stage2_26[1],stage2_25[3],stage2_24[3],stage2_23[4],stage2_22[7]}
   );
   gpc615_5 gpc843 (
      {stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18]},
      {stage1_25[0]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[0],stage2_26[2],stage2_25[4],stage2_24[4]}
   );
   gpc615_5 gpc844 (
      {stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage1_25[1]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[1],stage2_26[3],stage2_25[5],stage2_24[5]}
   );
   gpc615_5 gpc845 (
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28]},
      {stage1_25[2]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[2],stage2_26[4],stage2_25[6],stage2_24[6]}
   );
   gpc615_5 gpc846 (
      {stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6], stage1_25[7]},
      {stage1_26[18]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[3],stage2_27[3],stage2_26[5],stage2_25[7]}
   );
   gpc615_5 gpc847 (
      {stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12]},
      {stage1_26[19]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[4],stage2_27[4],stage2_26[6],stage2_25[8]}
   );
   gpc615_5 gpc848 (
      {stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage1_26[20]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[5],stage2_27[5],stage2_26[7],stage2_25[9]}
   );
   gpc615_5 gpc849 (
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22]},
      {stage1_26[21]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[6],stage2_27[6],stage2_26[8],stage2_25[10]}
   );
   gpc1343_5 gpc850 (
      {stage1_28[0], stage1_28[1], stage1_28[2]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3]},
      {stage1_30[0], stage1_30[1], stage1_30[2]},
      {stage1_31[0]},
      {stage2_32[0],stage2_31[0],stage2_30[0],stage2_29[4],stage2_28[7]}
   );
   gpc1343_5 gpc851 (
      {stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage1_29[4], stage1_29[5], stage1_29[6], stage1_29[7]},
      {stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage1_31[1]},
      {stage2_32[1],stage2_31[1],stage2_30[1],stage2_29[5],stage2_28[8]}
   );
   gpc1343_5 gpc852 (
      {stage1_28[6], stage1_28[7], stage1_28[8]},
      {stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage1_30[6], stage1_30[7], stage1_30[8]},
      {stage1_31[2]},
      {stage2_32[2],stage2_31[2],stage2_30[2],stage2_29[6],stage2_28[9]}
   );
   gpc606_5 gpc853 (
      {stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12], stage1_28[13], stage1_28[14]},
      {stage1_30[9], stage1_30[10], stage1_30[11], stage1_30[12], stage1_30[13], stage1_30[14]},
      {stage2_32[3],stage2_31[3],stage2_30[3],stage2_29[7],stage2_28[10]}
   );
   gpc615_5 gpc854 (
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16]},
      {stage1_30[15]},
      {stage1_31[3], stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8]},
      {stage2_33[0],stage2_32[4],stage2_31[4],stage2_30[4],stage2_29[8]}
   );
   gpc606_5 gpc855 (
      {stage1_30[16], stage1_30[17], stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[1],stage2_32[5],stage2_31[5],stage2_30[5]}
   );
   gpc606_5 gpc856 (
      {stage1_30[22], stage1_30[23], stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[2],stage2_32[6],stage2_31[6],stage2_30[6]}
   );
   gpc615_5 gpc857 (
      {stage1_30[28], stage1_30[29], stage1_30[30], stage1_30[31], stage1_30[32]},
      {stage1_31[9]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[3],stage2_32[7],stage2_31[7],stage2_30[7]}
   );
   gpc606_5 gpc858 (
      {stage1_31[10], stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[3],stage2_33[4],stage2_32[8],stage2_31[8]}
   );
   gpc606_5 gpc859 (
      {stage1_31[16], stage1_31[17], stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[4],stage2_33[5],stage2_32[9],stage2_31[9]}
   );
   gpc606_5 gpc860 (
      {stage1_31[22], stage1_31[23], stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[5],stage2_33[6],stage2_32[10],stage2_31[10]}
   );
   gpc606_5 gpc861 (
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[0],stage2_35[3],stage2_34[6],stage2_33[7]}
   );
   gpc606_5 gpc862 (
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[1],stage2_35[4],stage2_34[7],stage2_33[8]}
   );
   gpc606_5 gpc863 (
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[2],stage2_35[5],stage2_34[8],stage2_33[9]}
   );
   gpc615_5 gpc864 (
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40]},
      {stage1_34[0]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[3],stage2_35[6],stage2_34[9],stage2_33[10]}
   );
   gpc615_5 gpc865 (
      {stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage1_35[24]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[4],stage2_36[4],stage2_35[7],stage2_34[10]}
   );
   gpc615_5 gpc866 (
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10]},
      {stage1_35[25]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[5],stage2_36[5],stage2_35[8],stage2_34[11]}
   );
   gpc615_5 gpc867 (
      {stage1_34[11], stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15]},
      {stage1_35[26]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[6],stage2_36[6],stage2_35[9],stage2_34[12]}
   );
   gpc615_5 gpc868 (
      {stage1_36[18], stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22]},
      {stage1_37[0]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[0],stage2_38[3],stage2_37[7],stage2_36[7]}
   );
   gpc606_5 gpc869 (
      {stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5], stage1_37[6]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[1],stage2_39[1],stage2_38[4],stage2_37[8]}
   );
   gpc606_5 gpc870 (
      {stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11], stage1_37[12]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[2],stage2_39[2],stage2_38[5],stage2_37[9]}
   );
   gpc606_5 gpc871 (
      {stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17], stage1_37[18]},
      {stage1_39[12], stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17]},
      {stage2_41[2],stage2_40[3],stage2_39[3],stage2_38[6],stage2_37[10]}
   );
   gpc615_5 gpc872 (
      {stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10]},
      {stage1_39[18]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[3],stage2_40[4],stage2_39[4],stage2_38[7]}
   );
   gpc615_5 gpc873 (
      {stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15]},
      {stage1_39[19]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[4],stage2_40[5],stage2_39[5],stage2_38[8]}
   );
   gpc615_5 gpc874 (
      {stage1_38[16], stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20]},
      {stage1_39[20]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[5],stage2_40[6],stage2_39[6],stage2_38[9]}
   );
   gpc1163_5 gpc875 (
      {stage1_40[18], stage1_40[19], stage1_40[20]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage1_42[0]},
      {stage1_43[0]},
      {stage2_44[0],stage2_43[0],stage2_42[3],stage2_41[6],stage2_40[7]}
   );
   gpc1163_5 gpc876 (
      {stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage1_42[1]},
      {stage1_43[1]},
      {stage2_44[1],stage2_43[1],stage2_42[4],stage2_41[7],stage2_40[8]}
   );
   gpc1163_5 gpc877 (
      {stage1_40[24], stage1_40[25], stage1_40[26]},
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage1_42[2]},
      {stage1_43[2]},
      {stage2_44[2],stage2_43[2],stage2_42[5],stage2_41[8],stage2_40[9]}
   );
   gpc606_5 gpc878 (
      {stage1_40[27], stage1_40[28], stage1_40[29], stage1_40[30], stage1_40[31], stage1_40[32]},
      {stage1_42[3], stage1_42[4], stage1_42[5], stage1_42[6], stage1_42[7], stage1_42[8]},
      {stage2_44[3],stage2_43[3],stage2_42[6],stage2_41[9],stage2_40[10]}
   );
   gpc606_5 gpc879 (
      {stage1_40[33], stage1_40[34], stage1_40[35], stage1_40[36], stage1_40[37], stage1_40[38]},
      {stage1_42[9], stage1_42[10], stage1_42[11], stage1_42[12], stage1_42[13], stage1_42[14]},
      {stage2_44[4],stage2_43[4],stage2_42[7],stage2_41[10],stage2_40[11]}
   );
   gpc606_5 gpc880 (
      {stage1_43[3], stage1_43[4], stage1_43[5], stage1_43[6], stage1_43[7], stage1_43[8]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[0],stage2_44[5],stage2_43[5]}
   );
   gpc606_5 gpc881 (
      {stage1_43[9], stage1_43[10], stage1_43[11], stage1_43[12], stage1_43[13], stage1_43[14]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[1],stage2_44[6],stage2_43[6]}
   );
   gpc606_5 gpc882 (
      {stage1_43[15], stage1_43[16], stage1_43[17], stage1_43[18], stage1_43[19], stage1_43[20]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[2],stage2_45[2],stage2_44[7],stage2_43[7]}
   );
   gpc606_5 gpc883 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[3],stage2_46[3],stage2_45[3],stage2_44[8]}
   );
   gpc606_5 gpc884 (
      {stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9], stage1_44[10], stage1_44[11]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[4],stage2_46[4],stage2_45[4],stage2_44[9]}
   );
   gpc606_5 gpc885 (
      {stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16], stage1_44[17]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage2_48[2],stage2_47[5],stage2_46[5],stage2_45[5],stage2_44[10]}
   );
   gpc615_5 gpc886 (
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22]},
      {stage1_46[18]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[3],stage2_47[6],stage2_46[6],stage2_45[6]}
   );
   gpc615_5 gpc887 (
      {stage1_45[23], stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27]},
      {stage1_46[19]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[4],stage2_47[7],stage2_46[7],stage2_45[7]}
   );
   gpc615_5 gpc888 (
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16]},
      {stage1_48[0]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[0],stage2_49[2],stage2_48[5],stage2_47[8]}
   );
   gpc615_5 gpc889 (
      {stage1_47[17], stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21]},
      {stage1_48[1]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[1],stage2_49[3],stage2_48[6],stage2_47[9]}
   );
   gpc606_5 gpc890 (
      {stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5], stage1_48[6], stage1_48[7]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[2],stage2_50[2],stage2_49[4],stage2_48[7]}
   );
   gpc606_5 gpc891 (
      {stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11], stage1_48[12], stage1_48[13]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[3],stage2_50[3],stage2_49[5],stage2_48[8]}
   );
   gpc2135_5 gpc892 (
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16]},
      {stage1_51[0], stage1_51[1], stage1_51[2]},
      {stage1_52[0]},
      {stage1_53[0], stage1_53[1]},
      {stage2_54[0],stage2_53[0],stage2_52[2],stage2_51[4],stage2_50[4]}
   );
   gpc2135_5 gpc893 (
      {stage1_50[17], stage1_50[18], stage1_50[19], stage1_50[20], stage1_50[21]},
      {stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage1_52[1]},
      {stage1_53[2], stage1_53[3]},
      {stage2_54[1],stage2_53[1],stage2_52[3],stage2_51[5],stage2_50[5]}
   );
   gpc2135_5 gpc894 (
      {stage1_50[22], stage1_50[23], stage1_50[24], stage1_50[25], stage1_50[26]},
      {stage1_51[6], stage1_51[7], stage1_51[8]},
      {stage1_52[2]},
      {stage1_53[4], stage1_53[5]},
      {stage2_54[2],stage2_53[2],stage2_52[4],stage2_51[6],stage2_50[6]}
   );
   gpc2135_5 gpc895 (
      {stage1_50[27], stage1_50[28], stage1_50[29], stage1_50[30], stage1_50[31]},
      {stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage1_52[3]},
      {stage1_53[6], stage1_53[7]},
      {stage2_54[3],stage2_53[3],stage2_52[5],stage2_51[7],stage2_50[7]}
   );
   gpc2135_5 gpc896 (
      {stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35], stage1_50[36]},
      {stage1_51[12], stage1_51[13], stage1_51[14]},
      {stage1_52[4]},
      {stage1_53[8], stage1_53[9]},
      {stage2_54[4],stage2_53[4],stage2_52[6],stage2_51[8],stage2_50[8]}
   );
   gpc615_5 gpc897 (
      {stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage1_51[15]},
      {stage1_52[5], stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10]},
      {stage2_54[5],stage2_53[5],stage2_52[7],stage2_51[9],stage2_50[9]}
   );
   gpc606_5 gpc898 (
      {stage1_51[16], stage1_51[17], stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21]},
      {stage1_53[10], stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15]},
      {stage2_55[0],stage2_54[6],stage2_53[6],stage2_52[8],stage2_51[10]}
   );
   gpc606_5 gpc899 (
      {stage1_51[22], stage1_51[23], stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27]},
      {stage1_53[16], stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21]},
      {stage2_55[1],stage2_54[7],stage2_53[7],stage2_52[9],stage2_51[11]}
   );
   gpc606_5 gpc900 (
      {stage1_51[28], stage1_51[29], stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33]},
      {stage1_53[22], stage1_53[23], stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27]},
      {stage2_55[2],stage2_54[8],stage2_53[8],stage2_52[10],stage2_51[12]}
   );
   gpc606_5 gpc901 (
      {stage1_51[34], stage1_51[35], stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39]},
      {stage1_53[28], stage1_53[29], stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33]},
      {stage2_55[3],stage2_54[9],stage2_53[9],stage2_52[11],stage2_51[13]}
   );
   gpc606_5 gpc902 (
      {stage1_51[40], stage1_51[41], stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45]},
      {stage1_53[34], stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39]},
      {stage2_55[4],stage2_54[10],stage2_53[10],stage2_52[12],stage2_51[14]}
   );
   gpc606_5 gpc903 (
      {stage1_52[11], stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[5],stage2_54[11],stage2_53[11],stage2_52[13]}
   );
   gpc615_5 gpc904 (
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10]},
      {stage1_55[0]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[0],stage2_56[1],stage2_55[6],stage2_54[12]}
   );
   gpc615_5 gpc905 (
      {stage1_54[11], stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15]},
      {stage1_55[1]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[1],stage2_56[2],stage2_55[7],stage2_54[13]}
   );
   gpc606_5 gpc906 (
      {stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5], stage1_55[6], stage1_55[7]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[2],stage2_57[2],stage2_56[3],stage2_55[8]}
   );
   gpc606_5 gpc907 (
      {stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11], stage1_55[12], stage1_55[13]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[3],stage2_57[3],stage2_56[4],stage2_55[9]}
   );
   gpc606_5 gpc908 (
      {stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17], stage1_55[18], stage1_55[19]},
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage2_59[2],stage2_58[4],stage2_57[4],stage2_56[5],stage2_55[10]}
   );
   gpc606_5 gpc909 (
      {stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23], stage1_55[24], stage1_55[25]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[3],stage2_58[5],stage2_57[5],stage2_56[6],stage2_55[11]}
   );
   gpc606_5 gpc910 (
      {stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29], stage1_55[30], stage1_55[31]},
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage2_59[4],stage2_58[6],stage2_57[6],stage2_56[7],stage2_55[12]}
   );
   gpc615_5 gpc911 (
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16]},
      {stage1_57[30]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[5],stage2_58[7],stage2_57[7],stage2_56[8]}
   );
   gpc606_5 gpc912 (
      {stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35], stage1_57[36]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[1],stage2_59[6],stage2_58[8],stage2_57[8]}
   );
   gpc135_4 gpc913 (
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10]},
      {stage1_60[0], stage1_60[1], stage1_60[2]},
      {stage1_61[0]},
      {stage2_62[0],stage2_61[1],stage2_60[2],stage2_59[7]}
   );
   gpc135_4 gpc914 (
      {stage1_59[11], stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15]},
      {stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage1_61[1]},
      {stage2_62[1],stage2_61[2],stage2_60[3],stage2_59[8]}
   );
   gpc135_4 gpc915 (
      {stage1_59[16], stage1_59[17], stage1_59[18], stage1_59[19], stage1_59[20]},
      {stage1_60[6], stage1_60[7], stage1_60[8]},
      {stage1_61[2]},
      {stage2_62[2],stage2_61[3],stage2_60[4],stage2_59[9]}
   );
   gpc135_4 gpc916 (
      {stage1_59[21], stage1_59[22], stage1_59[23], stage1_59[24], stage1_59[25]},
      {stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage1_61[3]},
      {stage2_62[3],stage2_61[4],stage2_60[5],stage2_59[10]}
   );
   gpc135_4 gpc917 (
      {stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29], stage1_59[30]},
      {stage1_60[12], stage1_60[13], stage1_60[14]},
      {stage1_61[4]},
      {stage2_62[4],stage2_61[5],stage2_60[6],stage2_59[11]}
   );
   gpc135_4 gpc918 (
      {stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], 1'b0},
      {stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage1_61[5]},
      {stage2_62[5],stage2_61[6],stage2_60[7],stage2_59[12]}
   );
   gpc606_5 gpc919 (
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[0],stage2_63[0],stage2_62[6],stage2_61[7]}
   );
   gpc606_5 gpc920 (
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage2_65[1],stage2_64[1],stage2_63[1],stage2_62[7],stage2_61[8]}
   );
   gpc1163_5 gpc921 (
      {stage1_62[0], stage1_62[1], stage1_62[2]},
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage1_64[0]},
      {stage1_65[0]},
      {stage2_66[0],stage2_65[2],stage2_64[2],stage2_63[2],stage2_62[8]}
   );
   gpc1163_5 gpc922 (
      {stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage1_63[18], stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage1_64[1]},
      {stage1_65[1]},
      {stage2_66[1],stage2_65[3],stage2_64[3],stage2_63[3],stage2_62[9]}
   );
   gpc606_5 gpc923 (
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage1_64[2], stage1_64[3], stage1_64[4], stage1_64[5], stage1_64[6], stage1_64[7]},
      {stage2_66[2],stage2_65[4],stage2_64[4],stage2_63[4],stage2_62[10]}
   );
   gpc606_5 gpc924 (
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage1_64[8], stage1_64[9], stage1_64[10], stage1_64[11], stage1_64[12], stage1_64[13]},
      {stage2_66[3],stage2_65[5],stage2_64[5],stage2_63[5],stage2_62[11]}
   );
   gpc1_1 gpc925 (
      {stage1_0[14]},
      {stage2_0[3]}
   );
   gpc1_1 gpc926 (
      {stage1_0[15]},
      {stage2_0[4]}
   );
   gpc1_1 gpc927 (
      {stage1_0[16]},
      {stage2_0[5]}
   );
   gpc1_1 gpc928 (
      {stage1_1[18]},
      {stage2_1[5]}
   );
   gpc1_1 gpc929 (
      {stage1_1[19]},
      {stage2_1[6]}
   );
   gpc1_1 gpc930 (
      {stage1_2[16]},
      {stage2_2[5]}
   );
   gpc1_1 gpc931 (
      {stage1_2[17]},
      {stage2_2[6]}
   );
   gpc1_1 gpc932 (
      {stage1_2[18]},
      {stage2_2[7]}
   );
   gpc1_1 gpc933 (
      {stage1_2[19]},
      {stage2_2[8]}
   );
   gpc1_1 gpc934 (
      {stage1_2[20]},
      {stage2_2[9]}
   );
   gpc1_1 gpc935 (
      {stage1_2[21]},
      {stage2_2[10]}
   );
   gpc1_1 gpc936 (
      {stage1_2[22]},
      {stage2_2[11]}
   );
   gpc1_1 gpc937 (
      {stage1_2[23]},
      {stage2_2[12]}
   );
   gpc1_1 gpc938 (
      {stage1_2[24]},
      {stage2_2[13]}
   );
   gpc1_1 gpc939 (
      {stage1_3[23]},
      {stage2_3[8]}
   );
   gpc1_1 gpc940 (
      {stage1_4[21]},
      {stage2_4[11]}
   );
   gpc1_1 gpc941 (
      {stage1_4[22]},
      {stage2_4[12]}
   );
   gpc1_1 gpc942 (
      {stage1_4[23]},
      {stage2_4[13]}
   );
   gpc1_1 gpc943 (
      {stage1_4[24]},
      {stage2_4[14]}
   );
   gpc1_1 gpc944 (
      {stage1_4[25]},
      {stage2_4[15]}
   );
   gpc1_1 gpc945 (
      {stage1_4[26]},
      {stage2_4[16]}
   );
   gpc1_1 gpc946 (
      {stage1_4[27]},
      {stage2_4[17]}
   );
   gpc1_1 gpc947 (
      {stage1_4[28]},
      {stage2_4[18]}
   );
   gpc1_1 gpc948 (
      {stage1_4[29]},
      {stage2_4[19]}
   );
   gpc1_1 gpc949 (
      {stage1_4[30]},
      {stage2_4[20]}
   );
   gpc1_1 gpc950 (
      {stage1_4[31]},
      {stage2_4[21]}
   );
   gpc1_1 gpc951 (
      {stage1_4[32]},
      {stage2_4[22]}
   );
   gpc1_1 gpc952 (
      {stage1_6[18]},
      {stage2_6[10]}
   );
   gpc1_1 gpc953 (
      {stage1_7[23]},
      {stage2_7[11]}
   );
   gpc1_1 gpc954 (
      {stage1_7[24]},
      {stage2_7[12]}
   );
   gpc1_1 gpc955 (
      {stage1_9[6]},
      {stage2_9[8]}
   );
   gpc1_1 gpc956 (
      {stage1_9[7]},
      {stage2_9[9]}
   );
   gpc1_1 gpc957 (
      {stage1_9[8]},
      {stage2_9[10]}
   );
   gpc1_1 gpc958 (
      {stage1_9[9]},
      {stage2_9[11]}
   );
   gpc1_1 gpc959 (
      {stage1_9[10]},
      {stage2_9[12]}
   );
   gpc1_1 gpc960 (
      {stage1_9[11]},
      {stage2_9[13]}
   );
   gpc1_1 gpc961 (
      {stage1_9[12]},
      {stage2_9[14]}
   );
   gpc1_1 gpc962 (
      {stage1_9[13]},
      {stage2_9[15]}
   );
   gpc1_1 gpc963 (
      {stage1_9[14]},
      {stage2_9[16]}
   );
   gpc1_1 gpc964 (
      {stage1_9[15]},
      {stage2_9[17]}
   );
   gpc1_1 gpc965 (
      {stage1_9[16]},
      {stage2_9[18]}
   );
   gpc1_1 gpc966 (
      {stage1_9[17]},
      {stage2_9[19]}
   );
   gpc1_1 gpc967 (
      {stage1_10[23]},
      {stage2_10[7]}
   );
   gpc1_1 gpc968 (
      {stage1_10[24]},
      {stage2_10[8]}
   );
   gpc1_1 gpc969 (
      {stage1_10[25]},
      {stage2_10[9]}
   );
   gpc1_1 gpc970 (
      {stage1_11[27]},
      {stage2_11[11]}
   );
   gpc1_1 gpc971 (
      {stage1_11[28]},
      {stage2_11[12]}
   );
   gpc1_1 gpc972 (
      {stage1_13[28]},
      {stage2_13[8]}
   );
   gpc1_1 gpc973 (
      {stage1_13[29]},
      {stage2_13[9]}
   );
   gpc1_1 gpc974 (
      {stage1_16[23]},
      {stage2_16[10]}
   );
   gpc1_1 gpc975 (
      {stage1_18[28]},
      {stage2_18[14]}
   );
   gpc1_1 gpc976 (
      {stage1_18[29]},
      {stage2_18[15]}
   );
   gpc1_1 gpc977 (
      {stage1_18[30]},
      {stage2_18[16]}
   );
   gpc1_1 gpc978 (
      {stage1_18[31]},
      {stage2_18[17]}
   );
   gpc1_1 gpc979 (
      {stage1_18[32]},
      {stage2_18[18]}
   );
   gpc1_1 gpc980 (
      {stage1_18[33]},
      {stage2_18[19]}
   );
   gpc1_1 gpc981 (
      {stage1_19[20]},
      {stage2_19[8]}
   );
   gpc1_1 gpc982 (
      {stage1_20[19]},
      {stage2_20[8]}
   );
   gpc1_1 gpc983 (
      {stage1_21[12]},
      {stage2_21[8]}
   );
   gpc1_1 gpc984 (
      {stage1_21[13]},
      {stage2_21[9]}
   );
   gpc1_1 gpc985 (
      {stage1_21[14]},
      {stage2_21[10]}
   );
   gpc1_1 gpc986 (
      {stage1_21[15]},
      {stage2_21[11]}
   );
   gpc1_1 gpc987 (
      {stage1_21[16]},
      {stage2_21[12]}
   );
   gpc1_1 gpc988 (
      {stage1_21[17]},
      {stage2_21[13]}
   );
   gpc1_1 gpc989 (
      {stage1_21[18]},
      {stage2_21[14]}
   );
   gpc1_1 gpc990 (
      {stage1_21[19]},
      {stage2_21[15]}
   );
   gpc1_1 gpc991 (
      {stage1_21[20]},
      {stage2_21[16]}
   );
   gpc1_1 gpc992 (
      {stage1_21[21]},
      {stage2_21[17]}
   );
   gpc1_1 gpc993 (
      {stage1_21[22]},
      {stage2_21[18]}
   );
   gpc1_1 gpc994 (
      {stage1_21[23]},
      {stage2_21[19]}
   );
   gpc1_1 gpc995 (
      {stage1_21[24]},
      {stage2_21[20]}
   );
   gpc1_1 gpc996 (
      {stage1_21[25]},
      {stage2_21[21]}
   );
   gpc1_1 gpc997 (
      {stage1_22[20]},
      {stage2_22[8]}
   );
   gpc1_1 gpc998 (
      {stage1_22[21]},
      {stage2_22[9]}
   );
   gpc1_1 gpc999 (
      {stage1_22[22]},
      {stage2_22[10]}
   );
   gpc1_1 gpc1000 (
      {stage1_23[6]},
      {stage2_23[5]}
   );
   gpc1_1 gpc1001 (
      {stage1_23[7]},
      {stage2_23[6]}
   );
   gpc1_1 gpc1002 (
      {stage1_23[8]},
      {stage2_23[7]}
   );
   gpc1_1 gpc1003 (
      {stage1_23[9]},
      {stage2_23[8]}
   );
   gpc1_1 gpc1004 (
      {stage1_23[10]},
      {stage2_23[9]}
   );
   gpc1_1 gpc1005 (
      {stage1_23[11]},
      {stage2_23[10]}
   );
   gpc1_1 gpc1006 (
      {stage1_23[12]},
      {stage2_23[11]}
   );
   gpc1_1 gpc1007 (
      {stage1_23[13]},
      {stage2_23[12]}
   );
   gpc1_1 gpc1008 (
      {stage1_23[14]},
      {stage2_23[13]}
   );
   gpc1_1 gpc1009 (
      {stage1_23[15]},
      {stage2_23[14]}
   );
   gpc1_1 gpc1010 (
      {stage1_23[16]},
      {stage2_23[15]}
   );
   gpc1_1 gpc1011 (
      {stage1_23[17]},
      {stage2_23[16]}
   );
   gpc1_1 gpc1012 (
      {stage1_23[18]},
      {stage2_23[17]}
   );
   gpc1_1 gpc1013 (
      {stage1_23[19]},
      {stage2_23[18]}
   );
   gpc1_1 gpc1014 (
      {stage1_23[20]},
      {stage2_23[19]}
   );
   gpc1_1 gpc1015 (
      {stage1_23[21]},
      {stage2_23[20]}
   );
   gpc1_1 gpc1016 (
      {stage1_24[29]},
      {stage2_24[7]}
   );
   gpc1_1 gpc1017 (
      {stage1_24[30]},
      {stage2_24[8]}
   );
   gpc1_1 gpc1018 (
      {stage1_24[31]},
      {stage2_24[9]}
   );
   gpc1_1 gpc1019 (
      {stage1_25[23]},
      {stage2_25[11]}
   );
   gpc1_1 gpc1020 (
      {stage1_25[24]},
      {stage2_25[12]}
   );
   gpc1_1 gpc1021 (
      {stage1_26[22]},
      {stage2_26[9]}
   );
   gpc1_1 gpc1022 (
      {stage1_26[23]},
      {stage2_26[10]}
   );
   gpc1_1 gpc1023 (
      {stage1_26[24]},
      {stage2_26[11]}
   );
   gpc1_1 gpc1024 (
      {stage1_26[25]},
      {stage2_26[12]}
   );
   gpc1_1 gpc1025 (
      {stage1_26[26]},
      {stage2_26[13]}
   );
   gpc1_1 gpc1026 (
      {stage1_26[27]},
      {stage2_26[14]}
   );
   gpc1_1 gpc1027 (
      {stage1_26[28]},
      {stage2_26[15]}
   );
   gpc1_1 gpc1028 (
      {stage1_26[29]},
      {stage2_26[16]}
   );
   gpc1_1 gpc1029 (
      {stage1_26[30]},
      {stage2_26[17]}
   );
   gpc1_1 gpc1030 (
      {stage1_26[31]},
      {stage2_26[18]}
   );
   gpc1_1 gpc1031 (
      {stage1_28[15]},
      {stage2_28[11]}
   );
   gpc1_1 gpc1032 (
      {stage1_28[16]},
      {stage2_28[12]}
   );
   gpc1_1 gpc1033 (
      {stage1_28[17]},
      {stage2_28[13]}
   );
   gpc1_1 gpc1034 (
      {stage1_29[17]},
      {stage2_29[9]}
   );
   gpc1_1 gpc1035 (
      {stage1_29[18]},
      {stage2_29[10]}
   );
   gpc1_1 gpc1036 (
      {stage1_29[19]},
      {stage2_29[11]}
   );
   gpc1_1 gpc1037 (
      {stage1_29[20]},
      {stage2_29[12]}
   );
   gpc1_1 gpc1038 (
      {stage1_29[21]},
      {stage2_29[13]}
   );
   gpc1_1 gpc1039 (
      {stage1_29[22]},
      {stage2_29[14]}
   );
   gpc1_1 gpc1040 (
      {stage1_29[23]},
      {stage2_29[15]}
   );
   gpc1_1 gpc1041 (
      {stage1_29[24]},
      {stage2_29[16]}
   );
   gpc1_1 gpc1042 (
      {stage1_29[25]},
      {stage2_29[17]}
   );
   gpc1_1 gpc1043 (
      {stage1_30[33]},
      {stage2_30[8]}
   );
   gpc1_1 gpc1044 (
      {stage1_30[34]},
      {stage2_30[9]}
   );
   gpc1_1 gpc1045 (
      {stage1_31[28]},
      {stage2_31[11]}
   );
   gpc1_1 gpc1046 (
      {stage1_31[29]},
      {stage2_31[12]}
   );
   gpc1_1 gpc1047 (
      {stage1_31[30]},
      {stage2_31[13]}
   );
   gpc1_1 gpc1048 (
      {stage1_31[31]},
      {stage2_31[14]}
   );
   gpc1_1 gpc1049 (
      {stage1_31[32]},
      {stage2_31[15]}
   );
   gpc1_1 gpc1050 (
      {stage1_31[33]},
      {stage2_31[16]}
   );
   gpc1_1 gpc1051 (
      {stage1_32[18]},
      {stage2_32[11]}
   );
   gpc1_1 gpc1052 (
      {stage1_33[41]},
      {stage2_33[11]}
   );
   gpc1_1 gpc1053 (
      {stage1_33[42]},
      {stage2_33[12]}
   );
   gpc1_1 gpc1054 (
      {stage1_33[43]},
      {stage2_33[13]}
   );
   gpc1_1 gpc1055 (
      {stage1_33[44]},
      {stage2_33[14]}
   );
   gpc1_1 gpc1056 (
      {stage1_33[45]},
      {stage2_33[15]}
   );
   gpc1_1 gpc1057 (
      {stage1_34[16]},
      {stage2_34[13]}
   );
   gpc1_1 gpc1058 (
      {stage1_34[17]},
      {stage2_34[14]}
   );
   gpc1_1 gpc1059 (
      {stage1_34[18]},
      {stage2_34[15]}
   );
   gpc1_1 gpc1060 (
      {stage1_35[27]},
      {stage2_35[10]}
   );
   gpc1_1 gpc1061 (
      {stage1_36[23]},
      {stage2_36[8]}
   );
   gpc1_1 gpc1062 (
      {stage1_36[24]},
      {stage2_36[9]}
   );
   gpc1_1 gpc1063 (
      {stage1_36[25]},
      {stage2_36[10]}
   );
   gpc1_1 gpc1064 (
      {stage1_36[26]},
      {stage2_36[11]}
   );
   gpc1_1 gpc1065 (
      {stage1_36[27]},
      {stage2_36[12]}
   );
   gpc1_1 gpc1066 (
      {stage1_36[28]},
      {stage2_36[13]}
   );
   gpc1_1 gpc1067 (
      {stage1_36[29]},
      {stage2_36[14]}
   );
   gpc1_1 gpc1068 (
      {stage1_36[30]},
      {stage2_36[15]}
   );
   gpc1_1 gpc1069 (
      {stage1_36[31]},
      {stage2_36[16]}
   );
   gpc1_1 gpc1070 (
      {stage1_36[32]},
      {stage2_36[17]}
   );
   gpc1_1 gpc1071 (
      {stage1_36[33]},
      {stage2_36[18]}
   );
   gpc1_1 gpc1072 (
      {stage1_37[19]},
      {stage2_37[11]}
   );
   gpc1_1 gpc1073 (
      {stage1_37[20]},
      {stage2_37[12]}
   );
   gpc1_1 gpc1074 (
      {stage1_37[21]},
      {stage2_37[13]}
   );
   gpc1_1 gpc1075 (
      {stage1_37[22]},
      {stage2_37[14]}
   );
   gpc1_1 gpc1076 (
      {stage1_37[23]},
      {stage2_37[15]}
   );
   gpc1_1 gpc1077 (
      {stage1_37[24]},
      {stage2_37[16]}
   );
   gpc1_1 gpc1078 (
      {stage1_38[21]},
      {stage2_38[10]}
   );
   gpc1_1 gpc1079 (
      {stage1_38[22]},
      {stage2_38[11]}
   );
   gpc1_1 gpc1080 (
      {stage1_38[23]},
      {stage2_38[12]}
   );
   gpc1_1 gpc1081 (
      {stage1_39[21]},
      {stage2_39[7]}
   );
   gpc1_1 gpc1082 (
      {stage1_39[22]},
      {stage2_39[8]}
   );
   gpc1_1 gpc1083 (
      {stage1_39[23]},
      {stage2_39[9]}
   );
   gpc1_1 gpc1084 (
      {stage1_39[24]},
      {stage2_39[10]}
   );
   gpc1_1 gpc1085 (
      {stage1_39[25]},
      {stage2_39[11]}
   );
   gpc1_1 gpc1086 (
      {stage1_39[26]},
      {stage2_39[12]}
   );
   gpc1_1 gpc1087 (
      {stage1_39[27]},
      {stage2_39[13]}
   );
   gpc1_1 gpc1088 (
      {stage1_39[28]},
      {stage2_39[14]}
   );
   gpc1_1 gpc1089 (
      {stage1_39[29]},
      {stage2_39[15]}
   );
   gpc1_1 gpc1090 (
      {stage1_39[30]},
      {stage2_39[16]}
   );
   gpc1_1 gpc1091 (
      {stage1_41[18]},
      {stage2_41[11]}
   );
   gpc1_1 gpc1092 (
      {stage1_41[19]},
      {stage2_41[12]}
   );
   gpc1_1 gpc1093 (
      {stage1_42[15]},
      {stage2_42[8]}
   );
   gpc1_1 gpc1094 (
      {stage1_42[16]},
      {stage2_42[9]}
   );
   gpc1_1 gpc1095 (
      {stage1_42[17]},
      {stage2_42[10]}
   );
   gpc1_1 gpc1096 (
      {stage1_42[18]},
      {stage2_42[11]}
   );
   gpc1_1 gpc1097 (
      {stage1_42[19]},
      {stage2_42[12]}
   );
   gpc1_1 gpc1098 (
      {stage1_42[20]},
      {stage2_42[13]}
   );
   gpc1_1 gpc1099 (
      {stage1_43[21]},
      {stage2_43[8]}
   );
   gpc1_1 gpc1100 (
      {stage1_43[22]},
      {stage2_43[9]}
   );
   gpc1_1 gpc1101 (
      {stage1_44[18]},
      {stage2_44[11]}
   );
   gpc1_1 gpc1102 (
      {stage1_44[19]},
      {stage2_44[12]}
   );
   gpc1_1 gpc1103 (
      {stage1_44[20]},
      {stage2_44[13]}
   );
   gpc1_1 gpc1104 (
      {stage1_44[21]},
      {stage2_44[14]}
   );
   gpc1_1 gpc1105 (
      {stage1_45[28]},
      {stage2_45[8]}
   );
   gpc1_1 gpc1106 (
      {stage1_45[29]},
      {stage2_45[9]}
   );
   gpc1_1 gpc1107 (
      {stage1_45[30]},
      {stage2_45[10]}
   );
   gpc1_1 gpc1108 (
      {stage1_45[31]},
      {stage2_45[11]}
   );
   gpc1_1 gpc1109 (
      {stage1_46[20]},
      {stage2_46[8]}
   );
   gpc1_1 gpc1110 (
      {stage1_46[21]},
      {stage2_46[9]}
   );
   gpc1_1 gpc1111 (
      {stage1_46[22]},
      {stage2_46[10]}
   );
   gpc1_1 gpc1112 (
      {stage1_46[23]},
      {stage2_46[11]}
   );
   gpc1_1 gpc1113 (
      {stage1_46[24]},
      {stage2_46[12]}
   );
   gpc1_1 gpc1114 (
      {stage1_46[25]},
      {stage2_46[13]}
   );
   gpc1_1 gpc1115 (
      {stage1_46[26]},
      {stage2_46[14]}
   );
   gpc1_1 gpc1116 (
      {stage1_46[27]},
      {stage2_46[15]}
   );
   gpc1_1 gpc1117 (
      {stage1_46[28]},
      {stage2_46[16]}
   );
   gpc1_1 gpc1118 (
      {stage1_46[29]},
      {stage2_46[17]}
   );
   gpc1_1 gpc1119 (
      {stage1_47[22]},
      {stage2_47[10]}
   );
   gpc1_1 gpc1120 (
      {stage1_47[23]},
      {stage2_47[11]}
   );
   gpc1_1 gpc1121 (
      {stage1_47[24]},
      {stage2_47[12]}
   );
   gpc1_1 gpc1122 (
      {stage1_47[25]},
      {stage2_47[13]}
   );
   gpc1_1 gpc1123 (
      {stage1_47[26]},
      {stage2_47[14]}
   );
   gpc1_1 gpc1124 (
      {stage1_47[27]},
      {stage2_47[15]}
   );
   gpc1_1 gpc1125 (
      {stage1_47[28]},
      {stage2_47[16]}
   );
   gpc1_1 gpc1126 (
      {stage1_47[29]},
      {stage2_47[17]}
   );
   gpc1_1 gpc1127 (
      {stage1_47[30]},
      {stage2_47[18]}
   );
   gpc1_1 gpc1128 (
      {stage1_47[31]},
      {stage2_47[19]}
   );
   gpc1_1 gpc1129 (
      {stage1_47[32]},
      {stage2_47[20]}
   );
   gpc1_1 gpc1130 (
      {stage1_47[33]},
      {stage2_47[21]}
   );
   gpc1_1 gpc1131 (
      {stage1_48[14]},
      {stage2_48[9]}
   );
   gpc1_1 gpc1132 (
      {stage1_48[15]},
      {stage2_48[10]}
   );
   gpc1_1 gpc1133 (
      {stage1_48[16]},
      {stage2_48[11]}
   );
   gpc1_1 gpc1134 (
      {stage1_48[17]},
      {stage2_48[12]}
   );
   gpc1_1 gpc1135 (
      {stage1_49[12]},
      {stage2_49[6]}
   );
   gpc1_1 gpc1136 (
      {stage1_49[13]},
      {stage2_49[7]}
   );
   gpc1_1 gpc1137 (
      {stage1_49[14]},
      {stage2_49[8]}
   );
   gpc1_1 gpc1138 (
      {stage1_49[15]},
      {stage2_49[9]}
   );
   gpc1_1 gpc1139 (
      {stage1_49[16]},
      {stage2_49[10]}
   );
   gpc1_1 gpc1140 (
      {stage1_49[17]},
      {stage2_49[11]}
   );
   gpc1_1 gpc1141 (
      {stage1_49[18]},
      {stage2_49[12]}
   );
   gpc1_1 gpc1142 (
      {stage1_49[19]},
      {stage2_49[13]}
   );
   gpc1_1 gpc1143 (
      {stage1_49[20]},
      {stage2_49[14]}
   );
   gpc1_1 gpc1144 (
      {stage1_49[21]},
      {stage2_49[15]}
   );
   gpc1_1 gpc1145 (
      {stage1_49[22]},
      {stage2_49[16]}
   );
   gpc1_1 gpc1146 (
      {stage1_49[23]},
      {stage2_49[17]}
   );
   gpc1_1 gpc1147 (
      {stage1_50[42]},
      {stage2_50[10]}
   );
   gpc1_1 gpc1148 (
      {stage1_51[46]},
      {stage2_51[15]}
   );
   gpc1_1 gpc1149 (
      {stage1_51[47]},
      {stage2_51[16]}
   );
   gpc1_1 gpc1150 (
      {stage1_52[17]},
      {stage2_52[14]}
   );
   gpc1_1 gpc1151 (
      {stage1_52[18]},
      {stage2_52[15]}
   );
   gpc1_1 gpc1152 (
      {stage1_52[19]},
      {stage2_52[16]}
   );
   gpc1_1 gpc1153 (
      {stage1_52[20]},
      {stage2_52[17]}
   );
   gpc1_1 gpc1154 (
      {stage1_52[21]},
      {stage2_52[18]}
   );
   gpc1_1 gpc1155 (
      {stage1_53[40]},
      {stage2_53[12]}
   );
   gpc1_1 gpc1156 (
      {stage1_54[16]},
      {stage2_54[14]}
   );
   gpc1_1 gpc1157 (
      {stage1_55[32]},
      {stage2_55[13]}
   );
   gpc1_1 gpc1158 (
      {stage1_55[33]},
      {stage2_55[14]}
   );
   gpc1_1 gpc1159 (
      {stage1_55[34]},
      {stage2_55[15]}
   );
   gpc1_1 gpc1160 (
      {stage1_55[35]},
      {stage2_55[16]}
   );
   gpc1_1 gpc1161 (
      {stage1_55[36]},
      {stage2_55[17]}
   );
   gpc1_1 gpc1162 (
      {stage1_55[37]},
      {stage2_55[18]}
   );
   gpc1_1 gpc1163 (
      {stage1_56[17]},
      {stage2_56[9]}
   );
   gpc1_1 gpc1164 (
      {stage1_56[18]},
      {stage2_56[10]}
   );
   gpc1_1 gpc1165 (
      {stage1_56[19]},
      {stage2_56[11]}
   );
   gpc1_1 gpc1166 (
      {stage1_56[20]},
      {stage2_56[12]}
   );
   gpc1_1 gpc1167 (
      {stage1_57[37]},
      {stage2_57[9]}
   );
   gpc1_1 gpc1168 (
      {stage1_57[38]},
      {stage2_57[10]}
   );
   gpc1_1 gpc1169 (
      {stage1_57[39]},
      {stage2_57[11]}
   );
   gpc1_1 gpc1170 (
      {stage1_57[40]},
      {stage2_57[12]}
   );
   gpc1_1 gpc1171 (
      {stage1_58[6]},
      {stage2_58[9]}
   );
   gpc1_1 gpc1172 (
      {stage1_58[7]},
      {stage2_58[10]}
   );
   gpc1_1 gpc1173 (
      {stage1_58[8]},
      {stage2_58[11]}
   );
   gpc1_1 gpc1174 (
      {stage1_58[9]},
      {stage2_58[12]}
   );
   gpc1_1 gpc1175 (
      {stage1_58[10]},
      {stage2_58[13]}
   );
   gpc1_1 gpc1176 (
      {stage1_58[11]},
      {stage2_58[14]}
   );
   gpc1_1 gpc1177 (
      {stage1_58[12]},
      {stage2_58[15]}
   );
   gpc1_1 gpc1178 (
      {stage1_58[13]},
      {stage2_58[16]}
   );
   gpc1_1 gpc1179 (
      {stage1_58[14]},
      {stage2_58[17]}
   );
   gpc1_1 gpc1180 (
      {stage1_60[18]},
      {stage2_60[8]}
   );
   gpc1_1 gpc1181 (
      {stage1_60[19]},
      {stage2_60[9]}
   );
   gpc1_1 gpc1182 (
      {stage1_60[20]},
      {stage2_60[10]}
   );
   gpc1_1 gpc1183 (
      {stage1_60[21]},
      {stage2_60[11]}
   );
   gpc1_1 gpc1184 (
      {stage1_60[22]},
      {stage2_60[12]}
   );
   gpc1_1 gpc1185 (
      {stage1_61[18]},
      {stage2_61[9]}
   );
   gpc1_1 gpc1186 (
      {stage1_61[19]},
      {stage2_61[10]}
   );
   gpc1_1 gpc1187 (
      {stage1_61[20]},
      {stage2_61[11]}
   );
   gpc1_1 gpc1188 (
      {stage1_62[18]},
      {stage2_62[12]}
   );
   gpc1_1 gpc1189 (
      {stage1_62[19]},
      {stage2_62[13]}
   );
   gpc1_1 gpc1190 (
      {stage1_62[20]},
      {stage2_62[14]}
   );
   gpc1_1 gpc1191 (
      {stage1_62[21]},
      {stage2_62[15]}
   );
   gpc1_1 gpc1192 (
      {stage1_62[22]},
      {stage2_62[16]}
   );
   gpc1_1 gpc1193 (
      {stage1_62[23]},
      {stage2_62[17]}
   );
   gpc1_1 gpc1194 (
      {stage1_63[24]},
      {stage2_63[6]}
   );
   gpc1_1 gpc1195 (
      {stage1_63[25]},
      {stage2_63[7]}
   );
   gpc1_1 gpc1196 (
      {stage1_63[26]},
      {stage2_63[8]}
   );
   gpc1_1 gpc1197 (
      {stage1_63[27]},
      {stage2_63[9]}
   );
   gpc1_1 gpc1198 (
      {stage1_63[28]},
      {stage2_63[10]}
   );
   gpc1_1 gpc1199 (
      {stage1_63[29]},
      {stage2_63[11]}
   );
   gpc1_1 gpc1200 (
      {stage1_63[30]},
      {stage2_63[12]}
   );
   gpc1_1 gpc1201 (
      {stage1_63[31]},
      {stage2_63[13]}
   );
   gpc1_1 gpc1202 (
      {stage1_63[32]},
      {stage2_63[14]}
   );
   gpc1_1 gpc1203 (
      {stage1_63[33]},
      {stage2_63[15]}
   );
   gpc1_1 gpc1204 (
      {stage1_63[34]},
      {stage2_63[16]}
   );
   gpc1_1 gpc1205 (
      {stage1_65[2]},
      {stage2_65[6]}
   );
   gpc1_1 gpc1206 (
      {stage1_65[3]},
      {stage2_65[7]}
   );
   gpc1_1 gpc1207 (
      {stage1_65[4]},
      {stage2_65[8]}
   );
   gpc1_1 gpc1208 (
      {stage1_65[5]},
      {stage2_65[9]}
   );
   gpc615_5 gpc1209 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc1210 (
      {stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc606_5 gpc1211 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc606_5 gpc1212 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[3]}
   );
   gpc2135_5 gpc1213 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4]},
      {stage2_6[6], stage2_6[7], stage2_6[8]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1]},
      {stage3_9[0],stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[3]}
   );
   gpc615_5 gpc1214 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6]},
      {stage2_9[0]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc1215 (
      {stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[2]}
   );
   gpc606_5 gpc1216 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[3]}
   );
   gpc615_5 gpc1217 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4]},
      {stage2_13[0]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[2],stage3_12[3]}
   );
   gpc615_5 gpc1218 (
      {stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9]},
      {stage2_13[1]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[1],stage3_14[1],stage3_13[3],stage3_12[4]}
   );
   gpc623_5 gpc1219 (
      {stage2_13[2], stage2_13[3], stage2_13[4]},
      {stage2_14[12], stage2_14[13]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[2],stage3_15[2],stage3_14[2],stage3_13[4]}
   );
   gpc623_5 gpc1220 (
      {stage2_13[5], stage2_13[6], stage2_13[7]},
      {stage2_14[14], 1'b0},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[3],stage3_15[3],stage3_14[3],stage3_13[5]}
   );
   gpc135_4 gpc1221 (
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4]},
      {stage2_17[0], stage2_17[1], stage2_17[2]},
      {stage2_18[0]},
      {stage3_19[0],stage3_18[0],stage3_17[2],stage3_16[4]}
   );
   gpc606_5 gpc1222 (
      {stage2_16[5], stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10]},
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage3_20[0],stage3_19[1],stage3_18[1],stage3_17[3],stage3_16[5]}
   );
   gpc606_5 gpc1223 (
      {stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6], stage2_17[7], stage2_17[8]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[2],stage3_18[2],stage3_17[4]}
   );
   gpc1406_5 gpc1224 (
      {stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3]},
      {stage2_21[0]},
      {stage3_22[0],stage3_21[1],stage3_20[2],stage3_19[3],stage3_18[3]}
   );
   gpc1406_5 gpc1225 (
      {stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18]},
      {stage2_20[4], stage2_20[5], stage2_20[6], stage2_20[7]},
      {stage2_21[1]},
      {stage3_22[1],stage3_21[2],stage3_20[3],stage3_19[4],stage3_18[4]}
   );
   gpc615_5 gpc1226 (
      {stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5], stage2_21[6]},
      {stage2_22[0]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[2],stage3_21[3]}
   );
   gpc615_5 gpc1227 (
      {stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_22[1]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[3],stage3_21[4]}
   );
   gpc615_5 gpc1228 (
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16]},
      {stage2_22[2]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[4],stage3_21[5]}
   );
   gpc1325_5 gpc1229 (
      {stage2_21[17], stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21]},
      {stage2_22[3], stage2_22[4]},
      {stage2_23[18], stage2_23[19], stage2_23[20]},
      {stage2_24[0]},
      {stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[5],stage3_21[6]}
   );
   gpc606_5 gpc1230 (
      {stage2_22[5], stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6]},
      {stage3_26[0],stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[6]}
   );
   gpc1343_5 gpc1231 (
      {stage2_24[7], stage2_24[8], stage2_24[9]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3]},
      {stage2_26[0], stage2_26[1], stage2_26[2]},
      {stage2_27[0]},
      {stage3_28[0],stage3_27[0],stage3_26[1],stage3_25[5],stage3_24[5]}
   );
   gpc1325_5 gpc1232 (
      {stage2_25[4], stage2_25[5], stage2_25[6], stage2_25[7], stage2_25[8]},
      {stage2_26[3], stage2_26[4]},
      {stage2_27[1], stage2_27[2], stage2_27[3]},
      {stage2_28[0]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[2],stage3_25[6]}
   );
   gpc1325_5 gpc1233 (
      {stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12], 1'b0},
      {stage2_26[5], stage2_26[6]},
      {stage2_27[4], stage2_27[5], stage2_27[6]},
      {stage2_28[1]},
      {stage3_29[1],stage3_28[2],stage3_27[2],stage3_26[3],stage3_25[7]}
   );
   gpc606_5 gpc1234 (
      {stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12]},
      {stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7]},
      {stage3_30[0],stage3_29[2],stage3_28[3],stage3_27[3],stage3_26[4]}
   );
   gpc606_5 gpc1235 (
      {stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18]},
      {stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage3_30[1],stage3_29[3],stage3_28[4],stage3_27[4],stage3_26[5]}
   );
   gpc606_5 gpc1236 (
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[0],stage3_31[0],stage3_30[2],stage3_29[4]}
   );
   gpc606_5 gpc1237 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[1],stage3_31[1],stage3_30[3],stage3_29[5]}
   );
   gpc615_5 gpc1238 (
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4]},
      {stage2_31[12]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[2],stage3_32[2],stage3_31[2],stage3_30[4]}
   );
   gpc615_5 gpc1239 (
      {stage2_30[5], stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9]},
      {stage2_31[13]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[3],stage3_32[3],stage3_31[3],stage3_30[5]}
   );
   gpc606_5 gpc1240 (
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[0],stage3_35[0],stage3_34[2],stage3_33[4]}
   );
   gpc606_5 gpc1241 (
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[1],stage3_36[1],stage3_35[1],stage3_34[3]}
   );
   gpc606_5 gpc1242 (
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[2],stage3_36[2],stage3_35[2],stage3_34[4]}
   );
   gpc615_5 gpc1243 (
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10]},
      {stage2_36[12]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[2],stage3_37[3],stage3_36[3],stage3_35[3]}
   );
   gpc615_5 gpc1244 (
      {stage2_36[13], stage2_36[14], stage2_36[15], stage2_36[16], stage2_36[17]},
      {stage2_37[6]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[1],stage3_38[3],stage3_37[4],stage3_36[4]}
   );
   gpc615_5 gpc1245 (
      {stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage2_38[6]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[1],stage3_39[2],stage3_38[4],stage3_37[5]}
   );
   gpc615_5 gpc1246 (
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16]},
      {stage2_38[7]},
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage3_41[1],stage3_40[2],stage3_39[3],stage3_38[5],stage3_37[6]}
   );
   gpc207_4 gpc1247 (
      {stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11], stage2_38[12], 1'b0, 1'b0},
      {stage2_40[0], stage2_40[1]},
      {stage3_41[2],stage3_40[3],stage3_39[4],stage3_38[6]}
   );
   gpc615_5 gpc1248 (
      {stage2_39[12], stage2_39[13], stage2_39[14], stage2_39[15], stage2_39[16]},
      {stage2_40[2]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[0],stage3_41[3],stage3_40[4],stage3_39[5]}
   );
   gpc606_5 gpc1249 (
      {stage2_40[3], stage2_40[4], stage2_40[5], stage2_40[6], stage2_40[7], stage2_40[8]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[1],stage3_42[1],stage3_41[4],stage3_40[5]}
   );
   gpc623_5 gpc1250 (
      {stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage2_41[6], stage2_41[7]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[2],stage3_42[2],stage3_41[5],stage3_40[6]}
   );
   gpc606_5 gpc1251 (
      {stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11], stage2_41[12], 1'b0},
      {stage2_43[0], stage2_43[1], stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5]},
      {stage3_45[0],stage3_44[2],stage3_43[3],stage3_42[3],stage3_41[6]}
   );
   gpc606_5 gpc1252 (
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[0],stage3_46[0],stage3_45[1],stage3_44[3]}
   );
   gpc606_5 gpc1253 (
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[1],stage3_46[1],stage3_45[2],stage3_44[4]}
   );
   gpc606_5 gpc1254 (
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[2],stage3_47[2],stage3_46[2],stage3_45[3]}
   );
   gpc606_5 gpc1255 (
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[3],stage3_47[3],stage3_46[3],stage3_45[4]}
   );
   gpc615_5 gpc1256 (
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16]},
      {stage2_47[12]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[2],stage3_48[4],stage3_47[4],stage3_46[4]}
   );
   gpc606_5 gpc1257 (
      {stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17], stage2_47[18]},
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5]},
      {stage3_51[0],stage3_50[1],stage3_49[3],stage3_48[5],stage3_47[5]}
   );
   gpc606_5 gpc1258 (
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage3_53[0],stage3_52[0],stage3_51[1],stage3_50[2],stage3_49[4]}
   );
   gpc606_5 gpc1259 (
      {stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17]},
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11]},
      {stage3_53[1],stage3_52[1],stage3_51[2],stage3_50[3],stage3_49[5]}
   );
   gpc615_5 gpc1260 (
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4]},
      {stage2_51[12]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[2],stage3_52[2],stage3_51[3],stage3_50[4]}
   );
   gpc606_5 gpc1261 (
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[0],stage3_54[1],stage3_53[3],stage3_52[3]}
   );
   gpc606_5 gpc1262 (
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[1],stage3_55[1],stage3_54[2],stage3_53[4]}
   );
   gpc606_5 gpc1263 (
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[2],stage3_55[2],stage3_54[3],stage3_53[5]}
   );
   gpc135_4 gpc1264 (
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10]},
      {stage2_55[12], stage2_55[13], stage2_55[14]},
      {stage2_56[0]},
      {stage3_57[2],stage3_56[3],stage3_55[3],stage3_54[4]}
   );
   gpc135_4 gpc1265 (
      {stage2_54[11], stage2_54[12], stage2_54[13], stage2_54[14], 1'b0},
      {stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage2_56[1]},
      {stage3_57[3],stage3_56[4],stage3_55[4],stage3_54[5]}
   );
   gpc606_5 gpc1266 (
      {stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5], stage2_56[6], stage2_56[7]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[0],stage3_57[4],stage3_56[5]}
   );
   gpc135_4 gpc1267 (
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4]},
      {stage2_58[6], stage2_58[7], stage2_58[8]},
      {stage2_59[0]},
      {stage3_60[1],stage3_59[1],stage3_58[1],stage3_57[5]}
   );
   gpc135_4 gpc1268 (
      {stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9]},
      {stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage2_59[1]},
      {stage3_60[2],stage3_59[2],stage3_58[2],stage3_57[6]}
   );
   gpc1163_5 gpc1269 (
      {stage2_57[10], stage2_57[11], stage2_57[12]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage2_59[2]},
      {stage2_60[0]},
      {stage3_61[0],stage3_60[3],stage3_59[3],stage3_58[3],stage3_57[7]}
   );
   gpc606_5 gpc1270 (
      {stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5], stage2_60[6]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[0],stage3_62[0],stage3_61[1],stage3_60[4]}
   );
   gpc606_5 gpc1271 (
      {stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11], stage2_60[12]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[1],stage3_62[1],stage3_61[2],stage3_60[5]}
   );
   gpc606_5 gpc1272 (
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[2],stage3_63[2],stage3_62[2],stage3_61[3]}
   );
   gpc606_5 gpc1273 (
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[1],stage3_64[3],stage3_63[3],stage3_62[3]}
   );
   gpc606_5 gpc1274 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage2_65[0], stage2_65[1], stage2_65[2], stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage3_67[0],stage3_66[1],stage3_65[2],stage3_64[4],stage3_63[4]}
   );
   gpc1_1 gpc1275 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc1276 (
      {stage2_2[12]},
      {stage3_2[3]}
   );
   gpc1_1 gpc1277 (
      {stage2_2[13]},
      {stage3_2[4]}
   );
   gpc1_1 gpc1278 (
      {stage2_3[6]},
      {stage3_3[3]}
   );
   gpc1_1 gpc1279 (
      {stage2_3[7]},
      {stage3_3[4]}
   );
   gpc1_1 gpc1280 (
      {stage2_3[8]},
      {stage3_3[5]}
   );
   gpc1_1 gpc1281 (
      {stage2_4[12]},
      {stage3_4[4]}
   );
   gpc1_1 gpc1282 (
      {stage2_4[13]},
      {stage3_4[5]}
   );
   gpc1_1 gpc1283 (
      {stage2_4[14]},
      {stage3_4[6]}
   );
   gpc1_1 gpc1284 (
      {stage2_4[15]},
      {stage3_4[7]}
   );
   gpc1_1 gpc1285 (
      {stage2_4[16]},
      {stage3_4[8]}
   );
   gpc1_1 gpc1286 (
      {stage2_4[17]},
      {stage3_4[9]}
   );
   gpc1_1 gpc1287 (
      {stage2_4[18]},
      {stage3_4[10]}
   );
   gpc1_1 gpc1288 (
      {stage2_4[19]},
      {stage3_4[11]}
   );
   gpc1_1 gpc1289 (
      {stage2_4[20]},
      {stage3_4[12]}
   );
   gpc1_1 gpc1290 (
      {stage2_4[21]},
      {stage3_4[13]}
   );
   gpc1_1 gpc1291 (
      {stage2_4[22]},
      {stage3_4[14]}
   );
   gpc1_1 gpc1292 (
      {stage2_5[5]},
      {stage3_5[4]}
   );
   gpc1_1 gpc1293 (
      {stage2_5[6]},
      {stage3_5[5]}
   );
   gpc1_1 gpc1294 (
      {stage2_5[7]},
      {stage3_5[6]}
   );
   gpc1_1 gpc1295 (
      {stage2_5[8]},
      {stage3_5[7]}
   );
   gpc1_1 gpc1296 (
      {stage2_5[9]},
      {stage3_5[8]}
   );
   gpc1_1 gpc1297 (
      {stage2_6[9]},
      {stage3_6[3]}
   );
   gpc1_1 gpc1298 (
      {stage2_6[10]},
      {stage3_6[4]}
   );
   gpc1_1 gpc1299 (
      {stage2_7[1]},
      {stage3_7[2]}
   );
   gpc1_1 gpc1300 (
      {stage2_7[2]},
      {stage3_7[3]}
   );
   gpc1_1 gpc1301 (
      {stage2_7[3]},
      {stage3_7[4]}
   );
   gpc1_1 gpc1302 (
      {stage2_7[4]},
      {stage3_7[5]}
   );
   gpc1_1 gpc1303 (
      {stage2_7[5]},
      {stage3_7[6]}
   );
   gpc1_1 gpc1304 (
      {stage2_7[6]},
      {stage3_7[7]}
   );
   gpc1_1 gpc1305 (
      {stage2_7[7]},
      {stage3_7[8]}
   );
   gpc1_1 gpc1306 (
      {stage2_7[8]},
      {stage3_7[9]}
   );
   gpc1_1 gpc1307 (
      {stage2_7[9]},
      {stage3_7[10]}
   );
   gpc1_1 gpc1308 (
      {stage2_7[10]},
      {stage3_7[11]}
   );
   gpc1_1 gpc1309 (
      {stage2_7[11]},
      {stage3_7[12]}
   );
   gpc1_1 gpc1310 (
      {stage2_7[12]},
      {stage3_7[13]}
   );
   gpc1_1 gpc1311 (
      {stage2_8[7]},
      {stage3_8[3]}
   );
   gpc1_1 gpc1312 (
      {stage2_8[8]},
      {stage3_8[4]}
   );
   gpc1_1 gpc1313 (
      {stage2_8[9]},
      {stage3_8[5]}
   );
   gpc1_1 gpc1314 (
      {stage2_8[10]},
      {stage3_8[6]}
   );
   gpc1_1 gpc1315 (
      {stage2_9[13]},
      {stage3_9[4]}
   );
   gpc1_1 gpc1316 (
      {stage2_9[14]},
      {stage3_9[5]}
   );
   gpc1_1 gpc1317 (
      {stage2_9[15]},
      {stage3_9[6]}
   );
   gpc1_1 gpc1318 (
      {stage2_9[16]},
      {stage3_9[7]}
   );
   gpc1_1 gpc1319 (
      {stage2_9[17]},
      {stage3_9[8]}
   );
   gpc1_1 gpc1320 (
      {stage2_9[18]},
      {stage3_9[9]}
   );
   gpc1_1 gpc1321 (
      {stage2_9[19]},
      {stage3_9[10]}
   );
   gpc1_1 gpc1322 (
      {stage2_10[6]},
      {stage3_10[3]}
   );
   gpc1_1 gpc1323 (
      {stage2_10[7]},
      {stage3_10[4]}
   );
   gpc1_1 gpc1324 (
      {stage2_10[8]},
      {stage3_10[5]}
   );
   gpc1_1 gpc1325 (
      {stage2_10[9]},
      {stage3_10[6]}
   );
   gpc1_1 gpc1326 (
      {stage2_11[12]},
      {stage3_11[3]}
   );
   gpc1_1 gpc1327 (
      {stage2_13[8]},
      {stage3_13[6]}
   );
   gpc1_1 gpc1328 (
      {stage2_13[9]},
      {stage3_13[7]}
   );
   gpc1_1 gpc1329 (
      {stage2_15[12]},
      {stage3_15[4]}
   );
   gpc1_1 gpc1330 (
      {stage2_15[13]},
      {stage3_15[5]}
   );
   gpc1_1 gpc1331 (
      {stage2_17[9]},
      {stage3_17[5]}
   );
   gpc1_1 gpc1332 (
      {stage2_17[10]},
      {stage3_17[6]}
   );
   gpc1_1 gpc1333 (
      {stage2_17[11]},
      {stage3_17[7]}
   );
   gpc1_1 gpc1334 (
      {stage2_18[19]},
      {stage3_18[5]}
   );
   gpc1_1 gpc1335 (
      {stage2_19[6]},
      {stage3_19[5]}
   );
   gpc1_1 gpc1336 (
      {stage2_19[7]},
      {stage3_19[6]}
   );
   gpc1_1 gpc1337 (
      {stage2_19[8]},
      {stage3_19[7]}
   );
   gpc1_1 gpc1338 (
      {stage2_20[8]},
      {stage3_20[4]}
   );
   gpc1_1 gpc1339 (
      {stage2_29[12]},
      {stage3_29[6]}
   );
   gpc1_1 gpc1340 (
      {stage2_29[13]},
      {stage3_29[7]}
   );
   gpc1_1 gpc1341 (
      {stage2_29[14]},
      {stage3_29[8]}
   );
   gpc1_1 gpc1342 (
      {stage2_29[15]},
      {stage3_29[9]}
   );
   gpc1_1 gpc1343 (
      {stage2_29[16]},
      {stage3_29[10]}
   );
   gpc1_1 gpc1344 (
      {stage2_29[17]},
      {stage3_29[11]}
   );
   gpc1_1 gpc1345 (
      {stage2_31[14]},
      {stage3_31[4]}
   );
   gpc1_1 gpc1346 (
      {stage2_31[15]},
      {stage3_31[5]}
   );
   gpc1_1 gpc1347 (
      {stage2_31[16]},
      {stage3_31[6]}
   );
   gpc1_1 gpc1348 (
      {stage2_33[6]},
      {stage3_33[5]}
   );
   gpc1_1 gpc1349 (
      {stage2_33[7]},
      {stage3_33[6]}
   );
   gpc1_1 gpc1350 (
      {stage2_33[8]},
      {stage3_33[7]}
   );
   gpc1_1 gpc1351 (
      {stage2_33[9]},
      {stage3_33[8]}
   );
   gpc1_1 gpc1352 (
      {stage2_33[10]},
      {stage3_33[9]}
   );
   gpc1_1 gpc1353 (
      {stage2_33[11]},
      {stage3_33[10]}
   );
   gpc1_1 gpc1354 (
      {stage2_33[12]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1355 (
      {stage2_33[13]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1356 (
      {stage2_33[14]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1357 (
      {stage2_33[15]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1358 (
      {stage2_34[12]},
      {stage3_34[5]}
   );
   gpc1_1 gpc1359 (
      {stage2_34[13]},
      {stage3_34[6]}
   );
   gpc1_1 gpc1360 (
      {stage2_34[14]},
      {stage3_34[7]}
   );
   gpc1_1 gpc1361 (
      {stage2_34[15]},
      {stage3_34[8]}
   );
   gpc1_1 gpc1362 (
      {stage2_36[18]},
      {stage3_36[5]}
   );
   gpc1_1 gpc1363 (
      {stage2_42[12]},
      {stage3_42[4]}
   );
   gpc1_1 gpc1364 (
      {stage2_42[13]},
      {stage3_42[5]}
   );
   gpc1_1 gpc1365 (
      {stage2_43[6]},
      {stage3_43[4]}
   );
   gpc1_1 gpc1366 (
      {stage2_43[7]},
      {stage3_43[5]}
   );
   gpc1_1 gpc1367 (
      {stage2_43[8]},
      {stage3_43[6]}
   );
   gpc1_1 gpc1368 (
      {stage2_43[9]},
      {stage3_43[7]}
   );
   gpc1_1 gpc1369 (
      {stage2_44[12]},
      {stage3_44[5]}
   );
   gpc1_1 gpc1370 (
      {stage2_44[13]},
      {stage3_44[6]}
   );
   gpc1_1 gpc1371 (
      {stage2_44[14]},
      {stage3_44[7]}
   );
   gpc1_1 gpc1372 (
      {stage2_46[17]},
      {stage3_46[5]}
   );
   gpc1_1 gpc1373 (
      {stage2_47[19]},
      {stage3_47[6]}
   );
   gpc1_1 gpc1374 (
      {stage2_47[20]},
      {stage3_47[7]}
   );
   gpc1_1 gpc1375 (
      {stage2_47[21]},
      {stage3_47[8]}
   );
   gpc1_1 gpc1376 (
      {stage2_48[6]},
      {stage3_48[6]}
   );
   gpc1_1 gpc1377 (
      {stage2_48[7]},
      {stage3_48[7]}
   );
   gpc1_1 gpc1378 (
      {stage2_48[8]},
      {stage3_48[8]}
   );
   gpc1_1 gpc1379 (
      {stage2_48[9]},
      {stage3_48[9]}
   );
   gpc1_1 gpc1380 (
      {stage2_48[10]},
      {stage3_48[10]}
   );
   gpc1_1 gpc1381 (
      {stage2_48[11]},
      {stage3_48[11]}
   );
   gpc1_1 gpc1382 (
      {stage2_48[12]},
      {stage3_48[12]}
   );
   gpc1_1 gpc1383 (
      {stage2_50[5]},
      {stage3_50[5]}
   );
   gpc1_1 gpc1384 (
      {stage2_50[6]},
      {stage3_50[6]}
   );
   gpc1_1 gpc1385 (
      {stage2_50[7]},
      {stage3_50[7]}
   );
   gpc1_1 gpc1386 (
      {stage2_50[8]},
      {stage3_50[8]}
   );
   gpc1_1 gpc1387 (
      {stage2_50[9]},
      {stage3_50[9]}
   );
   gpc1_1 gpc1388 (
      {stage2_50[10]},
      {stage3_50[10]}
   );
   gpc1_1 gpc1389 (
      {stage2_51[13]},
      {stage3_51[4]}
   );
   gpc1_1 gpc1390 (
      {stage2_51[14]},
      {stage3_51[5]}
   );
   gpc1_1 gpc1391 (
      {stage2_51[15]},
      {stage3_51[6]}
   );
   gpc1_1 gpc1392 (
      {stage2_51[16]},
      {stage3_51[7]}
   );
   gpc1_1 gpc1393 (
      {stage2_52[12]},
      {stage3_52[4]}
   );
   gpc1_1 gpc1394 (
      {stage2_52[13]},
      {stage3_52[5]}
   );
   gpc1_1 gpc1395 (
      {stage2_52[14]},
      {stage3_52[6]}
   );
   gpc1_1 gpc1396 (
      {stage2_52[15]},
      {stage3_52[7]}
   );
   gpc1_1 gpc1397 (
      {stage2_52[16]},
      {stage3_52[8]}
   );
   gpc1_1 gpc1398 (
      {stage2_52[17]},
      {stage3_52[9]}
   );
   gpc1_1 gpc1399 (
      {stage2_52[18]},
      {stage3_52[10]}
   );
   gpc1_1 gpc1400 (
      {stage2_53[12]},
      {stage3_53[6]}
   );
   gpc1_1 gpc1401 (
      {stage2_55[18]},
      {stage3_55[5]}
   );
   gpc1_1 gpc1402 (
      {stage2_56[8]},
      {stage3_56[6]}
   );
   gpc1_1 gpc1403 (
      {stage2_56[9]},
      {stage3_56[7]}
   );
   gpc1_1 gpc1404 (
      {stage2_56[10]},
      {stage3_56[8]}
   );
   gpc1_1 gpc1405 (
      {stage2_56[11]},
      {stage3_56[9]}
   );
   gpc1_1 gpc1406 (
      {stage2_56[12]},
      {stage3_56[10]}
   );
   gpc1_1 gpc1407 (
      {stage2_59[3]},
      {stage3_59[4]}
   );
   gpc1_1 gpc1408 (
      {stage2_59[4]},
      {stage3_59[5]}
   );
   gpc1_1 gpc1409 (
      {stage2_59[5]},
      {stage3_59[6]}
   );
   gpc1_1 gpc1410 (
      {stage2_59[6]},
      {stage3_59[7]}
   );
   gpc1_1 gpc1411 (
      {stage2_59[7]},
      {stage3_59[8]}
   );
   gpc1_1 gpc1412 (
      {stage2_59[8]},
      {stage3_59[9]}
   );
   gpc1_1 gpc1413 (
      {stage2_59[9]},
      {stage3_59[10]}
   );
   gpc1_1 gpc1414 (
      {stage2_59[10]},
      {stage3_59[11]}
   );
   gpc1_1 gpc1415 (
      {stage2_59[11]},
      {stage3_59[12]}
   );
   gpc1_1 gpc1416 (
      {stage2_59[12]},
      {stage3_59[13]}
   );
   gpc1_1 gpc1417 (
      {stage2_61[6]},
      {stage3_61[4]}
   );
   gpc1_1 gpc1418 (
      {stage2_61[7]},
      {stage3_61[5]}
   );
   gpc1_1 gpc1419 (
      {stage2_61[8]},
      {stage3_61[6]}
   );
   gpc1_1 gpc1420 (
      {stage2_61[9]},
      {stage3_61[7]}
   );
   gpc1_1 gpc1421 (
      {stage2_61[10]},
      {stage3_61[8]}
   );
   gpc1_1 gpc1422 (
      {stage2_61[11]},
      {stage3_61[9]}
   );
   gpc1_1 gpc1423 (
      {stage2_63[12]},
      {stage3_63[5]}
   );
   gpc1_1 gpc1424 (
      {stage2_63[13]},
      {stage3_63[6]}
   );
   gpc1_1 gpc1425 (
      {stage2_63[14]},
      {stage3_63[7]}
   );
   gpc1_1 gpc1426 (
      {stage2_63[15]},
      {stage3_63[8]}
   );
   gpc1_1 gpc1427 (
      {stage2_63[16]},
      {stage3_63[9]}
   );
   gpc1_1 gpc1428 (
      {stage2_65[6]},
      {stage3_65[3]}
   );
   gpc1_1 gpc1429 (
      {stage2_65[7]},
      {stage3_65[4]}
   );
   gpc1_1 gpc1430 (
      {stage2_65[8]},
      {stage3_65[5]}
   );
   gpc1_1 gpc1431 (
      {stage2_65[9]},
      {stage3_65[6]}
   );
   gpc1_1 gpc1432 (
      {stage2_66[0]},
      {stage3_66[2]}
   );
   gpc1_1 gpc1433 (
      {stage2_66[1]},
      {stage3_66[3]}
   );
   gpc1_1 gpc1434 (
      {stage2_66[2]},
      {stage3_66[4]}
   );
   gpc1_1 gpc1435 (
      {stage2_66[3]},
      {stage3_66[5]}
   );
   gpc615_5 gpc1436 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0]}
   );
   gpc615_5 gpc1437 (
      {stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage3_4[6]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[1],stage4_3[1]}
   );
   gpc2135_5 gpc1438 (
      {stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_5[6], stage3_5[7], stage3_5[8]},
      {stage3_6[0]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[2]}
   );
   gpc615_5 gpc1439 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], 1'b0},
      {stage3_7[2]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[2],stage4_6[3]}
   );
   gpc615_5 gpc1440 (
      {stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[3]}
   );
   gpc615_5 gpc1441 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12]},
      {1'b0},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], 1'b0},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[4]}
   );
   gpc7_3 gpc1442 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage4_12[0],stage4_11[2],stage4_10[3]}
   );
   gpc135_4 gpc1443 (
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], 1'b0},
      {stage3_12[0], stage3_12[1], stage3_12[2]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[1],stage4_11[3]}
   );
   gpc207_4 gpc1444 (
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7]},
      {stage3_15[0], stage3_15[1]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1]}
   );
   gpc1415_5 gpc1445 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], 1'b0},
      {stage3_15[2]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1],stage4_14[2]}
   );
   gpc117_4 gpc1446 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {stage3_18[0]},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[1]}
   );
   gpc1406_5 gpc1447 (
      {stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[0],stage4_20[1],stage4_19[1]}
   );
   gpc615_5 gpc1448 (
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[4]},
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5], stage3_22[6]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[1],stage4_20[2]}
   );
   gpc615_5 gpc1449 (
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[0],stage4_25[0],stage4_24[1],stage4_23[2]}
   );
   gpc15_3 gpc1450 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage3_25[6]},
      {stage4_26[1],stage4_25[1],stage4_24[2]}
   );
   gpc615_5 gpc1451 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4]},
      {stage3_27[0]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], 1'b0},
      {stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1],stage4_26[2]}
   );
   gpc1163_5 gpc1452 (
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[0]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[0],stage4_30[1],stage4_29[1]}
   );
   gpc606_5 gpc1453 (
      {stage3_29[3], stage3_29[4], stage3_29[5], stage3_29[6], stage3_29[7], stage3_29[8]},
      {stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5], stage3_31[6]},
      {stage4_33[1],stage4_32[1],stage4_31[1],stage4_30[2],stage4_29[2]}
   );
   gpc3_2 gpc1454 (
      {stage3_32[1], stage3_32[2], stage3_32[3]},
      {stage4_33[2],stage4_32[2]}
   );
   gpc2135_5 gpc1455 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4]},
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0]},
      {stage3_36[0], stage3_36[1]},
      {stage4_37[0],stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[3]}
   );
   gpc2135_5 gpc1456 (
      {stage3_33[5], stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9]},
      {stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage3_35[1]},
      {stage3_36[2], stage3_36[3]},
      {stage4_37[1],stage4_36[1],stage4_35[1],stage4_34[1],stage4_33[4]}
   );
   gpc2135_5 gpc1457 (
      {stage3_33[10], stage3_33[11], stage3_33[12], stage3_33[13], stage3_33[14]},
      {stage3_34[6], stage3_34[7], stage3_34[8]},
      {stage3_35[2]},
      {stage3_36[4], stage3_36[5]},
      {stage4_37[2],stage4_36[2],stage4_35[2],stage4_34[2],stage4_33[5]}
   );
   gpc615_5 gpc1458 (
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4]},
      {stage3_38[0]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[0],stage4_39[0],stage4_38[0],stage4_37[3]}
   );
   gpc2116_5 gpc1459 (
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage3_41[0]},
      {stage3_42[0]},
      {stage3_43[0], stage3_43[1]},
      {stage4_44[0],stage4_43[0],stage4_42[0],stage4_41[1],stage4_40[1]}
   );
   gpc207_4 gpc1460 (
      {stage3_41[1], stage3_41[2], stage3_41[3], stage3_41[4], stage3_41[5], stage3_41[6], 1'b0},
      {stage3_43[2], stage3_43[3]},
      {stage4_44[1],stage4_43[1],stage4_42[1],stage4_41[2]}
   );
   gpc2135_5 gpc1461 (
      {stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5]},
      {stage3_43[4], stage3_43[5], stage3_43[6]},
      {stage3_44[0]},
      {stage3_45[0], stage3_45[1]},
      {stage4_46[0],stage4_45[0],stage4_44[2],stage4_43[2],stage4_42[2]}
   );
   gpc2135_5 gpc1462 (
      {stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage3_45[2], stage3_45[3], stage3_45[4]},
      {stage3_46[0]},
      {stage3_47[0], stage3_47[1]},
      {stage4_48[0],stage4_47[0],stage4_46[1],stage4_45[1],stage4_44[3]}
   );
   gpc615_5 gpc1463 (
      {stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage3_47[2]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[1],stage4_47[1],stage4_46[2]}
   );
   gpc615_5 gpc1464 (
      {stage3_47[3], stage3_47[4], stage3_47[5], stage3_47[6], stage3_47[7]},
      {stage3_48[6]},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage4_51[0],stage4_50[1],stage4_49[1],stage4_48[2],stage4_47[2]}
   );
   gpc606_5 gpc1465 (
      {stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11], stage3_48[12]},
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage4_52[0],stage4_51[1],stage4_50[2],stage4_49[2],stage4_48[3]}
   );
   gpc615_5 gpc1466 (
      {stage3_50[6], stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10]},
      {stage3_51[0]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[0],stage4_52[1],stage4_51[2],stage4_50[3]}
   );
   gpc606_5 gpc1467 (
      {stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5], stage3_51[6]},
      {stage3_53[0], stage3_53[1], stage3_53[2], stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage4_55[0],stage4_54[1],stage4_53[1],stage4_52[2],stage4_51[3]}
   );
   gpc615_5 gpc1468 (
      {stage3_52[6], stage3_52[7], stage3_52[8], stage3_52[9], stage3_52[10]},
      {stage3_53[6]},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage4_56[0],stage4_55[1],stage4_54[2],stage4_53[2],stage4_52[3]}
   );
   gpc1343_5 gpc1469 (
      {stage3_55[0], stage3_55[1], stage3_55[2]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3]},
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[0]},
      {stage4_59[0],stage4_58[0],stage4_57[0],stage4_56[1],stage4_55[2]}
   );
   gpc1343_5 gpc1470 (
      {stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage3_56[4], stage3_56[5], stage3_56[6], stage3_56[7]},
      {stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_58[1]},
      {stage4_59[1],stage4_58[1],stage4_57[1],stage4_56[2],stage4_55[3]}
   );
   gpc623_5 gpc1471 (
      {stage3_57[6], stage3_57[7], 1'b0},
      {stage3_58[2], stage3_58[3]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[0],stage4_59[2],stage4_58[2],stage4_57[2]}
   );
   gpc606_5 gpc1472 (
      {stage3_59[6], stage3_59[7], stage3_59[8], stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {stage4_63[0],stage4_62[0],stage4_61[1],stage4_60[1],stage4_59[3]}
   );
   gpc117_4 gpc1473 (
      {stage3_60[0], stage3_60[1], stage3_60[2], stage3_60[3], stage3_60[4], stage3_60[5], 1'b0},
      {stage3_61[6]},
      {stage3_62[0]},
      {stage4_63[1],stage4_62[1],stage4_61[2],stage4_60[2]}
   );
   gpc2223_5 gpc1474 (
      {stage3_62[1], stage3_62[2], stage3_62[3]},
      {stage3_63[0], stage3_63[1]},
      {stage3_64[0], stage3_64[1]},
      {stage3_65[0], stage3_65[1]},
      {stage4_66[0],stage4_65[0],stage4_64[0],stage4_63[2],stage4_62[2]}
   );
   gpc606_5 gpc1475 (
      {stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5], stage3_63[6], stage3_63[7]},
      {stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5], stage3_65[6], 1'b0},
      {stage4_67[0],stage4_66[1],stage4_65[1],stage4_64[1],stage4_63[3]}
   );
   gpc606_5 gpc1476 (
      {stage3_64[2], stage3_64[3], stage3_64[4], 1'b0, 1'b0, 1'b0},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[1],stage4_66[2],stage4_65[2],stage4_64[2]}
   );
   gpc1_1 gpc1477 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc1478 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1479 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc1480 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc1481 (
      {stage3_4[12]},
      {stage4_4[3]}
   );
   gpc1_1 gpc1482 (
      {stage3_4[13]},
      {stage4_4[4]}
   );
   gpc1_1 gpc1483 (
      {stage3_4[14]},
      {stage4_4[5]}
   );
   gpc1_1 gpc1484 (
      {stage3_7[13]},
      {stage4_7[5]}
   );
   gpc1_1 gpc1485 (
      {stage3_12[3]},
      {stage4_12[2]}
   );
   gpc1_1 gpc1486 (
      {stage3_12[4]},
      {stage4_12[3]}
   );
   gpc1_1 gpc1487 (
      {stage3_15[3]},
      {stage4_15[2]}
   );
   gpc1_1 gpc1488 (
      {stage3_15[4]},
      {stage4_15[3]}
   );
   gpc1_1 gpc1489 (
      {stage3_15[5]},
      {stage4_15[4]}
   );
   gpc1_1 gpc1490 (
      {stage3_16[4]},
      {stage4_16[2]}
   );
   gpc1_1 gpc1491 (
      {stage3_16[5]},
      {stage4_16[3]}
   );
   gpc1_1 gpc1492 (
      {stage3_18[1]},
      {stage4_18[2]}
   );
   gpc1_1 gpc1493 (
      {stage3_18[2]},
      {stage4_18[3]}
   );
   gpc1_1 gpc1494 (
      {stage3_18[3]},
      {stage4_18[4]}
   );
   gpc1_1 gpc1495 (
      {stage3_18[4]},
      {stage4_18[5]}
   );
   gpc1_1 gpc1496 (
      {stage3_18[5]},
      {stage4_18[6]}
   );
   gpc1_1 gpc1497 (
      {stage3_19[7]},
      {stage4_19[2]}
   );
   gpc1_1 gpc1498 (
      {stage3_21[5]},
      {stage4_21[2]}
   );
   gpc1_1 gpc1499 (
      {stage3_21[6]},
      {stage4_21[3]}
   );
   gpc1_1 gpc1500 (
      {stage3_25[7]},
      {stage4_25[2]}
   );
   gpc1_1 gpc1501 (
      {stage3_26[5]},
      {stage4_26[3]}
   );
   gpc1_1 gpc1502 (
      {stage3_27[1]},
      {stage4_27[2]}
   );
   gpc1_1 gpc1503 (
      {stage3_27[2]},
      {stage4_27[3]}
   );
   gpc1_1 gpc1504 (
      {stage3_27[3]},
      {stage4_27[4]}
   );
   gpc1_1 gpc1505 (
      {stage3_27[4]},
      {stage4_27[5]}
   );
   gpc1_1 gpc1506 (
      {stage3_29[9]},
      {stage4_29[3]}
   );
   gpc1_1 gpc1507 (
      {stage3_29[10]},
      {stage4_29[4]}
   );
   gpc1_1 gpc1508 (
      {stage3_29[11]},
      {stage4_29[5]}
   );
   gpc1_1 gpc1509 (
      {stage3_35[3]},
      {stage4_35[3]}
   );
   gpc1_1 gpc1510 (
      {stage3_37[5]},
      {stage4_37[4]}
   );
   gpc1_1 gpc1511 (
      {stage3_37[6]},
      {stage4_37[5]}
   );
   gpc1_1 gpc1512 (
      {stage3_38[1]},
      {stage4_38[1]}
   );
   gpc1_1 gpc1513 (
      {stage3_38[2]},
      {stage4_38[2]}
   );
   gpc1_1 gpc1514 (
      {stage3_38[3]},
      {stage4_38[3]}
   );
   gpc1_1 gpc1515 (
      {stage3_38[4]},
      {stage4_38[4]}
   );
   gpc1_1 gpc1516 (
      {stage3_38[5]},
      {stage4_38[5]}
   );
   gpc1_1 gpc1517 (
      {stage3_38[6]},
      {stage4_38[6]}
   );
   gpc1_1 gpc1518 (
      {stage3_40[6]},
      {stage4_40[2]}
   );
   gpc1_1 gpc1519 (
      {stage3_43[7]},
      {stage4_43[3]}
   );
   gpc1_1 gpc1520 (
      {stage3_44[6]},
      {stage4_44[4]}
   );
   gpc1_1 gpc1521 (
      {stage3_44[7]},
      {stage4_44[5]}
   );
   gpc1_1 gpc1522 (
      {stage3_47[8]},
      {stage4_47[3]}
   );
   gpc1_1 gpc1523 (
      {stage3_51[7]},
      {stage4_51[4]}
   );
   gpc1_1 gpc1524 (
      {stage3_56[8]},
      {stage4_56[3]}
   );
   gpc1_1 gpc1525 (
      {stage3_56[9]},
      {stage4_56[4]}
   );
   gpc1_1 gpc1526 (
      {stage3_56[10]},
      {stage4_56[5]}
   );
   gpc1_1 gpc1527 (
      {stage3_59[12]},
      {stage4_59[4]}
   );
   gpc1_1 gpc1528 (
      {stage3_59[13]},
      {stage4_59[5]}
   );
   gpc1_1 gpc1529 (
      {stage3_61[7]},
      {stage4_61[3]}
   );
   gpc1_1 gpc1530 (
      {stage3_61[8]},
      {stage4_61[4]}
   );
   gpc1_1 gpc1531 (
      {stage3_61[9]},
      {stage4_61[5]}
   );
   gpc1_1 gpc1532 (
      {stage3_63[8]},
      {stage4_63[4]}
   );
   gpc1_1 gpc1533 (
      {stage3_63[9]},
      {stage4_63[5]}
   );
   gpc1_1 gpc1534 (
      {stage3_67[0]},
      {stage4_67[2]}
   );
   gpc207_4 gpc1535 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5], 1'b0},
      {stage4_6[0], stage4_6[1]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[0]}
   );
   gpc623_5 gpc1536 (
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[2], stage4_6[3]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[0],stage5_7[1],stage5_6[1],stage5_5[1]}
   );
   gpc135_4 gpc1537 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], 1'b0},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[1]}
   );
   gpc1343_5 gpc1538 (
      {stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3]},
      {stage4_12[0], stage4_12[1], stage4_12[2]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[0],stage5_12[0],stage5_11[1],stage5_10[1]}
   );
   gpc1343_5 gpc1539 (
      {stage4_14[0], stage4_14[1], stage4_14[2]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[1]}
   );
   gpc7_3 gpc1540 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage5_20[0],stage5_19[0],stage5_18[1]}
   );
   gpc1343_5 gpc1541 (
      {stage4_19[0], stage4_19[1], stage4_19[2]},
      {stage4_20[0], stage4_20[1], stage4_20[2], 1'b0},
      {stage4_21[0], stage4_21[1], stage4_21[2]},
      {stage4_22[0]},
      {stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[1]}
   );
   gpc23_3 gpc1542 (
      {stage4_23[0], stage4_23[1], stage4_23[2]},
      {stage4_24[0], stage4_24[1]},
      {stage5_25[0],stage5_24[0],stage5_23[1]}
   );
   gpc1343_5 gpc1543 (
      {stage4_24[2], 1'b0, 1'b0},
      {stage4_25[0], stage4_25[1], stage4_25[2], 1'b0},
      {stage4_26[0], stage4_26[1], stage4_26[2]},
      {stage4_27[0]},
      {stage5_28[0],stage5_27[0],stage5_26[0],stage5_25[1],stage5_24[1]}
   );
   gpc615_5 gpc1544 (
      {stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage4_28[0]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[1]}
   );
   gpc223_4 gpc1545 (
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[0], stage4_31[1]},
      {stage4_32[0], stage4_32[1]},
      {stage5_33[0],stage5_32[0],stage5_31[1],stage5_30[1]}
   );
   gpc606_5 gpc1546 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], 1'b0, 1'b0},
      {stage5_37[0],stage5_36[0],stage5_35[0],stage5_34[0],stage5_33[1]}
   );
   gpc3_2 gpc1547 (
      {stage4_34[0], stage4_34[1], stage4_34[2]},
      {stage5_35[1],stage5_34[1]}
   );
   gpc1163_5 gpc1548 (
      {stage4_36[0], stage4_36[1], stage4_36[2]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage4_38[0]},
      {stage4_39[0]},
      {stage5_40[0],stage5_39[0],stage5_38[0],stage5_37[1],stage5_36[1]}
   );
   gpc606_5 gpc1549 (
      {stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5], stage4_38[6]},
      {stage4_40[0], stage4_40[1], stage4_40[2], 1'b0, 1'b0, 1'b0},
      {stage5_42[0],stage5_41[0],stage5_40[1],stage5_39[1],stage5_38[1]}
   );
   gpc1343_5 gpc1550 (
      {stage4_41[0], stage4_41[1], stage4_41[2]},
      {stage4_42[0], stage4_42[1], stage4_42[2], 1'b0},
      {stage4_43[0], stage4_43[1], stage4_43[2]},
      {stage4_44[0]},
      {stage5_45[0],stage5_44[0],stage5_43[0],stage5_42[1],stage5_41[1]}
   );
   gpc135_4 gpc1551 (
      {stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage4_45[0], stage4_45[1], 1'b0},
      {stage4_46[0]},
      {stage5_47[0],stage5_46[0],stage5_45[1],stage5_44[1]}
   );
   gpc1343_5 gpc1552 (
      {stage4_46[1], stage4_46[2], 1'b0},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3]},
      {stage4_48[0], stage4_48[1], stage4_48[2]},
      {stage4_49[0]},
      {stage5_50[0],stage5_49[0],stage5_48[0],stage5_47[1],stage5_46[1]}
   );
   gpc1343_5 gpc1553 (
      {stage4_49[1], stage4_49[2], 1'b0},
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3]},
      {stage4_51[0], stage4_51[1], stage4_51[2]},
      {stage4_52[0]},
      {stage5_53[0],stage5_52[0],stage5_51[0],stage5_50[1],stage5_49[1]}
   );
   gpc1343_5 gpc1554 (
      {stage4_51[3], stage4_51[4], 1'b0},
      {stage4_52[1], stage4_52[2], stage4_52[3], 1'b0},
      {stage4_53[0], stage4_53[1], stage4_53[2]},
      {stage4_54[0]},
      {stage5_55[0],stage5_54[0],stage5_53[1],stage5_52[1],stage5_51[1]}
   );
   gpc1343_5 gpc1555 (
      {stage4_54[1], stage4_54[2], 1'b0},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3]},
      {stage4_56[0], stage4_56[1], stage4_56[2]},
      {stage4_57[0]},
      {stage5_58[0],stage5_57[0],stage5_56[0],stage5_55[1],stage5_54[1]}
   );
   gpc1343_5 gpc1556 (
      {stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage4_57[1], stage4_57[2], 1'b0, 1'b0},
      {stage4_58[0], stage4_58[1], stage4_58[2]},
      {stage4_59[0]},
      {stage5_60[0],stage5_59[0],stage5_58[1],stage5_57[1],stage5_56[1]}
   );
   gpc135_4 gpc1557 (
      {stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_60[0], stage4_60[1], stage4_60[2]},
      {stage4_61[0]},
      {stage5_62[0],stage5_61[0],stage5_60[1],stage5_59[1]}
   );
   gpc2135_5 gpc1558 (
      {stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2]},
      {stage4_63[0]},
      {stage4_64[0], stage4_64[1]},
      {stage5_65[0],stage5_64[0],stage5_63[0],stage5_62[1],stage5_61[1]}
   );
   gpc615_5 gpc1559 (
      {stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5]},
      {stage4_64[2]},
      {stage4_65[0], stage4_65[1], stage4_65[2], 1'b0, 1'b0, 1'b0},
      {stage5_67[0],stage5_66[0],stage5_65[1],stage5_64[1],stage5_63[1]}
   );
   gpc2135_5 gpc1560 (
      {stage4_66[0], stage4_66[1], stage4_66[2], 1'b0, 1'b0},
      {stage4_67[0], stage4_67[1], stage4_67[2]},
      {stage4_68[0]},
      {1'b0, 1'b0},
      {stage5_69[0],stage5_68[0],stage5_67[1],stage5_66[1]}
   );
   gpc1_1 gpc1561 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1562 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1563 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc1564 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1565 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc1566 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc1567 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc1568 (
      {stage4_12[3]},
      {stage5_12[1]}
   );
   gpc1_1 gpc1569 (
      {stage4_13[1]},
      {stage5_13[1]}
   );
   gpc1_1 gpc1570 (
      {stage4_15[4]},
      {stage5_15[1]}
   );
   gpc1_1 gpc1571 (
      {stage4_16[3]},
      {stage5_16[1]}
   );
   gpc1_1 gpc1572 (
      {stage4_17[1]},
      {stage5_17[1]}
   );
   gpc1_1 gpc1573 (
      {stage4_21[3]},
      {stage5_21[1]}
   );
   gpc1_1 gpc1574 (
      {stage4_22[1]},
      {stage5_22[1]}
   );
   gpc1_1 gpc1575 (
      {stage4_26[3]},
      {stage5_26[1]}
   );
   gpc1_1 gpc1576 (
      {stage4_32[2]},
      {stage5_32[1]}
   );
   gpc1_1 gpc1577 (
      {stage4_43[3]},
      {stage5_43[1]}
   );
   gpc1_1 gpc1578 (
      {stage4_48[3]},
      {stage5_48[1]}
   );
endmodule
module rowadder2_1_70(input [69:0] src0, input [69:0] src1, output [70:0] dst0);
    wire [69:0] gene;
    wire [69:0] prop;
    wire [71:0] out;
    wire [71:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_38_gene (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(gene[38])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_38_prop (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(prop[38])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_39_gene (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(gene[39])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_39_prop (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(prop[39])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_40_gene (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(gene[40])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_40_prop (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(prop[40])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_41_gene (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(gene[41])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_41_prop (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(prop[41])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_42_gene (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(gene[42])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_42_prop (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(prop[42])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_43_gene (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(gene[43])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_43_prop (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(prop[43])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_44_gene (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(gene[44])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_44_prop (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(prop[44])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_45_gene (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(gene[45])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_45_prop (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(prop[45])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_46_gene (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(gene[46])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_46_prop (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(prop[46])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_47_gene (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(gene[47])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_47_prop (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(prop[47])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_48_gene (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(gene[48])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_48_prop (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(prop[48])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_49_gene (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(gene[49])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_49_prop (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(prop[49])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_50_gene (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(gene[50])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_50_prop (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(prop[50])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_51_gene (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(gene[51])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_51_prop (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(prop[51])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_52_gene (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(gene[52])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_52_prop (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(prop[52])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_53_gene (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(gene[53])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_53_prop (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(prop[53])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_54_gene (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(gene[54])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_54_prop (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(prop[54])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_55_gene (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(gene[55])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_55_prop (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(prop[55])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_56_gene (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(gene[56])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_56_prop (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(prop[56])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_57_gene (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(gene[57])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_57_prop (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(prop[57])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_58_gene (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(gene[58])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_58_prop (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(prop[58])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_59_gene (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(gene[59])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_59_prop (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(prop[59])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_60_gene (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(gene[60])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_60_prop (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(prop[60])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_61_gene (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(gene[61])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_61_prop (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(prop[61])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_62_gene (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(gene[62])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_62_prop (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(prop[62])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_63_gene (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(gene[63])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_63_prop (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(prop[63])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_64_gene (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(gene[64])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_64_prop (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(prop[64])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_65_gene (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(gene[65])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_65_prop (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(prop[65])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_66_gene (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(gene[66])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_66_prop (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(prop[66])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_67_gene (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(gene[67])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_67_prop (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(prop[67])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_68_gene (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(gene[68])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_68_prop (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(prop[68])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_69_gene (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(gene[69])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_69_prop (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(prop[69])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI(gene[39:36]),
        .S(prop[39:36])
    );
    CARRY4 carry4_43_40 (
        .CO(carryout[43:40]),
        .O(out[43:40]),
        .CI(carryout[39]),
        .CYINIT(1'h0),
        .DI(gene[43:40]),
        .S(prop[43:40])
    );
    CARRY4 carry4_47_44 (
        .CO(carryout[47:44]),
        .O(out[47:44]),
        .CI(carryout[43]),
        .CYINIT(1'h0),
        .DI(gene[47:44]),
        .S(prop[47:44])
    );
    CARRY4 carry4_51_48 (
        .CO(carryout[51:48]),
        .O(out[51:48]),
        .CI(carryout[47]),
        .CYINIT(1'h0),
        .DI(gene[51:48]),
        .S(prop[51:48])
    );
    CARRY4 carry4_55_52 (
        .CO(carryout[55:52]),
        .O(out[55:52]),
        .CI(carryout[51]),
        .CYINIT(1'h0),
        .DI(gene[55:52]),
        .S(prop[55:52])
    );
    CARRY4 carry4_59_56 (
        .CO(carryout[59:56]),
        .O(out[59:56]),
        .CI(carryout[55]),
        .CYINIT(1'h0),
        .DI(gene[59:56]),
        .S(prop[59:56])
    );
    CARRY4 carry4_63_60 (
        .CO(carryout[63:60]),
        .O(out[63:60]),
        .CI(carryout[59]),
        .CYINIT(1'h0),
        .DI(gene[63:60]),
        .S(prop[63:60])
    );
    CARRY4 carry4_67_64 (
        .CO(carryout[67:64]),
        .O(out[67:64]),
        .CI(carryout[63]),
        .CYINIT(1'h0),
        .DI(gene[67:64]),
        .S(prop[67:64])
    );
    CARRY4 carry4_71_68 (
        .CO(carryout[71:68]),
        .O(out[71:68]),
        .CI(carryout[67]),
        .CYINIT(1'h0),
        .DI({2'h0, gene[69:68]}),
        .S({2'h0, prop[69:68]})
    );
    assign dst0 = {carryout[69], out[69:0]};
endmodule


module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    reg [53:0] src32;
    reg [53:0] src33;
    reg [53:0] src34;
    reg [53:0] src35;
    reg [53:0] src36;
    reg [53:0] src37;
    reg [53:0] src38;
    reg [53:0] src39;
    reg [53:0] src40;
    reg [53:0] src41;
    reg [53:0] src42;
    reg [53:0] src43;
    reg [53:0] src44;
    reg [53:0] src45;
    reg [53:0] src46;
    reg [53:0] src47;
    reg [53:0] src48;
    reg [53:0] src49;
    reg [53:0] src50;
    reg [53:0] src51;
    reg [53:0] src52;
    reg [53:0] src53;
    reg [53:0] src54;
    reg [53:0] src55;
    reg [53:0] src56;
    reg [53:0] src57;
    reg [53:0] src58;
    reg [53:0] src59;
    reg [53:0] src60;
    reg [53:0] src61;
    reg [53:0] src62;
    reg [53:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [69:0] srcsum;
    wire [69:0] dstsum;
    wire test;
    compressor2_1_54_64 compressor2_1_54_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9ff93e9e234da1e33d13352175cb3de1929d27f8f45951961a520693fff8c8ba7dbb7ad508b17c130bd497e2c69de8f747cfba8353ec17ffab6f27e23191e797d097921c3fcc2bdc0487c3739870adb0f30921ada3b480fe12fd723d431d86a4c8bbb7bf44144b86d2aa0c80e846457016e9fb8e921fdb4d24560a9bc748a524c86396dc3a444e7b662cefa547ed78c7bc1b8545baa05aa502875039031a431369636c7ab091cb94acc9679c71e23812867c39e7467adb59e11e3795a0550b482e90e717b165d2f397689c8d5efc38234485e39658fe6539d658af55f885c7d0147f79b362ebe76b578fcdc7fb3edb869c5547f2a4a106688bb27fb7225b07ef479525b6078f4c062080608b246fa93a4025878152c9d88cb7bbd734f23bfad474da35613c6b2201888f68041f5e2db4f9ad298742e14706f641e51e172e216fb0c67b83231876e6a728c50f1f9c4cd1393325333df18f507692e5faa5dc6d0a0fc9e653781904a3684634bf73b4336a4ea137b9e5fcde0e1b04847493f977423a6acb9a87c11c2500813b6e5e9b2ad793eb83a9e6bc946db44e4d83ce48b4da9a8a683d3bf950c87f0f55e14c2dc03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3462ed5584e6d7fa872b095d2f20b98059932a5a77d8d52c42ebf6b3fffe94a988445c8fbc9f21ff41b0aebb037cfe568643a804e12b1be6dad100cd7164f6fbdf9c064503b1c1eca04508b66722343582bac0489b6763e0f9bc5002d4406f1aa4cb5c491d8bb486254d1f64f4a283d9ba87ac20bb3d187fe9581c373785fd084b24f234f6da27b50ec621746a5c29e2728aedd1a248a45463a9c45860abd64c4038a1324d2866a0178a84cd837dc1c3f7349cbda13012513247996f2c3d8603426d90491ec7e478274e7162a29648cf26c772285f8ea65efa37ea96eadd998f4136e50ba7552720bbdedc0d50461738d6c49d69d21a6dec14e3f54da28bbbbeb032723b8d7b64d593fee6b3a80b7af887012416494bda295878f9732eb2183cd87f93b85b874e13ead0527d5a51a1b278f9737c3ed9011ef63b058c0797a8528221c8ddad922f7dd6cbed716e7f1cef6eec06f2eea3a145ee6fc8d1f167980c24f501475998c1d2bc607fe4b9dbca247f4ed3415f867dd5b7fadaaa4fbab0c912efdc466a329b99dc584f3bbe9b542c88a3c23221f387461f2b012495cbc7b69f2c13acd3821e9b540b060fd6316192;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h73cada2b90c9e261c2c228deab6fd820ac3c3676b52fcc0408f37e84a0233aa56ea52312d5da34e42a85da7f148039d0ad22430be47da01adf2e13ada30b1f139fb1cd221b04051e3ec9fe7ac91604474787fa89832dfe8a28690fc76b3f0e787b30ad783a4bca6f1440e2134cc385deaf8a4bd3eecea68e2f301b14e638909b76f444a6920588c8aabc045d2ae623f3035c0867936017157adae7298cd405ab74ce784f9660fccbf6b1edabd1d12b920a4a878b91e7ad3495d4c6e6d2951b375edf885fe33d9393a26cf67ba67e7ee915ce1cd3a729832bcf747273605ca97995f08a434ca3926e5ad24ddb3808a643a6626d2a05cf3ac45d780901e743e70e652df3adfc83cc50d9e82f9645ef508e50d49a87ef9fba3dfe30ff88ce68b3b7488e8fae5585b56085d812457659ce750675e5083534deecee32415fe6cdb7739b011c0957eea2dba68f50e35266b115213cbfd134b469fe39e56928e9bf221f7b2174cc724dec26801641a2d475db41d8b14ee87b8a3b71908f3ff1ff79cc6cea05e2521f7f917da1471440f1d0125afee1bf4f438d9cb78508004828e33ca73877eb3688a362c84cce85b848d26c81;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc4d152e6e0cb142bcafc73153761ec202d450124ad3fa00bb0ac90564544457c7a86dbeb41eb96f904c00d45ad640b11f4678f690a1cc4e001b51fd81d5862733f12bc28996593a5d56e51fccc27ea71eeb5776bdabfb1cd44bf95178407e97ca8dc8f39c6810013c18607813f869168fbdd5730fe39ee80c8e37185ce8659ccd1d42cfadc84d37235975da433c8ce6d30ed119c5ffb634c0951e245836966022274969013293668c820202d8089dfaa8d3c262ba793b0801a4aaf6b39ea60f605fb5287534b44063fbdeb056bfce5cf1cdbb735e49c42d69bbdafc987698fd5335042ecc0c9cfa2f9535c0f24cbdbe536ec5ce3f04d70dd8ad854ccc1a4ce7aa48c9aae496b106b8b2ba49bd112116c5a08ea5c65d2f0138e22437c148c13dca2905a40bff87093cecf6498079bb0cfc2ed27c73c175bb4edca1bb0ba06436359c3402b5f35814f80c2bfed787d810ccb7394699205e2f5addfab8a6791baf8d578b2210c7c224a76cbf2d726f7161017a630d69c3fcb48280fe2b9dd845b0ccb3b5947649d301bc0682e68b73e7384a380da8437300643525f54a650f60a48608bf35c3a0933460b7d2b376e6238a6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h7d5ca3f8462fab170cced99102f820d23773913c224aa84ee351851e5a2f685838c138340346039a7b6e30c01cf0ec05d1f11df53fdd3c9de1b6c82fd5dfb65e7e94c0d9042c9f2d10aff2e824830f5c5bcc8a8a87cb3090b47c188e0bc616027245807336b15503f632ceba1ee94d42821a5b1398a34ff1229b664633138829a666ae3af005d97ac04356009136af92188be34a60c4e71736c54c2d0a770e54de626e9931da4a0bfcd526b2dbe4edd1662a98e5cdaaa73b58ffc303569aae0149a7e6c0ad5e16c6605e2bf7481d69a8ac76ab34e02f967a33a965beab8be5267d22aba1991a52df9e0d317eb545e75dca2a4a699395f3af833ad70f22886a6aa5f0629d65d710bf4486ecd3a849336d96dd7178cb64db51b432f96066201662138cae69e5f70028cecdbffa30f8c921d667d385b2e61a8fe012e610d859cd54fe7dbdd30aedf5cec1fd4ec8bcc56b1ee5dcd7ce4fe1fbd4226f3e27f659a2a0913ba267f5642c6ba472ee72fbfe0244a8941908275540710787073997917b3c1887ec419109d651f60c43a91ebf25451c684b07ced6d50ba958da0514750584d2c0a629ae04e88d35c622af8f71829b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc99b4805872b0f96c8514a31deaf4302935edb5944173d76cd04bd62e23cadca62936ab0d3a0153e563badbd30116091f145c22069b27c7a6f7c5ec02df5f87a3430c5d60276a2243c45bc7833b286fa4893ac2baa4877b803246256c2aa2e46f5488904169c1ea00513598e008350bec3c3da8eb68fffa8d6a58cff7de4c012bc15a34fe8c56cd61431b3a0d5a576dbbaae326bb0975698f6fa5319e229a4f550baf796f4b5462573589ce202fac43e132f52a5e5c1172a5f0631565d71fc7c7529425a988f08a29d626b7849e7df9b197a844ca30d50cfaddef8e193255139cba8456088d002be0652b2cd16cb386c9fefac8d2a9e4123cb56c41ec7172e1f2bd0ad11b29aaee643a0c53b35dbcb3a58f7e0269958c44ded3f7d5794f266f9605e19a9d46956d9ef69c40e55c5bf7c4e8aed98de21000aa833dbdf7d1a6cd0891877fe79d2c109656c2e433d7bc3ed4f75ea047b67ede7a8510eac185946bcbf189cc0c94b69dd6d852cfef1637b199a708c6f5e8392eba61ebb7cab5dc372f1d337fc36a4812e4d1c71cda00b381e869ec8332021c05a0127704f70682d090ad564f23e2010c50a51d9ddf1ccb2b9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h606a2460d75284e075bbaf1268be3a5ec04d06ef6120e4e9a960356e56fafd89240927e726bc5bae8387dd78004531d804fee0f1e3fd5582d5d94b200ecd28cce486b8a1903fb6270278d76267826764525cc27b85f1a7798175bb0b60be18f52bd48a9d686b16f5250f87a6b3740340e2ac933f6741ab378b6ed2705841e091d1b7df9d2f16b7915ca75c05d700b5e5fe43edca3a97e400753241f77522d578c51d7964e30a76e17b193675d987faf64356e593e9e97636c3717d147e7dbfbd2c838deedffd862793fbcbf319822daaea140477b15eb2b2df6f4334ae000a45e03add78701769a1d97126a64161dd3e2f45db7976884ab5745e556b11005d2b89b16cff5da8ad59b6c58602744cc552879250954378df4377e0d01ecc258a8f06b9356ca23cb97f0bbf5bf17acb728982583c5680669d016cc823b3f0d5f7734761f79d86b46580f28a4b8d5d25f05898b6fe0ef9f864d9abea1581c8fcc3c45ec38cb18d1fb9b6f78b3f34a9e07541b27f0cb4cdad05985cce395ac63db46e30f1759bc5d8ecd6257e3d5fdabbd1aa1d063188f6d3b16ea8a891dc941214f78025ab7dc58c5e00ae27cfb36e5e434d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'haa43d0b043b49069294eff4282c8c4b9b24f6a76331147c2421456b20e6ffd5a1ae455501a963f803d681fb2e7700afeee69fc597b79133608e0c56225f15cce2eb55bb11311066334857332648f253cbd59fbdc2451df7c729296a144fd08fcce2c4dcfc2b0824909f2f42b508749fe890ff87d5d328f33675112f3ed74c0f7fffc844dc682e93c417265ff759594933693a23eccfb0943fcda175867c427f3d74fa75ff092f58874082557c53af5397d62752d69168482681e8af2670fc904f3cd91aa26e7b1a841106b88cb5e1c8c3f8d7c67b852dc88cd0605e5e0a4fb01726c4fffe84dfda9a4373f6f39c50cdbf18be339e45103176092d7ad81c7ee8c138fb2601ddea2d00eda5a21dd3022c67fa0a8c5f5c0582b5c51f356a5c56bab10f0caf9e2aa745fecd52a00fe1244ba6bb790049dad4a736c265960621574ce51d310c78553460d04522c300b7beafa9cf30440c009207aadf8797101345ed8bdd4b2d6a98594d4040e36b8437e9a53a5dfba64efb3882f6a5492e1008656e4addefa6e2f860a2340c30522751138d8e36ce8da374d0ff960b7dd07396c24730e3f664d68b0fa01e442e2a3b1a9ebb5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hbfea4c9a01c943ab393c9d0ef72485ad18016bc16f9c5cf53d9a8c2d37fb3525828b9d4e58b145464ebf7467c8d7dcf299747eca2bffcfeabf8f2588385f0146f81770b8f84744570cb9d51675661e40a36b9f61bb87f83ccdbe1066e3952b1676773da4f193dd5b8f57b7024cbf6124326c734ea79e642fe0092f372e3bb6a75303814cfb10f5113861ff274269547de847ebe33dff04b06959278a76a039f0fb274f1f5953cbee0f70f3804ae1d3ebb4dfb96a76789b5c41a6ce300d6763f27d2bb72b4d6bb0e04555d594cd77cbf4f7eb9f166d6e219700cb948875de04fdf12e0bb37a1cacf58e698236bb11a826b12213a4c18859f0dba3b8df2ba47d703eb63f9963eeda901a800fb48b4e0eaabfc356410c49b762e7aca0496180d5bcf538124bef40bc9ce7ed56a9a181f75f4f0374b0b3ab26df79e99c6ebaea70cde0c8a409eab0102899c63186dca4590a3282afe51f70e46b7470a261bb48e94a07179c1f39d7321402ded85529ae4274022f6f9713227e38c03a752b534a0467f15fc2012226909b00a45c57d3eaf0b93864363d9a048183e3b308298bc1ee9174ebc781bcf0b2f07e0a558624296603;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h71eef08b825579e518daa0e96e078b1df4eca2e79b664d4adbb513338ddcf4ad93677596ed965a21a6c95f452de3a946df5f633830c1d1c41799828b006278f2e8eb9aba7f0c6819d836d226d02f08902f6ddc7071ef53cc1c61d82145f35e40b70882e2fbd86983eeadf88bf38f08793dd8a068a07ffb9797561ab012a88c0d40cc50f3516d60780945dbefd6e00e1ffce45a8f259b6dbafd0438db892a0f5f2accfa358c26dc63ed75863b9738829b6128d2c4de21288db83064aeef2dcb77b2089fdf0e96e393a143fd4df0784b28b09c67cbbb189b7f0df4c688eb2fa1863840ba6f5d5411dbd461d49be0c54a5bda7e9994edb1f79b77d8ba8ffc10ad6e21d8a68479a5f6fcf25b37464679991eefd9701d3bca1b53ea35257b25eff4e854289faa70d1b721d4cf116df3b7d12340863c5d26616d8e466014bc128fa1dc366a393d0f63850422fe8e41565dec2982e05094031e04175da0300fd4dc705da0ac5ce2495b234cd00562fe6572e834c2146c9fe21f1c94c6cc5a375ec6b02eb65052bdfe76acb2fe9624ada3be79521d6d3514f5223edd0ee2613cec91a97f13904d8b2bf5a3af27c00bd86e732bbf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb4848df26cab1bd13ee4a7a29b020862458be18537f73244319e8f4216080b02ca644b725b82e479383df28da089256d7265c165ba37b351c50a3ad493f19bb1836b29c0e527b366105c90483925cc70d2add71f26b66969d61ea17bb07f7c93e3a449095dce0bce3b1889c54a440acd76181d99bd8955a7896c5fb1c4548ad423f4e513bf04fd9efdf289b00d9d59507970097247234778d73131a271be63c713b4eab7ea2f53b0a6aa2df6954cc94f5e0157aab62a89b7d85c023fbddc34d41f7f0f0972112c2bfee2b3c609b84fc52ef39664c25dc01842b1bbb831e57f621d021f1b8da0494621f185aa415b05b1cfcdbb6ffab7777fe89ddcc4354c72018cbbb0ac6088f3493ca8fea4fe82d873e04da5934105c4ae0fe09512530aab1f5d5ec803ee7a12928e62d15691d921201898645ba352922c0a3276b1b3c989fdacabce2780ce4c634620289a5328e966be4034c899674b29fe8ecc6a71984a05138d501bf0d151b2bd6c43fcfc4767a70a85a1f02f96d04fde76821c05abdfefae7be85db32a30a14c3168ea2810dca782eef7eb44115c16e7ee4e7fb2f05ab0f77b4c9cbadbe8b13a841aafc022bf0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hbdcbff480a2219c8d4c141127b51ce90649b944de7a530d0341248cadbf9238ffcbc588c56972f02d8cd7e8a35858e38d707de47bb0212912c870aec8ccdea7fa880830184ee6255f2d17fe6c11400dcd514ac59fd53f107a0801799e4f125a275b7b3bd4bced37e5fe3c3c6ca5eabffcb6a2a1a644e0598eb9d9e5194bf8e4705fd5b19f69b1378109c0074842fdffb8b92085182756aeb09e5f118967263f85e9af944671e99acfc8be740d549376beae7f1ce8e2717074462133ac6e2ec79ca682cdb2c74e1b229a35b1799c2bb38694115253fad1311ee2cff0c9a3b7dd14c89a9bf55146e56231d923dfe06af5bed4e19e90b5ae5bcd9295bba5472676902ac3c83a442153f130cba5038377a784a97b00fcb8c9540e0361db9098e287488df126aee84c8364f01e3e054c733b9b6404ec8cbcd133ec875a2f9289c3c8243686864a649678efb2bb83ec0a90757ff616cc0741143c48c9604fdd5519e1dd753ce81ebcb575fa9256fe57fe91e2f3098e745e49ca2a270155299b62f0d4df951afae35ceafe04b6438e2780c4ed7901bf3222f8648308afa6999d6adb82655f7015d5b5fc266d61c57ac6900e82f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he1eba7506a68057754b7f5cdb02a97140010322b4a6cd86bbc1c15b3a925914b84ce98b59ac685253fc42f828d4dd4a941cc9b4b0ff148d35cc2bbf787e3681320648c11c8074169d11f05c18a3927e7d8e3402cdfc8d3f86a2c6f30a0b18d6e428686d6a7c215737528500e003b95b5e05f6b7e692b93368d4a66278d7ca4ddc0f3a964be6348c2980703cfe9ac4b6694af472b036dfa9fa46ff62a1a0861db0c0d314eb49b380198ff7fef6f416320d2e508aaf3a357a58589321a9fa6168ff84beb6e3fbe6f7b12bcf956e21c5970e452ddec82949fef39ad51434b81703d536fc790743220be9dbadd5faa2b15b1f559043985794153fb83da85890e5e91ea2066952deefe70cd6cdac5e37971edb5b02cef8af5c96cc68e8ad202bc67a69d5a75e2bc545b2daafe8f7ec3a4986b51685e5fdc14aa037557ec67021028bc39847e022ebab537466f491b18941eb46d5699050148fe41ba5be60039917347541792f1a081b536e015061efbf676944291077fe4ba90a27286f5e08d0e8cfc23a89f83d858ac24531bb39de18b19232b1f3bafda8d35456100750275afb1b721dd80fceaf885697d0df47d7c9fd4e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc02a4042c5264a18cea1ca99b76e22ab74e6ce9bfb3528275928b36ff1a1c78703abdaf029973e7dc124d66b632cff50b8a5b4b008a7b858ceea94101deeb0176275c1fad45d03a405f2041f71a62afd9959babd5934bd907959bf369724dd3219356e7569c230b7c1985f756e09557c16964701a0620985137b0fbb9750f51db282ac18b7b827c741e8a0d445b30ae0ac1d3f1efa99b3e13721970f5576ad79321fe41c7103b7f8f943e80f24310b93e564cd459dfa751c98d4e8acf52bdd78a8bbd7bd3a8ddea90f3d356d8710d8586f2e9d1368646a99aa55a32bfc6945a35a8fdb8d9afb121e83eaaf8e7f49b60ed03b7e78fe7616cd051f3bc5dcd025530c3eaea6f25daa5e04939388564fcdde90f278f251c8a764cb61e7f6e5f99440eb2ba839ebe940be55902a02d5659db9358f150c46902a72ad0370d107fcfdfd157ecca3062947f1e2620edfccde0671c004fd69bbc970eabd1025030bc6a2821d850df26d2fee62f8004da90c53db6b0e6de69d443f64ad4e9f5283b00cb13cd4acedbf0c8525a7fa27401d9bd6fff1d74ad121013724da7c3e3f4a59dcc46b465d19b9c97931daefad1628e92f3a23;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf074e91eeeda696f79b193b4cc6d36caac738928b9a9716a5012bf31a90acb927d7f6a99cc4946ba15afae655729444167dcebe066d1f390e2d14d9ab29b64481b97c403800d816aeb6bac6baacc20cef84c1a3256ab1ac9621b7511954148cc152d715a95bf238619671258005a507aadbaa5d06181bfa0786fbd42ba14e38956ea4e1992e639a80e2fe16276dd87b55e4d5d64a5a7cc078da8f44af9abc5e5d94c9314ea727c0debc2b7baddbf73486a337642255699d3d1044b292b31a8390b92353e83ac8dbb63c0d1b6a01f43a84a1bd38d6039062f9e02412a4e9afb9af196727265e095720f739d3f72daac99cb6c0be10b55138f509bebb39acbc9a8aee123780a493e0fdab3edcd824b9383136ffb9b81819afe233a9cff5c332457ab8e8185a140773a7c79b5a72e2a3e2c727be372445b3ba18a0cb6e39f40c763263d1e294b0ae4644540e31ef633ceaa1cffaadb756c2c458390d6809358db5ab084f0e7f0734f10362cb997a41c6d84956a357029e9af902573ae0b78dd579c3ca8c0e0f4e1c8a92e7d0a922468bb2af2c0f0e616455edb7b9dc9a7c4615d74b7d1fc7e3342355d580a7f2a35b08ad3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hbc9171c36120b2216ee65f135c7a0bbfbbdb02f086c557bd792a60ee03fc4fcbef634ca67e7fb3eeeaa44b57291e9dc6c0a3cad5993a3581c87b93b1e03201eadfbeaf1dbc43c826dfb32bff11aa79b9b0f567ef1831a4f56716bfc14fca5b04658ff739868c125454a383df7f5029e1d5cd0f9a6be2088a2b4b04f4d9a6b78eb96684e01d57c61ecb3117569d9e228a4695e56a7e9f3e83335d50efac5473fab0d26159c5d3323c78152db1d72065f5d8a99fa192f28bba41cb74655e46c6359f3ddff75ee374f0f05b4cbe232b5aab3ffb511860dd862afb3dffda3ec817251e8c976d63b5dc72873fe22029199dbd900fba71f1e2b2bcf32003a52720cea6b8bf7d526b059244cd28c0310c6f85c705cd1ba79b00f0457f4cd57a1466a861dfb8d4770f612acc9ee04c41622497fb9c511c2f9527bda89079c1e32b18e85261919177b95574fac370af48f8554b4f9347aa9e79bb49f4d0cc18783ced9b425e9bdfe469de4eddb5f0dce6371bffc62837dc424c24cb7810cea5fbda2c8caf9ab56cdc4f4e961a0e50fb1c7476e571cd793f8a498d819bece708962b8d0e5f633a239982b2824ecca3a003d1df6b75;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h85e968135e2bc205988ebb1fc51b89e50131c08bcbe0d9bcd73496de446578f317d6907fbf7cd59748ff4c824aec7107039b7e11d04a5d3387992a30e2454b984369ffa124163e5bec0322264c16fa3110353987933faa14fdf249808d9cef4f15ffec455a6b4d3444b806bbd8c09c051a84f0a731b74379a3fd107aa9415466593225f43d5722188aa98ddcc74c757fb3263d9f7e243f85c5105b0370411a5532abb1bc66d9f7538aa500ec41d9db581dc752d75d2f31919757e7498c41ecff88e1108180c1ec538d6b9fbdea8d629e5e65a7d190a4a2df8557fb5fa5d6d065e294ad05d5201f3affa21e16ef3482ff20e9cd5e310ac063fa8787c6677bdd5a71c9ccf458a7fd8346f3740b2e1aba427cb104ed8afe5b09580f74aca732641aa5ff33a90a7641390f05686368799e1ebfd9b4ca3315ab63a1054e3d72a7bd33e40fc6b2ab62bdbc03d69c08bfbabf2246ef2ae2ba692dde0bc79a5a11240a1f2b6935664baf42be7bf9814fd891ae061c05f6ba1eb32954c35dd06d6fecf5250c3bcd1fcb2c11166dd27de45f0e7c278d865134c4568294b5a2e8f095cea74d5af75fe231d880f3d8f047fa0683a108;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3cee733d283f615d281d1a6b7ccd5ce0e4a5b7ddbd97095c6c7050304e46dd71366c4412ca5fb938f3a1907a4369951d883b7cbaf638d2c3e6b8911c443e8c5abb732d11a4278f2efd74fd078cbb825feb1c3a5622ddf7ee56c2847a671850c78fc81114fd35d4265b5e7f7fe3cef2c45c14782fc41abbb540079c5d015f651e57ce5f53a06b8b7672111701571abd1c0d8fcad9fbf9b4727852bece7681d95c42a4eded4bb919d77ee97ad6cc3871ade23047e97598e7267801d168f94aeea67e6899d5bb16975b32e8704212e14c7f94e87e19453373d8557b67c417ac3bc31a078aa714aaa518b50c316037b0ca231e0b51c071fdff6d7a491e8769f240f094a721697545077f36466e25f2d47c8b47103e466a35f69a1900b1c6cfd79f227d4afc21723c5df47928ef9f535730dd0701b2a24fb05cab9c8c4fc39f8f80e1e4e88515538183e25c9cfce97dab6b002736c9fcde24ea57f82635317c962f0acc8b04bb7002fe32955aa99d402c712d4438c25e729a92c8d9b40222e638c9040903aecf21e4ae4d8dcc745e2afbdc5f98623a59d08c10a4712a0a8de53ce927989c283108bdce55c625a385fc1e6b20;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc471e883dac233f25d99a5bb19e8df54e97668fe615800f75445f2ffc51fbacc31d6c860b2442544dab2c83e062b2cd4f3e69cae87bc92a400f29ce13a6c96085d715a5c5242912d53d0c9a660ef1cd0e53d523ab480212db3483a30f3b68b68a49531e9563ab13dffb21f73fe85ab9dd5f1162d53c7ba347bce6cf676a9b54f5b142e4011a7cbc946797c461cdbb8ada0b3fcd6d4f32966255365a69292c09493bdaf59bda422adf4c0e9bbed05e8f04867ef1c589b1d9a6c473b8330ed50b67213432884b28400b2ba573223bee39e5f807eccb4f3322c20fd894dd45e0052244ec59d9f6e9726ad1c320e73ccf89efb0b25bddc528498fc780eae30c2dfe231188177fd0464eed8a35a1dfb4dfd6ef8090d978111f3412b8e9b697d3e4ac1f67b9d0a9489bb7931e7a0d759369641b37e8c44a1df2100be2d9adb9daafcd5d80146b8713d3e6ce0a09e160855babd120d344f20a61256abbb6d445b888aeeed88d1eb933709dcb59c2dfc6db9486fbea64cb96bbfa6091773d6944a6ff81891f837e7e8662c900b8fa4133683a8fb163c4cdfdbd6168614437a6af7a4216926e65a2864bdbae6ea5f4d296fd59a9d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h804aa8a336578b855fdde089cc9adc735ea2ee8979dd1c8e377a6a1d359beb3642b2edec3878665acd21d5e77df49a18e7aaed6650a021a7c2527d6b809af5b10ad6694131485f0277e6680fd9ebd314fd58d59cfd44ab4396d54aff6b6debe8f0f91504d70f5e5814668a0a7d8944228e89e7e9300f6fec507df7e04a123730813d4b5d29594e82f73ef0b2a14c136d939f8bcc49e01e477724205275bd9fb8c684371a1b911dc3eb4c6e4b4d09976918f569f4abbf75036307871852eb5e573a79196923045ddd18c1d7b76454907af0311b51b53ac0a401c10596a47c96996e2ded6a85ce10f006aad4f141906a37143a35f54007ac856cf748f0c80689b737ce526901eeef9f66ef262a6540b65655adb70a4b8284f77a5e868436d5d4074bd7cdac13d8ff625d6f90417a8bb3db2060b558378230fdc0fe6f3ef7f955a7c91362120691981c281167e09d26fb584402b48a338650ae68e1c8b3468d9d793d4b510cc0303c7f120e8b7d6a2f266991bff9d79edf0fe7138983e2d02e13b0821d84b1700a0486df765628e8b5eb5ee079bcd70789d9a1594f3e1b737686745c5feed6cda5cc4cbb0bc3f4ff67a286;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf2d39b5f67aa867ce22d730464617eb48dd8c3033c213ffa901a803080db68dd526355b0ab9a305667f33a80a1f00b2ae872b58960fd1f05d3e837623f72bc6ce9d84218e79c8edead367c39844246ef7b8aa76fb4ea13cddf70461a6c20ef44966539bce4eccd3520f8b383bb5cbd2f4ae24781871d60280bf0aa313e11e7c8cf0653711553db0a849af4870a4968146f777f2e9b71101c930c12d4dce85be093a4bef41b1aed6c46b1f15d87d97dad85876656d396f9c991bc74595747a9a6972dfe644313a344e2786393638807bd85465fe182524326725f03f7e8be81facf272c5d683fa0815ef0e25bd1cd82d214b316d96fe004e16e2c5736234ef15b32c2028e959caacdeb58e16c16654ea57711cd21e2952fe952fbfab6d07cce1814c323fe9d00a0edce5f5b28ba845f21103408714393c0858522bc9681bfefb36349012e5611854b98333134402f30a1f279bf7fe157bb9e166ce6933878b1291fe1f6fea0c936f5db4304b6e84275b0902ba752cdc02afc1b452066f8ab6c0cbfab9c680338a744a1775f5bf0617f779faeb941bf0a95ff9e16b293fa6389ecfea5f0afb666a7e98093de7b221e0e32;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc2115824922bc22e5132cb384ee00a576c0aabeb231342476842019d74c77e380bae8ff4143a87535b1e61fca823193639c7cb97f560d85af3b981ecff83069f6571a1727023ae5a5686281cdf98b7dededaaf453470de1644abb3d99bea25d12393fd07066d38b435771cb061a72982dd7a65acacaa7342010e9361159893feabc0045ceb2bafd1ae7bf26350b185a0addb48df7c7d1557ee7a71a99404f75fa3a42c402f249f10295c0bcc4939361977a4951d2f36edabac2f4d4f13c6e0aef7f9b50e1b64ea5e9ede12f2295049325993d94da58f2271d743d185cf7254e8cd3214a125e30d9a4c5a50299e07230753bf2bfe790bc3ebde7fccf358e5a761969083b3cbce2c6d56c14baed53c0d5918761545a5809c9d6a59e76f3b1481164e6f812aebee7f34121cb25f6b6c08dfb0ee7f9fbb370a7f039906b89a2b1b4fd0537e55f51214c22b022633fb5b4c74dcd0cce0b72b0ac126c03f7462fc84d657b8271cde2ab50dfd4596a0fa65959cffa16e346cf15b31b476d2589cdd7dfac63aaf83cd188892235f16611e08702b7a222737b28ea4018f859a141faaad2d5d97dd60c2e0f56c14080882676fe884;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h577742ffdd086fbc0c9de33cc2e3357147571240543ddd274cfc9331352281646a579ed7450099a3bd1f850c736e3809e64bc849d09fba04a7d6905ee889b0d515b648772d5dd772d5ad29b86c437350cebd263dcbf111e32794f0fbfa46cedee01d3047df55156e7bce6b4edf189fdedf5c9945319cf3d38832c41583927a312f26b55bc1a600bc4420ef89b765e857d9cda1a56acf236ccb516a3e47cfa4de5f17da1aa235043f7572cf58ce2dfe28d92a270c1f838679be577d793f850dbb8486c756e15c0dd293449b212c6efcc5a299f7b483ae92e43dccd50db32ef8c70f56b385aeba652e248604cb9e8b7226ca7f7e556faaa335ceb88c12dad76d152db8b40e72c988fa8bb47163a8360259f4b7b2ff3bdde32bdeaeddca9cbe0520945511c68c46e3da486e2f1dd541d59613ccd927bf433c8fa53f8394c1e273d43fa4e1e752ed24c565fec815593381811134191977d33501649a9e08911e5080e4d47e2642e1f8740771702c0edeeeb20ff735dac53b76ec8d18400c1031c4963d7ce5de2b75d349494a0b93b5743fd81c92c242f75805669ed47879bde223b00f2641993c325b15909d7745a3154378;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h88234c2f991b49c813576dcb5ed7270a0fb33b1ae59269b151ce6009359239719ce0d5fde6f0aff22e45dd52ddacfb26c6c73af6e668932f897b277aaee8db7b6058388254624b746f5a2936ef1a76be94b7884a3bd0a86ea7963d62129e426b5368352a63b08d11f5481fe31e7175e559c3386701d1ec358633a85956909bdcc9d0d13578b2b1a6f167bde1886c154657eef60cd987cca51ebcca38880043895f74a2f705a332347ce98b3e2c1542be5aad2c023a9af3f2b17f83ddc878fd09d44b0ef85e39d337cb3ff888f7a2e4193f899b34d19664c06e4f26a4f74172e1be2a180b6365f5657d0fad4dac9fd2a5ba841d17d1b1ff8969ec8c9892c3c4ed7a1e51101139b2c1cac7c7ff113d372ca774b401b2a2d92d1d2c41e8d8e97abab7f0c79971ef3b0f2eee1401b05840f8b4a175e8fa8017f97f971ba569cdac6b2d68983929256aa916265ba9cea317b14f82d6d16b74330ccdcaabcd0a539d488001fefb79f7770822842523d36dfe49b5bd0dfc55d08287944a2d01e4341438ff1d43a6a1b1fb3832ff8d4c8e8ce26975e9a0abc73643fd6bb51ada047f43b56c0f364d9796d6e570f6209ce99056d8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9ac139e755dc1fc6378f2e8692b4201d8f632281204a6848734f0ee6ba3e4bcc87ab24c5601e3a191ec40ed1a8572d2347744fd3dd6d8e2c9102e703935c4d8b9d142b09aa6d49bb5a6bf92ffbd3126c62d0deca558dcdb397f4a82476ddc19973b63a9bcf10afb7c27acce15b92f336ec45ac7ce78ace3bef74299ce16a23789cf3f847afa40effc0a6b746dff710ea04e6c9e8fab90ad98b26b024f746cf8214c1e1e16ffc68c6b0bb2a16d3bcdba4d2785ddc9bbfec34a72d568e9b45c43f31f6ced481a8ec91b7adaeec06a298417f2cc9d16e825925eb4bde5492e167fa68f87a21c02cb1ab95ae20e5d2d1641286ef892e75b1e7d979f4de74972adb35a7e88012a499d3b448800849d0dfd63fa3328dc340d9e5039400d1f930bc382aa892eaf1359b489f769819d7690c35f4dc5a3536eafb0506df9872dc2b4f9703226aff5e2b810dd12fff3044445a3fa66ac60636eade57590a35443161b0330b0f55da9253724fca42a9333332febc5e4a48b29ca013f37948a22102c9425ce027d8bc558ce381ac8620752cc3e2553c7f7ca26130a51eee32c8baf6045c14bbc9f7e2d60bc95f631e5ff4a38513c1dd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc247b5a8f97dcb41115d4a7de6d847623a989ed669ecceb67a1b30d39ff9e092b1b1b8ecb4a91ab6197647e965f2928057932b5dbca2e78dde670ada0f02e6a1a23259fb43cff2688c37a210ff93ff6342e10ce04fb4c67d7b81ba50c5666dce89c147781d90066c951abf24cab1d6f716032c868a5ab77a672c4cfd0856779214cebf837f41d9baf0fe0dfabec22c9249cfa9c3b2b50ce9bfd2f60acfb43d77e70a698cc851387a785a3f784eae0e33bcfb25984d9185a60c73110c6de829d500c1a1f7b9f9fe50f273860f451a23e6876463c897d28fde0db0c4a64fd5868d989bcca53e570a5e9eea4aaf039780422293da20e3b2becce6b4df8b04aa8de3bff115e7eaa62745e84341493dca6a9089102c86dac8c7b3a729d285b9ac9d0fcd3be6478ce9dd989bb43df00d0f58f369fd977abb2a74ba7f76e1a58bb3e8c190ab2fed5f09a1fe59c44af65e170d1c1e17c82933a6302fbbbd4aefa4fb0c5547f48315f31edc4ffc00c2ebfd7ce4ef2b29330fda55d24ecadb60168e77b33dea5682c2b9492393230b2e04a404f788849a3f674b025a1ea5cd9a667c7dfd647142511cbb47b8fde820aa2df1c52790;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8ae42519d570526676632a865ced25e6b2c6de6a8fd90409101120772c8299e4023c1fd57b4347bcdc7f70b9dc8fd8bb04c6a5482a776e837b254d7bb404d3fdc79327d5554b59cf57ebff784747c2a0579a719ce1c482046711ebeda8f0630653128d9d0e70303558ae2d33052082db857e048c35412524d6cffd264863499c7a9a0e4a99c36a02ea487016384cba1dc4d1a7a7017736aea08607f66a8d5142fc803581a344d18e1c0fd9c648086d9fa1d0ca15d12eb7f4436516f2a5f144b46a1f160a1ac36b6de6d02d629c3408456dc21ad7c7d953b0761c7faa99f659e9c46bcc01f31fcd28d0ad9f9316a009b4a13ca23d1c12647e5779056def521900d0d493e08991d43fe2f8de04a907937719332bfd29eb274e5c7e50bf385844e5713beeecb4078dd1e9f86efcacd9bd285deb67b6ff7b6acb27666361bdd3aca324d09f04f2acd9541ccf4f2a08881d788df59c01710c20b5ff7327f33fd634836197469ef6e46f97d696c7c1ada4015cc7ac603f114f99f361a5281eb1436031daccd32e12c2308ff64f9d37a69503997c0f49459399a5be388167caf06419fdbcfcff9636c2c64675f1f1fd27fcc1c4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h5a0334ab3530aca103c3ca8ab6812faab9ace7adc184b6002b765717e9b91f83d51a092b08066c24bf106597f4d0beafea01eef29018158ca050b06e59dddf3cbd7545afa339602b40f18ee47e11ce0bf88a8797c7d5a8bc6804cb5b78ed07d5e0adc5f5d1e4ee4dd713f2899344dcde24f78291686a735e4aa8c6ea751d183c37c607c384c0644cdf424e1e49318876f0efa9ba4fa1930e961e7c38cb5927d5a2e969f64f7922e32d258b48cad7925c5b20b36a5d6ee9c92f39012d147fa463729fb59f1ce858e6f95a3a6d1eef90c4196163f050cb097e7bdd7058af74f411f5dcb4e27764837aa682183b48159e8905852acfb3b126339210033b74ad9a331714da860553b0f261937de74c8b1978cc76f5ba1fdc0f4ab8419c42e2d543aa78a4cb3d74e1c4096161d9e14c884c6d602ff01a473142a14ca00bb5d3e51588d601060612cdb0ccedc1215a73c1917cdffc25345e1e614a0ab361ddad3750920e5db37204f37ca2d7c674a4df25d3a5f667a68780cffa152a40e31c8fc2745de19b0e5091867ee0db023a7c4748a5092a332a3c21bfaca969ac11c2b070652c595489f9bfc31e051b9c6209ca3a81d5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3d65d31151a88bc79ab1d6007578e1bad5b5638bc180e59fdbf3fc23e34220014e0559a4d2998d11fc485ca2e9d2c6b518ccb75cb0e7c3cc806abc1caa7821487daab161b39cf1e2170d6205b2400d0a21dd06ddb6a4821d664a77346a84a5091687a061e25f71b74dab825ec6aafc61266a64c22e573c497f9e706eb01ea841c5d93998786f0da2ec82d0e4d350ddd584f4d01d191e895de84251e7ce438783b230d80550ffb4f320ddddfd6d176fce3cabaf05001861796bdcd3570e2964963d69918fb86b44f5ab3b52f10f4aceab57b056d841e9f6a92c4d5ed5c56b71a75cd1d455fff90de363e0c59ed5d4ef9d88798fc25ff1dda4c51d892ef15329ea2ee57af31cc3ed5828dd9f864a12d7b5a1e7e177f86d1a9769c87e4c1ede08d2c322428311e3aac12089e89094c814ca900e54f8fb3c1ee7a6ec4400c009d147629830791f751a1aa4a1205f2929ef297b0a57ff2fec7cb76cb71c67631f0f145a2812ea374c3743fc575bff156ba143054a284a8c5eda1f9ccc71ed0e6981811dde493c15072ece4d1d9e141630f654d5825d70f237a5a76c5ab6bd542c28d8dd836aa624ddf1079dd845fd85d91e5b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8c8b52eaba64d7f15b5641e7f4c63bada6460d5d24d874a9314fe8de667ca6b6919e38d5aedff324c88b3de5d9f60688f96a3ea8fead7ad04f631fa5ec6b3893b2aecc506d4365de2958115fc4e7e1b3b897d9db6f06239ba01bbdfa9c603b88b9cbafbd4d30f0cf0cd2521595757c530e57697739ff599e8d053fb3be2f482829ec3ad294d337a1604773262dad9c117d690b53e2f869a870c4e99cd48f77a64b9a80a24bc30152677df8860bfd45b159fa880734674bb24079ed6078015edb7d22cb36c26b57f0eeaf3e3339202b711097208318e2955c065ce21e599887e02072636cda55eb001f64d07818ce5a1cc5ef9f8318bb25f5a1ad0175f0987598c0e8107df50c1fbcfac83eb29a4bc36e012abe5f1376d93015c73989ccc43dd7bcdd73b228bc5bc1c245b7c4e5b2bd9db8d62aba61def89be582800538e2488f6438a4818cefe6eba9d06a9371e09e6f43c7bb51880759ec8b40784ad0f0e8db514df7d497884c9cc1a3bad07bcdce46316472b6cac9c66a41a773dbbe409f11a4a57d4b466af01e2b9b5586502a1a987d16d65e3503ce835993a4de9d22b655bea8800eff67467c32727a342cc0317c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9ea504315dc4e41d7727e12b3571f42aadf57c6cebdf0c4e3209218b567a9d5babecf2eb6b79b480e5e5b9b50d1138b3bbc474c654a62e2c6ddad9b51b64f8c9f3425c9962421614d264a2b66e845fd9bd7aea232e796b1e8987622005778f2ba9f401bf87f40003a3a4924fbcd6ecdc484ccaa741423319d2599d80fcee7ea728034d8ef2b9212577e827a5c482c709b1389dabf9d055099596a76e554d394eefd1d21216291ece4634709819d13ef91a983e607e65a4d085ba3ea6477fd80c3eb8d3ef6f3cddd91819acab70e15c06d56da433d3e777d8a00810406547df19aeca37c678d6cfccbb8afe9b20767a6987c45297e08d1f3e251fd6775a08203e57eed495e01695c6c73867f2f7b0a2c2dcb3b6f0c23aef9aa72cc57a8fd5330f5d38729bbaed656ae461b64589ac5dce23a7bec11d68836889d2ba36013962cb7ad33a6915aa48124b8c31deefbc4fd8f476fd56e8d3f097c8a3bf5385c9f86974555cb6a10fd36137c98c467290ef170bafd527de4945903b51cb02aaba86637e1d1db871130008f483c925f9da42bb77d09c28c606794799027fbb539ab1634dcccedc29af00a2222abd9dabb55975;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf42261f6af9ec8dd836563ca68302fc10866504650325f46b104ef5c6dd22b56041defb9206b053882cb24e17d8760edfae41fb9e8ff0448ed68d0e0c1b019d0935765ed388e035b86fef24537015f7d7d1adf813d9b8c9c76eab5dfdce62cbe33262011e022232e635bcd7166f4b7816fb650ab2f39467e82621291fcf39c7ebd1c58d773335386fb40b5f7ac723418e64f485ea26385bf1bb51500913836a4c17bc9bf61e624069cebfa1bfb7d45f78b93eb53594850b6f7d502441b02f68774729cb7766f3459e8aa6a943ec5d4596835443931b0b0c31d615632fe45dd0cc1dbca7152e3cced2d27c87e1209fc6bd0c42a748e55597a88964cdcc96333860a76ea62030c7953d915d1c724ff5b4823792ab755b9c6410823348ab2692e80a8d026577dc02143ef87a1e2d321eece503cb559b40e5fb298d12599b679fa6a0bbd8d6c4490eae2fc01625ac4e8f896c747aaf253e2a08b7ef25b7a21cd19ae3ef4b3ebcbac1721d95b75acf62c0db8f24e13dd9d6c38407c2b21ce9ba6e794d1449b50bfae49f0ca1b3603c6942ac13a7673d6829f1fa0f3ab8b154adab60181d36da66a47a331ea6aa1ea60b5f978;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h63996aff3d036374a2ff3e4266dfa47f720ca2130abeb2e3026d32679cf46d52e9082c775b97bdac943c750cbd73e427ae1f1eed3424a67e8fa32591af60e4891448e4636b6b17a340d645473caa2fd73c7c0708082e30f94bdc3a7a1592744049d297220ac6507673ac195db2eb8daccae887792de07157ddbfbedf518d3dc6b2b2aca26c9f2b3672e2a5d39ad78ba490bb7a9339d0a256b75af6c32b66a50bd9a93298cd3f329472756b67b2c30f387f392f0a2c235227ef083704aab001544901ce2d9622555318d481144b53cb3828f9e82201fb5a8ad447240c3355f9162cee22f03c899134b3fb2355daeeb8da817ce62ec05ca98edfc0fd41af0812a6ce58286bd8ba01554c35a9656a30d67eb11a62b9bbcd531f870e0f2eb65443068d3215cb1a481990eab305def01df8abf2fd3ff512b37062590849d9bb7ff17b2c743fcda3e4eb2098920a22ff050b6be0feb115806848cc6c0251296514e0376f30053b6baa105c81202e4084b3b235999550c5b20b215df30e488165a7af98de66674d37d8df59b1e9ead6b5484c67d5a3b4d6176b0f2fcd91e5ecd6fb2257d14ad667e094f170413f014901c8d5d4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd796659798b8dea1d2464a309b84801b94a7d29736c184296a605a21579afdbef9b4b47a035b3142158c7233f523a2c9ab106db2242f7a118cb34a4f3437309a7e4a9cbe9011760c7bdbe6b505fd02fb83a21e91ff3a0bb90dc8a3e1279729cf8914a3ad7631f4a36cb3e0ef3dc7a7c1626446061d9e341318790788f59d175a906441faa99e939bbb97a026edc909b73b3c74173fff8a01c70b75e8ace2b9cf3e670a022f61595cfe5035711a5b292d3b6557392548468576656ac4f64a48a52777e27e428872d618b5951e420ef538fd9dae218b2b6953926cde602199d8cc829a138aa9a9a4681abd1537d84630a2516e85597f79909279a84e17be70e4d9a16f194bffefe63894a2c62e36a89d1da32d9cb71d2ca8befb7c6f5ee80cc84cb73ba1b8563c172f10eed6cfc75e575f2ae2f4378dcb8a9f78d1041225325f799ec44145caf9fd198cdc09be169211dfcd811f7bd301f336d2319a35b1904d2f2b6ec820b09c7f4f3dfa82bd099a16d512ae2a0a9293d106e63da62cb8110d67b80f6dd079f5b85ac46be66980c887d717b14043cec928b33479f059688208ea32ac360594a1238e6c3077c8bee9b31b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h733e931f802704c2262db862be61880b1f3ab61e15d60b8ab1aa1de8118653ef749a427ac1b83d5d579dd19165880fc08537c77710b2dc3a18e2600b52699314da66f5174de42f82cb51870ed04edf52106bfd38ecd06778140e5728507ee9c6b2c18b41c5d5b94bcfc95d6db15147667ea15355f1ae7b12ce0c8a768e9935c206526e0d58aed9875d6a7347339b49e94b14fd7e2255ae4fe6f489526e3e2af36377b4b88104059bd7660ea4c7702553d51c096c24013fefb9768729553a1fb724ff08c8210e0ea6c0fb9293613af8ef60f7ff4529f1e23ab2e0abfe2b4219ac14aa4db32d499e0e98fdec96d2b221ba299e6f4ae5dd51b29c028127f80638f669e03ab4e4aa12c462e430b317ebc79a1d96c4924d22d9d8c84180990debc13ed3420dc11f947ef5803ec1e09308748be78ce467c3fd4dde906fd9fa4c080ca553ce76b3f6d560e0516540578a3c7b7d68976d597b4aa40d23b90aca6b9650bc27b4a3e9198a8803f141aac8df5f9953d89089928b1b21f423ceef56e6406a813b0150ae57653f15a55b210c09caf4456fc7c0544251d5cd7f544e24e04970281b0ba7df141f8a749ef2b9be0214d520;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h5498dadf5099ca8269234c470ebaa8e108d2260dbf1f904dc1c3aede5211ccc370edc7a913e1d3ad417d48cb4d519f0bf34004eab8b8dd319bfa57679f374553dcfb8401f29fcb10f6dbaae281ca1cb37b7c2f8ccd70326cb8ae571787397c5ec7828122bf67ce092e6c39edd2baa84af9a88a2ad2f6e09cbea09a6a292e297b17289ecceb58c28df291d3b05faf250f565833b1531e9b34458c82b39fb14c114f25eebee08cb9d6b291ec1229751b95cac81541346f73783012df1d520bb24a56da80fb1a2ea2c1ba388da15866751cf4638b2f45ff5e2211e22294934418fdf90291b6ad4d472f1f851b6d7612604c52b1e232e2f0d06222e93cf5014d0162051fa94768d31484963b44b6b5722714cf31bb6f25bb6f685bd3b2369a169f2e18b15c31a22acd58ac31395535173fa8f24951e5b31186a195555e4568c2b9e766e24825a7f7b4965b7c066d032183c5ad5060c77789ea81943db576e34f39be98acc3df2be10f8d6eb5133f8f9a3d63f6df505756dadf4f7deba05f9a8ccc37f5dc8e1fd57ed56213fb9f4323612da452e9e8ba5b788eaa39af78a1e70d82cf3e8b08ca9d0992239a55a8cd2c46c9a6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6f69462f9f023ce4e1c61f8ce404f95d952a056dad0f584f04815c8119b8bcadd5c523ab34e9fc3ef94039126b2da76100209bfdcf47ef1e5abf824f68e709b468c48dd2ddb5ac1fa9e16705502ef5f941f0145b727c9834b6e6bd6a38e34ca56c5ed0980bc55806053b299c64539966af818f7de44b38190bf491c33a7acd14c8a16f37dff62301680f47a2e69dcda4a491db7bb792f30ddd9930f399705146537330e77628bd31757b53da3ace1db4a4d1b4c534f8ac8e113b05eaf312b42dab8c5b15b408479d1baa5ee35737d93f2c965d88fb80cfaa35d2909e0455978b6b885d611e008a402472969dedd72088458e2581b51ad69d229e35b9330230e15603612b60a232ecdad23e5bca1aa1acbf1e801d2944ae9600697e6693481efceafe5fc7f925b4403d6ed67738f6d58200ca557fa813391483cf1b35d0a336300e3e8e12be741332cb75afa6c84e0bde6eb254a75de59030f8be814ac038884ea51dab15566155c91eb14a531cd0210d6b1cd587fa925a557ac026aea93b6d6f457840165609d1dcc3bb2c3e6bbfc1ffb18fa2d28126f2a09bf05598a0122eca0191899c9fd1b149ebd8697581d4f7f0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdcf9d764db35326840cb5c8305aec07bf9e114702141989c71e6d03414dd2ba9ea317e819a07fdc503d4a0f1d7d4b76535855f74ea5de3217a85a00a26d4466b1e638f910a0789a0fa005eb024fc8b55ce861f294ecc7241b4e06a723d0ccbe3c9409a9ef4949249281ea1dd0dc01546f16de0ac618d712067321a86f2a306f91b6e08367b02e0bec8125c9c9494ac582659a1114df36f607cb311f83d066b851628db50d117c770fede2738cacf0b74f92715e7a0e9100cbdbcea33e47d934663b25088106da414788c5d0b5fc657afb810f4db4928d3bf26cc474840e510588752455e5fe3db0ac9d05c7d6ff3e1c6d12104de92e3ec070c9118a5b76b74925fbd551cc6d5f82237eba6fa25cbef7d66582f19d3fbaf4c78333cfb41a35e5ca46dee7976bbd3fa6c2f92dff8cb104c7ba7fc8f9ec8f7324d392c60ca31361972cd64b7889039d5fe3aa8c81c05003182e03675658f03eeb617caaade04cf1ef5df9f8954a4652d58c75abde90145781fcd4e585736a4544f76a6f8bd15cfeba962e7858d952479bc5d5c787f204212adbb7d5cd5fee1c5bf3dec0781fdcfebe45134f3bff31db0ffe88ebd15af9ab5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8d07a46ed57a060e8657704667424b2de04ab2f007a97faecccd84a7c47b96c9600f7dd26022f28ae94dabf21e9ee8c7c048ad2a0c155d17db708eab51c8b376154929a638ca22e2f06c5a9d3fb8a8bc7f23d28e0b894b8309628503e59b2363a9dbd21efb0fd2a367a3c69fc9a7970d7a409657444db8d367866e75ee318747f265cf8062249574aace8cf2e67a2b0e27223c349c8a77870b5fc141763bf9ef8d884c10754f86f0cc0a55a0d675bd06ce18602b0d681b8e4dd3a019fadad765e680ff4c396dca2312159c6c809bde5b325eeb92793a2f7a0dfc200081c8e8708e5e0a2d2d3170a1b9063bbbe7f7c9ebc848701cb4f9c243e6d7bd62e73c624505e595a3d86b03a3f14b67ab2cecc6f0d7e1ed832f1a41d897c9cdcb92b75d2dd27905b8d68f8ec2f4d5c10179cbe8c0f48ffe0020f51d220e44b783d78b2cb900e359e3c771d1285e58e113ce1dec6bb4175bea5db8a7a571ea2c877d551739457687a5e0989a5607d5f1396ce72e72938d8c583d4b03608926de9c12beae0e62d0d791f13b139295eb56b9ab762dc5daa13d129468a9cab991dce8ebebd7e55199068e69e7b664f9a245e778e8f63e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h45eb0f235a2e5a25e87c3ffccdab06abdb18001da1094b27c2ba216647cb9d4eaa149d5057c8e2384cdc400392bb5df5851c31f271ccd7416937ccdf6e127be143663d0c73f3d6cb6cebbbdb16496faa9985b0c033fe83cd8bd703d0d23358627e28a5c399a3e5faf3ae8f602a79a875984f1f79038d5beb35a4347e1c1f59918ff4334cbbd9e24c6516b556eeeafd1396d9c404421421c7075c8f82bc0ebfe03442a083b04930b02c6d902e4306aec7c2cc55959363057bd7527af06b4202670e80d59d581a3fe41376783776b169e624f3aa38ef681961c22df4181f8923963f95e1a310927eb0c6d62facb3000700299e841889989b7aea78ea76d26d1b8b476e1d4cde7ad8e6deb6f8e1ace83d9ace939db5afa22d90f636f2fd05b903582ac8abd5e4dcc2350b91102bb377a665d083157017010293a0c2147911a37aeb76df4e004f838ab87746c87cfd4d3a0ef3c20d78c536f6252ddc19a6b891f3c4bd9b0f0ac396812bd271c219d4db560e49ce773c326ce6dedcc4268af133931d3cd20222ddf5d972a5ec13b890ac149b21ec5771412f26632d6a2e9cdb23c568ff1221f46bb10d0357ef3784039a4154;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h11e4777fb4dbe3c6da076f85e5e9505db770ab9920f7e8d1131fd11e6b8421fa0895e6e3cc43c4f5003a5497335ed6a3ea35d4aa2857f216f8b61914a91e2f1cfd277bdf1092866c5d340cbce6747e6104acc2f8ebfff7a1795d4dbe9177dc6fa61895557ae5ab2c30d1588c12aee7ecfa94a2dd1195843fdc54887ad75a437fb7cc19d6a8c4240140a73396dfda60936f2f4ebd6eccc6571d009cf0f57c0ef338df30d602c7c57b22aa5113df0383a1c15fc70ecadab8a15ce920bd81a3a793fec8704f318a960f8cd2f00d1146fcd9f36c0945c63259f740032af5595bc6d40c697f089ba9434cf18607f81b9854da3d6ff13f42bbf1720bcf21931ce9ba043710a528ea5ee39542624926c5be74ea3edd5db2ebb701bcda0ca632d96011da8a88ec427a708351d46b77a05177379eccb9407605df7e348468ede40097e4f481a5a12b167523a02fc4b0197ac33e55ad87307d4b66b0748711e1a4e35f4e722fc8eeb70c4d8b7244ec3a28c0de33d07479b8eef5d34eca8ffded1d7aa003dcb36791154b901115d640fac83d2b79737576e9c9ff5c2444fca254e46ee5baabc0bc3552e706ae6ceb5e5e931349f2b1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hbbe04afc056b2b2b18748405550484943a470ec02e2d69ec5df315f3523abf711ca45d65c287d9e44fe956bcdc55003d1debc055c19e15be6f4f46778208b0e336daf6c68a30dfeaf55d52cb3c754dcd829285e47064b02a652e966e63c034ae310ef225283bb45088757f9364b90ac57d7a0449566d0c9c5f9aecf6cfbf2f1ea699b72c84ff298e6c74a555d67aee5142a83c3df68e884e2354a261e8dd06cddc4abed8279a1b08aa828adf674b1b5743ea9555e9221b087562e7d7faff0b28270ea745aa467ed68d7742805bbbcb2d575cff0b30e9f076ea2f2116778f328f35142c223855a123518a105865c378b6439c28d35a349a074253a27d711bbda2b450bd7417f5b5aff23ad813a02f86048ddc2be5db9a549b2ab9b026047edbfb274b8c6bf3cef9933e8fe2af3f35fad422db0530da23ea46632470030eeaaad491d58dd1b97b06e2da832e620446c5c3f856a2f1bb8f51af0cd4a59ab42beb023419914ea4c07624e603e1ec74db27736bc0f9b3d35b6bd01a42e70cd49aba0407e000dde87b6f79b438d238b0b97d2a7e41f3b13ae162345de5a9ef243c72a22150c0dce67fb8f0c19a20d1ba8ccc2f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha852e745899d4287d118514712e472709fed97a141ff5be62b73fc8b37bbe1375539a67ab212b84f479d25c3c874f96eec6262e3e69e5105847d5d47e69cf1a39743f6c261bfa1e4371bb60ec96dccd9e3ac6c194d141c77af7fa3d016c195244ea72edf7c196574561822b4771b86b9514f899800a5624d87a06430857e05df9ce63be68b85ba5546631b07846bd6d7efd0d3c2927160bf66635542d8928e08c66912268ad66d64cea39e51bc2d1b0454b7e0e9447fa017f543b11832fd7f5ab9bcd07dfba9be21aadc158f289e073a463c2e2afa52a880f3566da84e8d1c237915e4d47d767d9ca4065224452f9eacdd3c819fcb777b6b0af43e04a7bc9f0473aad2922639389d3a51a97f2c91f199a9d934035ab25fbede65ee21cf181d5204d0bbed15ffa86855e0e693be5d3c9fb58ae7acf45e94f2893e7b7ab142caa6f6be16cd43c6cd415d6da413fc03a30ce48c6ed8d773813368f75ddece82880cf75166a98fca5001e8604f02e64d338000ae3c00d31d96a85627fd3b2cc3aecef3a29186a8dbae977fea9ef4dc8d7830daf08ceea21933662d27314557eb9608a7621096ef2c763752d0754165ce9906;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h1a1f768311169f733a3fd7224e2257d577a3f56acc6b62f62e5b95ab5ffcf64ba4c6dbb3545bb9cfb411cfac489913b553b7045823b3469bab5d8636db231a43cae9b02fc4acfe286bec23258452bc822e24c14843e66284d3e9290b4e385338b7c819e045764ea50ceb39e942980b9535935766b008657b4b0a25f70cdf18c5d92859a36dd9455cfa05bda92d6594042cf6659e0ecf1054811e7451bc385d114461faf5960cce2d977fd1c1ad7a3c2fa9e81c85239e8f93473928ce6984f25f05d5f7c28ece0096e1ed6c0c81992028551bcefbb43d639433442856ecc4b6986e9cfbd6793eaebd782d5ae3cb724521450f074ce8f299529b42a547d51a2ee9a437cfad0919e2069f43326ddf76b256509bc5912022713dbb1d1946999b8730eccd8a70efcd86d774b1bb617ddb670293bc369e2ed7ecf3f1a252821bd1104d0e7f6d1d85b96e0a25380f4b5b5edf4067bff8c3708b56c39339d539949de3782e5bae9b047dec8793007af07a66f7bbed67dd4d704acbafe000353d56e2ff23fab420a719eebbd3e09ce9b4809ca37227630e85462d259c503e8a6314231feba62d725b10f539b505a507ec27b7a031;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2e75adae6477ba67d211a3ce71d2bd1f442c0382770dbc863fb27732c9954c0fab91aa37fa3dec5d2cac9a92d292dc6aa1aaa1e5c3ecdf067c4093afdd6f28bc425f1357a34585b3ba0adbe3f34aea26d3c09721447afad06ab2c5167b288fd7d293ba48423ccc451533a6604ffcc8fa0bc7c0118dfa2b9d78dcfd442ac99fbb57be010372339623aeb2dde9fbfc3954899e53036e792b2c05ddf1f93c747e520b43bd3118039df610dcfb4e5973b24b30ccc6b9287e11b7dd031e68df2bdd72f63eb0cdb56f36c88dfcf42fb6239a2383686cff655479b13d065c9f1f34e67ef8ef36aaeecddf86afcb4a719fb69c09af924b6fa61f712036a4ec458fdee7499300317f611f7224fbd8bc0694d44245d1cbd8d434c03d5fb23ef91009facfbcdbbb82de3badb776dbfae0e2789222410735ad1dc696d264f22d41a7722b588a31c755eb28dc8dfd481e8c860782d3f08622d0b0f44b3ad6c71664d6847f4a9ad2cc8f06c5d81afd88617a1301c97030be02970a53954bfe65282cc7154c994c5bde4e6aaddfe42d6b9faac35f484ac301c927df6c85372eb7bc743ac061c881cf83560567b15da5b2229f81231fcef7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha16c36edc259842bca9467e30d6f466cdc8ae34fb7fceff7264b08aac39008b4744a969d7d70bc263f21167b9382f1e21a15402f4d1263ab1d1a064d162b986057d7d32cd841af55d603a6c277a39ae2dbf21dd2899f7774120dcdbf2602a10bd6d5275584fcacfeb5edef0305dc88e3818cb06d7ca150260a8d583268ed869c31734451edb17fb9409f62b7ccd7455773eb3410049b7c5ce30458f529a5facc99a3b7f1aae8ff3b4d96127c8c206f9a2c235ddae2fb2ca34a9abd7b0e73723e25fd1818c7d9c6ec6883da791c87d4e05a04bf81ddba95f00a2fbeaf1b12bd4ba71a372d3168ca200884cc89c780f3fe988beb97df16b759afd8f03d5836804f4cf8c1019ae7e75015a3d17c168a31aee133c67adcdf40d5d587cf095af6ba5df7ebf7cc0c97165c0590ba9b51577db67532726f957d20332affa3eeb0f01e27d723aa47c757f7ee8e330d6f74a7d0b2e29c26aadb5e1063c2a6e6fc736fff5502b675fc67e5cd13363b455347e38d0c6c7d36e724fbc0033587f125d40610884b0ed785e5e5fac3c0a319482794a787260068d98eb88ee38e103d843ce5939f8610af9b85ddb5858dd28b4a026a9c22;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9141ca96abe956e7df301f84673819ed457452c229bd66989ffc24c0ab175964607552544b0535f5249d86f1158686d202dfdd28995409bffcca4edf03a20c56742ee2f755f4f9874da17bcda96c9349548225e6a7c2a9c0e27fb631f1ae902621ecf3f495ca3ff0aef92138a4e0f8919ba443281eb37b9ffcb5d86289a0a83275bfeaa08667ce330d7ca738ae6b4910e0375daf0ee79e2383f3f8e4be79b827d72aaacf3c00513596bf1bdbb01505aff068ad728b62c2b1911b798ec44b5aeafe6fd83ab16ba13124039b0a3c75ea63abcb2c4acc573c3d8b760b84d2b1fb76716482b4dba0a45cf816424a862b79384f68533a0a59a266d53caee7f2fc76c1295c3b560ff82c57e32d53a013b8b53fc7ceadeef3614738eda15cdaf4432f1f0624fe79a7b20f959efe6590e070a02cb1cdbaa6c1c1f15815ab1b4a28a7a043019c5950f60490243d74d24aeaf78d8093c775e2e6c4bf8d0315a91d37a04521662a876356e87dd7d32765784e16ec8477f16fc57c6bde66658b5522045b16f2335f0a759289758ff15c7cdf44be54ecd245f5927272a63563280266f6ec46ab6f158e4cd22db40f3b5eca83fd6e9769;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h41e291dd90ac9f98c410f902a0235dc7c300da660a676e9a6e8eb2d5c74305ebf4993f63ee875c6132ca9b22d77c4bf4317a00c1ac269fdd67d1cdba8a51fb398f41f59716a37956fb849e7bfa9d1d84c2cfaeaffcb0fa3cfbb7ad950a62fd5226c7e1877cb995b289a7bfb9a3ac472cccada2dc253f866367f5ceba493d3ad43e1b0f554d8562a70a2b8c3f5a30949fbb6feb30f797a52f5a887adaa85e62b1e9720f6a8314ec814ca704e1e0721406d1a40c0c5f8365f410fefc7c3cfc0097a15ce96ca4925baadae90aa6fd1452993c608bfaab0a23b183d06e24f7cf240c396d4907903879b3969870f392b7a253fed510ab6600407b0ef88b6ec1d240bfbc299de6daba04c5c04536557db34fde836c20cdfdadb9b18b36d950430823fba11af22a35ee095e5e8eadc00d92ce9fe5340143f6a7e23524454649a1967ee6dd1b9b7e4b88cdc4c8663f4a9cf07f13050cbeba1fd33d7a416e3b4615fb5909f6394f848e0245dd8b073f543ec9116537b77dde9fe3e8bada143b7d251489439761510a5b41ac3933864715fbafdced3b354a168fd29434ec29c5e3ab39d4e19c4db3d688dd063fe30eb0a393fb5935;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h124c058661a37de444064ce29d41254fee5be8310ce6816be4d8336fbd2208ceaac587080bbdd12ffff2917be368707128f11f4af5253aff61fcf33b84b6ff868ee6c5dc24bdf3b797522d147b9aad11c1d48db3d21caabf31953341b1f3f6fe50f2ddcf036e93d7df36979b5330359c49d21e5391922c5e9fe51fdd964568544401751d0df91667b0c1f1c825eb8fb6d4a8f900a2556ae8f443ad571e32f70bdaeaaa04259860091ff84e6774acb241eb6223bb5194f8056ed0c527bfb71f3b860329de92491bfe30b360a7a138e85e03049d246a3895d56c2a7495a8ed9d463ac69a7c61dc27aeefa53e4d9a57304387e694eb6a34763d0178ccec9d52bbab6ff12182191d560037106b0c693c6c37a816b518f0ce42490dcc73ae1b7e6eac1da2da86aab110858bb56d8627cd900abde1c567981be6552b385394d484ed3eeb99aca84729a4cecc7572509d9aa54d9e8fe74e972ff3ae69d125a8f8ea5496eca95c526de6c77bffe4ecec87cc3991d11cd37a4ecef28a3ce1c3cd5f8e7e8726011ed8cae9a07e88728e230a281086e5524d4fd9ba4d40b3c94a1a816b92a04c4999b632b61859f9901acd61cefbf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h1bed8e66fedb14935dfbe4baf1c8e6f8813602ce150580b148167da94ef45b8140227482fa0b92490df123e237a790c01414a48125e040b974881b3f6b4a52dac6d9deed2b502e55af4d36e5c623ac17045d346d02c9f1c887ffd086e12719ee2a4275889bb215a94321ea6ba6f84b85542b18b2f078920fe66e191429fcb03d13f5b44bb09541dddb885ab300b084986bce4d2f0b995b2230fa514e94a4c4b1b0719bb3f2cfe0160f1f43efafa9ee913c81e89fcb1c8e8932da439c64b244c5ce263e041bc90d28ec303120441b99ccbea8f44f2d3166ba039999fe3f9bb7b597ed3a6e36346dd3fc237c5299a2aa57ea343784653f8e4be5044be63129b67a1af9582d01a5a46bf87e9afe156d12a1d2e5e2d4145f2f2ceab19fc120bbc451ae3b227fb6cd38aa3d1fe820c508bf5f71afd9745a526995da241c0bcb40c312f644d2ebb9ae1ba5a8c4b3a377fd7c7eb3b08f87d620e8bdfc503d242bef0c0739fa85e6632ed506d10d80e2912be265d572dc3a2d9fd701c555e53ce98b9f6b1d4d51951cb2356a49b607799ef8fd19a0f5c1954e62ffc4d7cd2b1e9fdbb088068103f58d8ae1e718ff3c40977b41e8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h33f5fa81eca0caded1ba93a7c3c4dd1c592df850024d68a665d876af954b880ccefb23dd2e86f3e206f2c01aa4ecccec97adde713fc6f2d1ba766de8c41eb298f866a5894c29e10bd24c39bb989e6ee451ce7ac0040d01c7e12136bf28ca7f5fe0c6006507fae99bd08a59d0f37135ccc23e3b5c9fd812a4c32ecbc1305a0c4d3a3a64a1a1297c1a6f2115f12d9524f6322da744f7930ab1889aa5b49895fc2974ef093c62989cdbb1cab148c1053ee3876d9d7b4d200d36abd892348750f763717f22fef5710d4b77ab9e86813eba7dced396e6b7753e4ce4deec5b75c4f437425418316eed0d0c892d003fe0f8b4ec4c889d01e1df5c4909a6cbd7035bfdbb4a3722d2ed88722cddd2cafd4c3ff374260109ddf63f5560fefa0ecf86affa2f4a10abc1d8bc983548588f50a33641ad031a14d9c7ffbcb01f31a3505c2e431bdf6898c04e47c1d51f3a825032b46f0383e1dfd4de772b5ea950cc12cf40bcd9de8a42fa676336e980b7c7c5b61e700cd5233708a4119a9e9f295bd2f3f715aa65cb486982bd10028a362b6173ac09ed59d25e85f097db8c45dd3ec0d9e1942975256baa3a19d99f5bcd2f6b06d288f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h626acb3545cd478d3b9c256f31b0e785f7b42fd1c9cf60b3e8b1f33b223cfff2509ecad8a10c0c46ca0f9ca2aaf5a17e54577ec7118a3784b49a2e1e38ab8cc9fcd5d33a89b533c85915ede48b8ec41989bb3d15d8f05414fdf363b42b6fe866887fa2a777bed5e7c3ad39919f1fa8c69b58f9798d54c43c69daf92da91d1708a8dfeb9a68873291219cce812314113b9faa1d25a68457afe6aa09b87c6906c2a95d4a587c61fa993052e9e968496f82a1280453c8fa82049d774ee76445088bf6dbc9c8d7a70650ba98cc483919418f2809143df13ef9f6faeaa04e844d2b50a6c093ed8c94001bc3910d7d0ce4ae822b5664c5a81be43ddd6ed8b5ee5f9fbd4609beac48e30c4af0090b9a0df5a07d953654c76679f0f7a20f9deb0404242629acc899b44159b30c6420181d1cf3c99b9178f152571f28a63e8e7016cb44bc77d722ffbac0ede47399efa2b6334db64f381fd64540d105fa854c9e4e81320e9f6905999e1168da4d670d5cfc1c7cc18329bba6dc11ea269797b786bcbadaafe069494a9e67ccc77413c1228156dd3b282dacbde86be1e6d260d96b6b3841fd72dfe477aed12756ba7210ebcd26c15c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h85f06d54e84696d00b1d13753a3e12cf9352281762dbb41367d73b26aa8f074a79f68dea425bd74f7947cc41d4663bdb72bd1b71214fd877a1d8169089de865a26c5c619a01a4c3f449861a6aabd4e05d7e2435edaf3e34f17bab126ef9286bde66a29de65c8fbc633f3a07c56d15cca8bd3ba3fffa9a8b287dc574d5336561d25e332de3f065586aad4165e6022b2ab02679e0eb59a38f11af77580cc77ebb48e122a37b9bcd31429cff20a18ae64a6a2a7b32c43fa7928c1b0af83526bb6b1902a44a4b53a002e69427374e8cf1500afe651c4ee3b929fa7ee33e06430629ae4b802387244377b0d328a28168805d55211d1a2b58ad88e91dccb31cf236213c87796691dda388547edebaf1460245f71355c0e1c96fb883b002bf8f3fe53fb7d947b594800762fd757d183a685ca35768bde3bf6614c52b92d4bd60283ee83177664fd1b52cfb91ba2a71a321b52ad75c3b0c3f5d67766d34eecf3ebbaf9bf2734f526a4c6060be4c1e73ef938290eba2c7ebdf35d09a2c5b43f3d9f178f78b40f2a89707050d494b3f227cbecf54771fe48bf18e54b634f6cc789561d559adc0a901b0b23a692f1492c72689555bb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h4c3cba78a46f95167569f0eec2defc2b66d79b06a7396de308ec5e4b374910c405e79484ecec62c99f0ab157b16228d67ea3dc74858cb4981eaa59cdf08c2fa40ccd5cf98b3a48a0e222cf1f9c3001670e3f764c2ab0f3f71f99c8561430cae838da1339d705d8bd9c0e2fa9ab58a01d45382e065a681c3247ade108f1318ec50133805162619a3cd6424c738e43e148477d1c29610f4582aac83180a7b3da6e5274df463078a22203892d73d9f5ae991a45d6d14ec3ed7b5e45cb51f2267740163e58145345e027be88b639f34c52723ae79d088cb2ada6738e00c8979c521acec92bdfb7a4962cc7621789148476f968af2b16e4cd4448834556b534575d628a551d45d16ab5c2a51270c884ca4448d0eb4877c64aa9fa6cecc1ffa6f200d63a30d36e261531438e6515e943cc6892abb7941c611200d4f2c0e8f1bfda134a7d2039f4712a7d6e51cfcde99f524ddcacce5a8f65de16c8176d56a490ec48202b64bb6911b5a252a5e44e4f92c99c4876cb8c8805034d06507b9c94ecb84e58766c785df203625e490dd2959e9dcfbdab0114cea2ce8db3686379735aa4631babd8c619896011d222b2ea3078b7510d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h511c580d0f2e10d18b1446a8e09d4b67f6cba4f02c169d2a2c2248a206f1caef1c20ff7d13a6e31138b8168765dd10a183bb78af4331fcbcb8f16594762aa5cfbf7f9e3b72d87aab882ad45c2478778b9f96922dd1e6eff34e43b20d6cc8b3283332903366dc6a71dfc000de27ea5d722afc93fc394151c55140a9fa8309ebcea782d26d08b331ab7254a925cf1e128aca84b7b8b9a9bd9529fb5b859a468a0d639151bfe713079510ef20900e0025ac957cc54e2c681ce470379691d0fa1b772c43d368a6d7e836a9fabacaa42f979e2f646f6154bf6306dd90a1fe8d2e6b8dae9f27d723800e54304400583f5ec31aa93ae21959f4f91d3adc3ac40642c7cbde6b14173703dd1d715c06828582a88ff37046ad204964059a216ee907b9faf970f2b2ad0e60cc56986f455ce3101233e822530839a3264a50db37eabf36a3841fdae4fcb9185bcabff6168866bf77acd92c00ae5035e4f0f6999b2db95f62582a848bb682aa71df2295d7a45b7c43efdb6e37a8bc9a6b1eb2a31550f2c0a1b729c359107e5b3c226841d9888b5d057be02c0a5bb755dc55fe1937abb7e692a030210666e8989ee8f798a6a9e302d60;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h5536c5ab9c1ed8f3e4a2204c31bbb9bc1414c47fca35783c46e3b906a93047b9f6189547c8afd363562dd241388fd415cc1e8ce64a91c07c722d577164a628b8f5ee88082fa79dbed7fa8916d00eaa874e123cf3e3c7e74d4d7696b03d168f53f081be84015ea8217d78acf4024ca0acdf759f852ea7cd791223b6eea52884a76e6dec98ee6b9734bff8cba48f5a5c486dccbbbc41dfb3bc78528b94c6d109ae05b81832b9db51a74e6a328b523f8f66b61e01b750a980f84087865d32a93cf2aa99cc1c6093021d3b7c804fe2adb52807204e935b15ad48aab7b5ad598f4743f9c8a1125f602c59b733084e11a83810fe4274bde8b18d19f103eab6eb2fcac5901330ce9441cbe2316e28dff468fb1d8fae1f4a11a941540915b360d4faab9a23e1f4e4f59d083dbdc6fe5357bc6ecb3f92c16862997b5edf41ba56d187e5b91bb3b9607f733b8bf03659488259a44b53c6eacd112e74f6f7a5b58de6fc1c6fbd381ef5658254f49920b966c6aa15ac51863388ad87de5918b982439c224822595be521ab931b568d570477006b8b0fa818cc10ef6bbec319323764b1c42337943f8f552024949abf831e74def1b5c6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he6723983ba464d0ceb671d535c37df1bd58d4aa088b4339369a0f4326eff96be94d65b2b872d652a7ce19c0903c96c381c26f5e30749027f66daf663a6f642982215f2355bf576b42a21d4a313495fa9d4c8106939bb34708d64dc27fa28eefb077acf930f84e7aa9d46bef2c36029ccafd913cee2c9a37486815dec4ec4af9222d80d1bfce39f825b2e3b8fb145d3a6cfaf0afb9b2fa0ff97ae462143e542714041e0fbec614b72841753fd4b9b593beaac17b3203e06cde107385756a2f1536914bcbc321649861b9980bd50c0087ee0ae68277786f0f4b24e1c49faf779634299776114cbde16d279cb1e7a100d22011e9ceb8ecdc1770e1b0bbd1cd3cda7724ea2950cc8bca093c885faab68f0a8d9f996a6c764eb7e70aeb64f2203a9831e069382214451dffca45511c4b85fe77e17dfc06a65d4ce9f07e7f616c6cedb5153d6cc6de1f99396c0f2f11b0769329a0d6428ab310f6a02c6005b13da474db83ded29659a442813a823402c990168588f641a46982d222c4c93aa8adccb4ffc1f0392d35b47aca9d75778d153718e8bbaafe06de67b5d021b557d3c20c504aa6c9194d94b764192635eb172f32ea3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h27d1871dd01e30dda79ca7188decd7b2cdb4cbdbeab84a92f62f27a472f586faefc360941d70f36f78a180983c92651deaa825a374bcd3e0de4d4cf6e31c0c130f9bb0fc91e378fdb6a6edee1f20c62f09818337bc8f6074a17b06abc3f94de59eeeaaf840ddb62a11c9c40812ce16585ed3df638f69e4ff450ff77211e9cc24c11a3d59c0db487e3abdf1ec59c48723f6660e7a5d06a4c6fc5465bbe68f21bfeb8ad302644b6c6c0d0a099ae8fb979fac9d3bd0a6ea88df57bbd193ef2d999e5921aef7fd1d4996aa1dbeab1989b43709c7d7be8a80ac973656c4a9164b2e54bd2f00de8e8d0c52d0e60e52a96dbc6f95dc8cc4bbae07a980498d94f53fb208929f4823af76b2f4cbd49a904ba7495de25e75ca05627436eb0d6210b328496c7bfeadb1160978d02315773fc68cbf3ff9ea7a03f4de3a36c5976a1ce1bf0917791b6ae9d5907cbf4df8e8c10f6eeb7a4d7bc1e9e75b4fafc44445be980e003d14ed456b00811305f85ed130d5e90221829eab38bc52f04be2871b98d0aa870f5ae871c279edb76411c7754157946127d8003390b66e5f1bef4fede61b6d5e68f241798dcbaeda9bd233732dc9d137fb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h400bcc50c00bb108b73131fb766faaaa8c084569d04a6b4fbfa9435b0650d3a3282fb49b994306ad08d47b40eff5f073c00cb0dbd33e87f16c6e6a463ddc0bae332de3fa27d7c1f2ea8bd15ea1b765fb234e910ab1cddfc5c47374b4001ea6281ea19d154594c4b963e9f6963395e06acb81ba5ad7425d12e4142c082e88288c9d998b4c599bfc86241517a873c4cfa42f2d4db93a81c88801cc33585a4dd52b8659925b5dc6c9db00d3b4cf90d21e13cd02846ef1fa7614c5cb2ca8161debf1ff3475d5cd16a923deb294e8245ddf280d59e1237defbb15b4edb4e30586cdbeb32f33b29a745d382f4dd80e21f94d8ef6c5b0e0fd9b7b66b7ee6460e5c2c46cce8f3edc19a0040a1255ee4a6d9167d201ebb480f6064bb3df7b1e7c7b6e8366981f3becc3bf92de9bd191317a1532cdd52801ca40f727d982311eabc2d1cd9d3ee49405c96f418e5b4e1b5a8b626d2e8d2f11db101eef4d2da947b9a4db36b43de2cbf34b0ca197e0c2af116318eb478c79fe69c5c44a13b3fe4384ae93ee1c60b5bfbf730e9b97e0d4b7d21e7ed1bc5e47d83467a9fa2d8ea85a710954389012e4d2e015381dfdab5ead83aa7a2401;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd369992b95178f431b324a29215a9ac5c3c645df617bbd4c5a446b91dbfe3d89eccc7ae1f3bd757942bf3046a58081d42734528fc84cab012a0ef0f3179e3d98bb4d78c6c6c32cbde5fff86103058128b7472f1951183cf4e363863d04d4dcb9b270d29e8b033d883c1f5ece843a476f5e5e781bba4c3a92f56f674cdfbb5b1793aa19e472cd27bebca3aa62619ffe929db35818790fa74e8f8be43e614ea6f949cadecd35f44d61a69ae6c5181f8bb6b2752b1d475f99b45daa21969b06a4b50136d4ea576042af44306dcfa6e7c4ca1f1391af24f4ca9c54efe723c195de3265fbed52ab52e9ffd0898c68b5556804119bf88618cf2580bfe543eb5c4d69b7274007c5b2ed141fd104d169316caca311b52b8ad3e7db40888e834d6eab8ce6a00069a3857d1dba9295f5c30604a6aab3daee4ee34e7e376ce7359835a2cd35f2b620d137e559ce5376de7fc8d4812c41fb01c70d6245bdb8dadaa43c12af55bcf1b699e3ea47a1a572ec2c3eefd807e6234b271f481c03d938bae81508445989a6cb47261836e9290ec406145d2989ea53bd18a9fb0c96fbb1b3ec5ccd14ab7af96b65336f236cd8794b79b31e6cfc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8b11497757f5d714e559e78c8bfaf70a9df7945ee535f8958a7745e2076e42bb0a1cea6922aa1062aa162495586c5dd32d995ffe2a028c27115e14e4cd7497c1c23f32e5110a1b97646a3f7f878e77e8219c5efefb7ebe61745ccd1c5c02c38ffeca6d27780118516ac7c76a9bb2b294a034000f9c03185f30462d2c2f499e316aca3991639c32795002983886c4594f2a534f198696b8385b7181611ecb191840bd3c01432416758279f1d44a6f3391751806480193e8fc69097a06dbe1905a60a89e45c9568c20515a7a277355894cb8ce6b838b719cbb9c538a517340eb54eb24493b48fe6f299d947122251939f5c0cbaa3203ee3975898fa33e75154a76645ed5d4d1cc375cfd1795272dfc50cafc94bb4eb71ccd66fc917aeee79a6d8ddd27dbb83430aa4a87bbc30ca1f0d63c05aad2e3f313fd20abb4ff69a91c80a11fa2cb0bfb9cf4eb2ef17cbc845bfc905442b041ae280f4b15ca29349730486afff9dbcd1cb93f1080c8013c5c4a24a4e85e082da9d9e582a62199da3a848c094e9903e80d462e38812e3d9b71afc03d74efd4ab07c8793923fca9c37f733d4eb9fa6cbe9070c36ec948a517970d3459;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hcc61b7b39ef8d5ffa6d76ea1abfcb45276164b7708b6f1013663ee402cd651df805049c633f4ecea92badaddbeb33723bf94f1ac945f601284c9a0e019fd2db1c0529e3d9758d902e2525caf3da6afae6c8689df951758825d4ec75ebe96943b376f1eed3c69dfb0b04ad6bba02f7442cf9eee4b40c481dbb9250f006483fec6a3e5786787f64464537555d6fae23a6f0e9a99464fbeceba86562d61d08d1bf5f73e7271572b75bab679b9310eba40e91554c0f0c7e1c9ae217aca0067293ea682bd69ead84cdd44118260e9b312de717cf4e4e9eecf5ea900140a4afce64b569f616c33fd8f262c908717ccb7fbca1d7fbbbb275ec91f1fd05a4177dbc0ad91b93f2a32c728dee51114d0c2ac4d4a311c4af80a0a9a8bd42105a977e9ee707d86a4c9d71764cd78f4e09573e3a53b906872b1d0a459b7a33a33d32b7c2c650ef21d87be4cfd37f4e0792b0f15b6dde8a0367e208f88ae6bf9c2472daa6a5a3432b5e613f728d87a7e11dcab7090048642afe273ee1b9d6ac64607cec8601d25de8aaed3bba5b7c3c4b5c9d4edb5ff03ff019ff128767b86c281b1953f972bd6b7d1210dde2d13c53669884ad5ad4952;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd1bbb7138dd34294ef7ca79b67103d716c266a1ad1909b15c3bc169e1a387190203cd0888c0164590b6db9e1af8694a97c0b961f5903abef85af12fc98abe878ef4cd41a06cdb7254e816ba3e554055c8487e2711815d23c26383656abaa37ef772e8f0c114f4727247cd5a136c4f9d7efef2e513c5e3b8bb7ff6a701bf12d77aef68a92d93d6a9447ffdffdb16efaba5140d654b2cb375f791df30b7cdd24cefa1a624e3cebf779dbd727b152398c0dd578baf56bebf6ea65017b90894730742665c0bf330c974c9ac2915805537014d289f6bc094bcfb94a79f78696c5f55a7ec47c16fe3c86e1ed701f6479c14e5cfefaf09d0afdc16348269579fc27d3d313b5c76ee1efa88c6cc04edaf1288d1d7e31abbb753ad6f7babb0f632d4e24e5cbe2d6d47811fbd85d2f7b3c6df8a2a6c05612b85bf40e3df37535c2b9df53c59929b0e21d3f5197a79afb2d8f2aafc262f304332a13fd15dbb04a6e54d64ad12e9c93ea3b06c29c498336b465297c5a20c804f6a621f94c3558b3db231928a2de309bfd7352e65873520dad653640a6d3c42a9466c706a94e0e4370930fa78df2faad7a95825b162cfc472143f85c4a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he543696e9789d263bb60079268ad7535b2b46ad77789602e2a621e4241d3503a03c023e845d48c3b549c9842b800221aae3a39f4f0a08cb76e61899ef25963166b97435c6cc429a703fd891edc07f86a78d280a9b5c9aef56da172cbca6274222df2cff2b7faf4da6a06575fc1f7ea481eb8d7fcec54ca131dedc59a8735a84339ed8d9cdaa2c8a2f4984ab667b27648de28ecd44f7bd9219f7b8a166209d597aebb951b3d84d5fe8d8cbdbbdfeb6640e8384d87dad2ba3be6a883f131bfed4f7810b6d4fd41dbf14518bb46c00fb2fb19782667268d32f51f7932040f22afce96cc88de47dd6d83355ebbed8f643c29fec062d9e057b92aa3d42418657bce810a0d13b8b17d1e7c36a5db41a5912f413a7c0ee83577a1d8ad72d9b4ea3cfde5207b94eb14193f76a4a93d646ab946ba0540fc83925d3e9377ea9eaa9261dba3785768f9c3fddeac2100e514f0351dc8c7dc0617055d033e0b0028ab65111d5fdf2befb984ef8c02bd6c787660bcae7705cab019ceb176ee056a94bde0fd0e64d3d056e6a0a4e64a1310462f872e64a4055ce404c31c458f313006401a6c289992b8def321a547a98737cbeb74eaeab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h16b431e1f00010c1dbc34afd60c1a4de17b1940e8870f46ee8890eee8645d4bbac743d9141ea6d32f7a218247c1d6f30ad3902d040245ed1cdf0afbf25ffb14c40421740cd661426d1a193d432680ac128c297087af66e83884072bdffac38f9a9c53cc074e660527ede4573310f83b8ed0f1fd0208c5986c1d992bf451374c0bb6ccb270024f6f57ac86c3ad9fb43722a65ba81b8529b2dd8cd5d4d8267b5873c4169718eedef33ae789aeefc9347204e77047c1f5b8a92b97b652098c67dd563e961ee7457c9840b20b5459ab201a8770e8df2175dd532f45e3941f74405e9845e4af81ab3d9b871eb05d15e3efbe6556929d42751801ebbfa7e1192069a84cbac5022cfca92c40f939ad4d4ac3219a36c49dd5faecf6f57d779b58a14afbf259944202f2a85b43fc67ffcb459ce2c991af8156e338f0709f3d36a2508b08a486d3137c5b4d440b79dc3a7c6db0fb48de16ff1454bb026cd915ca2ac5b280bc94ec1b26d1d1be45a42798e92d9f3155622dc24cecf55ba9839c3ddc8071f273c5b3ff336fe44bd48d580373caa56e145875f6c303cf0f4dd508f93cba2aaabb186316201051e9ca4e527fdf405bbb0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h671bd7f5026722bb44206e25b999d28eaa5b36a8ed0309b1611d387f080bbee493fbc7fa355ea88685987f4ce928b6ac260ac8380037055f1d63a23e6ba7023d1dbc60632349de4c39bd59ba1f3f30fc9d0a57233954db923842581d3c81a7effe259fcbf5962c11598b7cc83ea2948d26586ef9d1f8b19f9048a0cdef7ebab04f8a95cda060b31a4ab2c1ca55f38f9c7c7f711e5d15d3eee75bee0eb7198a115d69fb2f2918a5c5095d63a16aad3c9f1adafd06ab0a3cc8947e6d0dd98831c6195e3b37b7f02dabbd436dfb3f7c67bfb9f72f519ac87acd34c7c485697bad79c7ba0641a4c8e65c6be4a6bc9be6870860e2c4e94d681da20d1b0176dec47d064482dac9c1439301591a14eae78534427b01f1e19796621de26244e7f007e6614a92c1a8f4e7756c627a0e71901278d14c45a66dd7b23cabe9a3f8eef9e5c586165688acc5c47012d9975de66ab8ed209248294de6a7d001b279545ae8abce84eb54acab135480ecec0acb95de8d62879fb1bcd3e40ab486e01e716e6176238a7ea94ff01ca183f14de2af994dc5010a2d4f238cf7a1e4bbe011776af7b543f7cec98279ff2b387182a3cbc5d0abfa43;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf9f465204f6a2fdefee8c092840e126508707b5aaa706bab509777c91c10cbfac270d7b9a984b4cb141d7cd1344853e2193a3fc2794edd57c45dd425c8b8a8086bff3036ec2e285e12fd354c6e004b8c74cde2805e223848950bae621eb701b31e236d6fd7482e2ee11386743124a3513f003b2e7bc0659fae472d51c52f8a5f9b3c3bfb50e61ac12ec2b2e6970c720296bc8c7cf1a57a6ca3c04a0f03c494f4d4c322bb547b5712fed9c19aaa61f0f5ddd26976c239dbe17368150a976aeaf896d592822f765cb5e3af9c3ac2986d564f76d06c790c2cb08a66a58499d7d9a019fb299ef2e8da79f3c5039a500f2579104a0886bcf5db393daa451a533b0186bead0816c6a5a682145e8f318d2326d5e723494e118107a0addc1fabc4367482141aa302b2e413370c2b0692ef66acddf88968c0da62568161732a550a23d70d8bce1952b4f815afa8a7e5962b6ffe0c95b5f2337982eaa467117b476c77ccbf353dd6d9b6a2e845d3dfae6d325ee9fda67e95ef28d49312ddbee870cabd37cfd6068b4611fd66afbb0600b5fef13aee65544ddbb829be9222fda538bdbaefaaf0c7d4c084c48af0eb37439c7671dd92;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h670b92e29fb0fe05704abd77509075d947e0f2b4a6df038b2df3c2757726abd45ea65cd717f632907f50cc2e29539bbb22fa5af50d5c6be53718ab879bbd6bca5ac551b9b54fdb48952436fcee5cd9551cb33a73d2f98783d66f0f205d82923de02a1d8cb2d1fb26ebbf30421ecd617d0257ca66933f994497722eff1d901bc943c68194632cace820cde0e0d4cd0e09f2ea7525ec8a4cdd42afb8d586d6bcc42f19320a175017aadf4c2ab1e59d0b99d630141363d4c149ad49f117b9c183712086809d189f52db106f028c368503a9f1c428a31624bba649a14029d7f44011678b1df5490d514e14f54ed4cc40d51fa2fe4aed30af2c9ab4896e26bba987100e64af20e86726c594959ceecf086c65f9f768b8aa4af0a48562ae9b53e6a4285a133d18f1282204f422a194a5b1f8cb0d8c6005157b9fe2e6286f936bde38eb6782e74c694e9a4f178eb20b22d205d5c2fc8de384cb3ccf6e110ef8e1d2ea84d78c28f02511e32504444a37fd040141bd44dee55e665ee0fa0a80045321dd1da7534a4771c730f1bf6ba0cd29aa495256396b86227f4a09b1c465314c3fdde07ab7251099020933b3f08accfbbe30bf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb8885b7835453a5dd11ff6d3c86bf120d5692d874bf2e7656638547a6fbee0b13f6b8b5d919b5c1a3d139b5c4af2f939cd393a613f8208b16a54f456038fedc712aa9083936e9693b081ec4370bb9b185f0101ae6ec5ba7d9d098eaa10484f4d65507471ef66d612cde24de9b45fdf45fa4d80d1a403754de943c4fa13159d670f60e081a71b1f31422bdf6980a2320046187b344d4e3fccdc2fa72fe0881488fbb159d3996af0136b056662724079458b7de6a20eb34f310eb40ac543b2fc0d846df66d3735f4252c82dee16c2d4afc1519e96de965628b9afcd13496a25973886d46505b7530e1779e1935ee938bba3daca3e29ed4bb83ccc9b46b67c54337d1ec9ce75a6990a43524ffdb23bff873e49f5969fe5a54c245b436285d208e54016aaebed0b369c4599cba7aeab49c73427a3c6557a61d8f585e15deffe0a91b3417727ab7108b5c54f34850b84c1251a51da11f041f47e2f8542d84d265e55fbd0438d3598efba203373126024ab2ed5cbbf486eccb6cd5d60ea33b75d7a6e320938016f943a09b4b645711d7e5aaf25327f3ac8b629c39916b4dd90426f2f03b16eaab962a2049873061ad059f1a9b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hfa000f37b8f389d05770180b2c6ffe5bc7b211e3e4a02fda28f50c628f1ef3879929f3662d7d893993c00e15e48e26e71a2337a761aa5991223467d5b7ef5b740001c5182bcc549f038083d2e0f1f130b54c186d3840ea6b1bd0f2cdd7d3cd3e0a466b5401c127d882314f331eab3d9edfcf5ab1ea53444ff8c36465d69953f4db5f5c16951734be34beef5d2d8e9d070e77bd1305bfe3a2751a1b32a4c4f981d6f781970c9ee657a46fcb305e94add2470ba1a13b6c094782e0eaf36c91e9da32dc74acb0b18878419e7e50aba2a65f3e7e3c67d1f3f236345421859cefabf382c538bb56a225ecad97e201e28de1d379c93980ea27b67d04699810c6b360a081b66c6c36e4a981480b6cce25f4bfd1a388c410948d250fe0e69eae7c7f2a33bcd58e53c443e8d421a39be86ad52dab5e622d5b6cb1fd50a9ab6969fdc2a3c226b7fd49c5be4c862561baef714ac91aa901066e2594aa980e07867e9efd20e3549adef92fc6927a96fd8bf2ebe9fac981e3d65ba01709a6d5186f4b0aff604235e6ffce77e0c4214f74200f8a5e8269b0e092250cb877265a830b2b5f884abac0526da5f594f1fa21c725d406fd073b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd9f7d6e10f4f2d92f1ce43be6035127c26d8858b97860b1c9dc1b33bd923832d32a08718d1c2ec0bdd1906648bf672c5471fde5f018e03f2c562f5191dccfd2a2f355d855eb5545e366bf8cdda69ce776bf26d7e5967f5a40cdd37addb6b666f16bf627de2fc6fbfbe35e1db2ff06558a0bf133a27c4b4c358493c8fd4d3dfaca35ce19c7a4b55a5138621072816a35b3fce0e35fac92a6501fdb7614b7cdf7bb2adb29680eb3c9055b882a8253798a008e4af20ed31a797cf02dec1fe38dee1fc68b085251b1ce4ce8aaabafb9421754477eacbd971e9dc2a5bd6dfe791e882e7651a50b09cd8e46e942dfcd4f9a3ce1d6efd319b27b2ecaf87ff3e526c2cac0be1b125bb1a8bf08802ff7e47fde864c4ea6e57a254d2aa6d33e6ed830141f3202bdbdda5a482131fc83a8f882685d01560cfca924992a27c22e1df0d1ba28f183a4d32a764de1a4e20f30fb40b367bc5216316e188881489a33354b7439f5b2cf8231df94b49a61b2e5dfd602a096c60b68887aebfae5dc03319519e651d696f9f6838d9fc3a8db0abf058f9922ede2ab2e1517a5afda8147990b2974abf5fb13df75da64eed3d0384f290587382a1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf3fa649dc035dbaf9fcc6e6180b681456262afde7650d97525be744eeec32d16f3c1b522adedfd31ad69881ff4e6c577d839be6611cf3a03367ce08ff26cd8eb6117412e7e2114d4c969282e55091b093e8e067a5f8a202b5b081add1b85e8eba5e74c2221e5c1f511ed97c86320cd3ffaf456213ed4cfa069c42c77305b63721c8db53b04c3198e7d291d32ffe59bda882857799b2c71b96d18abffd66bd289017eb219945ffe2ee57cdd75a7c9de967b2f8b9b3f2dbd802b52d60cc0a6f9facc892ebbde80639c546f69775d18e70eedcfab06ea3fc3471a253e06ec79662d28845d3ea1ff11c2e43166e329519b6b27b50b11d17bb2b6c99a629a8ac9f7b5ae667eb770430819c7cc2f60d9a925ec3c5c373b9aec8dd14818178ab15aeb6147d94f54abffc94080464f2b1c162d27faeb3c580bcf231ed91c4b21510511a0ec2fa3afe1551e9fbbe36b031b5ec06b46a30d5ff38e7170d5ae5af803be6d42ba2be9f64d468859c371c65663205b652636eac2c3349bc7fff4280f58f33288fff57a923278d3cd9ffc2de6d3b680d1894f36249bc6d61f984250882d54dab03ae3d4fcfcf373b6f34306628265640e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'had15149d6835a1046180f28aa4d354db8c1a4ee213cfd21d59fe3d93d893b0bdf75dd9feec712df48c7571ab468c81675c9d334a83dec30ba586ea2253fa49797253958d07dd362c0ee27088a3a0d6dd9e4d92a04acd3f02e0cd51d042f2d7ef7810bb7c070f5275e72d03a5a2d39ab779867d7ff7c6d5db6cf60bf2b1693523d05ab7bcebf6701025949302dbbdbdd1eb82bb45867f64d16a3ff2ad03343d0931e60acd2bba13f36f0a3e4549a1dfc48694c64648f7af0cf8794112a244b5f33569151662456e5543a738264e573051bcbccb705de308e0a28d4fa082e1a6c19d91dc95a04165dcfba6ad942cbd1481ec8f466498ad62cfc255321eed8a08bb18a43624da77362a10850264b198515e43f31b6485b8317e811a5feef9340098297e59cf079a2115a0a23488e34d1488bf053cf25371e427bacc9497603862013b73abeeae02535d1bede8dd2f4faa202e6f3315b379f062ce394d64632330a48b33c2867abfdae8e1fac9191591d7054e85e0f75ac035ea28c7461552845b474ae074d2773d32035944a6254d0a52de2940329939695253efecaeaebf0735922291691617a9b2453c2ec18c09101e5f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hda430a65b56519b60e514473f48434b5a4913047d45c667c6821e486d4480b309a121daba6e6ed52392650e8ef466fdacc0cca5bce22526486aa611ee598bee99b20e0e287049a64e8e7f144a43c5cf4ed5c5ce098e992a5127af98548fd07316ec0afd9d0c3ead5c8186618601bf2cfe3d58e4179c08db617d6834a56a8197ddef17e911b9e386713ec988a22face149aba6e99fedd9453858644e2e898ce52bd7cc55891dc94e40835a5e32397b14f4a0960c03819761dbfd50656f4881dcccdfab9fc4f4f6069b58adab314c33d233d45d36d8ed430a13181af004f8a8e5544df94d86552cb6acfef5bc9224ff50a1b8a50635e6da60b7b181154417602171993f1538dd091648e369348e9def8496d6d9db584685554cba559cf59d020e6345043135645a1ccec4540573d61e6819aa3f98026e569fdc04dab671d7ba99cc709d68514c21415c5aa615efeec15b8416e40113066926d14bb8d5723c1907cf90e46c91353437c45728020350c2cb01607813673785887e2fafc7a20434635385aa00d6d98cb65e2401a6db52f90b7e5396b36f73f632ab396fe61ad8a08f3a17f064d4983be1976e4e048fa72747f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6532e899b2aea61f4ff837273b1d452c988b7193bf047d22a6989ae235460ced5c5dda57e4ce70eff067244d0d1a361f0c81e9c7384d7e62b434156f4d6e5429a35e42f86fb8ec58906e5c76ba705f96e46bc09343ccf6873514997a87f1712745edfe3d13ede347fcda7bb0690cbb2295f5b6e66f5e509be94f444c8495e6624a87ed2c7307c5f47ad3cb5bce8e83e69d36c656b6d2943aa11b9bb262b5fde44a0bef7ccde99ea7b762e1f6f86935c93a975c7156fe7f3dae89759687482636e87e36fa4fd89bdba317f47f37f7049d3b6def15a967bb121081ef1cf325732a781c8bf2bb59d8bd8b72917da2cb20ee72e0c03e115c1564998a6e358c2e23210bd984a9ce059c647c06d1f161668d6ac4fdf31ace80af8fa24e96abf1e3f4c49991a0fda224901e2663fa3525fe7da42c7161252cb302ea4ba02beda78fb889fbecdd0b3e1ae3e3a9ec1ec55214a763251ec4d5c2b8072799db4108cc01b34b0307c2605a56d23dbba2df5c7e0f39829e165a34c17d5681aae764ad7a0d6089f714a660957d1ccd6d327c1bd5ba6d654bfe221345c24feabb545b96e50dd3c4642a76b23f232d4dfd97b603109ac57d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h4d242c817315d14e9092e9a03528d9ccd0275f4f1f1568e12ed0a4449bb7cb67d187668d743a7abc9f02c11f80017f5f114c78a294b0991d920788a1d523293e5f81c7c476bca8c60ebde6ba35fc9792bda83a63e71ad4a127562e4ebdad59a485e12c7cd6393d79b4f58905532351bdf5dbf1cf47ceb903edfb69010e462b1d3516d0a1ca48567e1062fd2fb16c2914d79d99974a1fa18bd57134635707ce9601bb096411d124ed4eecb1c700717cd6fc96ca41ad601a1c875e19ddbaf835ad5f2e8446e378800803cf208f3c9bbe539da62500566b155c42d9b129a64a478fde2c665a8523b08a83517eacc4c8dbaaeab8e425b9c3d5bec17326ceffa4c53cbefbc300eb8763e1caa57de4a41fcb99d9f823205fb53bc0402ba91aa05c400ed90ea5243d6ab898ce2b578bbf45aa376bc89732bd9acd5f26e72ffcc8a1358d22bb27933b6415235716830c537a47dc24a62165b409df2fc521b37248844fad60781d3c52cbd4ca61596ced77e1c377eb9fee4124dc9f2226cbcaa319055bb9b073123216d4157c33555d4d071c4d84f8222d0c239027324c7a1e55f805eff52f6d471fce0f190a74b1bfabf3239a49;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hfcc5eec583f275157d6772a45c355196969087636b3e6a01dc7edf6961287acf56a6896619e795787f9a23fceb539ada4b233bb4147cd2cf9a9db4a955962a590ba4325bf473e368b9120060eb5a150dcb836d5578347c28fba69fbe8d8766a32a2419e1faaa8162c361b80a75cafbf2fc5e7900e1518d770c1c39ae63c9341ec8fd237efafda4bc00a2f7875227dc75c08967cb52c457a7c0a191e1590adb44a50a6fc9107c8bc7a379a75a8b6ca90dd352ccc75719b9193a3c519cc12c20ca5f90cb05985d98460ed803b1d422c628cd546b2bd81675037dd20843eec096c4b701bfed17d003f5dfb857573fe3c6dbbdd00212a21509a1bfc3b7e86426944e1122928ad244c2b9f457b601ca86c38037b2b0b40a5e4e1174170c412a1471a765210518ac40698bf8a5d10389aa4bbc5a596f7b8a7d4a260d3ff7f1678322e8ff4485a71900828289d7458e8a97b5f6a6aa594da033260f2d4bf5f714642ddf432666e81accfabc9247c71156d1e398e2ae2f686b1a6eb146eee05b76faae7a07281dbd414225872ddea9012fbc25b50e3a37ac19efb2fb4707e3be4a5c7f07e4c0007abe139fd98db12b12cd890eca;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h53863db83ec475ffe7134d56de0b200b4bf5b9d252ce181a4e440d278f24d36ec0fc71fa425067847fabf03f8d8e1cfa1d17adcf14c757d4102ff14484447f387750673f8f2bb63817b7e252ffff8a4b1ada463e1cffa85918e76045c237447d2ce5bd33a8e3d099c4f75edabba190ccb01249196990aaf150b742eb87fa57a158e82942e8a0a3c8b7613925aaebdf038839b16c8236c88581b6604672d0290a10161229630d1a6876988bdf8f199d4c241b2500becc878da5331f15cfe3a5ac1f68e21cb2f78ad6478184ccad24c6ba38489facae4ce81c51c6a6e753ace2d144cdeca2f4c2c3f7468351b771e96a055e8ed4ce44ebc5632292d424f4bcd6bbdb38bb10a46cc2466ae4e33bf7b159e85312575c594b63721fad081b90caf1fc761e46fcf21255fa030ff68fbd774bf9f0c54899eabee729ea2d2f2564badb4a04e12f1ad0d9ba52d40e88adf3d69a809945979f83ac1670a965c19200121f66129b1a77138a345996d9cb4cc14df902afd4702aafa44f6a4583066771dfb781aab8484a7e6682f9c1f3c1f7fa29275967c8eceeb962c2016013dc5a34ea09c71377ae4de1fd63bc0cee0bc1cb6b7191;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb6ceecc27e6c5087573cd9efea028189ae60dcf5f15190b821dca74f86705409aa78151d97256ed492b611301976f0a6ba3bf700123fc9a920d347c0d5905aa8d4a6f29155c1666024fbe6e4b142a405ef61569216e598b13edf41863732a9ffb72b10247a682fe2f91089d151dea0ede2611e03fa2ff6a13527bb7b8c41213b9fbfff84b864556fc590024c829087730fcaf8692c9e262cc714f2ef37e3334083736cf95dab5c0b099e8eb996e227a6d5b846fc02fe09f00b40c818ed6370d31a24e0fda7a78bd0a7f4a1bb8e5837b3a217853034cadb613f8f3c6e412c3946c315f3034cc913e44e87258062d5de5bc0a843cf5afd661194b3d1a83025b524f3ce286924f724e27dde7aec0acd98d4d02939b7d6c2325dea1983f81955bb52768311fef982c9f2c3ee3a2473aa90f893e7a4f503762ce06a3767ba31305a4ce6476f2fda8c6a2bc0109aa03c911594a6515e804753759e49f5a8761b907909d45118c977317cb495a2348db89a6a18a625fa783e22ac50900c86ecc172fdcac0094097930bd21a8f99ab10a3b7dc31f94660849dd4f0b3045707e3309abed8cb3c1ba48415c31c383d1dfb56ba2058;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3fc966dcbdb0571a23f698ef72389f4c2cc4e9ffc1db76697f6848fc5ea402479a2debdecca8718b287b7733f672eedc33e7f7b71072b65064ea615e7e913b93acca44d57006ded1d03c9a0c5728168addbc002bc210f93e135d8847919eb26699488cef55cf1693b7de79acd91ee58c9713e82246e187b003e6f395af4ff2bd675b75d9f0545b2241ba007d31332220d154d2c965de6eb86b51ef29071c9ceaaf386f291a511421a7d34a1ddce4caba7f7318149bf9eaadd16fada82849704090c746a2bebb2218c87944e276876d74144e85937526c7c4b37791f015e428c3397904ceefa928bdd9c6f78d07298352512247fa12817ce7cc40fe224e8ed478149ce2354f731ae995338f55f0bbfd8f551ad72aee1b276ce4edeab5a8828a83d5bc0e6b61c90bddb252642f8903e58b3efdf0c59602f13cc53fb231701210eadf2d08341f6d9001d73aa77c633bd6861c904620d46f019289ed4000a63488935fcc56fa88973973a77b015e129dec069d7f3bc8dbfb09cea52e28f622b613d880c92468e30b18502af01ee05d7d3cffe50b94d4ce9de2d5cd2a4456b5ca5d9b140a750d621fe0f89fa9277ff9475dc2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9634f052f06a7200b1f084f5f3cca4e50957ad00fc5badc417e1f9ab7162e17f0028b70ccafef8c94a0b79f995a5cae6fff495a0864ba18029be54719ef5e01c869a0eb8ebc0b1f5912e930a0edc69f4d1b440e52b068e2835b4df74ea8de2034cf8bde82ec9d3c3954a57bdece3811896bd3de8aae1b16197d3bbdfa5650d5206683f88a22100e1024136979f6d490d3334ce8acaa55cc8268a0263b117ea3d0918a5316cac1a34b579d34ec31f4582986b99ecb116cf466c53e4b396ab0a8fae775bfafec04053154b30104be7410fe815cc71be3199c952a680432611e05ac290cc8101b344469ed7e54f0c0143eb42de5157bdc8b356e8b294600dc67bc96c833c7fdc583ddadf7d93c150897a69343c78feedb3658ea607523013a73900ba8b30ed1bdd367078e52fb43fc90c3c906e490d2077104327f7a380e2317ae6031cf0646592b2721ace1162640e20cb0413cb7a84105c725314782d5cb9a9fc0eb94d9f21eb4ca464ccb46c8c724335e34437cf1fe13ea4679b79c5c1c173102b99273eee06f21c5e8ec732f69021894a64f4314f8ca707e290efe3a8c3c0449d216c53e06f7ed1e4c60d5b2632ee4d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he97481a4cdf5d29afa12d4a1c78c8ff64a112549299ae533ca89f4c76848380db64d592e618a86a24bebfb7ca24a591ca7dea93c5d5f12e9a371e4734e0374924c22d8218dd623a30167febecdb05a4b714d1f5c8c197834bac1bc0f85f4afe0f5dca565186d5187167d40c25bbc3edd5d193ac004c2c23942fb26dda675ec501f4a25b44c7cf68e1eea8f030031b2210f2700b025aad54d60f8af89affff81b19727ed3c593a6b325d6f2de0f5fc3fcbd47d99265d87546abab81af430ac008f317ae4e9114c089c554167242857cba590026af1a97facefa245ad6692d9e308ee3892c8ab2c787b1124334004e360413a2f94b50c5c982c7fe1b228d636ba08e4eb2954d1b632b76dc7fcbc561206948abdfff23b29a354baf0960117da25cdc739af41e5e7a8bb39ce2aff6d5db682349c1c3314b4710c50e238aeb14ec50599fb4ad03f220f2e83c62492b05e5a16c4277371c9a906ddaa6ae3b192a25ccc1eb2ef89e9836988cb4f6f7ffe8ea298881eb708ee40de5b68bc782d83396d31b758cacf71403f2737a01dda6910af1aaf17fc15a83471000e21fe6edcd9342bea76f3b62735332c018aef87a2cdabe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2df00983a919fc37c6245771c6340e2b9c81920ef2c1d272b05a2a86d422b16ccf6cbef07c18f4ee005629f6e75e37ba6e81219bc1028ba609ac077d21a743e378570417adb91ec97c0b74d48eff6fb9362804e4bee8314069276ccf8178b6019174bf426928678ea96254fbefcff9753e5356b9193091bb1e70ba2c2db16f1b1fbaf2b7a4ed69c950e4e9d60b56f6e0e5fc6f70046bb1c306987baf8b49ef58a9810e62b4a25581a27df670e0d6859d9de4a148e97d51b327c6cb6c3ea37fa976d9d05c293e331bb9c7bc4504481a9468954912e4884deea099cb4ee7284fbb3bb4ef7572596060a35a472a8c60ac09b1c887775ad8daa444051ed7c8464b0ce433242bfc5ca0cb05d0e1825e72e7804cde2e3054fc2ee384c491b1e53ac19f94add8d5712c37e2092e3ced966dc1bc58a1214dfd9b27d9db61f05b1dcc77cb7f6026f38325a0b06ed5ed341b928167da6d472e55ed27dd17b6d0f4a921e5135d0d9c9f273672d709bafbcc28943fea2994ca023ea51e7c5cec0adc45b47f3297efad7a7c94229f9faec264818c0bee286b503a1f9e1d8b79b6dcee78d5c0c5a7c54ca45043966d154d6ec016a7ecc1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h5e1ad69cc22a75fc30b38f299af5b7e9820f785520bb4f77b588f2dc30b55afb9050d4954767cf50a2f97db58fa4bee7b84d60d6508ce5883b5c211ff707cbb658eedddce40dea7fc24afeeb7ffcc2213f13e77e15eeaa7057a59820265bbad29bd2181cd5da86a63dfb67de0f4581167454de95affdd0111fc95148fb7c5544fdd93a38c3d0df01ad90315ed6031b36004c7c4fa4db9aece747d73ff4a18a9a3b691a8c16dcf95d6a94cdb0a6f424c18df2bc8937a913af6b750e664fcd711531d20f849412b229fdc2a3c45e6720504e348dad74230b1ff76862a8e752b0d1333e2ad64890a7a2ab142a98347371d6ef1a17f8a9663216b881c9a04821fe2dbcbb307d94af1ec9f715b6bb9c8dc2d90b28042795c16f59951fd0c2890bbcd11bd71c7054b7b5a8468ba32dd2ae6eddee1ee05ac725fff886adfa32b5ba77d0f857d12365d8472ba6c04e13f6840509a218d6280a2fba13c5537b088247c5a006dd722ba51799883eaa1161cdb474a5d2ce2c548f5f8579d3a3a34a5720c01befdcac689f4ef22b9edd74edba85ba19fb91ccad86ce9e83aa33eb1c0cc0f467af39eaa14ee7fa0df3dbabf4a194dd2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8d0a1fbcfa63465bb550d7c6b0ca686bb2160db384b5c26f31672ee6a28489fb2c3579b6593a9cad198de81e8846dd8ef486b4c01e70b1d7502c48cd45af47b4b396d80c0bbe3e62fe7c3fbd07925403d5e5212319253c6297ead18c89012b8d52721b7021cb63be860dbee1aa2266a9372a351eada3b8de85a15dc6c2b4401ef752c02b4b08b186d50e03c73bf6b01545c7b63dae2e6188c444a40dfb46f1f213473057791d5fbd9145ac12b9f5d642c6101096dae5c8453b4cc306f9d255940c3cc344755b953882e390f7a3391a73230baff26e6d52691f4b67ff9c915fd7ccf5bb61963a6ea819e634e5d58f81924f890d7b03e83c33909acf7d535bbadb0c51e5e5d9418a4fd324b234ec5ee86dd7545853532cf436e22ac62dd705d9b35e217f307401c1cd98068a1641e7d4cbbba8ecdc43b4990f77620e82f9d4a27076ded658363b9d310513f83264bcfdb3c1070404b84e9add3c7df873f3b41811df28ac2764707f9e9039bfc4c2f1ea13b07e916522d6cac737ffbe0de9315d09fb48abee4998d2ed120af391fa542f45274fbd762a3b906a8d8e2a79f6a659f6098b8d071fe8fd8b8513fd62709190c5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha31e26804cd53b9832ebbca0f9a9bb2e4806c969ab0a6e6bf5b861d5ae515b3e258d1e9e4882586ceb5d6bacc02c9d429a4be6e383e1837092719688957ebbd74991100d7628c772ceba20757396ab3bcef267e0b3e4c19726a327553050f5f2a1e4d0ff2ef0d8914db128768877805ec70748307dc0881bb4a81c027068037aa5f7352ce1aab2570f4bf811d1666c087e8f292647a92748fa244a18004ddc384c3da3f713cc02931334ac392fa438fe58c05c2b65b587688b68ff31b321a9bac6e4c732f8b48404c3627f1527abb74c28a2c2123401110a4be1108dd0f9b46a237deb6acbe0f2b9bc94b36356f6a2e99105f561e4bc98b42447672fd4683bfdc94ed63a0a4ecff6c355bd67cbbffae1ec0afc800daea915c2715fa57aed92df4834752598ed6f5bc7856780918ac141858147b0fed6d8137c3caea300452523a72585195c5377757e198dfba67d1ab8b70bf3a926fd2bb4e16a02be7ba316a946b7f1852b1b973cabd3b7685f28db7b064ec92ecc84e8e953ea0450faf53594498020cf1894409154c78e7a973aac9da637776c7bd9b2fcbc280686205b62186d9a5bae024dcc6c1516d950b5879fe2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hff6264ea4cfe03d82224bccffdda97974f9b43d0a1ca003c20f8e6a66e49e576fef66a447f12517a9946ddb97475863f2dc38bb89e6b61641fdb877ab66c9c38ec6c1a691664e174fc994f3acafea33974b97ef0432ed7e97df5f158e800acd4b2a86f0a1c3148fb49d80afbd51e3a0cb3140e0dc050067da852f3e61edfe6ea8e91055867628a9945fd0d1dd84e2bb1d97cc41a72e4b1d0b33bf35aca8ec19eb42b028fc6ec33e98ae83e9bd65ce9bc9e3a43b94d5a767f186316887e9382e464ceff177a9c2083abe09a1065701b136ac965a6c6c0079b99551d5cc4664167aa1fb7d4942a3fb9c4ea65d7006a65d9ca0a4aa6e1ad43e030b7fecb6e2e6409694a71cb200551aa225721f95c689bc823916ac2860e0f6a550f354e7b72d1f9b227b59560559360b529165b49926bdc20ca7823bfed1e1ba92fa2db5e8e39601feeda3949bfbd54ffd0d3098575881bb1abdd00fcc21cf2f413752b802dddd874246e00449d91d4861867ab84567d9b9c465a41b860bb4335343ddc6a995558daf55b693c1fddadfc657021fb8306502ad5ee204f10e143b83742c4c0aba1456de824ad5e08a7a2270168f7b0db6fc5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc3f0f626090843a1b2c98ba7e7137c93518226ec9b1f244cebe1f570309246b1d0f4a72fabe1a0d361f648049ee957a53768779d08de0885c5d1a59d50a0ff78261ae308b3de23d1e308e55e9080666dc926ce203844ab0bbc66c81f0017d28b7ef419b8d2f4fa793530ae1ce9395c3a1b099971eae6ee5496961ff24ba724bd78e52ab7c58157cb64090dcdacba0b5dad12963a73d4dfe8f2f395231cb878d5ce998057fe4b5eade7103e76c986551cf138f5dd115dc57093c551582795eff74a92247bab6ae7a1833366fd53dc193fd63a04653e62283f5852a1d180f73e3c8a9bdc9fa5352494b096e348516f0ce3654845d2e5c7f2c3dba41ce5f1256018169dc52cad148d002792b831cea4a73402347eb7e1d80112eb76693a96eab061cf653f7f2d531d040e1f8298e3b85b6145bbf93b9031c1be8c8ea8c42d56954db430b4bcee49d3a7c14703f0ab9cbe982aaf0d36886488d93dc01071a7c86e830950d09f7b5e20820752a626971fef811d470e67508a470cfb0936c514ef18824898af74013071c6aa37b6407c8678d9f170b87781c3e4fb9495501520d46c1514535fa759ccbb335a10c5225108d299;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h37fa95c048dc872c54dc4cec7d6936f04ea6f91aefca47d0ada77db902c1dd17a17deacc47436f437d16c411179c2878285d5fcbf0a508aabd9fb006a360d6c674879a67067763111fd8ded1d0b6c5365dba34b8f259707892bbce9c63332cf0713d64e10bb46746fe2e610cf0bf13f94eb2aac719a4602913c23934f525fa09e6889cbc8286eecda2064b256c730f085e928f26ec12b9e733ecfb30bdb1a509e042aea5db6b5609f74745484c4270c63d0d938fb444ad7c17552b2c729b7d32a8a9d71698613f140fa0501b7aa5531b2986d3ef63d29617efffd1cb2127368bfd833f4dbfc0d5221635d01fd4e07c04bb4aaf59ad55becc6f6335d8f8f64f240dcd84fd76b66d7591daccab26b0c5470a6251dae919cf6921b966649a14cfa0c723ca36d0614b0ae204a70de1a065f3a1e3d147d75d86242c86f34ccda96d9563b6f5f9fe6b000ab56caa8506d3942144105993066626ed6cb0984628d85ada9ba54e0c1ab558788e1a33bbe6ecab065f93d2e654d6994e81a3ae00cc41650d5100e7bf5c095ff919b47a586b16e33190cfe4251e3ed4da24924a1173900ee357e4b57aca487b80b11a3de30a518ade;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd331d801b921437709e97bf8fa773bae2c7a9ac31d987865a55f0a10d39c82e018a8bd83968fe3672cd8efaf6d7e35f72d478f4348c3174d0da3845576cb1ac46cb70b06ad7a28140984943f86593aacf895d194e45b048bb09a05845200b8dcd8b352db6bbb3da4a8ecdb946f50ae5e3be1d6651b79ea380275179f3014402022b6cdacb96e8dcb804eb1be1b24ba646b9aaf752ed3fe9c7b2554244a695da9bfd5d816a8cd187a9329d12bf57f2ad69dcacd8ef6e45c2aa2e18d78e00b45d6ab896c7b0036c127d51e3a368387f75059a6807b1116363fb7ed92967a44b3d2c653363e5977edd16513b7fa3ac911f5605a3d36c04db4d23905867b7815b0fa196bb300baa6eee03a89ccbab43c8dca25e29fc74c6dca3e3eae7bf4ffc83a0979ea674b36fdfeb66f8f3621c4412e4383b63e12e19832d00a9ab3aa97712f342a6c59d0f2ae74c166cc42eac9c14eceadd9fd31eb8825b2da2382a1e7250e44702499909b9e6bc13dd57700e09150d2d2ceaab5421b0d86e426944388377d1b77df5d87f74c2aa63eaf8ddbcca5e642707d5720564e971e6a5d3661789ae1450552a035a298ada395050905a5c632d2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd71a7d6145b573a6f1ca6e0e352920bd2d9946a797698a41cb02f79c837221723d024223b2a8b1bdba94e4b2d5c7c6302059731a25727163bec7475625ff64d0b8008b6754b925bb015ceaa087d438dce1539e26737ec721cdc3a6ce5edbe72b1d162dd4381e97dbcb75df5f0c1e558352d098abf686e2d7b6862103c996c0dbdc917437b5047ae7daa9fd22db77c51e4778c38a05e18ffd313cae09809eef90c301817d54d460ace16887ec1b4f155d63953115c9a81df417daab7fbfbe9b972aaa149691138efc91c81c04d9d862e0dcdb240c3af339a8914ea6298bdbfa8dd49bf3f12a4608de21090d50b0763e27a526a75916eaa0686e5832c40432265f1c8c9e064d80f7b0b3600583712b50303c2ae50b49fabe93f0003f91df21ba666b243d9cb3932b47c820a4ad4ab826d7c47a38d9b467e4e1bf7c6da6903fdda363c76dce1b861646729352234945a7c4d5d8f963b31b8342f1b20e6712cead40fa9b9fc23c8120671b554070532c1f262bc8513ef8d11c906af0e224bcbf68bd23162c07afb9a243e98bd57a7c4cf1cf737693b8e06199fa1b78b5c8a55559c42db0fb957af1f4b6fe2405b77ceffeac;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h7a885cdf37493e900b3abb33ba9f6899e9178dd28acac70fe87b261a497beaa9e8eedc698fd9866f877409c0579f393359213b0046c1e05e17be055bf2b392563773288c9f2cb472a3f602c08c81ec7da0bb85fcc3174279f77c37245e6351b7d5599a95f2566359a8f00c760446ebc78524916f80f3ee0eadf9944a7c07a04dbb0d9649bf2e2f709526fec98765557bf5ae0f95c3ffabc1ac8e03fb5e761328e183469760042daf14d8da0528705f156c415ba5dbb819eb14a29731eb7966a641f2579524196b9d9f96dc073c19b3d6d719d813a4799657cb622e13d39f2cc9a2532b4976284a3eee27cb9e609aa3207613184f0877535a23edc23e80f7fc5cb274ac2883ae2870de6866dc0f57bda671654a3609234a42cf458cd1c6b2ee82166080f40c38c220c16b93242f134b5cb755cf27a8fec87380b399b38639aba295e49d0afc48903a60583cb2ff805a88346c9784d8507b637cdfcac5b0986978fba3d20731845adccb8472eb4a0094b00adc943f1b2e9afee52a24ca46fc4fa306c3c54a0f728593dba65613956a0c106f09e58b249e1e8f34f21000bec040242d9f9569be574f0710cabe4f89d3f8c3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h311beee547183b033b6f0797941a60a03b8ca90ecc408a76cf7cd85ce0ee3fec9b04b04b2f604de93d8a6cbb1dbc869dbd139803c98f78e755d44f2a214cd75841f9f3a7076964cc1ce379a6245130eb2d981aaa7b5d52d8725d447b28fa3199d870a77ee4909676d8d6b7898b30ce6bbfd94d85de4dbb7b865e3d239c055379a1a24a546601a5174a9ee9e00238984139af4dcdc6174d8030f3290c7974398b0c7850399f5b54d5cb7f2405716ab7761966c02cb8318a11e7d97efa56823210b13f00dc78cbb0209176f099fccd76eb928a0ab2d8c7ff3e18d64264b64e0dcdeb43f3f9f954220befb9e981b4d965819bcc7941002b89233984a68b76aad3f216b9f4d995dbc0fda828d1b70818f6c9f9dbb77e9b5282fc62ecd2c18e71c443d9dad918c7e6c1546910ce83491e4bbbb42137bcdc8f71d047f5196ee9430fd9e9b9edad8ca1cf9a7539e897c290035bbc5a28155b5c26446106a918ddac91960324c22a0b7ae780d23149721de694adf4b1406e499b71863de1160c423a76655cd972affc9672ba9fa8b50431aab12f09128dec1a820e39b3b0161d257b0fd021631b2ea5ebbadd84b0746f218ebb20;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h83847f56429f1b43a4c2f1a723095679ab70ecfd95c439b83fc10a18e1ac55535957545ed150904cae4714e2ae1b80101d2f1f778372f1cb117e717be668b3314df66f43928d9a5d05d484a37d620bd18ab6737de6f36234fdeb5614f29bcbd56bc7d8d44139ec78b6299db57445a83c720932ec86f2419d976f6a30876a336209415f1eda67586edd33b57c887448b8400e828f42311da1a2b1a80f0e421fc38294353e69dd2350b0fbe3a0fc81cede7ff54c736ca3e8892f81513138e1553222c684a939a10c1ddaf9b70d3f73e14c1ffbc46991b0a0564cb64a6ba14c4cf3ba71b1022d530b2380b8368afe7092e1429097acb2295c5b4dd3470b43f3e89d278152326d254215113507f2c8ba445b704e0351d4c4c3ce3ca0c6d3a18a6cf20f7f9e8d532c591e965c5203ffc7c7949b476f346f822185b2db8ac8d5d89142f14114883f9d072004d258b983b150e9f3b800bfc4a1d046445bd81c9b1e3f41ccafe2140f69ca34fbc5ea2a89e0789c16b356f05d8bba93b18c762101dcb146648353a29cc2135dc213283be936a8158bf2269f0750505a381baa293bc9c8b3687956800cd3c84fc24293d0cdfa8f9f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9a156153e9bd3c6a65115d846925dfe09923fd053d6a2f1e88f9291159b8c66154aa5e749186ef78c24b7650fb44d03fa5dd01440ec66c709a556098552969a5fcccf697525f6d3667ecf82cff5a8e3d3144bdeaf6cd951c4164d032f08447727458310e646b229560686aa8850c4ccf5d118791ad4dc5bfef42da157d7c55a5fec07e81404b7d7b7b78ce6da9e7cbd526de55dd7a49b5f5d92f5a27c673ce845fd60380d6e7a17175f711f8e29e947ee8b4cc050a609a942605507e1c22827e3245a3cd98ad09ac58959993a85b383f16b89fee989bf5bd27aeddf3c97109232b3289c57cdbc20380d445fb1d95de8f58ff08370d0b14133da178c5a18899af3768c80bf4bbbf3918478261fab89d1fcbc3e639e0773ea78257e0a7f0b6f23010b0c635822fcca3793527a03f6f8b530eafc8bd82ab540af713d64efd678bf175808e90e6c1a75dc87a0a6d2a5850f4966a651e67c5b96f17985f4bb1c2f00b6de207c870cf76894376ff4af58121ff9cb98c5343f04ba0651179b1ea55b0b357672747118509cf7d9bdd1157146e195978c0fa06b73578e9d452fef2c96c4fd40736948b3c7628027e783e98b794b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'haff75d58e58ba2242d23d6de2936c07f1d7b6d4e7a97c7bbcb88055ccda8978f4c0f06b51d1154a20bcb8aa63373044bfed47590ab79017a1020b237df8137aad16c7ce512ec006e80d26b4ec023bbb829fad0327016a74e993f23fcaa112f2fd3031e434ba1fe383af2a6bbe807d0cde3b23c4b5a943c33248ec1ba1cdfc122949aa09854e90879654ca54af91b0274d16637fd32b0b3c7909d9ba50f4fe0e39499409b9eeb7971d05f397e44ecf0c80cdd8b458fc35c6acfe961d89f9f30488bd469d911b2795b725fb24427e74db88b94971d6dfced322d26c665413468427c3fadfc3d72738d1db83a83fb6c6469d7fe79c48a68bdac3d025afd2ff8f8f861ee58029daeb5edd9f7f227fae373061f216b542c61d531cfb69f0766765aaf7a4e27678aaae22bf137dddd40f56c727cb5ccb4d510e08f8136cc8f301343c3a95e95cfa1983bcfd1f00bb4fc7ce8eab9836948e44e8776932b6238368e0d8c7f6ceefa1b2b71f624e9b43091f78e937b43e9b523b9f99935e8b14c47e684a97da9e6c37cd814a3a7ccb9e9a71d8dd7c706c46eab229c11df4764fa68be9b4a839e2ed9c05ed264fc066d01e88ca55e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd262d9d61cbcccd852995d4b300abd2f655239fcf55e726e2e1e8d3c118c7ccf9a628cdf73c2e91621ae8d6e466c68c9d5682c59acbc3fff0db4dfec23301ed0ecb17dafc179acee6e2b5f9adc7bf90e753afca72a6b4117844aa579e32c95d832b6fdde0c43792ae772ba08fb7b9e2f6ca599d95f810c4611f9dbc46c1914733800fc18df8936e255bc4efcf1b7e208d2e1404d4e233e21298e48ebe14478c252545a883141abd07c65545fe2e72469feafa2cfc067054ffbc4ba1ba41f3d555a0c83e1b30c9d5106e0bda69afe1fc7eec013e3b1bed63eeb988549e739f6126b7b4454a6017569f11431e6ff7cd2addd56230ec28ea21e9f6620c9c17be6cbdd30de9ea2af34d315003ffa3b3b5ef262cd24818a68bb84fe4ee5bde764c800a2744e41f6d4fa8a93e2248893705243feb28cc9c2f849e8213c859d5b3cc9b2d4a36371bdd3063b037caae7fafa80a01e548c287e2e456ee4de5cfc8fba32adc319d4e02b632101a8d7db7dc1363804adf7506c1f5044314d1e1367bc6dda65f69d169845d8a205fb385824470055c0dd9707e863b5933de305164ea493a7544702b5e24e102da4accc554aff5a820d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hcc678294a9ac647c48d68d49194c53e4f7879b58410c28134d671dd5d88f4396d17ee0de1f6c1390540b477aac879ebdc237b7b86572a3d2805ac4c8b69b417667226600fd1e2e67ebe147d6ccffe08ec7c681baaa53b5d75ac2a586be27a7a73768d823e7a801afaf098b54bf77a484d8b6897203638bb251125d37e68110e694f0cbd6cf3bf3c3981586057d84330df6447481d9e21184d6c26ad07361bba8af729f74daa25b9c04a8b9d9693eeb0733a6df23566a09a341b94f176a3d989398c5b8bb59a362f62afb4e14c118583b597fa987e41df00ee71b254657c4bcebc471ef0c2b1d90f74abb86f445f526dcf955978097004aab6ca62cbaa17bb4949b65cacec0e59f4c58ac2764b1b0f7dbbfda71d5d52007db89b895c2b5da84b12e5c9d7dac5eaa92554f523d065c52937bbe4a0efbed2fe8f694eef1a5e8a1cadc754f9f113636ac1f4d9dfa24be818b698713e216a1ff5743b4f8541946e8d74adf8bec7950ea4150478481cf39dcd793e6ad321a314f9d61897b58bd799700ab89a948345450880c53a0d9653ee869df36afa5a55a64015a95f3475cc1800ee9a59d4be303f952260019a29bf3eee8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb40fe3310d47a1b3b445b3993ba99b347269684720ff2dddfccefcbdb46a378162401bfebfc5fd92340d874286122b07357415b6e9556a50286f33fbea0d9c3214403a5ad06d2aab8753743d72fc209bec147af3b9a89d8c6955899c7c7a0b67f9dfca09aa141725163d6292a817ee75b5201703fb9eacbafaa7bdd78427704ea46d559fa2854134bc59421038117f27bc1d92b559b2775f2368e5618206aba98d8d2664e97bb57b1916dd93c2f871faa3291bccd20c6b11d5dcdd85a22fa0902adfd8b71141ecb0526d650854ac42aee8fe36bced83498fd570984ce6760f79f2e10e594eb426cacb92c874654931c8197d7a2290de0bbcc4bdd9020fbaba3123cd2b88a94569e3a52ca8a9c356adea9800dc8360354b0d5d0ce0035f73fca68aa998b0c41477e1c5eeb3867f0a20e9c55909cb44b0982bfd764b5d6bbfa5776cc9c5eae9fee4648e3f0dbbd9a7ec45089a8152442594077ee49a879ef881a69b07d6ced41aa957007984dd8869a76cf725584cc11a00693ed31a144fd14db4cb42c1e8068aa43511771994ac74e006a2cd721f521e1c83cd9bcae375019032ec1142f2d4c597febfccd71d7b6bae17;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h91dd44ac20eda81a7be97ef5e817a4aa7664be1c924803f6ee250b87fa42902ae53e7abeea8603470d71ffbd9d25f39e12ee5ea0d924ed358f31749f974f3f11d94307db13851f5daa5cbff9c439f416318bf2aaea77fddffb7fea483434f58d0d8da754661b5e5d1d993aff81745e63bc672a04d7cb13c2e0a7af8413291532f5a07fe49f4b2f14ca22d89543257a97c1a193d7c53d7df08036bdff99a75eacf8f8549d2e200edd33e5a6b1e78cb07f6760b54332f0d42a970d61f80d29caa00467cdce760310169039fd6d63414bdd175e14622560b7d45d4538f0eb71eb72c2dd9e9cda0d26e821a1178e54e7fe2134ef4ad54868a2636dda8ce27e6908f2f66593385d4f4146838c65c442b3b2bff7f5acb3c1064d15c74c35a8dab0cc88dfa799656ff9707cb6f54152e09f27ec068388d67a1f04c8e7ff3310b6b7f9861565054305b5346dbbb2fc38938ce9e6a8b3600506270ee3ac56a1a21658c9ed7a20ccedba6f69f213a0fdb4345f588a6a7f9a38b533ec580a14c607f2bcf688700e7fe0f66392b1d33e66cee6fff02d9bd6edbfaf8fdc78931191f7fc0717bb692ac664cf93d23547a58b6accb4fb7b;
        #1
        $finish();
    end
endmodule
