module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [25:0] src27;
    reg [24:0] src28;
    reg [23:0] src29;
    reg [22:0] src30;
    reg [21:0] src31;
    reg [20:0] src32;
    reg [19:0] src33;
    reg [18:0] src34;
    reg [17:0] src35;
    reg [16:0] src36;
    reg [15:0] src37;
    reg [14:0] src38;
    reg [13:0] src39;
    reg [12:0] src40;
    reg [11:0] src41;
    reg [10:0] src42;
    reg [9:0] src43;
    reg [8:0] src44;
    reg [7:0] src45;
    reg [6:0] src46;
    reg [5:0] src47;
    reg [4:0] src48;
    reg [3:0] src49;
    reg [2:0] src50;
    reg [1:0] src51;
    reg [0:0] src52;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [53:0] srcsum;
    wire [53:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3])<<49) + ((src50[0] + src50[1] + src50[2])<<50) + ((src51[0] + src51[1])<<51) + ((src52[0])<<52);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf5d17fb1de37789ee08f04b6d8adc6029cd08676eccdd2a193b34b1afdd6b455b496366dc9e537a49b11524dddd69b76062e632d2ffe4437ed83b136e3f825f95377c7ae83a8b0aca040c60ce6c08eef607c220ace98e7de70af6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hac85acb57bcd5186eb32dcb48c7987bc94e9210a799dd1a1bc7fddf93d86262b8c698f180c0d964c2c235ac51a47f567e49d667e8ffbbefe67f0e51a7271108bfbc7e8779625da9368dd91dd5310e398ac28ee1e357aa1ae8f3d51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147ad707cb3eafc82e5b35879946a00f4b81cdf042bc5347846baf4a5087a025784fa69627477c1a5e5b9ef2cf9215ec4a5459939796b0a04cf489144e0f17948b9d43f855442f4786f17b24dfa7d37fd4799bba03cf30d4887686a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c77d95f50e9dd486e83dd4d0a24f3b29681f12c031ba8a72b02fb560d241fecc4a5deb06a493fe0cb806851e663dfbaf9f48d0e76cfc7759dba9a19f4e1b9ad6469d438a8cbdb1127360e7600a7aba769d06241bf9c1b95de4659;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ae06c56ea7994c9fbb2ac47adfcae0866e30b769491cbc9b53118561b4527fcae8ea4fca0b2e7603041adccaf90cfbfff9302130e7b72e1f994d14c46a2244655380054575f2ed3bcc3d2e4b7f0d15390f640069f9f4f5f890431;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156b569d365a85bd6645d45f9f47a9628ae0b7a72c12bad5f9972b909411adf02e04f5ec3da9d1894e12465e67373b52a73961694f98995919dfb218b9a85e5049be0a9028af125e57b91bbfbfd07d6031b0e1c9ae2192b05d4c5ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fce5b5e1ee52b583419aa595fe6c73fdc999c8d37c84e3ad1cf12882f8eeaaa042aefa05aba5dbd685a0e11115bfa9c982274227420782d6b5cc80dcf4515a50a2eeb59202670e4314d062e71bd2a240afd980c878c8c95d8a737;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b09c735e7ef1ec4bcdbfbf4bf31541d34db1a857626186b3de148563f79abf6b7f7bee41e9a23c1d08f2b1cdfc872218c0613af92dbada1cdf70c0ecd6da2a9abc0ecef39d8fa47ab05e77624b64a0f6f7a6bf51a052492852a97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d295fa2dd1ec648985ca4f7488e541a5659878c2c515073f57265145388714c1c9012b362f84f2a7226d3a0f321297cd26417935a378cf3d574454df78b6b2aa2ae1bafed2def8fc5949055e075ae741b075f1a49069c91de985bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f2c0303185182c8a35dd67339f3b0308c59a4c0f8007e5340ebbc6009ed10bf1ef3a0c283ee0960ea20a9a9a965a3ade1fff952d56fe5d7879c56f556df90f2aa7803d075dda6cb95f625eb4af3ee854cb14cb6f5c48afc12ea27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b33c68e0d43fcbdbfeeb794e86839fc050d8ef21104ed06a73f856fb2149f01a961e9e9e0a180456f17704395f9325a29a1bcd8355484690ef32fe260b1c8f3cde3c87218b58a1b9274bdaf07aa5e8b8120aa2e414e6bea8f5536;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3bc8c51110a9ddf5488deec0121d4076002a8cc59b093666331435f2bf628fbdd32301625f1a0ee960c3fa24e6c57f602cd8d47fa43e5cd146e1b4b1f83f668417f073914ee1d8aa0126e0872f6bbe64cba8255fcdaa978261a0b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc71442161156b6aefa45d3c8b9c8fb47a577ee0a5150b1382bc8dd35758117a6fb2f5cd2d2de85c92a4a86d089f2d190fb1651f5ef729054bebf43b113ea45b2ad5f53cb8bdc6fce270ffc2e0d313f55c45a7ea34b3bc82da8fefb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b4ddcfea3aa298ee05fdb5c5a4926b4507e1de5c46096fe945df26bd245129f53595f742d751aa8330cdb2c9c7b7bae0b7fe990ebfe546d3bef4eee553a90a892dd26b21ffc99c5e1db18ec5ef6a540e4f05d7e713765fa1e267c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169c2a5677bb32bd47fa02353dc854e2ea7fadfb7e301cd6860b20ed02b151b867841ec23426f60f885603f13f58c2744cc527d3022f93edce9db2aeb1c4e21e8a40e6d8810f90bad3ad51ba135b772fbe497c901372af89c6bb851;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h704356ba7f8deab1a57a279d2a0888703d88308f24573356707fa32d64150f1a32d55bf8aa53db0e479bb473306a28490cb4764c0e1a430293bd2ef5e3c593e29ce67bf7bf8e317ea19992e60563afe293a0cf222fbf32b747657c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h66d7bc70b68c65ce9ef707628f2ee13edcc6cbc47131dc64e9c11ee976498cbb0733141b981c2d13b28b1b28a5db90034815fd791c9f08f0c7e662c9f076a9bdc2c489d0d3f6089a4945666e6b6b6a7f6b87daa536f3988500ea06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d669efc1c2eff2586322e186ad7246004783f8db07c4729d302b70382235e8b38fe8368671ff8e06f0d07c619e81ec32de836d8c6270d3f5534d6a848f84796070d68d7c09a8af5d1c0919cbd9d5a5700bf0f9ae358b84f39aa38;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h109a3a755090735b6a3f4ab1835f136ec3e732d58d5a20327a2f54860032c3978ee7304bf4db64dad02208d697121b9dd92de5e7cb076b82eeaf371c52c7906e0574e8fd2da880fdbf4480d4800b218db6a4c52eb2d7ed341587509;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14395059bf74749ec0f48fcffd6835dc18d5f90efe38bf48a0f0aaf30df21145d52eafb855f35a0bcdc2a8e14e8e373d3c552e7ca5e7502c37324957d47c10104073a7d11fabd44a54fa426596c14111e888a9e2d23d14d85396397;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9af5320612f4c9a78a0aa71845d2ea2036a9603062a4f06c8b61e415e8c707e2a53d641af54c4b062e90fa53cc041c91c48f94830fa348656945b88e22e2c164d4cbea76cb20b18e6c3aee03f2b5b631003ab9cad84192d365045e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1505de29a9796cd859a78e42fe3cf79a0a251475da7604943e4221d27dc08b5bc275713b61b726efd438eca839fbca24eebcc41168f23d55731b1fcbd86f6f17d19dc2f7326ab85dcfd32374a2763d41704e6c7b4c9b40f9f85b44f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7671df2bc84764475756ae6793dee3b5a46b84f3aaf60289f845e61c1f42bea16c2a96f442173dabeef784a79fee931f868cc6f39f32078cde54acf909c6d3c0a06028b0684da2d256fde4bddd8f7fa6677cae20d83e038c555dde;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c3fba36882ff4ec78dd98a49a8d5004bb94d30a257bc5d1c490acee22a915416c93e571c51332e839500d66b235ce6cad049418a468aa4698098c58db101099a37ea66d5f1690a80aef02043b09af5ec87ab0f49a581212217f49;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd82eb0f2f945c5015c22825e78368d28dced64e65ed47d83ef4a34be5cc3b8ed86692c8fc3d48a1c2684408c3d0077f904a2df16d126a1c1fcf95252e4ef0bfd428d16356c86061d7e46044af122112b089b3026ee98d8d284c0b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c221339796c1485b742aba8b7c20219bafdbc5529b9d1207bebe9fed3ab06d7ec0455fc09c06ce335c0689f36cee45b6346ffe514afd14a8736c7650d97e73f4906b25adfb8fe263c0e54750e70da016c7b2ed172aa0b34b477721;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b0a440b6317f5f1750b529a863e124c0f72c9370fd77bbab055a882bac989db53c75f87b73e27518e529dbaa1a205983e83e7fb786e86a9268d0d851113307345d797ed474071a45a4cfd82076bd4ad5859eea07f9ee5d33d464d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40a783e6ccd0c0f6ecc5a7a84d72d95ed36bfa9538b7611755ef24b0ad47fe2b48279dbbe664644c18b8af1b21cbc3a28c9cb2a0e1d07b2529d9814b35c5df27e07657bb023694fda8cf390559180bc704e9db1e369413eb5ea3d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17eb974620e35385bc3dbc95d60b2cc1c98b26613fa3b2031aead109b4015e6d81b8c136a59ba389e36a3d4a2e7272a8cf04a88f85bfa900f88b98b8ceb136119759c85ebdf7cfb30d67442ef7016da98761808a54adcbf496de327;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b6563017c0650f8cec632849c8fa70cbd2a74a36b3532bc8f02ce32c6ef54b754efcca03dbe19401f0f7b4d14f74af58a68ad260bf43f774030dff045ddc625adcb7353ddbe9c5ddbc95f24f977980ca7678d3dc6c9597a6a80ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1171d964ea5857268ae18f218260c36969023f53c0d680c4a9f689f03981bdff1b94ce2a12260306162e8064db0d45e4682010a7c93575c6d1c89283042954938a5501beeb4cd8c7a995f76d50d0178f94549d81424af7041f1dd97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c54b0981759b9b7428cef344ddb4d482b7d1bb1db80c0485baf839d8b1d874f708b72be455e6af97e6ab09e93a4fba2febe115b4da4ff2fa30c2c5c4e2b7802f7fa10de9eb4abd082fe881a9d081f9ce11bfcf67475572d02bac2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9433999f19994f2c9fd86289b98dc7e8b47840958744aebf3ef1ed98417c37d19ea1e8818e9ad60a7fbe9cad051213d3ab5428627ecfa7d0a468d7c846f3329816a9a899ccaa704291f1662785119556aa338245bec9110eaf3fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174e4035bde1cb6bc5c46eba9f5c98265f4dc3c9786f677b5c80e731e5263a4ac4effabb6b3ed134ded567d1cb04671d367f742cff8028e0d6bf5d031ebb176345374e0e94eb58e54e2636c81e467bb4da32146cc10ddcf14d0f4d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1433aff045e6fc16ecbdccdd23e7c9dfc5544fedac9989e304f2791daf6fffbc7478fe0a4354cc4b7e0f39a0d6ce8842df6c77623ab99d5ca20a2d66d1b20ee39101cf320a4e64c036bf88c78ff22ebea3e3bec8b4afa4517d58946;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79761c7528787f064da1b3cdbf21339e8d595d60f5ed95c382fb00ae85a63bda7b8a66850a0e6f57644e2b522414547b9d7bb58ca66b1db16e404166689be429eb809d7ba2b87c49df6dfdef290486d5caeb0ac3d13acdbf6fafbf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff39bd8f825c630d90f791528493d22a6ebc327e97981425746ea6633fc96aaf78f09c43e395a2dc339f08bd33d17b829eb6c79f27df5ff483b6af5db80d621a72592906158b4d42b9b9f4686130bd2bb089d31d9ba0bb5f32fd58;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb9acc9c6e77f7401721f07b8830dd890ca3f36190ab3abad58bd298c3ea70fd016341d7909e673530f22a084e1b864067b494352542d205c01468548f6ddc836083cd04ba7175f3be0ff7115389df156997a27f1dc959386cd19e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8759a218b0a75cef005d9265c0415fd199af66a6fbc2bd01c221571d5fddabf61a2f6c237440e910246295dbfe9d7daa55ced183cd57dfeee7eff6d3effee18228bd7ed2752487deb44efc7855fa786dcaf013d5c1e5e0ad4c4d84;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2df40b9d117e4f7db4bd31379b74dc396f49bdd9bd674290e0af8fe4765e39773ff6a050ee96020e87ac970604328c86a89bb28456dd6c30bf02208b58312fde0e6c28dc0eed6ab030b00426d61d7ed5e84688bfe062a9af29e66b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b319aa52588fb49389ac28685471ed612347345ea30bad01fec4a5c0b4b9f539febaaf261c386edff69ba47801c77a84e9a6d5c9df8c0bd2cca9a6681438e50e86ea6bd069b17f4cfb361ef50b9ff9efc1076b91cc9adcf8365318;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h124b7123319c57e2906d1e165c7a8a81756d39db52ec4edbe6ac5a5d64f7c5f622a548d14b8788aa52f0753a34f1af4b6d9aa4e1cbe2b11a8ea602e5caf74db026d47714f0748a452301bdc4e91abec5c7cd15f0a0763796d334aff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1760e14221a91bac4f6f84d9442aedd096d28bd711e251e3f2ae5052587c858ee64ad96c3e5c46ac727c27a9331126b86f773c71b898523d31918d5c7dbf14f38c69d1abc3ab77b509880c6eb87f67810946f3214dc65521978f178;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb8b336c9ba20d6708155e9f443e2db580c4e476672fe9c067aa1fba9ec48acddc37f56f257debb589f404818f6d714e68214e0858deb1264cd9e9423bc9be427f6aa63641c9a4bb9dc0b6e9d8b4c69e8615af52e3664f717c23cad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf44da6b22c490514ea2aba5bfd33f7bf80762f31e97330ffd7fc7430e0c167ba3cff1eef990d498a433ccfb43443d4a16a8dab43dbd81a96ee2bede070f5e7fd19fa5518b59879828e4a6d9ab032d641666fd3e9b6a6d08ccc0fea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36540a7f088a8be5ad87b662d8362a56bbd72fda4dc5b4eae7f31d2ea67d3bc16c87888ec3c921f3d83905be2fc1bb811985d4cde56ff3dae4f1a24f4ea94d2e9dba8a2ecfaee0788477f386c9bbb5cac805d33db4e49d59c0dd16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h39e95f4092630cfa93d06f23380b4f13b5988b01f3028f5ea410c6ae56ee5638360790e990e21ad170327c7f30199e305633b392e79e95049eb15a7acdc3a00d95269afdbeb6c0861c07448c4575f06d4cdaf183f7eb55db6882b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2bdd4aec0ba8c2a2d56ee54ddddfd7fbc43f5a349c4a635bd83c1b757e4e20350daf17b018de643af839079f5a155ecc21c17a5b757b6f393ebc78b81473538eac88c6577f508c879cf2e52995639f2297c2120e82f99132df80;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ed72321ebf288445c376a7febb0d99f56d43fbc7fc73d99da59cfaccf9d8be5a5cf6146a041ab9bf253cfc7300ce2728f3f8b8f961389f599ad30e3ecabd087943c5a8241e514f1d39cd3e1dc7c76c1d05d4bb4aa864126652529;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec4ee5fe203324dfdf9ccd9b6b3ed185f013ccb50951a8f3c1c52aee26816930f09c8db59bad2c4062e143d7740dedde228809d4a096939613f036e0fb5b0c03cf23296092e1a0c5e40f4ab184e6742bb043399a20e361b2e589af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb84bb3fae16373e3adbd0db1bd3375d6dbd0a8cf715065d420d990837006b4284efe595d023fcc589d7ae74b6a7f31af696817afc4a49a9364cfe7708735ce53dd421137ceb2b5a2ca51bcac312389c29cdff1fb07e62c68a88d4a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d303d89ec942450033488dfb49c4a12c1e9474abb1cb50f687307a53fff518878bc10400ba152ba0a4913ae47f5f9be76747e1370a20f5b7284a63d0a4895d7d6504d215e8a23af66c2b0bf841a94f21e7cba5bcd40c00f4aaa28;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9ae932283f5198df66e6e8d9bb1a1eb550e7c2762586ca84e6c18588e26205dbfab97426f309b09c0a9b88a51248ba2b9bdcea40ba803cbc748f654d77afa832326863937e165aaf27ae757f86b1cb7248c4392ec3499f7943249;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1acf48017a29a02534ca2d846d8599da6d22292fce98a30aede5ac537f5a857cda3e7f46cc992de12d26da2d90e00377cccc93cc538a1b72de362f6ff64c7e64fae9359362d3b280b01b1a21078046ff15ad0da4ba23f2890fbe0fe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9b4b048bdce53afe1b5dab849631aac50a74256f35828950acbc78f0aabea276ac18d2f45a32bef7a9e89d7cb84252b433b80cd6bb584043ed220808c933026824851d147217f60ebeec6e74ebdeef9904839d90fae65d81f70ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1d3076dd848c97b01b6432715f7cc4ad8ac9b2c3ceda83d37bf857d7dba3a1248e7c63393855647c0c6291460b81c4e4e62dd808fea3521d7ddfb2eb2e439969953da17fbb6f4586ff51e5b40ac99e2a31b3174fa6e78a175809;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1f0647f85080e7cb0b8eebfe2ce5c7900dcd6dc83d18e21be8f40ba6451f9edd25ac92cd38d8c699917898b81b4d117b3a61776644035de38bae6009454a5d5d49741196e829cdcccfae8ce15c06ae616b9dd0dfb91c1726e81a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a873a5486ed8dcfd3e1a8f7c2424221fe4a2dba9d6ade6f4fe7598b7aae84bce7de95bd3785c841ec954b152b0f3d84d7934135b2f10850db161ec44222201ba27efe167475a5c47ab1dd5fdff30c9faa4edb28d0920bf1a10fe68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e43b56623e2801d4665695dd8cbeb8d4fa48372e827372b1133c70d45bbdb51b823661cbee09d430cc249affcb9706221225c61599cc77a9478078d3e5ce34946c3ea77b1805c121b2631809c590a6546077804a6d8552b85bc1ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4f5f165ee9a2b18a05966304d085809493457c7dce817a752eef3d0852b35f6e4018af20770245d907a2871f46e5edf54a77985eb6b07e7e9d915316f03118c66e819379802c7f10d36eb5187ff9b1ffaf7b87d387edfd25ac047;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c06f185332b2a2cc1724951b7efd5ee4913d3205e95cbeb2899993df7d8af1bb93e1eb4fb7e0a080b776b0348621624f8e81f8b60a1107bc90a9b4b9b2260bce0adf66baebb024ba822d075133f81d8ec3f40786fcdc367487df8e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d3facf2227684472f2dde18fab85a80234a18fec173d89fa68a37e13eabb1bda90990e879a265b08af83efa3f45c53c839f633777a66e20aab1c579b4cf2c20f77781a71f4aebc3dfebfcf18a33776f57b16cec55c70d16784997;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11501a60f6a5af197b908aa495642517cf30573d62583019f60ed57c08ceb8c0c9cd282897f351f8be8b57ecb08d57a79fb10a0a0f98846683ad41daa4d413dc2337e24024c8fed92a04566c3713942d13bbfeec9a4ae6210685900;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a0ec7f0e75d592f7f296379f9d3c6e49bc5b816008c7fc23c869c1fe482a98482a5d0e74d7759e3f3543354538780f374d3b2a12cc8695311395175c477af5b55dccb5997be156bba155b960456d203b086f8d10c5c44573b09d9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d5dbe3e5cc97c210cf3111da46f8db4eeb0b5fe816750306595a8b3b8c5d1183dce3be133f8ca092458d16fde481bd0b15f14f79bfb1bcf3f5cc7395443bc628e6dc2e10a61b6eb06eca477c598e42fe1441edf64afea71ae3914;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15dba2c54929d86f3102776c393ae456cc259c02fa293459501ad06386f0c9f5fd957237520fe37d16f6ad5a3bffb80ae05cd06bf8b8209659962d442da46be7d0fdfcf433af5b2ac8a755ce93443ef0dabcd36d3bbb5fab93c2d23;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aaab33bd67cedf5a62fee13a2b0382db8dd7df97917874617166f285290c4f51ef4e79a5923e6b7f5a85d42de1c712dc3e1e35af9bb0a19f66c85af34e0159c4fce64782e06fea00717df4a17246b18571862fb7af05c6b450108b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1450d7adb43fc2a2dbd4ab6ed8d9a4dc4d00cbfffc37ad0837077b5fcff6761d943c38cd59a6758644fd0ddd876a6d2281d71121dd83e3a091a23c41ea7a5aff5cdd2189aeb95eb38381b541aa81aabf68965cf20a6b6f054527109;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd09b33b6b06de1fdfc060b84bbe7c7d936053e2253b20026d52040e0bcd98d5b695b1b59031f2e1b1c0b86137b5e38ce7a207cc87b36ab732f1e5c6ae8e5bd681a8475bec90aa3f03cf78973ee44070c6c7eb327218048953ad2b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ba5b99252d40471904b1cd7538ebe482b8cf674e367d0140a2b34a6f20f88a7be835039ce2911ab516c22a91290e2b6b7b271ca587892f1183332b14eab90ef5697cdf51ce287dda6a0ea2205fbb5123aec6a3379dc8f68c0878f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0622b6139919308043dd71bdc594f7de236f634a971b8be08727c8703c7c25a15e86dc127bbbbf348ff56169d0c75c33cbfe02a745a220b94d17e5df96a73ca3a642dc3578b98ee94a1c3953c8fab1b6942f525d17627643cb6b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114e7fa73eed7779e578cd01690d15d2a99ee06873191f4a292ff7c02f332c0126dced6ab84956578010c005b7d37cd8acaf41b0c6f7cd0a3a14eff9d3ec7c98efb2cda3a3f194c418686a7ffe64d00bd7a0fa58f041605d34e4e23;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14846bfa1d9daa09b65193307ec43eec54f7eb3c65abcdebeec9695a463b58dae877295c59d5a3db6a3e69ee6a14cbca01452265ea63241c9e0172030ca1b64c609b53d7e2237e82bb3bda60264a11fc8ded6c1eb6e0eb4644c71b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff5304468126607c219d614654cb8546fca234541f96b83a8d96c55f410f4e02782debe152338b2eaa8ff0655efb216f477e64b724a5f7cd9800ba7a00b6a358e32cbe9e4a22b473052dec77733cdedaf7256445698fcbea56e1b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80aab09a7e0af216415c4b9fb613ec86a2851991e38fc3b182cf1888bfc2a9898c5c5c320a5968e40eb6c12cc1326cc9ccdacbc5bbd016df2301d57fa1950b8313dbc949936b0afa37022ac871b53293f342a098bfaf6452fb6683;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1ba963fda18f224b863af46aeecc185e2de40c2bccafefa263da45c8e5ad2f3c8c28bf7a3dfa0c0daf9ff713eccd12912ee855aa753aecc9189a409954038e9092416a0a3ae3d0448a550711e8047909bc7b3b435d032721302a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148002924da3c377b45713c1923244714906d6faff9b2d79b1a4351452e24920e246761037c6b5aef6c59d79eb4b6dcd7e4a2981f4a81ebb59474d10caf88463baaabc2cb5e72e743129e817d883372e5448080488fc17db06fb008;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9be3fecfd6ffdf7c87129f9f5604e0cc7e034969c8e74713ac538e0c06635fea7dd6a9757ff5d7376e9e499e419106e7bdb1341df3f261fad90d51ecb84f54ccd206c9631459b941762a90a59809b398dea37ec30eb13e488ecd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a78c84fa0daa8fa1c03659d984a30afa32a8dda2e7e60de6b35a2b42ef51b227b7ae670af37107aaf6d18e17404591e066108a2079ca36011afa061e556789880893c430b01d72e9cd80f561a9f210d440777dfc6eaf87c048e941;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda6882574f1fc6dc257102623833e4a1b3ce86c579e672dfcd1fede406dc79c168c0d7765ce56d920f9c8ded1588df4707e8d7d6e8cdefbfcf92abcf60c002b3ed5bb6ac51ad8128c77ca906bb8a3f480a37bb50ed3148843a32de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a63b88998b185ab6d0bf40bd2f546fa77c7b3ccf8eca9831469cbd33367eeb702c32471c0695516641f3b56fa7810afd5aabccbcb8150284d38ac339f743ad6bfe6917eef9c74463e82818ca1b423039ae7bfbb2079d13cf8837b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f789115f852dec724f6741e683da8b2f2e92bdda3a6737b948288815070ea36c35f346a99f36c95d7af6ac02bff3d794c3be185a6283479535dd4b0777ed9110a0c8747bb7cab3122be446f69166306979cff4723ee1f8e92ac5a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143ccde8c55eb1bbdcd29a64b950bf03a32d199d25b68f557b5f7d16d89ce07f864f01d49cf7c768f0c471dc93d9ccf51abf6a0fbd47b73e6bfc5b7c6dbca6faded5a59c2e444c9c56827e77639cfffa3365e478983e112f6701d38;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1260f06aa03beb4f6811eacb204b9e2778418c78da6d5849d5adba427279155f3e5ba9dbd6e534e0c77240f450e6d482c803001e40137549d355b21a7e15538c530aa4f6cda1f44f86e6258a32f9ae3b38b640e1ee3c0b646fe99d0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1377c529fa8a5c991f3ac3dfacbedcb9d2f68586cb02eea363bf4f26f665e1b2475cc0fb8db5a669e78e4055c30d9c588a336fd12bf362ac7349fcfd427b1bda0b8af4135658af980c60f7f35782df10e32d95e8bb47b190612448a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cb453816dcaa44da6647c82b46948929facb87e591028f444a250f5b9a32e99b8f36a138554ba2543bd1b6f0b8fc6459cd806bfdaa9e5def572360796d61be578d78c597017c16533a1f4dcaa800ec9a01bc58f1d31c2f1c65b6d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6a53712aa7bcb64c303f8c4eccc2af82c106dea48cbeb9cb1ad39bd45c10d2c74536cb4d40e0f49591abe66e76e91a5a286f6421eb960ecb7b660098650bb253c1907d01d56808b4dbc338d8f05ea057a032d1de8e483235db5ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168776e78e3e4473b4a1c0b5ab81ed5f98de0613623aa208936dd425ea6c04d11439742d89f702b00e9a98df6b4704765e4b0112d6f34a395ed77faf86c227fbc75bbcaad8439b7cac5e7c675913dd4816612632066bf282fc11735;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c58563cb70f5e452ea3ea702215b51f63562d3efd332e8f197d89e5af358a7ac75b92b5cac1242c95fd88b3b8387cf34e102a9fe1fab9ea756fb694d52dcd34be36728c91185603be1b1149d8977ed0750f99acff90eb9fce50d6c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4e9265b42acc0fccd11a69d8db2a04019fe50906a0a1e039149fdf1a19c9ef3402a8a08584e48b10953fb91a3bba3f63f84d91efa8ae08be4d7d09ced9e48abe18b5540c39c4e26f50f37ad725f9dbcf87404379c4a20b09032be;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87c146c01600d806f8b4b11158fb776129f5d40b3e4ebf27f5155c7612ee4f6095ee9fdfe7ff19fe748e8c01f69c3d3bdf9182c02b44a8125870a0dd089fbf9b328767edab4fc2b678688010a4c259a7b71a747efa899d2291037;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d157e128f95eac65012ceb1ab5cd2c10cc47fca74cb6df356cf79aed29987284247e122b526530c61f644cd96a8ecf1608993f4eb36094292dc8eb19c3d920bdcce6733b061bf76d994206dd5b00f988aba118453d827345955c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d544a4b95eed8b3e9bf567f03d4aa24cd4af3cbef14637fd0d544abcb4dfbccf7ae67f57ebf69c14aede4cb5bc01b194486fd86666c3a7ce29e0dc43654d1dcf6113cccb2f4097fa27fed73731b68b314c5df9e29ec9e41b10e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3fdf7d9fb1f55371cb045293a25d55cb4819d23296c48fca8bc53759ecf0810cd87d3531fb47acec09443fd3be6684986d5a2975d3a562d2adbecad9d0274ffb1479b5d0c44d503ec9f9eb95b41f1bdd60ad6b9ecaf48cdfed3ba7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he81ed7ca3f1885a276535233ad707f98f02a4713aaaa659cdd2487a51c2ffba330e98d658dfef250b37549df4d255675ff9c319c7dd06c29a693c683eb2aef3f3ae882d0b759f25de2d29341627920014c9166b8a24cac3f8e52b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136b07f1f231905b2c04e76aee277e34b6bb2eab7eedb8d0389eea1ebcc62f0afb16fd5ce16958002c4941415f627496ae78028f499c72eb498971694fd46bde30e9c991349601340a18720be2b077e26bdfdb02481f0c95e0d5712;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a25f53a6708cb37d25d4e13879bd5ac5e05b687b97f75efa324579bb34ee74fe20974340f0dd6086ef04dc0530d5423856c76f9f2e8ed14877212449c9e64acd54074cb02b890f83ce1b80729fb83e5c579420c99ae8160aa3738;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa16c097ffd16cddd6894f1032021b46325b4a330c2d89b6f20fe5b69d57997483b200c29b1a0e66457097e6e6001b9f952ba73c3a5dc7f427b42994b0b4a9b85a1713a0c0ba1488a3a576eb86c2eaef19c2a0f615bd8c32d59525;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4847ecac198692e04770f78230905188cd22f71f1faa6c5db1993b0b6607715ea1fe70f289c72eed3db94fe2f6a85a7505f87a5374dccc05c7142ceae257bc357fc695c03aedb8f2b289d93c0c8994db39e236426735064e5c6bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b592b860ea52e725899924c317e2cfef72f68d16bd9de7eecd342446f27387fb2bd406ed93c9ea0a0a659021084941124d12c243db1f747ce103e1951b73738ffaa176a8a06d973ce12df2ea3d55966b4118ffb39dc4f745f0e230;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5b9891bd6b90be1a8fe87f86972e44d08c1415085eac823b768ceb4d8c94a801a7b7a7aad02e034c7ca7d63c09c843205a20b67fdf674e34f3fda44a7e7e2f03f11bcad54ea8dcc557f8976d641f4b679294288e59241decef82f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h572e5c137ba18d3ccbcdafae0794204358da96fbe3a719d5068ce44041943fc1abf7d8fda11a05091a36b5c8632b23fe6d6fec6203b141c1db3ad79688146f6d56ce1f35c907d91b8a310ef84521a8f83fc14c4b1b16c5b48d3aba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144e9fe9bca930dcf8975617ef5e5a9782b71a1ec8b73a3d36b61be748d6914ade669141f55e532898e10d22f9e8d277683ade6255e03fa172b0b3bef65e5264f5ca4ab6a07642d7c25b7445f5b1011fb6aeff0ab4921a0db8197e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab44c2f49e06ff28946ea2789b276e7ed7fd97c7d2b821a7244fd4ff4b3f00db5e0d5a90590fea344adbeb70c55ba0389e36a5576b4ef89220de854dae2f5880171bc7fa975218b09ebcadbadd8a55afaa0745934e7bbcf27f4554;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ed282b2dfc5c6a1935968d7f576c59777c233bd3b11040dd00700ab5c998726fdffa4d40c19af80fa3780ef43cff435041b447ca5db0af42eb9217186f3dde79d41ff1d6071648287cd6f2eef083dc078366771874f6c0ffed620;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b06a762b6cb449fe914f232b3b13498b66a67070f91ed3cae64477bb83cfb54ca2cc604c0f6cb52c3d14a23f2f7c3b2a418a4f78509f1d7d3040e60a4c43744a38ced382f300553b0d7b548ca7ecc613ab82c2a6f3327fb39dc4dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b06aae53cb34e488f4e4876511dddae1b9737db596ba1d8861ddd2559072b5bf4b456d8e860408a1bb323c541567256f830e7a75d7efcf3b2debb616ec7adc7ce7a280315b2fa5b4c407f7ac2981b869dd16346255b7b4842f409;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5902980694489661c1f730af2d921675f182f9c735458c49300d67fbd13ef0c6e65189c96b28811bb8fe67dcbac1f034b404bfd4a9e1e5b688d939e348a826819ec867c2083cc4e0775d4da4a3bbc5bab5fdbed23dfb23ffc14b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d25b07beeea998fefde328a4cab76a238d4b727afb4e4c0d8526beafa7f97b92e31c50acdadfdcabefb7543b7032d3da4a0c4055c06efc5a630559d95688e941bf5a05a8a45d53e02393548da580954a5dd9c18e10a00df2ed54c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf11ffd8b6ed172642131750c5e168a9852787aa05f1e548a531ea7ad59eb6072998d0b8107e224c82a0069c340a16e5456423d8c6c583759fe76745249bd430fee286063b8263c78847f24d2c06e13da20a133b940a2013f455698;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160643e149869a45389aa3b28913ac9ad8a47e7b318bce351e58d2609c4be0c836027b9a1430eae4d376af7453127eb7326e4e4d88fbb6c6b7ee3935d460f7b20ea9da5d5d8ae5cc2fc93c5290f47842c9bcd4d8425b6882172d874;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2b1f7fb7b5b8cd9ae1b9520c15003518bf55d14cc9e0f5cd5f65cfc05a0ae29815685101bcf2a5989b1eb8e649227130bc12cd8d53bbe0a70138b66515f0b79baf160a7cdb8294afb99340c6dd42a83f81633fdc5ea43a2703a287;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2b3b1d7a808d16495f2b7d83addf8f25be53a4f0f272986650967ad0a4211d5bcafdbc49cf9c17739cd3534977e3a3fe06d681f3dbbebc401d179b828f4ceb5776e107c3d034a8aa3c28204a9cd161ab7d7034894784f7fcc4ddbb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h349d9ab3604353cf0ac9b6be6c82618008a51dc297eade176936a4de8da928b405a9c4a1fb503112fcd8973b6fe31b2cadefebf84ed20e4450f2880b31adb4a2dc3566dfeb34df75122748b076f8a632acc16fed78df85ad59018c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16cce0d86022416dbd0a0ad32f91b41b961fe4b461c957bf6eb1cf300d8f7f0fac4b78033bae989e573c0a0618a91d9199398522112408cf2dc16899e44d96f59313285d6e0e9f25af60cb5b22c9c5bb6909f47b4043607ffb0a05d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd28c4e4dbd393f53948169c66bfbf786616da8413179a5dc3a54c85d07ecf39a8215d6f3e2078544db61a1beaa79ce35d1ac5b3948637311e5d7c926c8f19386aa134422d4251cd39e54e8e697a4061bec5d32e249aab3165e883a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h425b8af8fa6b8469177beaccce07edef1b1d9152dcf6b1f8f36887a882295ebabfc57f5bcf81261642fd6309a7cb97d30ab3a6167cc704e6c9de6e770011f9fa0119d102e4e8f34508c68b14b15c921082fba79b331bd957f54042;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e30257f98899fb161a87a56a763628b693f49f066ee3ff1b16708aa2b046d95a40631c468e610a36b0d32d64ef7613893113cd4d9a079aff311ef4039b6c98e10e0fd11c41b9fbe926c0baac293f700c246ff6c192194f7571f61a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b51410e6aa66be1da1c4b9e750ab5a39d988fe0fded358b4c59521edafdc8d2ba4f23418e6e2c29c0f4c6273add4402d4f0ceba69fb503cd83e17fe65c4c08e426544619293ea9fd08239440459512afc6b822079d49b480a26dec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab30afb6b7e2aa6561fc42acfcfcba345853bca574c59aa9150fafd2beb758f2b3743cf31388dfc940f15fa6ff8853eba8f1792a6f703f9e3c9b1a7257147a2b58a6342ff55f89a513d74f6863ad5573b1dcf3d4302171985ac968;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177d08cdc01eb0e942385a5ae06b4b5daf26f791542e49bdabf16061283613d11722ca7a3df814277a0f7d74867e6cf7738d93fa2d8fddc1f309b7705340b1a935321f9b49bcaf979af4d5fa3a3c1bd0465ef23d0968d0aae340019;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h918710407132592642836c654f8acb9ffe4a9769fce3116fdc80d4e6d60b52b590280ac4843e301ab89784cb2278ac62116c4197941b2b7b9be670ecfb849e9e9d6d39f2e2885a269ceb72b64590a1f96db55d82f888b7175b1b86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha09e66d8390d2e4b09d081e6941afa63970385d0dff2f28f9cfa4b38a3418eff76f3f0d566f669f789b7156919fddf98f3f5ece2ba7f7ef831666114dadb7bf75903d448038ea778932edd4f683a80baaeaaad4091a2a4d233cc6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b7393e7888794494ce04faf1b2c97464385ad6b221602c3eb6a6e7da0dc5301ac05f46f9059959e8df71705d6b2d535d06da2ccf04b883f9e54a87979be8c989d7838911e3c7d35dc96fdb0a43a09936f03991ca6d90904f2a96f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8e3cfd3decca21d22b5360acf4328899337afaa9633dff1f22785c99d1e7dfe6e076443928f9f0fbf668815fd71c13803d2e4d2e9f1907499ff5b503205c081c1b08fb82eaf18739402dda929c4592225d596bd5c5b8ddc327604;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7126a876ff3465a93519ad3e4bb8d82df2d133eae407217e757472b327a54cf41b5532c7889dff3d0afc1d183e22aea2509772e7b9e19cc1d31b118f7f0cc4211f00b2cdf6be0139a39edefc511091dd3061ceb2e0e4c009cb4ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123191963abae05615220a4a48039bf83c2253656894de888ef26aee6fe1dfffab40424d60e71cf148198d07f6eeea22916866edb9e8faa844572ff665cf310f540acd6fae12386ce4cc6afab232db78ae8edcba44b3abc13756cc0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5426deb5a8bcb7a592dcb86bc7bc75d12cfb9fdf8fcc2fc2547c80e0e7e98728a1b38abc85bd394bdc2a8b42a05f4f5cd9295107c4508c8b74ffe4615f69d08d0c8aadf45f55a3826813e453c2ad56c9e530959810f0fbf887f85;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2de259dfa0cbd89c7a98a8c784707e7b7bed6bde871177b9eacda49c004f4963acf380a3d4c38fcf4db6c5ee6808549bf4f3ab4731b1cd9207791f5cbab7c7ed818a2dad97b3157d4e1b91066583f25488269f5022fbded78cee0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa01f672d6d7f932456ac4c025dd3f16fda2ab713908157d66cdae41e84c299c61aabab19804b961d19ed6f2f48b73ab03e4a4f6ca9040172f696145c4850f6cab1169800716ffd229b73f10dfb646ed0b8955fb98f4ad203e79e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c537257ba9d18cb3d7077ff42c1762d6ad993b966e241d405be562a9475edae58770a145a35820a02b5b77c0838fc7cf1a6640052fe1757a4ea26c04e4171020e1b7b5427f63e7d12b9565a2b79f6cb09b29ef896abd4369a428b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf1fd6dedb546c45a10bd12cb2d22ae29ba569fd43fb917d1e9c3f18d8a654db30f4ff1df942c1cc10313f1dad56d67936ea140bc74dd3e73633df63cdd1c95da1387c1a4af53c409c9d39fb6681421f599d79ca4d8b185706ab50;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec6759d5374f35b0e05f97949f9a95a00509fe7225935e586776592e66724205377b51ac807b88b2f0422f0cbc123da09ceaf5b1c066341779714e27c22a1d4fede1b07a489cafbea797e69a5ecc0182281858cb142d3e6540684c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1fb3bfbaa1d6f797de113c7db841f1cf31c06b79062a6f4cced9dd54141a0bfca5025fae9bb2153ed694ec07c6d6dc7b560c6017f2a93bac6ed81644d95400f5e3f9b05f0f080211190f463ab0802b322355ebed1ba7e2c5bb3cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d8bdc49e9b7158644f8ba005192e05a11c3e237d43b791446d6ef9226c955807ca71785628dc598533357cb5a8db047c26e0b7143d2bdb8f7b2d28ba3c1a7d358c0b4a02b1668f0148ffe60cced58bbf614cb3987ec000577265a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3c8787d73175b490187016ab6245b10dd7d260496d9d7b30694b247c8b7f211d16248b9a81037e6b2bd91309e3e0bb3fb6cfb5470c512d4dcf852948764758352cc64eab207870fc633367c177f622866e876cc77a49653de52e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc924f313c3828dc0bacd89b21eb07b2228af62c3f095ebf52a3ce92028d9cd10e641cabd9955aec78a30263c8ff3780dc69d38167752ce9e782dea4694e26c1565a7cfb26bbc7666d210fdae1f685e508cd13c0f95662b14dc49e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b306d1d4abd977efd3f340696713b5470e45ce7e946199895b4a3ee4d3f3e3608b1567127380967fb659bbc3f3b73b9f4eba209274974a00b298a000ee0faa660a5a3cf787689481c65599c782f07487d234b08c8f155a9b3074a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95600ae701ff0c88b8a86383f01c99d70a280d469c8e5e40916e5280864a607230cc4345ddd8fd75a88228dadadd043a83c18c83fc42aa90db49d868226e98be321ba19089a2a02784a91138f792b778d6b137bb0df5d72869a477;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef985bb69bcec3cf1656cffccf98bdeb0172175a462e0f1098f704d45e5aad67074a3a98b51796261aaff6b39184aab09c9a0036bc51120672c7d6b376e453e4f3e8f8b6a12e5781a5954ce6aa234f7e3c7868a9014281eebb8094;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc9fac97f11ad664792fd00a3f7725f515641c41c59fe2f30d75d04e54c27a171619422362321c1f898a2357f6201eb120a82de77d73025b3803477a5a034e86965f01cb37742bdd0a5cc370e835bfd9a997a7ef6167a81a7756e8a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87cffd27f0517219db047659c17faf99372ce3a232b2ea7d0ab1db10e8c830368a91532b73236ca413a505875417890331dfe21e93ceb9808e45a3549599e8394a12e605163f3a6caf2efce1a7a2eaa0b623ac3dae3863f7d8a65c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e7c0f8174c596b3d7e74abd03297165afbe2103594b1fda3ace10e21dd4a884aca96c37cef4347cdcb971f64ecaa8eb6ddd70d722c71f78663900037da75df18f283a5c59cde6e2819b635c38996665ac6b1b402ca12af606c0f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h726214c783c4db4e39684cddc9ac951d0fb40f4b922d32ddcfeaa17a632f6baf49c58410cc599b7afe0d08d36ce2a19ea7d8074c68727dfe556eb1ff2719983f6265e3ed826a9aed5dc4682b72a8cf50c852c5fbeb5ed0c1d19cf6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed907eecc4ce7b08a334703c2df5bec3d7f1e47e8657961ffceb143ad0d5e11dd14fe18d06d6302ecd75e10bf25c3e2ca52f08a7b8c07a87d7a076d8fc4df1cd7d147e001462f8a57cf793d3fcccb0e26a43d5cd3f25adb36e4ef2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0015be9ab916345150b5055220defa1d309e58a6be3cf55368bcfb27144344514417916aef1e7b6f97f2f7458d54e2c6e3fedbcb711b0f1621490f7dd7de2ae7c2a97ea21afc004ab8ded434ddd65ccf6930eac1781633132d6fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd17b2c2a78b52e248fc978fc28554a6daa42b9ae9984b3fc552d7958d7d80da818bd474b51eafd6b59c70135f91f0fa6aa85eb493aaac9cb0298924272c6e4276eef15218e102c5f1ba5b12ef1c315085d565d37fd8b722025ed6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd183ef1db4b435f0e86af3e3d04427d048264197a6ba4898cd26d613ac2b4806934368127fc8b78a7b6d3918ed70ba03576005eb6f678984d63e1c7b4e12e4b0fe8c326d27560da99505cb09f24e1e17e8457e8ff46592e145a2a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33ea53214a708170489f163c2c7b18164a6d7cfbb9d5c702930694763543c8e2e2b6e4b668a94725b6818eefb95d2acfe450b04d6cd1cb91fdb195133491044d5734f1a02fa694a181c4d9efd32c6da2ad7ae165bc7a688006937f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h118814bdf1d42d18449b15aad1b3363e80833c878d69f925d7299a38126051cad5d6ab30e43d26a06cd2577cff889f5ced6aba1818faa1684c6cae8152e3dac038865dbd019f3bddf7e38e49367f8e395e89d4d2877813e011bd4d9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee018e48169038efe251c3094c0b763514c0804b8c748a2410cdd5af2ff1f8f3833c583479aaec0a4bf80474c441dd9d21c62fdada4c1fbd8130c3efb580cb17382502b2d6eedaed4948cfa59a64c41cb5acf2a43af0cda7c81e15;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b424b3b0d483a924bb320da78ade33bebfa6230088637221c8ffb919fc612491ada9ee567f77ff3ecdedfb7e633f8d6ebb39024ae1aca836da3f9dd51823e5fbe660cb25e25c7994030d5d2b443f883cc1bda8012a20c00df839b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1160392717f8e3073389a17793f43971a62e624c5f91b2d7559082cbb6434c82685fba3ba9d7b983b64ffd553d0d002b2d37a0f7c558f7cd38bd8634909b1daafb7d2eb3d9748871d9efa3631543fbb72c76a385f62bd4b1cbfd829;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d92b0ecfa31665b231ce3e32cf01c5ab77540f4ec8586ee89f7fc19e983c22b9c55fc74dc50cfb1b475975eb5f8035aae1b515be46ab076e31467ad05e7503e116e7f12f26739c85db631e31fe053659c525c416de767115aec2d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47c563c7afdb94c2a53783612c561e4cbd1b4e9cbbb03afefa1617d2694abe941a437130c4e24d9e63e4cfd904da90138148c1a4e3afb26cae449a096b4d796a62f8d51cdb9d43661547deb38797e53e0ebc6f3348755383dd289e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de92b79754519572b7cfefc013bd2e4d34789078050768ee06fa7049cb14282175aaa53e1366c03375e9eeb299cf1f3a07e50bb4ebac91108b6f22369f7c4fb5ca0c599a4cd7062bcd83ae41c9958c5b4fe88d0348cedbfa9a759;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f83dd20b2db16f15ea14b344d91e7d80fec564fa4f6d69153fdfa5828a15d7a1b0a12875bba4cbcf56dec69677f9e9112b02013610c33c125ed626f020c6780741747318fd3b11e71205d123e9ff34dc35f5edc1fadb602bd2adf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce35291e90a5827f1f945c870db3e03db9335ada57d57fc416b3187009f998347ed786211bda4945431f1821096bfd5770d2a291a093c378595f11e3f13823cdd58d22933071c922cd4ac2b5bf7e7b60e1be10b942fa26cd61fa07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ed0993e34d48269c88f1bccb4c5953e6bce0c9fb0ff04fb43ec219769629fd86d92d1ac17126fa4bd41b8700c5d03c5ed5da597c742de500dc259cb01780bedb5df5cbe44488d4a872651c203e1f1d9f61a8a86d7f6d867545dda;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1971be48b6ec4e4ead5fd6ac823a717a56104341052acf96ee3667f18b3d7e863f544e9533e9aef46fafde1b5c8624902dc307ba219378f0d1b515220221247c8408fcd6627e56824e3a340be0458fbd2be48cc5f178a73a1caf918;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63854d769aad8d06b43f3481c69c757e065a8a3cc62ff8f0d8012395c8621ea2e47e7fcf6ff2c1eccf38f36c380ea0cc9d68315f9918ae4af4b014a20cfee3608d24f91f82e73ffad0c01a5b82e2ddf6dfd89a9499d5fe9fdc5b0c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h45800ffffb2a466ae90ae9fcb396cb21f01476e23f94a0ed3e64e33395203048a9684f7c08b306a24e4dae836559f77807a4218e09ec153de9c7f0348c303f1887b9f2934283325a589510446e2ea291ed8b7dad7c90d73c76381e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158fd134ed2ce1dfc21d6982e3b06ff1971f317c74314b1e1a6d5688cc95af234316ebfddb36221fdd10a69626fc2c927a8337bd6755216b6d67718b87139675ed888a6fa0b08e458b02db138d6be6280c45b0cb2a40a934867d715;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdeeb1eca89ec8b281f3852066e4f433221e105cc61ab95b0ae6a286a4ac5fa8abffb36803fea2907afd50f3da05980596e9be947efe5b914eb761d1c2151fd5f947696336ef4d8497477812452249d2f54ddd5d8467558525c85e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148e71b6fdb8d23f8c3eeb36b91b5cdc6bb654c57f9166cc9230f70045830e84f49480662e524a89c5c8f0834f27e1778aa514cc6ccf3c1cbf24c1fb8340de3e66feb529a4c85fae4405bb3bed650f10e26e8338ba118c540e61688;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6039fe861da8c8f03b038e82aaaa1d7c8bcda35b7f951e554df600c6fbbb5cda1086efb492d2e327744983af25e626d693380c0c0baa2c05fc3ec0795ac67721d0a86fc607309ee00347988c916eeaf9187a1d19843ecdd71ff2c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2a6650ae6d2d956d06c6398bd5573b115a5e87c261c67adff28d7bf3d328653d0aaa4669f46abdf1d02bbade7c896be8049a33c938377b0a319962d4ab232888956aa748c4486cee8c503ac03b3d44354e924c7040437d7696384d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f33ae8f5a7ac65f409709b8bd8aefa36ec025e66de8076d56c79232ec0820d0bb5c719e6c1d7709b54b08dee9b4de862dede600ac8d1163e79ad63d240c5a3e7114cc7829c3927eb27b64db55f7222894cf6af804b0d0749f9a7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b16128fde15825a212b9c4e0542beb104e34939816a3aefed1c9e75f6831351218fd106d865270e45a360201d3d669c0ef7452d63f2d9047939dd788de06e9d26e08f71bb66f54b958a62adfacd9b64e5a0983c08d31c39c40abb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1514255629e7a7ca4c1e65a0b248bdd7c903e0b4e30afb30e20844b4051063ecea54ef2523c5e90e0c6338b87d8edd1146b7bc8db4d167553a0e191a953fb3f483d2b88cbb6073b1c36a090e1d71f6ce6d625a308ea14738f9f21d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7dbd0ac2f3b06a8425da1f7a2da3dbf3c2ac918e9d77bd299b525e93fcc031521d30c2323c380863105b85bee668133dd6e42a333082551953de0ed95b3456778d1d2f2195418704b847c3641f1a83c56e199d8cbba2d585600e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106c5cd224727e0d3014da86f5128f064ab5cbb1280a24210afba3e315ad76b3e520dc702d014af12e06cc2d30f796d6b5a6f220df7dc3f4989a162c133194b0fd4c2c321587aaa39fb6f90c742fab931ee38946062c400cf0ce723;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7fd990f8432ac438a2ed7260919227702ae41a8840db536d2f02f6681ad0b7a94d8161064a8da87ea7794fc8642917cd414b79c1ea1754193a72cd9a9c098a74500546397abdef69523b256896976448469799c4144e1c2dd6149;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa0370539be1b94dac608dc7c82a5ee94e3c329b5dd618a5a26f1f914c0307402fc7b1a1089191a030339b86e9b5d4b5c22dc03dc53be21de8942674108e3eed04ed02586eb09ccdc393fdab6020214e866f05655754f6829442ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b96af0b1e147afe2ed9bd90c73a88a05e2eda219b667ec5ce2bbf90fb2f971b14284aad50537edb5a0cdbbcfcdf37e9f3d522255dda1e07a47a1b4c19f300c9d39f5a180b426cb86723ae366eda0a880c3c5258c6e085a80030e4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2755e8d586c9845d92506244568b2aca5b11b7cf8e35ad6eefa943d5a9bd805530567b0c827e2475757a3f612ed79717c80ed8169c19c840000447fc315457e41e8a37a301856f1068ae6742de4154d1c67173000ff02566165a25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8872c40f3aa92c5b05ade71762af81be023122f56afc1bd1c677ec00fac5f8f1e05512fec7186e78748e07b9c5e7c056b9cbec46c6efa48b3135330d6016329d274f87ae67ca943c25f26893e88ab55a214c6b0ad3a01c5e42258c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha0481a59e77b025c537f161868f9b0fe791c5e4aac4fd40c4ddbc75250b6cb8215fa9b434ef4603ed0cab1523a13bf25bd017685c0d6e39c54c9b47c311d1f0608f87080e7aaa4e7f12e7e7a48b893bbb458fb73646fc53715b97b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa4d3969793754b5776a4374c9bdf6827d536d90d3061d9b7d067947715c2d4511cdc105190860483495a9824c98537f93bf887875fde69727eca638a8b6f9291071c3f9c98e1e96f4f3bca1686ad3123cc9ce61ce1ae2018835cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6afffead907fbcfe3af2c6df764f5445483e72d1a5d4a57375d80ae439d53fecd2869bf895b8455a5665a830416221d1dd46c83603a9847fc24649af29c1ad54a89e5b5632d6928ae4640353f8a9a92ac7e1f60e8b02cdd2372f80;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he38beb75137682c06c66bf5145854957c3af2aebc0efe65c15e194881f700e7e4d047ec234ac6c6ba6f59ed04507ba25e1de58d5df6a6db24658dfd7e532bf4db116f211b24616a681d305fe07f7dc8f4a65f9d5c7e9a792cd9e1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc217653ab306455f413c42810613cb919849eed03c4a3c58e1ab457fa78212d7a4cc3603115319ade70cbed6e6ae9e4f7275b04168e9fb4213279a59552c9b8d99da1a392db093b873b3622fc3b7a35b0faca0d16e2ed722b6ac8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2bfbff00ed99a3a6669e570ca15049d2d83b33ebc19d46be0fbebfe1222b2b18412cd4ee2380ff59471ac901ffc2168f45d6d498f0af31e1733309d3a74077d73f25e98a6cf8106ba44b998194dcd6bf361104235efab23e98511;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197083e4e3d767e5f825a76bc4c4c237d142d19e8fed5a20cbd12cc9432aa38c706b3e70159dd8d1e41c6a0e5a07839ab97ae72941b2f2e27b39478ba7ab15faa2e499bda0937f358fff77ca6864451a565701b74108f01f4ea9e24;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18777179870ac39146f311e3fb09cdc6aaf610781816154d851dd51937e5d52e54125216b3b6af0546226e3d57c96746ef4719aa06046d10a3593ea441eba2723a9a7d26403bf8f87a8132f9f5415621cfdb52158297451001f1d74;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173f886c4104e6385f3a5d5bddc47e89ab0582195049a47c79d13a9029f4871464f977483275167e728508b5deb7975d358ff6677d0ce2a8f3da0d3ea91c7c913001b9d73cc9340f897fa2a5ce295a274b7620ca67cccf95c19e921;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb008e66a5166bb9da9931f37e319be38dd2452fabc3b06273048e23c93f4fd727647408182824f69108c440b2a3ebffc590e305892abbcd1b8f16835f83721cfd74f45345474829424db631d3aec75d7bdce68683b57c0b3f93874;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1add4e6e37b6535c6036ecc8fd4ec2ed87fd79ac7b1a56d5f4a4f7e2acb473f8b97751180586970278bbb9491ef77c969ee5cf49e92bc3c38520510a65b85b34a0fec8ec72cddbb08dbe674407c8175ca29f2d0d7f4ed4fb8dd355b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5684459fc3c586d90be93517f1b88ca79ed1cbddbf84fc0b09dc2a2183edca73e0fcb62cef41c0ef884e47edcc44c780b2281f07bf9f0127375a3c524dad1c059e169b031109d741536dc009b020c0646c9f2471efad1ea069ae9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he675535b2c79ff309244a06847dd0862be601f96641d097a356bbb1b3c685eab1f098e4e2c0f6dd057f06107cf4b8226ed84fc1adac1e06921664f71656d11dc6f1f71235ab20b9f410e2279eed29319805e76bb2d8f1b9bedb09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155f4560be4ab2901efb92bc669e91954f0f3255472d8cec75cbfdb3498b8870d65754cad6687e2c0f3ad52fde4f98be22a97407a726bef353ccdbb44e568383a9a0184c11bdc9a83c1d10c3d7b244118cd73664bbb23fec07ebc9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2be75238a1fa0411614b6f42a8844ad8a749e718a8361805a2cbfb16458a41e450ff25858552d34bd3213c2e5ed26423846f1084ed1939e29b3590a37e60e6f06bb22cfd8250833b96e4a6ea54048c702e5ce90bc4e0fd4627069;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40e69918b76b09a560cbe44104305459ba8f3dab2f624b53a199bc3f988f48ddc10ca1be207c48c73d8703b66b41b0154449d465464e3c90810dcded0540397c061fae71b07c12825cad809421a82b9a60c396b1f6ed240c10ee21;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b0181c20b3c4a1f9f506b9809c8bbd8a65050d822fdd07dfbd63a2031469bdc75c985f64468cd89d23ad745d85dd38976c7b91ed218f832b6fe1d1d08c94285a0a78e90a64765404683f08cbee06affae6c5b30a1bc5910b3273d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78d106f7ceed81302445f4771a77faeb019c01d9bc9ba9062465992fb60c64516f592b0e94865375715e5f056347ea97fc96cc4e9fd48bdce91ffd5754b39df48ccfe9f104e8789e49725c6b471b7768a1403e7905b0a8fa5ea6ad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb2dd6dd1715e917547bfb74afbbdce490f9cfb3f385f88729731cb47944c5c036e40cf70bf715fed860edd9f4c9854ac50be0df50b43ad183c269bf92338421d425ae3b4ca35b370107611c20a27a2b5e27b3f2cc427f50a2d1de4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eced434357fa6c72d01a7c8b5da9ae1d971fe4fdcefeadd9f8ee9156302bee954d0de69998dff801c8ec046a044c51a2eaeafc8450b51a1693ff002aaff39b97d5a8bbe257fa4962cdc70ca25ecd2bed10c63d2171249675da974e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c20f4f57310f7695ff32b37ec048f11b3dfa409669ed3b7482990db48a18c8c9731ed8a06859df689339cc34f2402e44a2c1a1dc10d70b6a799139d179afb560d89246333328ae76435dfdb1168fe3f57683f445672c49e3b3929;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1823c05f2a03a9040d1842024a4e1b786e8024d576c97403feac19ea9f65680d8d733831a25c69fc0c99be2723f3899c0fb523652cc41b6821175784955bd3a90499cb401dbba50197aeaa59283ee9f9c8182e63fa0e26cf02385c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc26656f8a542597160e5065dd2ce373448188e291ca6df69671a6795e9930efdacb61add99d20b26858bfdd97cd79588e435a5c273ab6a31c57e1bf55f389f2b1619c90d71194611c5afeb967b25e66daa633f7cc4bda4b0588c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h128116eeb55279e77d1e9d457e4db2a1b3de5cd6df7bc5388d8fc3693cee30285e5b0aa088eab3e2cc69121f7b88f484340ef7a3c8337b3c464cb280c623c2dd6447fa3860d9396ac43355f2aa6410a38579198ebe588e4438b1111;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2b944343d23bd951f0c7a82ee288fb1c7282c9689680a7e9993750242c32d692b2a61dcee4f92bbb5167ace439f0031d0de93deacedb917455053fa6af88a87e6f41451969a160fb535cd9b7b738b072734b72256c8baa1af3851;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c7c24f68c459f2fae4e657e19455b12bcb0f0f16fd2c9e16b9dc010c9cfd84ce8ce826133412500559fe59a67e7209a1a52226fb0cac41090e3c7540afc092e4c1086be9b024c3dd59004662dade17976ff9cb89eae158bc66bbd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab40df89ce23761177eadaf468c0f745fe7ad2cd1bc8aa3c5b98280ec682e491f42fc054fe4e841887b61a136a506ba502066f446e16acc15fbede0040d6762f2484372a5a9b2ab6745fc9595c56783b00968de63651763a3c1bbc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6688b100aadabff31a9683b7493cf92e16039953155f6f68a2421a21e533bd280cc1d268b0a5f054798eec8317eacdf61b638b885296f8a749d745db4b27f38452e87774fe5d8cffee58c2e4fd36157a0c61d3482e6ca7ca4ecbdc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156f1780e168678e86a800478c2ba9d9c2aede4451d4e9240df0ad53226bfa927126e53413c6bf2f99703d5ed4b56cc601f243ffddcdd6171530dd2c3bd5f29b2fb64c3efce4807f8de727481b258fa609d96f7243a84d6851693ad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114c11b8a7f4ae87c9b4018e9913aa0a53215ef9562f074f029acd484723016db3ead94df71d3d456665fc3da828edb7ed1df6c8a5a740c10867eec3764ce94c0711f842c4f61287197aef07ba256ed13c273585abf0e659bd0b6db;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd528482b1bd44f31dfc71a9cdca4b0a968bcbaaf29555370379adc2cd39b081203e53aaf5daa3ef3fe89ad862f1c039da3c767ee1feab499487c58902431e766152c985c27c822c5318848ef1ecd894796e380773c1b42a4fa4b77;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2e8a6bdb3aac01bbcd0fc799228d2aa8a6496c8d5343f7838be6b16345be0af9f0434f336168ea243d6235b1e61e98824fec3c54038cd5efe4aaa8e23c4399dfd2d3086ca2f020f9a972f3f5b0ebed25a59e14945e428aa0b968b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5c6497b7ad1273e58a781ae2e786199b30938a3f55c47c48a73658efc1c74e25959cbd88e4a3f9677fb12a122ed7d04f8cbc2dc2357b80265cde042f29b1136cedcf235a2f6c33dfd213eb87ed49916998160175dc9aae3fd1fd19;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1779dc5f2e13ad8f60764355a67051de0bdf8c449710fcccdf4d2159e40107d25fce0428b4764e082f135b46eeda39443044f1e2d20133fba4086816ddc497a6f5dbf7160cca5340b7b091c2c9c306fdebb816aaa830b15151972fe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d43f232c0c9b46369a390cd577b57dc9df3482a9c726095d6a27dbc25fe03b99aec5a3259afc376e95cb85bea05ace5f57b8e68ede559f6b00434da1df136c4f5fcc4c7625ca0202f97f2f7d8fa2eb9642d0b4715de8b53931d2fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136205899524ddf82a7d441a3210c07395ca6a0cad033df2611cfc7ee5751a9bd2f478fa72103ed09b2c25ca2457cee610da09d91cc53f9f1f081b2bba08811f891b90c4405462b24e6094a73591f8d7cf62c65db1a3aacd2060b1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h52197b52cd4b8446a1ee056cb5a40df2a600f1a97144f085fed385bef8fc83f768e9983f6d6e487eed4cd5d111d27c37c39b67da182a3e34b6a1723eac91baedd3dee5281d58ecda01aed5ff16f31ab981da6739368c0ad7e4bc8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6221c4905883a0758d3818602f97aa395daeecb29bc4f55542798cb3075faa50c41e0904ed10617da9eb1bda649ce1bbefada51ab0c8c0ffc722e3c6ad0537b074979304ee93ee14a266ec94c607ee286b8c5d2001686bbb4d0688;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h198ae406c0f631081d23d3c1efa1f744f80da0d1d95ded8fb929f8572ad51cf5b1d9dc6614ec57f7ff932a8bccc583bff0ebcecb92c9be3221e5965528ca28dbfd1a671f5f392d9c0072b47d434c872fce789fdf7ee33f593eecdc9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ff211df2f65d7a3ffee462594660032f35c24e96691d073ceeb33b6c8a93ab990acc593b5a5060cbc3d8d1caddf331e670248244e0675bd5ad594bd28a987f4581db5eb6a55119489117d4122381e450eb7c2cfdc6d6f2144c351;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3bbdb12559dd5e0024494518ebd81cf1fabc8401211a36f778133c36ba772ad3842ef200e6007528738b584407de9edc3248a611e2a8f786231b79281b7db20b522b3a389f099f2cdf3d5774f291e2420686627b0b76a98fb365a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc881baf29ad386e2500b4027d41d965eece96f8ec0389acbd3caf7341773912276cb882c706dacfdec7c2676ed77c9db2b1521d358e927f758a3390d0d6cc82519346c0f7aabb3cf8e59bd551fb08a6b1af611f773fd96e58ffece;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90784d639f6bce67004febe0acc4eef987c58d9d271de740d38c33ae7e4151a375efeb7ebd68c817d2f400ad477981b7a40320a8fa3cbd1be370468395f87916b5c4fc0b772a70f1db4f05a3afaca011f239af93890811e7b87af3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b474c1f12e99fbdfd120a128907a094d7e5b5a8b833bfabea09156d7653d9603ba34bf22a9d61dc657dc0ea031c355a6eec5ff23c83d4ca27b046eaf2d4dc1e982e5a52608aa435d4fe9486dcdd72367a955bf53659e07ac7ade4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af539382a3f06f23929f13940d8344780d06a8b56921826386762038be62151be82d9fcf4794b6f1bb365f12192e457f1e2ba8b844c524d1a90f55794cd98671166a452b2842e3fedc7af191529f3d9d773cc58705065469615a64;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40b54871d6c6d86d17c8f9426377dac6f14b06ec9160d167f54ff5aeec5c6ec983a8441c79902312a4544d6f5996ba26da71327f2f318f683ce492791957030508d22e5108ebc20d69d643c4fdad79f7fb33e2865144237aac2943;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcca9fc044faca2435c43a73290824fd9a71b1655f3d291533c04bb939df88d9307ae744108c2742da0da3c06519b3efa629efb4f722a67717c5baa14d7f52577fcbf1919730d05426bb42c1e9da7732b941cedf32895b34a287af5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3bb5e34c88b54fdb9de13c789d2ae2b0207f13304129b23a6a0c9967adc2de403ff8bc9c8dad37fb471ea0a6f9ab25df1fcff45269e85f1dd70ca9a567f4a3091d85922be299eabd78dee78797dbb3d6cd639a942fecee3a9f9127;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a15a9e6b6a2f71bd9733f2d76d3df690837641e20a76b7d717d68e47a930f10ccc4fb761cb7015171588f242fb5cc33a14f930a3eb76724ab1d720e30c9297fbe2ae903ee4d95b45d8b40a5b7cc327bb7f7b31b0292ce936766b67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1034f294987dd36156fbdd23dc8e255a54f3af5ed6b91d015c7cae450f85be624570f4979781d2f1f1ce025bdf4a5c3caa336422a8a483d50f4c95ba8ec3af526ec96c843f40adf6fa9caa1b37cd8b94f5f8f7e0f939991a23c2f86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53401033d1262a94c104f48e1d0dca8021fc0dd7a35e4a5e5ff5b79e72e17438f439d0f892ffd30d359d77390dcf22b84d43005a780946b0392af6b480b6b1b0883e9faccc20c34d71c2fc5ed80f26fb7b4e18ecbdbd26e55d093a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h154394b22e95b2bbff4f9d691182b505e994e0a1d0a143daf8a0f7b9a6ea6cff3dc777934c8c2415cc510cda2f3db253899a7dce96bf3a551a5ce03c0f62651c11ac92d105fb4907e239916718872b1ae000b0f4aaae9a6eec6ee60;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda8ead2f5adf51eae1b1fd6612e8797a2f53dfcd42e9628266de524b5d82faa81c4d6b1712afe18ee5eb54c2fb9d19b84fe2987f7601527bbfd0c72317e2c79b51b1e37a5ba3e1aa1ac6131691faedaddfd4fc7884549cd209afff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h134420903faf218eec92365123397dd0d78edb7d7422e8df8f97ac0154cf6be3030e0c5c9d1cfddb67844723af7f4ccaba2778e47bf963936d137c50309d4d5ff9fc34b9165a7504da56a90aa67cb29ef9f65be98c52fbd0a765af5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h532d75c8a40b5c28aacbc34f2a095ccf5228dc8c9528920ee28c5bf549ea5d9ba2f23305de8091487e9cd8a8b3afc1e2e9155d625297d25e4c9bd51054b572f43d3e0be7a8a3c2ca22d7067d79d265671397fbf7bc5f912df8232f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41e6223b397aff1a3a773d6e52897d63d09d77a2636740b91d2e9ccbeb518141b5b0bf2b777c57c3f573ed8738f4d86b20966126252079cb739223728639098a7b23dba49857ada102bd723e75b9d8fe1cccb616708364372738f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c404022e2a6ad6294c68fea458aaf444bf500438b821fd84ea9597ade2f4aa17a55ed605a896036ed8793600f7f35512b33942d5400931a67780e9d5eb15de1e1a4621655a65ffc1a1a2805a5487d533c3d44e3d2731883afe646d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h118a86d07f33cb4fca67fd2a7a8f0202320a17eeca97cd0e23a265d94d2f129559bb07dab02f4ab688c423367eb47b7bf05e8725e7ec540ded411abfe02979e3e1eb013f1cc7fd1c9b98a9ab1f2ee7c1d2ff78964f10b371f614e14;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4183ee7bb060a0dff1f835543965fe02792c3b4351dabbdefcfdd4126fbc377a603e04de172057b0446e72f9f3fe0928c21c1096a1f557b4683c039c1dd3bdeeea7f805aa10e10c656b15da938bc1cfa2382210839632dd1131ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144d8ea4e21fb0aa4f4ea1362e7e67d6369ff0642ea2b9175a89368bd81a51279a7389ec11444273e8594bd7d6fa38f34c55b6bcf30736100589294e71240072c5f731a96152fd714c3da23243ddd5fa636a37b91a7fa8cc317b563;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d165ea5040a1f3a935d89b02b9f2bb86c617b1a2fceeda12042afa1e3501f3baeca5b2b6d34051eade724119efcad70ce86bee57a8812e056f8af6b7226d7a17666d3a505c0e771c256eb46a1a32743fd9e726e6393efca059e662;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha67291e4c35324353700b8138b127f8fd61685595b55ff4a8243498b0e3b529745a159118ffef95bfdffb72c6d0a293f66ce3fe5eece989e31519914896b3d7a1ef811f7cd827bb2bddf7c5a6ecf8dea8d49f7dd0eb19f87be0f90;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1219de411ba7cedd0247eed053dd3d03bbb1d53994e61dbd78f2113b0bbbbdf8f5605a722dea5a80fd1ef7ece3b83227056175deaddbe50a6f619a4544bbcc15bd28b2b6d837b7094957f8dd01f9249a51599b88b180b43f181d1bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h995886eaaf1d890a60110c913698cafb8f3aa8064bdd38b79efa15bacd5e373c80695acbf12bfc5c92434b10804979d8c752d5929f624369613529d30b955933d2630085dd22730a6e0a0d4de55437810bf5afac97095edb53ab25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76f5890489e99a80eacff7b0fe892bc7040b1916c0a1fca3daac9453fd86aaef0eba900d2f078cffa2ecf6131f25bfeea8eb460302c9f52d6587a1673a7f955b1473de3130d0c608a941a129151cbec00a692496d1ca8e1d25ab25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c9d0fc4fb12116364db5f015c4fc8179682a61bc26ef89f1c6292da0031636b8a03a90c070c5be55521fe5f3ef0a6464e48e59ef02973a0b799e57fae1371e19389f4f8fc7b79c1e65043cfe7c34f80b6da172e0bf087ee9d99e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6362393f7a0e90e4aa9975e8d69620f13c0ff51fbb6404aff09ff19658e0074718f988e9b043ed22848163d9fa043e32c0d41e0a95732a27993d437d2043775a5d44e593cc3e74d1aaa818279c1ef07958e81f6ba3738f3286df13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he96919748f68fd53b2ea7f5a44a1f2bdcc4bff8f19d2b0dfb36b3583e51bb935dfc2a7f0975574e7108ad02905d7f5eb5e390ffa8c24cd47c56e5737ff7e0aae83d52ea00b3de0c042d7d373b830c62ef62ec42dac1969165ac222;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a566dc8fd6a6234e2d7229365d14c2d07a00ab3153d7bd4d470cc203439b928169e03c3f6879bb6b0e466e2be06bebf87eb9ab9512152ab1456995ad90ca7a3d9a19f30116c67135878a45da19c756a4f78c7708e46212f50d13e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cab5e42d47f80e75e2884f973d4c48204b6649b855a77c30c0293b3df09a6515c3f9a6a342d0e7ffb2c17b9008485d803ebabde1407be18eeac8aaa1d3313c134087aaa6b662fc5fcb2eebfb7e8eb47788701e42e6a203ef032c8a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h285e61164968e18f5bbcb6ecb155f4e307d0ec89547039c2f246b97d6f347cea5e6c14e701726a72699e407603207d84c1137d97638729bedd97cbd133a6b8abc4d15fd4a674c7f1ceef1b9821b57fa03571e70b8c8c1fdc6eef44;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc6403e601acdbcdbc1afad5ad33938c7c5cb0daa3dfc4cf91d5e9cd0637ea5cc84abf37b95353abe0672532573aa193b8dfe3896dda47969b985e6f57b2c2d51d9afbfe8452c2b248570de2d3e7756b39b071c03962d4edc8d4997;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf301bf6cc4ffff23f69d35ac5a8cc8d7c71350aa8726d5b5c576b5614e234f93da326eb494f585d330a69f48f0476a5b116006c2f97325cc6fd606b9c878afd894e1e57f04c3c1b57b027112085bf35ad3d1a7477df188baa6a66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17827252f3de23a3fd631f81888b2457a20b3103053e368c55f9432fbb9dc50fe8997f84eb3a7de9182e8b69319e36cf3ef8319254d3984c14d0daed683a6e5abc6d94c75db30a3560f8d45bd63a4fbd1c398af2cc2b1a589c6e1a7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1664f614cff878855a847cd2daf2a6b38959bfffcf0d8ac39824a811e150addda8e51bf9e47194f7b8ad26e8ca6efd67724963671311f6f08c34aa1bbbed2870ec680ece1bc244c5f3f5d7ddd4b2c7b717a157f22fdba532ff576b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hacada758862a95a5fbadc591c0e88f3c5f32f72a0c35307a49428c5ec56f01510c6d5332466919488ee9a610b73fbf8040c81cd16c3167b3f03a3d800eda34c0dc702334bc006ef68383fa194dc7ad01f4c81ade7da0d2b78bcf07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25d32a1b78925a025a7c1868f9b0dbd8bce85d425a267fafd29a4dccc6d1764009afa82106b70a5938c34aa9e089874343a53674a7b4a8d0b7538b0adb0c66317d5b15132c7de25685385dda4ea31a913318b37bb0a5bc868821c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ada3d583fc22f6b3652953db9d49f104b647299e5cb9a7782143774d3f8b4722709c0b73b06dfc87b9f2996987b77db58c205dcc3235d37f6e5fd7bcc5e673f0526dabe1628fc3f61fbe5fc52074c7ea03e5a55fb53062a986299;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11516704579b9e701f7576aa992377e5318d1733c3c193401a6a27b9cbc68e3e500f9af9f829486791f9179f37e01070d85124e2254257d9deb57192d058c9f472bafbc347a4eafb29580fe9501ad812f6b30f14750c1e2ebd68e68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99207ce48b8909c4aa415d03b7a0ce19a6d341c41d0c12f5418e2d3b9984b6e0c4d5d1fa1837e56a436cc251e3f0060611b4c699ccf009d19f2789b5ce01834eb726d8576b6c2b026a09dd093893b29bddee0a90d261e2a840f38d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179b08d9ccd9d1c450fde3ad3e093101ee38fa1fe20e147067e9c78716f3744e3c577bd49178ebefcd3f5f2e8d3270dc6918260ccf838b0e05d3d14f4def50e5b316ce87c1bbb162b583f83457fcd259b5744b0bd8e9a29510f0de1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b2733c54ac3ff4c6e7efe4807eec0576c03fc113a23f131e6daf90beedaed7592af18ce7a5c9a073e92b3871288c9395accb0f719ca0f9f22edb6eef32830661f59d26889a85f6fe1b1fc9bdbed7ea70a914a42008d32843f4544;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194caa41e3c85d8717a586290e558ec6629c0fac0c77d642a0304b752785fb5007952c3c3a3a721d47f4b6ac7829b042d36962acb28ed464bd55685a8c89bf4de6621f52f96fad6889487726c029ce37c619dc88cbe1c8707685062;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115ef02f381ca7f7ef5807c189d0c7792386a7acfcc2d3e6c4c7ae1854c89adf8f769627c79e74d17a17dca1a011315574f2ef7d71a32c86cdff7d39ab22dfbce857ed8b72c09855f84dc11944a92234193e3e00e88dd7ae8b8f074;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180c25c0da166612a5f71eee465b021e94c7bbc942264bad7613350a6335fefe0b52a4240ae668d48d17b22c39224559a18615845173fafd3be7c00a01018af9f8b0c71eb1c49f0303f2620ca2b3f91bef77c48d935432dcb028dac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d63f409f83458bb2fea3f813e2bf1aec0647cb9cccce0230dae62ee8fedb9d7036ee07e72c94b349aa339c37ee3311cc04e531444ad45f89691fd01519d810f8cf93639052088d086256e88ccba6b196a55d003d5baca1f9eb3c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11844764a42fb7f5ec13916641780cb41bfdfe6356c7eff0349caf32eed088e0bcda87436d3ea69de346f5971d8a4f791f927964e825a2348535d4e47730512015f3822ff00668b0995c292a5fcff51ece8cf4f6f7de63e83547422;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62e32997c9bfcc0cbea3fde5443f64974448f6fbabe9192019fc738d94ae4cca5e14ba1f1169e4f6e3fbd3a33b557df8249368c60fb84be0e6bac805ca8f64cee3ded5ac549e309cc4df916b3129c80a0227caa24c5a55aa5f34;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1d4f4a93dc89afd76d8cc8734ccde630b6d8e29af377d251e21ce496921fa61b809273176093de034a224da33e9d008ef867be4a153c1f7a83968a6f07e6b3d95d0f1d9263bd40da2d3249846542740f711a4eef23f73413561a5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h873ce6ba623006c72ff4f75fe710c4b010367c3c40a9d60b4d4db493a6cd278611484cd91decb4ff2a6fd6e1c8e6c48c8e5858d359813d8c565f3ce0ec8dc991136219602ee896bdcd5c6f4c3575427629edff59ddf205e9d8493a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1821284d99be146b765297f5f1b14d225b62c991f40b6a28932d46d968555b01483f707c1724a7ad217b471a8f0e4a085d82225f43ec6c576bfe394deaf25c11c6383bae2da68742171c48553286d4bd6b3273a034036167b9d1199;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d9a3dcedde261d70344e535d02660df3eece8651a9fee7993a8eaa91aa2ed40b8ac4f4b61d32f310c0257c1a5e8c915bcc22b15eb2fbf958a01bfe2f8da511546fa2c05026cbd787bb3debe78bcb80c4b82c70dfcd17bbc3ff1fe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2baed1c4a991d64174ca66ef111ec81b57bd4c3592ae5f44f5eeed77018debb000577e5121d37401149944417bdfb534a2bfff3b7fd98434947dba924bf64cb5841102de4ace3a594b360618ffc8ce5bc759202d52639325a9343a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172630943f70afe23883fc5fcb99d3530fb61b31c20bb6e0d0bb52137b433ac103919b8fda41b29ef8a8337f83d27fe25929ab9f2f76123c10c788f9cf18e619a17b858e6f47ecb32c8a14cdea965aaf00b7c960a05f4b704dce0dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72007119ca6a7261f76f576a2f62ecfab47c0ec7808b2a8e90a1f32de8bd542659d4dc7ff762454d45c78988c139d89d4390e41bf5dac2bf1130e25a620bce15017412c9d2141ce1ec9df7a4c3c2d73553f3650a54f59beac4cdd2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37d1e315b17c4288829920e5c5bcfe5275ea2c1fe78adcc431dee4f616af99daa4c51e8d3b7acb20147a7aa099ad5e84d83b7d7f23d4c54eb570dc5ed6bcb43550793d38fa196b6ade4ffab2fa9b82e72bdff9f9f8134ab821441a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3aff4fd3851847a79a0ecccda3baef8b9fbf48ec6df688a16edd2058f3d0bb4d07f431c0be492b3c36533408f4fc5b531acf0a97825b9fdfe935a6886be6f9d22707b4e3132bc1162faaef1c0ca31293b7edf4b5c4348e028c3227;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8d52a09197cec769450305a89394eae2928327832928fa9856ad34e766f9ebead7d9bb398d52e29f71970c571e5d74f923c264c749a89cdcff8d8c2f603782ab36120b157be87cc12c0292c06d5d261f7322ac6728534ec6a0b64;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16741dc008baa49adfc6e81ba066d3dadeaaa3c127c1379eb322f40b30f0a01c3ea3db1b9452fcd432d9b7ab77c7075973fe86be33fdd3e0c311d0b5439c30ae82b106855fd619dfbf57930b8f8792f83993e665d2964e49bee7376;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f3ae53af0928aad98d254d78ab4f55bfe17f490b2c2d282ffc59924ee41ec416ee632ca032a22b2ef163d12b1a7d518dcbd741a80496a5afd5879ac9ae1de94d865a1bd871769be37b94d61f024b98b8ae436029075e65405b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116f12b2d131b610e5452bf6d0831d6c848e31b5b18d45b250f5adaf61e06dace493b90b75819daa690f05d076239239ee3cb3a093594576d36f367b3c3057ff3544fa81a13691a0ec9f5786c21236d37c031d0a37561e62a160ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0a78964dd78d0dbf288d77aba44cd3aa3b14f7c18a343b9daac37778591a00912eb9306b42ef8ab3e51a53058265b20a306687865a676bbbc70ae6a39a38b551ce5f530a62650bab60cadeeb496cf0b7285b3d840a5c0689684d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc127e487d1a3db1aa727635b6f4c29c4e34c00d2742919a641ff56cad14ec4dc0bb0513da6b1756bcb98bd97cec52902776bb0eb6af87d1ccb56351c68a0fbcd7da21f03a0102ff648f815cdbae550e3477ec5de1f45148172292;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa112d404dc42f693864ee3cdf3f4e46fe839fe29e578e9500ed4bd07a5709b634e63414c751ccef5aaa2e8ed1a9fd1a7aa01095023a0f889b6fbee774380749f025d2f1726417872d37e66cc3db1d6c0c32d0686f101e3f2ae524;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1390e50369e96207dd7a2e0ee46b7e29cbea59a92b188b1e21d968d194ebb2230df5e2dfbda54cd913bfbcec1d811af0883b5eb8f68c2b8f1a2066e7591c9118591f22eaa0892e0cd863d0957558564aa9848d9e7229ab2e9cba110;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd90fff01dc473246b0983c68103c3c97d2dc8f098b4a3eecb53797f3679ccfd7b0d174aa30ffdd8ce5f8d4860aa2dee0b0ccd3ac151df8c3bd4ff1c58b617bd8037285b6c6a2e8933ae17742e1ae30c25f967c4f37b57dc88ca161;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc4d54053cd291d1c4c02fb18348fb65ec418f41405128e65aca216fb059f340b0dc4044fe97b99344a6f0591f67229d5b7d17f1441f5db9f7b4fea6e00777d4d65f7fc6962314fd0210d3ccf31a4e0508a80b27daa45a921fd3d0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h922f7d589692525bec2e18d7988b559b33f305ff30c942003fea464a1f6f971e7fb5f27b54cdb7b47a32d0d2efe5403108c77dbb13487f4beed9eaa2a5ceba654e818499d2b7c561d2ecffcb6005dc49638c14171317baeb7fda46;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc3a57863cd290c127af82d388b9f72db833484b9e265a46c9b7c938ffe7379f114ca70fd1585d8a7f35246268894bb91be0bc972c91a270b29af7595fab3d7634564626fc2327820bbc779be0ff646942b1c5fce244096a45eb645;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f9a37f110d8b7619dca1c52b5e656a1993dc6130c936187bba95663fc57b872e080f0ed6f0f48a31a7429a9bb52047d0ad45bddb02d99a64ddab80c35402b99b61a82eaa4a5374e6d956c8c8d7075f95567194c0dcf020bd6e3b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176d06f78caf52ce7323ebe5a4a853ec3ffbd67db0e184c2cdafe70eb1019e0de983fd433d363a640d9d6ceb3397c560b360a9bdf51bc0f05fb4296570c80af6626bc784e93503d3adc2a99a76b06638617623cbb84db6c55b131d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0917813a50a880ed273dd4f50aa08a07caf6adae83a62a20b738adbfa02ce94bb432713c13802eb0b7ac7e62954f7bd3e4713c5225944ce98159f45ecf8450f4081d988b061dd4912e0bb1b88135bc5689fa933303edaece02ad3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1117e090886ca003327352b8972e19d57a1b1dc624220ec7ed11b234f642a0d4482b2ab3761b8a5d04ce63725d55e25a5a7665dcf15f0013bd7483a0e31c4f15f5e5092da230abe6e9c998123ea6b79c21c77146135c45b16fe4363;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4fd29733f480a3420098a70d9ec44774d8840566531828f7c254600dc777dcfde1429b7135453c0b03d022136a4bbecbb105dbb35cfe074e6e4c3a4cfcb56896329ad4de23b2b367d74ced98a3765febf27c3ede2eb45b51ad295;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b57c45495d4b4595f889123fb5bc24a53c9baa3a1924cfe41d06711e93b6608914086dc3289602c6f70fa6d5ff1cf895736a7ead3dd747ef3d19c3a85b11c05e4414504152bc3c6ad0220d0d095147aef4596ebe24476ed5d20f1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0c2f5a7a8a72f5e58d6d5a6835b4b1ba7eee69d18ef662d678fab63f7684226cb4c3d7e5fe4d44782d64a1ac264b7cb46677da8387fe31d14babd5a787b7c34af37bb6b5a909f5653b5e4891df5c93cb441b43de33d3d300406c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h580ce561daf2d28cee4aa2fc17d15117df22d15ac46604215b90a5f0441f1905185d8a4418677d73ccb74174cdbcf69b448aee2c3d89676c4b93a0db463955810fbd6736813b20ddb09d4f567297e9ed8bf79d99d24702949f1c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4230796984266d1717bb8b219ab20cf586427bcc8941a68892d356de194e2e2aa34cbf2eec616919728c5ce8cce1f3e640d538fc39e8bf3d9a1130843ae14a0eb88a152b19b1f8c9b8b5794d52f5d8e45888edfc93be80e4b82196;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf28dd0bfecdb512c84662ba5899c0f3c46af8b6a6de9a50fd9c89fef166bb3b72a50734239a74735de0b8d68def053a9ebefa5ec218ad1c8612f2844a9b996ce3306822d7e01e5c512cc7db16300dc6e58cdbbb6e6bd3798fe9fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce6892e4bcbb3fba69234b16cd9ea822a210c8801d011f0063fe454ab26f0119d7ae6466b30a2927e60d222f106ab1a493bf210017dc6198e287f3f737b5deb3f66115f23f8561f751bf17c2ff9d2e3d05013d917bdab9c4a9a70e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eac93247206633024aefc84ca03313e08a83146e10a3448ebaf461ea7cc5260959ee2f6ff41eb7cf44454a2af6f87befc5a3ebef8aac5a8f0891b1e092bbe9416530af8bdd31ac700c5fa46ce4f82d419eeb424e38b3e81846452a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h582c28af8960418c3f4a1e9a7485677c32a74c0ff27e16bf4936644492c102a0836b3905842aac2323f125b320832f5d117c0d15ec3dc73e4e03b1a594635f12cd7efb7c8af517c8e52d0bdfa5deb7c12fc701f010c44a22ee085c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79e0bc742f0c55f59f68d1f887097b3f1ff6eb2cacea562b6c6cc0f049a0b4597360a48ee4be7bc4a53dbc5e171b56dfa1390d632f496bc971da71c95d994ceb45235c48705aee6331390f32fdfb35100cb655cbdc7df392b076f9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23b6697293eb0e352ac142067fc736e67861c2edcd6d51dd2352dc3102c162e63bb77e5e719676dea6d581ae232dc4f15b700fc217071169b849a99952e96a0e7a50f2676812242dab9432f5f87d242137578da1fdbcb649411bb1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76c39435d268aa037980c4dc7fee8e2187ca07489ef4fb7b0f69590fb19fdf77e9b002ecbd9358abda97bcef4dece9d1b1874ad8ddaf812e53deece2bd318bc389298dc489f4e8a78d043bbd6b9d676662c9b36c4e60d1d18542ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefb0032c530954aba28236b017e7a7d0f6c3ba592697c8151af41d07c52048ef359cf591ee67330f66aeb9ffef746fe2e445d0fed4fac5401dabe512f2c959399e65c564664a5661b0e95e3d36389687504c03a3b93579cb840426;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2a887408f4b4bb201c456731e26c1956c7968ebeae8898e5cae41e8d97f9e53298c1230ddd4b1bfc31419018686bc1de8c3c57c22f2bc6f2c60f5f2d7f75ee9e97ef233864cb81b3f2afb8612737e0d1640541ada0046aa9f04a44;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d4b18319dff9f84d08cabbcf980017b403929fe465428b8da7126fd42ac9a3fb771b81b528209340f1b7c7bb476fdb51960145db0001e3ed9944e0259784911313e7ea1fc211f439a27037f9d37c303f2d88f8e6adf4a496d7556;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7b73098b528d8e023691bce99669dcaecb30836afe3dd9cf40e39dc925923e7d4284109014b9ec37e802ebe064e0dd360ac5ac732e1ff87ff697a0399b3019f15ea1dbcdbbb4d9c2fda26727556c252dd67c8cafcf340f0f30756;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d4ae232a18bda757860dc96402f25fa492abe75cf89b29a377960cf58aa572fa7872b7854c83ea956099b1d19b50b7c752b080bb5308381cb27c34dd0d050b38c4239807bb25a2e1e5da525f6b0fd4cc721b43fad281bc97236a7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16155654b7118e98c06da07370bafd22f790c28e05c75bd7b0e822f2dcaa425d2f93527d64d9e66108771a8d9e233ff35bd56939b625a9b9e603a7b8a2f45923d1b59087a7c934999a2be68437d6bb275a36e28b59e13510a01def7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdbdf8d0e3cbd87ede03f5919408bf572a9197708a45fcfb62b3b8259d7ad2a6a8bed990356d0026b8aa9d953397b5fe37b8c66b51c1ef35ba158112aa7346969a6524593228e9d370f81c8cfa031b5338e4b52604d1665753d08d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10bc79dfd5ff84a7a9785c05806312db39f9153cc44ef9daf38fa455166e71416be933f9be9d736295d119597245dacefe65638906458cc691bf0f3123001823e9730bed7067773c6ac66b9fbaab2925b44f16c454f9212943fed04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24d13287392a5d4a2346ccabe9eef3faa7613108e7af198c25738b83c6ac3d93515ff129dc0edcc0e41cae58aa1ceb06c56fea4d22fbc9f0f7eac0512d46c89bb22b3f16819c933de9eb04dec53caeb69112e6e658dac1cbfd0d18;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h382ea3f72cb6607e304a71cca3b8adae22dd405c827d58dcdbf6b18903da4526f908596953ad36b23dcfae3397edba8468eeba0458a6bf972e4a79db3a628ebbaf4d3e19ac96566e583880cf9b82e253d668e58d41b40c561ae22f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h494fab09cf473ec0f24d8d5ba88f398328f70b45f6683641f2ecc142cfe3ea6755376c0e2194316eff0368e1b7e1a034c7460e28ab6d773439b84a326d049fa78ecd93c5f1f8c2efa69242e3767e74839e09db9ed58c3c8bc9ff03;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he357b87d2244bc2f3ece4d1def02bda6bc387d535ee71be25348ae0b144bf4512f39d905eeb0ccb2fd7db3c1f303b35a2f8a39fe1b6fbee2c0d2811da43a9c8e45f74a4a06c88cae8bd73240733b779ca67140e021d2a69c785a64;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da37ff7a8b09680df8a6f802b197701283195809eec9e708162769bccec3ed6ab60144347cd61363aefcc77e510b94c2499378b3c03d7d8f63ebd9f274aad15a92aac6ff56b97301442be3feee0f77d5b671989e9ea1720b5441e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h689882c5de8bd6f71c0fcf4ccf75fb3b99984e6bf5233c76ee84c42a61b8fa7789aa513910b0e0fac1a77e0a60347a1d346e07582f8ad0e9b395036a9e2c66c6aeda334e7d45617b518b6a41f4c3f320b26c566682fb6aa014f014;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85b90188a13d0eb54a099c4c0e6e5420334745805cbf7fbcddc951330932f8e4f94e50a8bfa4c6c67e52d555f34fd74c23e744c13d3043ae200732475c1dc44e5b962733394dd400b448fcdfd44bad214b72791830473e18456088;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ea0c51ee86045f14dae631e8e61349cdce48e9a481f6925a0acb1124fac36bc731878773327d4d0cd14dfc710baef7a3cdfebb91eddcc020d2629723a14af64ca54f5909768cf9735eeadde0acab33a323cf44ad0bdd86d04c1d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he20d0f9b795ec42dd25484c39ce4c7d54e9a8dbe8d337b3079466c353b070c78fba8954a3e722f9d712c4eaaf6032ead5fb0021d10092cecddc235553d8140e6ef49b149415ab5b4ceded8c8cf35e66e25c8864377b21fc867598b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h128da73049a2551f575529a1f05a10f7ab59ca15395f8f17fa4ed27e1edf407cb5fab214c7309027acc7576defe18800ccb6d20433931eb7ef8d768ea22f7a96ffde79b457051dd3a6fa64d3cf53889e11445106073e539c4598e4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha146bdb4c106ce6070bed7d984b71bfeaa5b7fdff47a8cedffeca4f6ca469623193601af124d592bbfc2dc750ddd2dd9131c1daad2f1d3eeb10e20315fbc7ce7b19395c8a6056e4235c858d1c993442ce3024fb768f4122197684f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8e74cf8fbd4843b8a7aacd0fe339db0394bdc48c1ff18337955975054c80b0b742383006111b549d4f1ee7f6bf4bda1a032ee6ea20b5a576eeadf872bf3132c0ff75dd55a6269192bf86e4052facd3c23eb6405af89511e2ea217;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4b16bf22fed5de81a587758bb49a9fe2deea2266502f4439bfc44c72a250507b85b996fbd67d1332499cbf715dd4f34fdd72eed9a0b07b7295ff831c839880b43dcb960e9ff0e9a1695f4ac825f9900c28408323503fe4ed7baf8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c0597f0a76e0f60e8a7f3243b32593688b98e324a548078ec7f696782740cabff12823951ee43422d5c01312b2298085b15263089ecebd5811fc935e7e76d2d1e5e615a4e7616a3e9f0a1e9f04fd3bb4c8139fbcdf17773c34e94;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dcee204d7a64339b682a5ec9e7c481296387c77ec35b5c30fbb75d8793a82b006d30e8dfff836542e947be162cf8170698822f830a09d0d5b5a10ee20c2af41e233e5e8d6ff069009655a98269909e0fbb2d0aca50e9435363e66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ac5cdbfcff03b1ce61a466e290f011d6261f2d2219fe2462327986c57710dbd3adb86e964b517584f7a7d15a2e7d7f0979c7b49128ee95dcceb68e2fa60b09735a88cb639edde575a106d4729c13a8d44fd588931db9b02ff7a79;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8d7e57735fa2c2db5ee652882f420f2475bfd29f304303b0800d94bb9e27f5e96380a49f3e9548713f9c368d922df76b7830025961247da558677525974909c4e3e0081b028cf7ca97b1b4f0832e0f3bf2baefc29dcc0fc32208;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8c6afbf3c31a012026d2b0a82cd000c49a1daebd1d5692237cc16ca3164399bfdb439e24cbcde4619185f1cf74eed1588f2fe3c191f067766936b58dd90301f1cfefaeeb5b7c22517b068ad2360a51c1352883fe414f79cc18bd5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h766d40c10494404fe378a031e7c1b919c7fabe75b20cc37b3b4234dbe45d944cbc2a7fe961bb6a8eb6d3a9489bbad1d12f6caf3b0b6efdfc583fe3169b3f801dad58a860b1f3fd5b507ed56a0b14736414c4cd8e926b635c9dec25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18848575946bf69b68bfc15813d93895eb43638bd57002aa130d092ff0b977710a95fdb983447033b91b3773d6a1c9aa92294d88f7edd8623c91af3fd402cc1c8e2c7595992b2fa7825d89227509cf08234cea7f9b48c521016d6bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19cc42cc74f9c812eb85b935ecf69f3a389cda8a02de4104f3ad50ba969896bfbced30b2744cf061d886178a93cfd57a49a30fd6f4cb9c7039d375a96b00cfc6120b91f51390b3f8f486b55291a75084aebf578c0ef17f75842533c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec90aac4b9b3997330271371932e801d9e9fb60204f6974cde792d8c67e4879ca76fe24e2440f1fbf580e51e0d31654bb716dcf966b36ed09eaf9356835f898acb0e373f003c5bfa1aca7bd6b1d4e29292132092468399068eedbc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf0282bbdab5ce72f34a5522e0bca4d3302f749c1fc3c3d30586dc859e317c641fadd778f55a517110262615c01ed36bbd1a4533e8fd3586b04d32412c136a8526b45d78076b511ddf70d9a392c7aafd297983f796ff42cc709e7d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h590b90cc7e694bc47bb0b2bd3661606567c43a235b3544cc1e2130edaba655ff62613515181a7873854559408d80bf23b4a60aae32fc18cf78794db0546e291c120b3500f1534dcd7b23397d422f1717460a87b701196f969e28f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13e8a09f0fe94cd3a3894c74aaf1a7bca1e33e4201fafb766ddb4360f7e6ae73cec3cfc1a82049be88481c14320d578f74aa1ff31eaa4bac8a1a02fb8ad9ee2ba66246cbbe7f6313f7935f1e29d1258514614d3347ac7990ad23703;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1490e50d0637a45916ffb3c36825e727b4ceba2ecd919c8f5fcf1a84e4a4400a5bb57505af7239374ed8d1db1baf25ee17fa78681c81209dff9d482f33063f0da763b6e4d99baa0152bf0f08d081e5d3a3220f9ff57f7ea200b2c3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1365c15d2ec7a55c32b2d5b8c4b85ab822d2d64abdab0d17d8fc0e172828327412336f5f7aedc57be4f6a932ad019c32cd48d9539bcb895243de1132c57972871b202a7b2fafef82d7c403b3307bd13c6455936b755b2f1b898d901;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2807b3f5313868eb97010118c222abfba41d911959c45be693fbd88fbf93e95a33604bfce189bb278e92814c56e0e16761b42fc55f4d61e910ceb0b92dc0b5350a10766ce9e9bb4c9b112458fdfdec2cf2707ef9c701541255108;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9a6644c38d1f69249ee367f46cc1addd56afea0044c33448f356ce073f2181263dbb9f7c0269f28bdda28f8e029f7825531ba662fbc509daaf696917b14f1ce7cb7e61d9aae254c88b0cdc8c5f956b19b0ec18c841f387743d973;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3116741bbbbe300372a76bf7f58a8a6e648e9988112a816eac2287dc1dbfe8e04931b57e1a7bf9c6bdfb965ff652f48ea71bfb6a159e672aa8e14247f064ac41bf7942a9b9ca7441fe3ce83eda12fc891d7879cc4991b6f82d9cfa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h191f7d10e49f8fa31c4dcbfb3d4d2b3f4a0467301b4267e605e7114cb4d5caec75e73d60a84b3afb5a3529d887878c6352b8826e12f91c89d06aadd06f4f61988754bdd2ed0d99f40e1aa1155ea80e7e95a501a51a6a6702f29b3fe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdcefba54f241a44972b0b4f64df6669cd221e6bac9b04866f634b8e8d1883a7a3b7903af570a10357be497eff14d77ce568bc54e306112fd37d1ccd1c8ffa98893a1e7e5eb440201788b74fa854981f29d47f038bedbed512141d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1afb2309ccef84b74cd4a46ebaf678c624566d93f4a1e1d2eeca3a5b73e40593365023fe0505c8242e8aacd5b32f5bf9d13ec93b8727a2fff876de3ca18209c84db5ac1b9ac577a269c77a19a979ba4aa76cc1d294b12490893563e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h100e395c2c5687450f5e02485a4a0411bee2958d653f1aab9aa1f4f6a5487ef8636c5a82d123bf29a298a8e36b640b05d188ed2ae560a4f030d09e454fe693e6926a8aca052e4b7964ba8a5bf9b07d5d5171789b9729dbe1c1bbd8e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h159c996176ce8106d3ee111061c27e4133e08ba7b41f87ed2a521ee376264b98ec94751da2337432299faca3517b3d73ba3ac08aeed871d30f6658c52aa9c66d5799f42d301f2cff2fb682d7100a4e05dc25967b60f6b9b867d7a9c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15652bcfe5b22af499d08761d79f74883f2c36ead513162e0929fc26ff6cc5fcf400948dd3e3021a970114a6ce8bfd412ccd87e11297751428615b30eb7ccb752468d8dee3eada799fbd51ad836a7d68f33d6a2a7d9b1fb8f6037ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1883358a3389942ce3b1e0dd0f2023dfce414213d3129bcd3fda59d87abd4156112a9552e8edb0d8b225debbccf630d6262f2ff47c63f99e0c56cc872df12f45229c06d3f16b78c2f7440b95075aecb4336dfa43421e0aded5a2da2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab755a144bc5eec4d9799f93de5299ce942cbd9ccbca92e537b82e0faec895439c3fd9cc5ab76d7e8b9dc0f5f70239221e75d497736afb8b2543cc218a17529a215df2b5d7a2b939a29fa69b86537c5b284a63c593d396032db430;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168dd7738e1368f462f7d2cc0f5f44805f8a56ebfd8eedd5306c4895556fb0fc5543cc69ba125d6f4cd798722ee4f4b9dbefb332ec17ef40a3c4b9db80ed8c5371f297a3a067649d89e684ea758824aadde561a69d26a83893dbe5a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78563eda381eeb3d20b6061c36d80137e44139355c147b1c263b543d6e06fe5db79979930b6cd509a6547133f0fa10c4174c439d4c1cd04f539c6c4708d5d09dd6141383913aeb2e77b18899b52181a6a596c815efcbb02127f8d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ca1ae34673846d4d2f0f2063a91a3eeeeb619828fe64a61104ecc45c337600f01886b92f141e47bdbbe3294064b3d0df60570c44e051b5e930a60921d61bfbe5ac6010c73a2929cae33b3e8fed6fd2b356fd069114b2b87ff7300;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8beb8d775fae510ece3f71a8d79a5b93510807a2ee84229c6a26ed321d7473b191fffbcc8ca2b12d99a19170706645f30e325f429743e646b9fc8497155d1bd6b7d80360d205a4f86a031fda06d1da3a457ba08801ac7b2f39218;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c475acf8ddbc104beac16ae7835b634a42a4c2f55391ff85d2058337b0b3cae36bc9f04cb11d217edd359e80478902559551a98748e76ec8f573058f297af8047e460fbfb307d321a68fca557d5469e63189987193d69959e1f94c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1492cb7e54dc92e970c4671913572797ddd3c8e9c51f0c10b1611d13f169fc98d73be0983b5162b242f8a73652631f1b853c5a3cbf6f887d06b8ae43bc1799551d552a7d168e6f9aa9e49e2f8f5e82fafe5b3dc3b2a9bbf3457172b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8d6e2a15dfedb37b04e30ecc72db784698e7c0519ecbe7989b5c5287a780cd44aeb4f31a7bb43e0c69a45071206cb6c13266590ba3a3dbb93b0253285111ca07a81bc520c2dd258e01fc16ac8caf5fec44d034beed8424bbf760e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h135f5770ca9331a753915c3d9dfcbadd3552093b67ed3c84a3d58255eb502548b64ac0ff3df0f6e02ba4805c0c033655311d0d9786743ef029b1388fa155e0882b7f9d2b2e70e17ed3d31036e0ce142334b6287f21958e6785a5c65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h901bbe8e7e83f72b39b332af54100d6453208fd416f7c8c2f7e4f193d4088d7471e7722a4dfbbee8b8f369779d31a27cdc7421117374bb0afd7550255be6ff671c1e99e652ad5db23b931ca0baafd143634011d14b27158f567ff7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf15af3260d8f9fb1cfd1a8e65f6922297af8eced597951c9db4f68f2bf45f652c8f4588a0e6d73b316ac6be024303c3f7db7e9968f6420e962c50649b8343fe9e25d730ecc43a44be83814f40b70893fc8df226fbef3c4813f8668;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11feac3687a0a6d17e6e44c9b63756af8bcafeb9a96f15ea41f3731580d7b33be2feb2949cc0735d85839cc7edef071b724a5c2a3b14321b51c03490a0d6a1f460b5b980e80a6bd16b835b94233d86a9ae47a73640d7b608b2ffdb5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7384ec95206115ae1c2f661678f31cd4e09a6c59b06ff995da27dd9096827785d20a222571954a1cc31cc633ebc9ab5fa42b1e21e5e511fd9243a0e17747ade4aa545c4db0f90901c8bdf80af490859d8fdc6ded0a931b8cfc41b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f921c4a49f4b328739960c8555d44f2dcc44c84cde40eeb7e1ac4e8bf482a9cab79ba63c13a1cb73d6a2ef434d1899137fd5353eda8fc00317abf5e4a88910930b65c373a2f3658421a2eb00d5495d6f2cba6c61aab6f69997d75;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b46cc09ac8e19b4c87b99aac2e534db9b1d60bddd6a2129fa6e5add8fdc2a0541dcbbb53a2da8cefd9fbb352a1322d0807cb69f4ffdcd6efad4c6fb1671fda4b2b9f9801d8312a110ac3ef0e75fb9e4228af1ec429ba6f1889713;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196ef83ef150040f06b7571889aec2e30a6c323b702261cc8d623ea55035b315f81b1bc39102f198ec0496f462b9758315879c60c883dcd1c4c0dc8e6a6bea0ecb41320d24c3b908c7de0a57bf7ff8dd18dd43f3621184a38e55c91;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176a3135957c53ec04bc7b9949217fd6e803239a76ad2b1712064f4abb2037fd2a0da6ee26e4a7dabcc4587739e25f84a129018df907322611b84354d7bb459f51991bb93d6b9ecc5ce53ea699072ace8c3fccba6e8fcc418f6a312;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h738b0e94c0b22e7a226f1ace8ad9244b866faa15590995ef7de73b856dce62ed3b35042867da8dffc418a82cc2d4888fc8323f538c8de87f0fc471fec3d4147e2e9868d46a649a9f3cbc0e5a91440e1f526474612108930680cf06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ddc417438fb37fae90e60863cb140165cd494dcb5f8fb5cb7abfe3996dbe3e0a1d69caec12bf8b96213fa8bf6c4ab841d66622bfc756f13a0c61a5453a984d3da406c3be945e267b15920bcba043e9d6e0246d8939cb5a290f564e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1b27ea28c76da1b2e4ac5aabfa93b30aad008a26f8718233464f4e7e7210e545d47d88ef90dc2d78f93d7ba62f026b1c46b00142883fa4a9e5e82b0e756ce38dd8c9abe8c5e5921a7ed26087cc0f20140fc2abaf4f1ac3132ceea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cc1f0006fa17f5e92614e1b1e54a334ff0d5a1285ce2ce35e9de002675fc10eb6aff68026926d3e857adcb8b7de51d1462aee891948877c8920375bee3c4c11a89035dbc54b26442d0a505654b6ee38122ff2b88afc5453f0d8fe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f98f28dcd3565575c4434601ac7ef602cdf971bfe8343fe6dd06529ec5383d4f231693654cd42200fb8db0d661ec748217c462106e4537ac5c052c64936a55643ff2c0518a5a64ae3be6f5109d96e4cc3f5bfa7279cb631cbc9928;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb3d18b511fd8bcfb5ea7513c0e304005e826c2d74969dbc927a78a5188043c97c2dcbcdb5b54b3f685d9a93e5134a5dfd4ff5bd20837f5ed4469fa2dad7bb9a2b3efef94fa7df73adb7c1412a29b6c28e0fd395b5fba6f1aee51da;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d82a31b4286e53d4e831f413595218371f38f491a53349c120b34d0a6a2e9be162688d6e46c0b9e73017fd5cd7926e729863ef27b51fa2df1fa78bf94009e976ebcfffc95f4d66d2b9913093c030c33f48e303841203ad114bae1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f267874d039333ede98d375af6e71f37d17de243c256c250f4731e4ba55f1d6958a0b6dee9fce171d67489b2820a95876138dafdb026cc25a181f9f7faf5e2f6eb0003a10e7a5930791b842ca171e67df54816976f631d0224567c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd5496e3083131bfcae54279dfcc5dab48c1b90194b77b421e4697ce1fd4fd7812d9daa11e6e8b6402d6b42c45f05a38a1e2c3808da1ef61b25abe190fd225faff882500286f369881c9adafde6880e93750dad2b4e12d2c7b66520;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89eee1b6b2ac608a87dbcea5d2bab79b6b4a82f51cb6a125729814de82d23a60a011d05c41cf88ee3e9cc446a05ffc1ac6db8539515d4ab52e33572428187e0b771b4b279ffd55ff49ec4db7873f863a6cef7b297093c246df9041;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2af1e2b11bc8026ac4e4a25c5e8f92b579ed6623596b9d505f2cda0f922e247fea00c56c11241cef5762dcd971782e603561665893994d33a390e79658677d53d75619d36ad7c7e03c478a4d2ec21e906dfa7a664865e09f17178c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h101dd90e234c52c07227b2f32dd66c06db834a74d5f6ec3fa859a388837035ef3bb996d0549ff73db659335c5965b54c76bb39bd34b1e411470ea1f46873a2a492c6995fae698c9c696a38afb7615d2413fa0022d67552a6d57e10c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e556e7b0fea48911a80fff256e04eed5333074a4905a6add86834867b426a1c0566dcd94438c1762ed58314a6dfda91a46c76f70fedad6a8c63b046c21c4cc201d0b98f29ab3f0367ca8c0c91b528f0cf76949bdda9e1791390f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10145e032df1c69da16e2fc2c162bbaae76e63492b33505cb69952192276d1486f5891e6bbaeb1c347a7938638d1ae6d872fa1064c4eb335075315f346e7058b0d6f890eadfb70a370842f3bc52111b4f2d016455a96b39df9744e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3558dde1bab26d994c7b941ef0cd5c1cd6348a4fb2e568a140cf8a3912250f5a45f20482431d114e417876b77afafaca408a07c449e1245c28ef89dd1fb20d01e723a079ae6a6590d65dfb5a687b6c8dbc71aaaeee2d62cbee8b57;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h826928e40fa958f522a5756890daa0edecee308a6269502c5195873bfda69ff2df41728d88aa47fbb41c47d4b1a1e00377aabcb8df98fa189172db53f9f71cfc6584a77f2b1f71da8d57e61edf5782cd7c67465db9a483b33e14bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c6f0b83bf6e8ed879fc69a55b464e3155c78539bf517a72fba288e8e9725b5d9112e7a3368eb12d376a26e12c29ff8817d65fd536e5dee9904a314c39b03afa471792f1d2681a90a191e686b9b52ce7a3d79cf1d566b9c9bdd225;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e3a1a1b90ef7ac05dd0937686292ae79aef8a8cd8ccc05ec4142a8c612100ce8a500566c5fef5d4f5971354c4014d585509730a20661fccde405cd9fb09b889374a32017bfcbdee513aa48e6094caa0facb40f4bf706033536e20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h257dbe50f48a07c447d4ffb10cc6059d8c4ca5e1137750ef3f291986a99958f2dd5d6c7764989aa8dbd52f50fe7e383a7e26baa7268207953a7967be1ecbe1945a2513ccff39b9dbb814d54bf311de302b7dd1c2b807a25bca0c05;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h236077dfe033c33b318148a6f63c2a60d619041b4dcdd2029dee9ccf4ead252f0e1e9eadb111d321110ce1ff0eb54f91422673ae532f315c012933d38b0cc9730978f802acabd70cf4eb3f1bedbfdd2244ad16def154b829f62fca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1471c95978e84aeca9cb1244a79dbe4010ecda4e8d14fe37e981bbd02036446d493f2d865908188a91930f6d2f9a2c789ac37445a3733ebd7f3f4cbf13464f721151d0a98d9c63f1b545d5f03836601920d8811cd6f4fac33dc1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f05056771b479f55a3a7f775c25954a26b90c64a8321f03e8d68d17abaaf65ddc41563b15698942416d4cb39ca86fcbee28321bf1cc39095fcd91d8509e28927bef11f05d054642047ff6f72958dd32811cdc109c1836535078044;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc281572b3fd56dbfb7112e372e34168a2882750759f390f8c3053fa3dde4f4f6ac0052c904541106ebe18cdd2e0dc6d45c132766ebd83fe891db89652b5c49a1acd84318d5636c55cead1b487433917efae0d8c3546ee1265b1ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a78351d8fda6a3248612b216c6c110b6d15059b392aac7a357ca1dd31001106f4348531933bfd08407fc45669f0a69c5a055f86c972073312b803395c922d6597f85e495284d4555402fe751c37a15030ac7879c859968d53742c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197cd1a93e26adaae9c7cb692405a7bb165d5914a2f76fd377e691d5f8eb2723fe17b59f428150f6880c71a87863eb69c382e1e149a18093bbc61350c9f32a329b45283b8c3a22cae79b6cea309b5d40167d21860b7b9eca33799ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f4ebb9ad47328ada2c987750ecc82c2226e7fd173743a7f9d4f1d43a2e5c5642bfaf9c72c30f59550277c0669c165cd7ae02e12d059d39980e6cd9f5a4802aa5575393653d4a258b395b484b2e0cfa48bc587dc77af0b8005f3627;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5969b68f11ff79cddf9deaeec651a0f9358f1ed52ecf71b1a2dc555264576aea741162881c6c73e8e024e493a5ea2160e1ba05dbb435b0d6d7583edd1d3798c4f0ceeffc936d1317305b4c4a22225c8697aecc851fc6b9de022e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1628f275a8444ec7f0cea43666d8a07fef119cf9909fbec03b7f89e1acfe178da4f25aafb58f3d414d95ab958abee853da8cabcd84ca87f48c4c66b950352e4170c29800a4826ead63777f3d4ca004679b4a10848b15fc98b563829;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c60893727a2cff85f7818ea47ba6ba073f67a013707195df4118599a1a84b04a36880bd8e89d64fe7605bf08c7f09708775511f19e1d696d2b31ccf57dc7429210eb6f2778927c588f990ac20a48135c70d17cd87bdb17a5c1cf1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a9f604eb96c15dd3e475be057e6c1964cbbfde58071850a2dc857c61fc2f62e50cd1f69b079b6877286c8352088bc861a1d29d545da9a456fa2195e160fadb3ff78d1430b6b98d0bc508b2f59b19bd6c2671881c4a953d8d6babb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1894dd15d17649a4bdc257ae22dbbfa6bba85b2fee4e32f169c9059fdb95d5088647f536b6dc216d3d44708e5ad7441ab2f440429c5d203f0ef3d188e327cf4a175b36d328122f17b445c3415ac9efb2907afdf4689655cda6f39ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb2da1f6592fef9e10cce61748c376ee7dab81c2253d02e2e6a85cf64c3a8f54f18028f1af62b1f2deef1689c236c01e8ed74be12aaa91a9848769925352185d0e0bbc217e2c24b212b137926f842dd4c7b32f6c254db82032dfa51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c05c75d244c6403171cf2a9406e2871169fa3f18aa0fd43d7dfa3437ae33f1590aea4ae0f86f36439ec818628a0733df53e217fed5544528f0808de7a1573f49541ff4782f5efb63c9654c529f16341d928ee81c40294101099777;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h154fa8a4da7cd1a5673d4d716ddff951b3546f2b4ca6318617e586541cf517cfcf7270eb95d98214856ce3a8f4a0991310acc462633cb0ba3d52ba728e4d888175090b284f522aef34e61d0dbfc97cb4c4f016bcd9169f312ddef5b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9301ba3bb92c71a6720a92072799cbc2a1348bfa265ba599798671b754027bf652ea6313f9b29ccf232dff367db0a8165fcde259f6fcbdfcc3d646e519af767947be3381a49821bc4550a72d2a2b750acc23590d7ebb87dbfa069c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a84e7325b2c98da9cb0280b39b1a1ceb534224f2656b3e023d29eb97e16317590729e2353c0381486bdb140846a316fd3759463dce70a4790751d022c7ed1ec4a9216b8ab36a533ce4db1f0aaf19c85adb03ad0ad7ec95ddb5a5a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c86cad4bd055d592d59c9c51845d194269c441b99d35aaf4dd645aeec815d1f14352963777a95bbfa0446dcdc00c641c4ff09e555e02057586fb78a8daddd03bf9993b6bd3931eb3d042a82eeb540a8f08e9a97e73467a8db4ec4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1313bfc3740df4996378ad0daed789ea9e83e03dbf1061b0fae8340969175c50bcdb0c8372120fd21c23109ca18d641b399cf34b6fc415371dd269ffd968915c06af2058d1aefb54a2aa26990a6d7fa5902d5183c5f75b55ad16d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf22418145f2ea7d7602562c8ea094930f7c4ca51cd3cbced8537eec202ae653ff596340cb06380e978878528dd33e231d34f37490b54930331fa016731568a2ca236feea8efbde28773040a23453d73e028e2142a46c2484aff505;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14365c997e1400aaf9dae01187dc86673e00ee4db7a96dd1f320a02ea1eaea2266f49d3f7a7c0036f9f1b96a36058c5ef96537bd428057563c309a70bb2a252e13b5c35fc9b570957097018e25ac87087d05b4a92c73b90d6034227;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170924d28b9c867e239ce93346eb510256ee9acdfbcc70c528a4211946304967539b6337832d4443570f710429d296b71d27f7c4831ad074d504fa5c76484ccd412764667efeff11ec55f191dbe8490c828cfb2aa3ef5c89325ee13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58788fae10c6e735119f0579b073af39c8fdac1da04b8ebc62309950023b24878cd1b7536499e4acf7bcd2d1fde8b5b371a01db10d642cd3886449c03a1df37b3f1940249183349a54c7ae3d82bed2666b8b01fc39df66ed7aede1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121abf57370cb6eb0b6e1f52de395cbec608a1ab0109e44e469839dd825c4a8a9548460c6fa4127f812a26460728098b90de79c67c1af82370aeff3ccc4b217c7ec5dfeda31d6fd57e23d6bd1958dda77125ddc8369899cc17122c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c22bd149f768950ea96a3bab6f909a7fdcaf469153f7cf8121becf67723aa8f263f7622a84c481d61beb6c1f682be12be63387caf09f027afd13e7dea16d51b628fdd815d91e6a0c84acbb81419d18c291d1b1b1fa65fccbe9ba5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f7a5b576beefb8910d0ebada9589b27f4cb2c41e2c975287669c96ef6a2b9bdfc03fce1a1f062c8530033d0a44eb9106c043d2c3faf1a9dd9b95faa2cb8456563c87e276290b78c3f6b4554e9b4437643ac728e5c1cf3ec2c27c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0c783a96c1d395c72d2986e86e69f9467652588bf1af6fec62cf70e9d5d9d893b765b2efec3cdfb85700700eab7f6294c89037b48937cc41d465b38fe24063b2db7d675fbc406b93ebe9cb3b3998fb9c1abe915442b1cc0e28549;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf60f8dd8280d4a81653df9ce93e9ff702d26d75b46e3261a8ed87ee39ec9628eb5ebc9e01140f0511bfe26cc93bd39522ccd88e29e4a1ae388dc1a108592c32fd628e09691677809fbf1991ef6a5f68b17ea3c66c534a6d2e0b6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c8128c0a64eeed746894e094dd3a9e8ece2f6eb448757a8910cff22d9a9e91cbe015c77375422cc8bdacb2fa3f9158aad0fea573039c6f45b71363f19a19ec4e26b94602938469b4923a2436bed95347e867b58bef8b8c066d9e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdcd53c7db50eaba94ab2c57188c0dc001db52424aa423f4c8595efa8409cacac361e155da3e64deb2aa8729fe64fc9b39034d7dce54a6886431ff767d063543515fa2bcefd6ee2f405d41cce650ff025e31eeee2d6550bdba0d940;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa71e7eeb52dd3cc45042db5fe3d8bd558d75fef3852aa6ea691d3036cbc0471ceba5fb4f1cca71df6f5d320598e4d6f3eabed4116bd4a43441bf8b4b0258d7b5ec19973d829eab17da19bd1410fdac544e04ba045c1e298a917f0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17106cd5ba97799359d6766644a7ea9e25cfc5c8182ec0b4769c712373eacce4196785c3567b88288afd03d0e657af0c700d815bcc2c0d0586ba1d44e059a9f6a3b57ecfea058d877c6d3fa325017f2c2fb4f777132a8d208db3bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9232d8fe98f229fce448ecf0592b86538098bf505e64b511c1a7191fe2410ead3f650f8e53f08dc9312e286cc188a22f51ed6cb82525846138c98daf5b3e129cbbf6fb3d97ac1f21da6bec1c2becd07ef76046a2a04a043303882;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf66991cba805e0ea699c3f604b1bc52b72fbff3b5008144cc0f360e7b1e939a3c60c38087caad8d594ec88fdb59aece16c4317e43c6caba53bc559b442c8ee8bf201c244245e92e710917e533a5351bfbb649d680486f9d3110eba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h163b904c44d5d28a458981534a58140548fef33e32230b5da54949aa77a988ba761388a86773758489e153378aab2fe832939d587b19e6791501aa556b47a97d6ba84e340ff98ff387542774eb2acddaa796b589a9951f3f4cacd51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1becc9a59ee37d6053022092a30b4f50582260503d60fc09fa666a52d4e0690fb393945f194dab9b880e16dd6233a62a9967911afe154d8ad4b2dd16ccde5635766b23f37e310e4b45f8acceda6dbcc26d423102d88a00f70ab49b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193426565e45e623f935eef6cbf8dce97219dafaa108592d307e15f231258f385a235eaff9f19a1173d35e68e0eab2a03b886fa5ba32a84a8e8b753e767d2e5ef6223d049babf0a7509a0e4ea78797a50aa57cf3c97f6373eb0e0ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17290127c6c2a6a9a0446cc8a2a8431ebb89935c6e3e30d567ca2c147353e05d689fc132b9b6947c29062ed7b79773982433b6bf06b94ef0bfb720f457cd431524acfbcfeff38bd1ac8664f992cfdb1f8e6e88411ceb166d28e1e9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce1908d4a9c218f9bf94a15f3748b7504c0f597cbd77b1d8e908d1443e709343a938ba228acb8f736bfcfb7914d7c915fad419d9e67869c404b45aaf72e502906fbc286b1e0c277f2d46fa84ff51b4f3e71c9c0bd8f8d4f83abf6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5286133b6ae004a28bc868278ada5eddf0d1432f7a910fe65a8da94ed63d266b00d65e006e7429cef47340c584608f1c598b39851d18387de5148e3b433796cd03129ae25d840b392f4215fd7dd3055035bc5d5dead11bb2af084b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fc2a91a69a61ba0bd7d84d69212b80645a4da943b6b0d86c8ff6e0cc6ed9d91184d036ffd44f78af6e69157964c3cf1f7cde642cab758066a97c9ebf19f4225327172fbbb947281a1f4d6372ff41130977cde08a10cd77c713e67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35fabc67219f167afffb82f523031a50d588a7d012fbca89f508ce65794cc7b10b79c72da6ce860ab7c6e6b8f8b6edd460b278705b75fdf74661755d6d5fe3d3e772003c504d7598eb777918f9490ca99444619ebb479682f4e9bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c5232a4ca224f951e37daf431e6986c4534ba0f4f5a6f3d3432c165fe512373c5c9752b580750aec9d4d65078fd84a1b51264979f9bb24632624ad6fe7895cf98c90f365529cae076f5ff559593c812f55a6ded0504635b75f7d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h307704534050b401116421baa95d128efb18ba13f43da084a994f92aefc0d0771daa64455a102810f3235f5826cd88c1eb3e9c2161e047007510514fb6753aa9753ec9f90a3ddb89484110cbb7cee5904e0753a383430c986cfd3d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f852d82461df77e39e6076dd6a549ef6701f84311d04f6a63b3ecad4348c8fb006288f5c4dd050ec12f2db9061769db959720ffb25f19610ab8472b79a00a6416eb431008f6aed8cbad8aaf8d34944904161347f2cd0304627bfd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9dd93cc5d5a8484ab057f431dd9dff3cafa0f2a76a199bbf540e71ce9b63d13dbfd8fefe33a66a895cc157c4c1d493b4e7a6439f83d32ae4496b399d8abf8dde1c7633101098ae5cfc069aa5731b199d30d2f8a61a55c7ee22db5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdcf5c9aef62420452020629b1bf81df799982c00557da2dd3f4fd174bc17b5ac6d124da1364978e6bca1b7d8bc3d510f43a0bb3885db0a87f7e6430c16988e5329b0771c945546c1590c36b0e2a590c465d566261b99758605003a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc54f4a69203e10dd8b059aa01c22e655d671e883988ab5b956c43b655211b0cee1d50c2ab11fe08f7aad1cd588159e4e73530e3fc2ff099c0144254171c594aa495e4e10f9771fa63bf0e36f43e0bb6f63695513111b4d4f0e1365;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h205e05ac9156c0df30d0c07d8a9dba7915d99ccd069d41d573f5e9c8209698d4978c6b4aa782e88f073084a5468f1853b07341a919c32560a756efd0929f05083bdaeddcfd79a7938f0ec600d0a4f7a10821c26cba39f095888b97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h159794e5719c4bb2ca0352583c28f422715d9d1c92298efb67320f1ba9e4c78ea9e74b68ea2df84ad631fd9cee7a95be9fe314fd5bb357891c7ada7ca348275cbd9304f4714fba64e1a956b5d37be7b6f1e5847f29569caf1fd6227;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fbf9ba4601c914add989b239f9f84b2e4349e813ac72a5ff15a47f8adcd0703384e64ccbf691e6ce8fc2df61c0c7cf563b8565a34695d3e2d64b25f41b471c4a56c01aa69d052388e3b74d9ed634e7de4a6058f4fc18d78de8c74f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3a5e22c916d08fef839695542ccf4086492ba972b5e8288e45e2868e6107914cd65542a14f6cd86ce88534334654e098326e76616dc63dcaa4a5c4531e5d6dd6c6ba34df679bb20431bf4c6a6e9908ae851a00260faac3de721098;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad36355a424b1ca15a4f4cfe049e212bdf6846cea84ef482ec7894d9cb5b16a500432a4ca48c66111df20bb45add91dd4c5e46d0a458ed9d7344cd7228ce701d17d036a7d6258fbd43ad7bf44c5831a69a8b1b11882df965befd65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5d48899026675dd6b78c485b7c09a4d36e7196e0dca591d51338284d15ea91c4a257e8d5df76543c13eeb5da6aac4b7cc279c194b348bdfd5b2ee0f3d78c05ce651d99a441f3a6827d99320d1f5471b66dbbb92bae11ffe8649f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0e598082a195d568b0555db0bfac1a0f9acb19b236ceac34c16c0d03d2bf3e783e245155c06fc5579a28db5d237bc6709c60b8cc483b61994312626fa8bfec0f92f7c40a7ec451e5ce08b6ec7e44ee462e10e78b874771a2d3629;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38721e397ea2b7fad4cf48828d2c10e2917e75edbab2774dd3248fd313005eca309cbd99bc742b8332489cb47cf758f6efaa334a8035d589061c9d8a42e04ab23bf59253f6432c8d7eb14f89f949160ea6a5849a3d984e4e409d8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd97011ba130bf9771625727f276f419d5f891bd02f75a64d3e6586b39c90b38660174cbfcfe2827d88aea2ed9e557836de1b025cce1144acbda1b58af83665c31af9e175f92a40babec19e6011fcc151dcf2276134a182098d01c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c98cf055abe87bb5ef16e900fc194073644356ec054e721f285cd4e3bf8f8943eaaa635093d29a0147539848eae89b065eb9f66bbe005ffbb3ada100335d7391cadb3379f27098b46cc31e9cf2192df041983a517adb283f8ddd7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha0884da9c538eaebf4ef21ade8068f67a69036b3b1adc196e52151b1cb5a40d9849e5091225c2262cc76407a70e42321a9a61c9bd1bbca060e3f9024ede0d7b42080ee67da3c5092277d7f3b884bdc50d84380c2303dd0f4adb0f0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d8a0b67ed58c70e096b70ae632825b4be89ea362089ef18f8ef9f0fbe2fc5f997c2b9f2a0033aeb59be94703810438b23cb86bcb17c9efc9b96da5748ecf39e0e6333be1c50ca6c97623874ce69cfe69bd923ee6a8d41a995bdf85;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182842b31505e7d51f3a3dc9b47c8cb4b5b5b3e2059629343a97be6f01fab837c9f383daa4921f35e20110809f31e8da72f85bafaccd750df9349fb2007dee430c6512626046c12771c8483d50ed02d7f5b91f7d37cd11442c091f9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h775c3bd1aec6b26193b07175424e2006baa9404c2d56032b0f29c005e90fc160f0b59fc4aa77ba096e3dbc7280fc748a4389ddfe15a2a96a815f6b0c632db61aff5396a12d53784c8809161bf89baae4771f3faf4b4baea5fc5a71;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1219ae408fa58836657ea7cb03530ec929833e78760fc85652444842a1105ee2f014d8fd47d2c4fa524033ec687b175fad820157dd1afb218ce13b2dd1b6492d310348bd749568abae571947d8d220fe068dbdb823f311b57ccb368;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1815cc3474c0914d6ea6deaebaf205cf2010e184a3620480a74101554efac2ff5fa1eb38d31db40cb3720df72350f4c26cf6d55efd793100aecbbad7f413c7675db51a64181c7cba24ba1ed3ea06e5eed1450c86c28104e49d034c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf5d109ca6f9c538975186353e229b18bd9a8ec13b3604350c15c34505f23698503a6fd408b4ce1cbd8123c5f2637d783cad2f199f043ea43e0dcd23daf7ed3f6c40322f48202d5d4a064ffb7b24595a9e3858fd47c502490bf3b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c7b3cd54af2786bd59220c0b3dae5d8dfaa1c9d88d6e3165020fa6467a66113ce68f9affcaf8348c29300d10ee2443e0db139610ef820fc2036e416902ac8c739d1cd1b272fddbe8cfb0c8faf3e6ef0e23149e8968eff5dd84c210;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1f895dc821cd2a3281112af7072717e50de949a32711b48a181fc34059a7e1cfd966d4e0690c7b152a0902fa7d93f2608ff4f48ce1c952d1d954edb5f5e22c5784beb29853b575bee684c07dc1d399ede09cb7b08e5e9bee42c96;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38a8d6829afa4e17b39dab7e025f0c9b737bee5fcc4568d079ba117bf785c3890401cd42c8f16efdcbd8771566f09f9d3cc79277bbfe4e075bfa726a0be5da9655e8bd67180b3dad2233d7f13e47fe4fb2477601315e6745fe9dc2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5bcb3455766d5a008879ea65030eb93f326545cad5a0e2f0ce9d682299c3d65503807f4f0723f6a296356b65ee0dc5913051ef5705cb84592ca9d12a93cba0eae827e866a4c691cf549a450d5922dee77f9cd754a82e08c27d699c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3cabde87c48e22c57e3ccb85b59ce0547f1ae0d83ba0894fa89a72e3b434a913aa18b5de5a6bf02efbb8895c9ee2c3feb557e1514a8daca7ab671b3ff34bd758268e58bdb47932e401e33e44d03491a85fe1e3ba156885de5026bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h747c495f0110815c100ef0216ccce8d8b86816e2d5a1dda2ffa72fc32d222027f94bacf6c154005b5cfeb94c3ceece6d42a39f2e388382f2c58702e306239f3e682a12e7c608a7117e603c9150f120a550d91b160d8d173ad3fad4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c31e5d6ce1fd784128ee6c1729555f10a89b9e3b883865b0a15c69f7dcd0dd83843eef3c93013b3a5923b017e1e2997dd980fa67a311e2da04b1054e68ee00da29e4f9d5017c96cd4fefe73c0746d8e309275592656217d4efed08;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bd2b1129c94018953daa9097747936c016772c324369ed7bd7229c5530850340bfa47e0a3e77bd7342bc33a14f77ac7a51cbf5bc1b134eaae4cf1d7d58262647004d41f7d8bab1b704a014baaa04bf65d1f71e3a44bb09a3ad4488;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78abadc61e899c44650d25b7e245992627e64466374bcfa981aa2edc7dba7ecfa1f12a5f39d0981790f35aed1c28fb0577857ff950ba0cae8c2d2af9e353cfd7b08beb93d61b9d06fbe270801b4f84f9ad6f38f0fb8733597832af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3975cdf4ad017f5e2e63a7419e723c9f770b904cf77461b113a956f529ecd6068094e76e8c8ce21f4346f88a8dc647f48a7ab90c47cb17fb6e6b30db4729626054b5286f0979da43de9b76c1d6b4091dfee703f7703a444bec6d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6fd20aecd3020afb27af42fea3e118873ddda1c23e0c89b299e323817d5bd92d03c6b6979b4c9bd73177aaeeb133bdb356c08c1b83d598f6c56aaca6947f5c8756b1e8f690d3de70406f7a766fa4f7b6866c13266077263b8deb9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff818436cf3f07bbcc5da0b06f293fa220b13495c9db010a797ee17672d6ef016c02511d407e23ee357bf18b127daf1b82c036fdae3920224cedb0176462438edb4f3d8e72319dd1ef28f36d050cc426ddc24caa978a3eb3174714;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114cb1c61ebf830fd063b278675a2e0abebe5fe51f073d0f4e2f8427694aa5e5bdfadf93693a445f1525a8d32e4df85078216f42f88de97ca3d92cfbc41138932ee68871ba6195f2f4e5786fda16cf0075b835397b08c1d65907013;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d3e16e9337388a3df95d428b10fc828a7581e9d9b90ba1a9c221efce141cc337024187000bd9a07d2138b1c65cf6175de254cddec2508640b3cbaf93f803e5fa70731dad1e7878fcbac662a0e32469e363579686e95991f953cad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9f6fd18f46fd225312b7c77ce9f2fa4ccf88b8e855cab7c6f3e1aaccdd4dd4d92e30d8d08aaae0a68e5ddd1a20d30c8851a33e88865a616972603faf06f85c85884d5da86da86e1035fc91056af47faf56982133ad58eb0edd3af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c9d3daafec34629df9d3d103ff82c4be54394cab21356a838c57d1f0e1c516ff71bec8b87375bcd2928dc6f0cde05bce80719e4bcdf30dc520340ae579095d8e8dc0694fd8061164ec396c715af085b199276f8ab0bf3fec772faf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15685c284d39a671703959329971c2940b86375ff88c90b0715760e0383517913cd6645cccc5ed73b4add3bc0d17379fd52640cda373d87dade9aab494e5b6f6c36403c7515b3d5dfa5e704ed31c9ca4cc31b406eee034c0a1d6543;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa8b24dab636aed5870ae863d4801a0bda02d5cc75d5818989e54f2538d6c21b0ed80841d5b2ca0dc1f6e456260d90919023846233b0daf12b609291f676e95a2c5e51ba2089f0381956271ebd172ef54bd541fdf2692dbce16a2f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc38693c719015f953c13273ddc6ee11b163fca360fe6b437c79216e4786b9bb21bd861636a330f1fbff33efbbc0fa85bf9826a24629a796b23f96459254f625af4b6bae1407fc4be0df0e7c61e2f2beb055e6f19e9a02d5d26bcc4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35267dc7d10fd790ce059b4ed8366abd0243e4c28768a0da838fba029f60676adf98ed2ad48fb8e1e953a45b69cca3560055f29930df962ae02d990b15729810d7232815e2307015e3daceffbbe2e80e4c9885d9ef730a3d8dd5d9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43df447a0b49d096073a27dff21fe3b44d51f1c05544feb0889ff150e5cff3c12cd6651a043b8f12c45ad91c3858c1c9be6ce645c738edb430943f32bb7e935b0e87e72368eaaf5ae5be45b0d46e9d1e4ea56df61f71f95844f25c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e5d5e4ac8c7421bb787413962d23159727ca83b98f50c38901cc0d359f1a68192551b3f31c990ac4765504ad6f3668da24d88fe4c17616072259241330ca02a8381cdf5314611b04b6c0e9267162761126da569b22ada648b256b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hadf99616da0f296bf9e576706bdb29826d8451b60a5f8ab74d96521bff8a29d3325838ae3686d638a25f55c4ca3606d6be168f1a767b6b8374356fb1827f6369ac31941ae568a1b53102f19f19d104634fcdb03e4fc36483c95edb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13fa6daeed3733e9be642309bc0e514472843c51e2c58173d6173aed273826b2dd475e2ea9f3616550819e3939a6a716bf28b8e9cefff168552c03bb55806774740a6adb855e1be31dfb27143acbad06f878bfd8b0ba838b561a1ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7760dbc101921ff39b55fd5e18e139d6cb11724c6cd93e929e5a2e4d6f20c1f4d4afd53908f8ddce032356343b4391ce522d17054b9add186f212e09225057e4e348a69853510caeac5558ad946d5b4a0ee7b6d8abf75f629d560;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c2402bfd4c215ed98a5bb9ee01b5d740623203bf44acad803b249f86b663da00b24e30a2d208c7f3dd297c689517cffbd7ac45cd1d96d52835711d258a5289becef48f6034d29453d5f1351d72aac189a59e47aaa2d2e2890aa686;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he74d18c9358ad4e5ab439fd9105c558f6706e9840df391309c4573e7ed6ef9d8cdcfba4a509d9507ca814290fd1f82711cf70132330611542d6a30fe0a0eb1a37df3a9dab70a0a9a0cfc301baeb5262dd73fabfd9e360dcb55d589;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc0244fa303f3b12ccd7ff6195fa8348a6dfe373e28865b4f31594b1038ada4a8bbd71e5b82800b005a629fbb0bbea2b9d6e1825617fc7b9b9faf900da9958170210c9077d622758255655fec80bc27960e416f0d80f77641882f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24e8c1adeb2bd4d175054247f92ed6f52580f7ec10f5d32a0d5f070f3fa94884fceb2798b1edbd7443980e608176dbe5eacfa658b4e4ebb3e469178dddacbe1cba6e338be8c4dc086b64b35471bd69d71ab998dc41125eb1cc8773;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd6fcc1dc8421dfee2c42de3d4cca21ef045db428b489893cef2b1d7310643dffe9133e219092b14e875d9f07b7801a1d39825762b6044895a47994fba7aa2219b57a1c3f9d90151e0bd0af21b6691f66aa3050207e249d9789e32b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16dc18456d9d8cb5e84746f1501fe4b9de2fa789b4440cc836a076a35be0198fc6c1f442040071e72e9ae2fe90b67202750c1b3dbd85a65a7d6c4c4f879e8be579f4169d7c8fe0b1b7583c481d61ad731353497a383d7453f45cc99;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116738d6308f4f0491d08d125a45d75f73cb10ce59e5ab61a981c6f8a6ce0cf3a4e391de98fe2d5cbe3ebf5dc39b5346d1767376d53586c185c10f68d4ff4d6c2742101efa9077c82c20eae12eac8f73a6d0b35153cacf3c55694d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e1a744a0a2ac757705db99f6ed7c613668cc567736dd1c3eeaac0c70ad15954cbcb5600f9ebe3fb672133c5eb31d8add350cece2e56fe544202cd8a86896034924a1e2a40eba6e45de5015549206ce557b7f3c76e73ec8b9b75b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3b266e0e848c3a0f1abedc215f00792afb569fe1f833a0fa5ca1f07a3f6d0d7cb0f7f12aad5afc6e80f3f0abf030e52f869941648ca64caa34c6aade289d0f540ae07d31ee8c52d87cadd8a1a764679ccb55f524970356e5cdf83;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11431ecd9f0d0b2c4d68893a8da80609acbb02f89e7ee2d182dda902137f559605338eb881dcba9e4de7cfa6e75e075b836a803699b5b2d508a0b1ae76f89cd471680f88758426e88a1e37f40339ffa266f2e7213e300d2c2656d64;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h754b236bcfd2f7a552bc2591d27de6e99fbbd4d75472e7b5eff4b14be4b0a315d2eeaecf8bbbb0bafbaac8806ad944784499599bf91da4d7928a64bd9772a1225594792556276f1ad1296d1fde08dd38ed7e73c4dadbfede22580a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfec1dbfbb8146f02d77805e0f64aab6c3f3349e38330df5c927e19594f3d7d7f7a3bea6f42cd0070cd1fb4bfabf2054415b4058ec3265356f1f428e9cf3afa38f712e9641040eaa8409e00872495d5e11f5dda1e12846567051ca0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfbb90311536b60420425614309dbc390a4559bf2a2009c09925d0243d9be5838dded5134e78c2388b3b9e8ff0d9e7fcf418d3fdb7d73daa51f360b6f73d4a2f17b70b1ed07330813084136878ccbc45ed0693f891b4c7f0b8ad857;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5d60af45aade17cce924093b127e2f871f6502d3636d9e75ab7f38edef3e24f85cd4e1f831b0f0f2d2e2daaf09b249cd08aa49e701460fb0b712b1da454ee7e2031dc47b5d1c5cd1ab874dbbfabec7e8f645c8c9c501bc999ffae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78616f25a0753da616301ffbbfede3bd4241a786137a13d1fbfee84e18c4cb6642b6c4314b61ab32802d4be388f69961b1fac66246afe21176220106abd5050a22b97efaea50ba39e868b52fc1b537f9be05e01433c9de4f54b230;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb1ad917ab78b901fabb897417c5b4fd7eb2766783003dfcfde2b321644b6c9c1d1ee3281798f52bd00e8bd8a11d1912358a05570030552849499be793006d246779f030709fb7d76808bfebd73feb6f7ad438c780ab285306118d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfb7bfe639a9ba116649057b113fea15606c9c79092907989c58547c7c1c93c6b2af9590209877ad18ee1cdfc2b6892244349361a7a7cbd23c10d39aba76c7a3cdda505bbbff2acffe311590b93c59bf14e821cb4082571b71bb751;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha381b864c783c5722afc67947d5a4eff3257797c58c79c39745e5d85913209c6e769e80f348f369b50d075a1dfd253f87723bff2ab245538e02c343181168ae3450de0c9a5bdbe350a1c3f78ea5fcac7e49dfde7a76ff851940a5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7532e3ce02a621acd079392180badc592b2e574e695450813c231e3d4d6d585e9165ee3d60ae5294f7433bbac36148e65311506f70e73125cc3fbdb402a74b28f11f672367934831144e60c547a799381da54847df0ab8f750d5e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5eef5ce2654993dce807965e956826b27656a4918683e20fc8395f58a2a481b3e9972cd73db60194a7c69f05902f7c6d87b7dce43de2d3b6742f1102ef4e9b3960097626a52413ddbd2740bc86089b152d6d3a671e3f1df916ebe4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97d0f22d89bbe3983c15ffb80dfb2579071068bfce3897291597244d3933cb131520acd42b696f946224098d87abc16a6e740ab63da37ced8325513edb7ca56972ea7730e0c005d5b096b5f90f1b4cd893fb9e7db0172c0087e743;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b547764dcd08354e91011ebeb51495bae2a0c45b059a78d4f1573e29a8b6e71e6d6849a9fbdaaf2bae94d05a095587bc18689ee2c182f29c22c75eafc229ba3d6252f9fa9b4d7c8451f4759fde1fcd6171cdf4172961d742e18a9c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfbe43f1f5ec183714cc21603afc1c5033c5cc9b7fee5e790a08956200e93154b821c43d8487d70b20aa5ceb403152d59372f60576faafdb0b2387d356f8adb918d386b43027a8b6f2372174509e77f4035043d8e73a85c78cd0923;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf0249b9d94b859780f3e66a76df3826dec9c14cd9ef533292bddee436e2dbddb0be471f04e8039de7d0f16c1ddd13e82fd8cff8d75e799782b78e3870210baa8580a8317a3d169660e791c739387f5e2bd1fd7d8cdab1768e39252;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c6c29f8837ba6d9de7d5d5dc4b9fda3172cd0b66d6ae619d32560c9649cde9510101c8b1817761ba9227bbd18919ce938edcc5b34c735e612de39eda4bdaa866444e140f50c5a703c5486c908ceb24ef821aca903c520636fd52e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf2414bbddc66134d885a37cb7889321fbd7aacf77297b30e8b42e60e3a27c691d2112f58705a1107bb82ce6a0e719ddc1d1c22b15c45fdc2633f2d08d223e47ffaf4fbbd1d550b5b7fefdbcac88a8ac6bc637de8e439e66da484d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130620f4a6b0a7ef14a35282f950d0c2254a23b7175618ac9bf951fb7f32174658656edaf5a8bba8ec81cc3f913e2c3e9d7ff56bcc980f6d775c0f5bbe0fdefc460a266e06946ff7feab3702ad57f8be2403922ad931aa08511cd88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be5c2a45e32b9655bdb4be0c6f76653cbfba8fa0f51457eff718f3ee2202b3ab7e445594791cf99eb78ec8b751421001d1e760687216baf023eb88854ca9a64e5a4806d7264836ea334ea4716486914458121d6f64f1ff92ad4520;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1852ec75e350c76bb1b25de7f7a31347f2e4fcffd6cbbde1d4aab74c904dce85c4d185b767165754c6bb10113cf16d2abb1cc3b1f2dc0cd4fd68d541fd7e777ae260d9f76b134b2120f0b0ec7bb867fbec1ef2c3f4f68fe41776c5f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106b240c3f6420df5930fb6906bbdb4bc16041f3d4eb485e10e10adb8f5c40f134f878f16a24fee266d47179ac274d5c158e213e8b02baa93929caccd1beedc4f9c1b8f75457891547ed51f580ce189f421a61d0329909372d4b380;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153e64971797459b7df33c783796ed34ce9930343ce048bfa543e76f89570126cbbb14992c85df9bdc84083d524df872a093fd02375515e6bffa9989e929f41cd383aa7a71bd1625753b43ef731ff5577315a23bb277a56a1d7e061;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h181b1ca6b6f61d09c9371e959419217729f0aaba285aaeb6124d85aadebd27dac75686bdc03dc40b7fa18a0a9b7651d1332fab085f566de8c6a8b865e43d083abef4ba7b51731e0780f5c149e2d2ded6df8f06cd1e2babf4aea28f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ff55ba77d89b209d117828f2ae9309fb96f102e6b33f4f28953170dc376c49da28e92a3381d79c3b931a1f590788aad1f9fdbe1aeeccb544d37e821b0ed68ff79ce045813321609c4654cdd7d31b111e3fdeac5995599b5cb5d98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h349b7c2121563d8af0b752b7e64e9aa9c5be2fff2dc2f8a7e5c7f83c59f00d4a90a44be023115d58c388c4733c314a855ab45739b961609e749566edaabc69eb0b502d37c809ec58515907c394ca4d338deddc2d14c0a34c391053;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5b0bd0e0a1b97cd44802cfc1639b16e7d45c907c920894d0f8f0ef0d477f0ff410c1d370571accb47cb13591df9991d82a90368b974380bc93d53687f91fde19678cc3080aa0f921707dc684cbc350210b869f3fe1a539951ac9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76c8187f2a4597bcfec96579b78ed46468e5b1bb53adaa4e07463cf961612bd35d7df73a4704603cc8d2f0dbc2584f3c9e04c4299836ddff2eb40d51727acfacfc2517d1ec75db819ed4d208a0e5dc274c783e5eb909e33fa84d22;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8ec7ef60f04cd5986439e7f0ad65cc895f7a8376cdb8137c6f9c33a5023a1b455697f4bd00b84cc0c287c0d199a1d982bb5c271441d8a649c504b9ef2c48e34d4fe558ae0bf0efcc159aa3e1a4939034c330cf8afe2c6191e6df5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a28d81e162cb727cf816ccf63987e2168cdd7318879eb47cefab236807d1d08744cf82d1782e2dcbf78830b8aada765f04eba4f7b414e5cb05189e1259723a9386d08633da390f38d4845495f51bc9bbb9db038c02e34da28fedc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8792b3bb15f5aed2be461cfd8568bc3e8569b39849b1e5aa7eb458538d3b0cf53c579d096b5c3d0cf7fc644f5ec617215c58e553ded5613c61c8193d4a396166bdce48bcc99652de746c2134e0a7ee7c3953f63b34cee52a97fb5b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af52e8415c933f222d7bdb347706746beef89c5c19505a93b889331a3e6712ccaddc93b8b7e43df944ef1ca2ae81bdfebe33b1b87a5aab472219601ad535930b58fcc604c40b67efc5a20a0bccc580fb7318cef9342a424f1b1d45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8890497c4d77d171e4663f133767194c4a249fa82a4da7a5d110d2f4d7e7db02c4c8551911923c091613f602a37946a41fe87fde641525b269a7109fbbaf624f8d4fd08cc310030aa50b0cd5207ce7a5453ba0183b0357cb33d741;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h936af7fe138cdfb36aa612a1ad4f7b94a4903f45d44362b9e41ee61df2d0c8310de68705d70bc7f47d9176ede8e2d6635c925caa1304f8da82c0367698cda8ceb9c9fe804d8fbba585d9c8ebeb478d195bc90286477f2ecc972003;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ce219f415a5ff463e661a60668969a619551459246cb66559e5fc6a1f5e2890620a3c792a90983b0c4f4340a48dd16c6566b7b26a9a1cdf6002f2380b5455bc0ca5878aad2aa2c70d2b360d69cb967159eec91795a6296acb2084;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1390f929c9e2a7e646e0f734421536ba05407d2ca19f263c696597884fdede270646336caa3a7f91a4aa79a106c9fb601253025e7a459e8bb3fd7c36f7d2fc8940f4ddedc9d72cc196f181fbf8209f2612df37d80fc30a0e157b513;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d01db631f0ce82f1fe09dff619c394f2fff9b01b5ff1dfc635128899cc05d4233c53836e651bbb71daee68cde968da8b4705887961b2ace817a4597a1bee5189138dd3dd97f677178c04fe647ec46d817ad09ef1145bad63339ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d06ae0841c66073a53ec4bc93af10f4b1f34eeeb753c3cdd5f69d02827b0ba3aef77235fd191cfae346fddf6b31cb45cc41368532e0719b5c3c64a5cfc04996b8f0d9d65200c4dbf09c6a3a08fd5d251d0386eeefd18cc62476062;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h82f68368e2ec82f6f55236f2f64df3dc3d25e7a7ac12b1318f2e784ac2803eceb6ee97016a8376fb8fe80983b8f10e088a6c3574814b24e953a3a5ca096cc72b2f2ffcfae07fea415f1278ea6a92290fbdf096050bd34a46ac9652;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e00cdf0146ba337a5d64711490bb79d920dc8f0d071319c99d9c94f5d98b89d7a03e25f3806ea29ccf63964651a96f0fe7a2cb2d0599c09310b07d1cf37f806af60da665f53bc2f07dbcf77748cb69b6feac7990c98f2bcc00dcc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104d4c622d237471e500ab050f0e6e510649d5d9e3951e107bce4a0ce7781f44977f8b48b08204f6cf89b51d6ddd94216d0558d7f631ca6652541c3a993895f0aaea673f4f7dd8335a6e5f7388053b17cc023684fd83a7b8d857277;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7ee52fffcf88da51e34b4be18d69fd8d791b2f90551143515da9f34c5bd61050150ab759fff0c8e1746df4db8046c09efba885425fbbca5315fa01612af58550c0a0d57cc80390fe2fd6f9c3ceb28fbcc85ca38bd154932d9ea1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e09b5c1d7bd2ddc3e0c067299bb94416fad72373703409ee98bd1cc4691bab5c1f7a41b41630ff573ebbbdc445ac699ba2370e951b2b5a6226e2ae43b4c4a944177a45525331d0c9d01123249ac8912d688c99e9e2144b832c7bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h149db145c60d61a6aa893e3bbd27a0421346d0f6fbda1bc677a5de0300dd970120be9a5ddffa9ae03264a849399e9bd5b4143e8b9b57d55eade39aef23eed88f3b8dbc0d714cd350fcdbd98ab18e6080f09ebbfd780e3cd21b76353;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f445eaf7f3daaa856b86f15a18565b76010a2f2d354d1ce688a04a05e3954fbc7992d9b2729185e3984dcf950bd11007d1c2b7fc6c8726aba7bc48677e4aa5a369e4af6f5dd59419d99a68bb135870ac1854c94062756c2041706;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf323dd6964d692ca369227f22a0953fe74ef3ccfe22a25139a3e49ddd5d76221b59d350708516f02569de3cdc694605bb69302b453677de51d9667a7787ec230acbbdde3ec73ac8a46fe857d2a228d557908aa69565886bf257acb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0284d893deef4a980091a59b6839356150b4cbd40379e7e770146a0cfdc7fd3a9ac7bbcfb13d4102842570e5518fa0219a9dfdb3bbaf539897ce992779773325d9977b1d745f8f5ab7199440fc09824359d5eb88023d6277f141a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ac69b0d21a0c782aa70fb02a6a653f6fb8f3d701c22bf9dddca9c0bfb3f898a6494e00cab2787e910fe95a7ca42965dd94e7cdb1c2c3054a96821c7856c1a8e830d934ee72450a8d78ca5848fe16663f61029cfeb3c28688b6b677;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1773907278b3a39c6cf9fec562cc2e9619ef173fffa47549da04e6d6416b40048ba7da7009321294e78773133680460fa231051e644bca4d84fa1eecafd722da3cfbbb00baf4518f071dde7cefa69e8ba079cf739d73eb80cf37f05;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb89b57441408c44b470d58b1d9f1213260055cd2d4bb26615f88c519be1fbd3a268fe71d1293e5c6e9a14cb9129c1442ec05e8691b398cd96cc76108ea3d9fa76f8af70473143757247664e76c7c6ad49e0dc4c7161e4d774ac944;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1098fa7e10efbe5de6e8ad5f428d194e779167d75e2acb8bcc28e35746bf69b14c5bf86c7cd0af02e1aaa397e3404f48eb780765dd0a87bf86a9816aa7e99ac956902960b99cb8e907452a25c74e8ba9cab2521522c7636b7dead9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167331c63eac7ffb09c48c017c9cf074d0f401c6477df8538162e33ee150f4ef662438e88e38e84b99c91a924e3ccb3dbbc875ab27fd652f3bd1e47d390bb5d9632086ea6bce6cbc39020c334f2777b56fd4df0e59cca997fe4262f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ed18146cba224ace198479daf2e659ad7a5ca15db6eee5138c4c85f518889314937d49efd0a3c3df5a7d561697cae1c4ed45fd05d87dc4a2cd1d40d668c0e206d27ab9f5eb8d517677bf95ad172483f1f658fce0df0d562b2a5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6bcd6ad6958c3359ff08281f6a56b5f2e6b424968305a69fc9bed7d027c4c432dbd42c0cee1d46d3e6d8cc74d1fc23168fbd22b8c8ec13a15e4bf62f87b66ed343b10821fcd2c163cf78d186e5d5e271a54442e93f1f80acc63870;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1756538ec63c85faaaf40e1ffaccbd69d47a488895271213a252bfc0e2b6bb2385778bdec8cc4c4615ca37c524c20de5690770a7de4756f5258ae8f7032c42d582956471df6bcce369c5d76e8049b3bf6b4a2d2c3e0966c59f7600c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f606f6bdad284127626eac09d081a5980c2719e2c08607c30d04061947132eaa9a3eb446ea5b71340ff465a4ad674807b63a80b06b289712c1a1223464d35ac4d9ba40ef35097577e386fab986e58ebf042690dde6b70e201357e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130e4bc7521c5737d5d41d730b7b8ab24402b2b33be2cd75b2f5ae550feef1e3d0dec625b27aed2351d5d669db815291952a1ac7e0453c342ef435c73d751f2337ca10e2585c6cd0e7695b2f274c23e5ae013a4c75ec8592f0d893d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fef308e77853eb368cb4b22627c406c40d9ac5567972f1a47fb0ade388c951ab2d6e8939a75abe8973c9e4bb0695da72f0a48932d1c487f45bd72f24a66828ae037baed57bdc3514dd6d6b08e0b2983c93880af3280df586004e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heaee999786b044ef10a97623d85832d03cba362027b065521942029865fafcdf4085c84fb662e5024c2a72fe3ed970351597b7b82dfdb4f2ff2871dc39e5998114d2f4118cbeff0206ea5f6034170ccf4dc356308882fc26f5939f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b06ec97c26f1532cd9c3e7190964f94a162b2ef816c109350e5d9655468b3e44f097e3a5a04c4da943d7c28be60e9b0272d8a2755e7c35e91a9febd0d81274bd3e86aa44d5615b2a6a443181decf77b6b3e7dad2b0eb1055ca2c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7c6f1c4ca1717289da772968161a7bfbb2b10b2445def5f9e3670b7144a068040f23cbf02374e375cfbc9818dc6b1f7e16ef7f5e06cf4c92de41efef9149bca5e29c55a5352d970023c35824d9f2645122bc027c61540d0e0f662;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115591846e04acecb3f9a6dbfb904350d02faf093d9b30100b8e8887cabe33372e42e4de83484bd500bf87804a57366596d25b87b83d02f37cf2ff3c31a1a8de7de6a69634d28991054357dcf6ebf7249ac3934a741a71f4d27de1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e557f83192674da7dc7237ba7ad13e76108ab1028464c7ef3e819eb758b582b8bea73667ad5251cc80d6a86901883e6afe5f4df3ebb6803ed0c4a217624cc0c6b29604bdf3a9d85bdba637f74481ddf86030bd518e5bfa3bd3672;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb25e843a77fd5a5f794ea60a648703115468b1003f6ad3f6364f2756411fde809f70fed041f17e5715fbb9ae4094e820c0550a7df9f97e2e2daf683ca4231cecbb8a11609f81204d93045df9c7f334bed7d2db18fa4dca93f1c651;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0cebb7be6b63ba402b1fdbf3eb80bf5bd2d760523ead9d2c608668a37beb9dfd0acbe33804149f2cfe78aaf42577726e3bac5c4c829e29e571c04b947c706b7bf70b1e16e051534265db5ae14bf81abb1e47c45d15fcacb9bc687;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16cc39de1ab6ac02ef06e8d5e0c78168640a9ae8a723a8b11366e02e64599bf0db295678b270301c8b6fb5213ec5ac510cf1926e51dcd7306d5893b24ef783223232fed11d2c91040938a1de90019c7f0963a9be028f71cb5241433;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ba914d2dd8d60c324768c296a77b3b33b44137eef2a4227160b7b003b9fd92896b20d7ddbf49fe4c6cf76630ecc73f189ab3e654d97ddc322bd0a597802849d41fa2dd48fc951ee16a851105c88cdc8db767da71840bcbb14f7ee0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h820e7938bd07e13bb65861f8594a1b9deb9bdb88404eff5b88b07007c0d06276d62c4742f394851e54928582ff4c0d06f44a694580c6440bc758d7561fd8702ab31251bd3584b62f08e2b57803580802b9ae884e5bf162f63fd730;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ac54661f15465cb778bbe14ca8bf1a33fa1738df62691bfdc2703712770249a18fe8c98f64bccf9aa376553b986ce605a3661a9300770c768ae821855507877abf735476617b37a723e078ca03514a11cc652085e3f0f6c61f593;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef050c5035827c3d9e47ee80c0549dfff0eb86f12129ff25066753a1fdf1c212b3b14fadb791fd5154d3697c62729f36c7aefcafc6931bb6a7fed05365023bbdfa96f405308560cb9fcaa8cf3729fae305726dfbeb2ab13e792f1f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123f370de03d070eec3c46ff3f36a5e07f5343b8e8a6c7adb6d59b2dd56e9f3ffb742ab7418df711e6e77bc1c568faf6dc2c38d619cd5c176d089ad72768d070962671bee0c3b1de61e24562fb53ef83470f951eb367868e87b3c72;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38852e89e957db35c0c54669f071c168ac6c6dce9deacd30d852063d6130051db912ee8167101f48e8ccfadf878635de2b0e72fa97f77ab54530c15bd482b9136a38b5cd5ac1c15cd29f762a70b69937157bb09a450c40ba81e33f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146d17e1883a756ea6cf61411bf9515e23a055ea43031508643f3dc8ad9ef77c0cbfd3cd498787fdb83567b9b078ed58b2c3645076b6c08214f7a33b994e35ed4bedca8996988f8d2b5e7ab27f0c3600dd8929e2ac05cef4e303319;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f0eadd7f7e05f8d9545a8ad3787b06950cd3574e1593ab8322d729ede43e6aed59b1278fa58fcc5958ab3af573ac9ed68b548b831900c19e162aed9524edf5e8182271b5e7e124c0fff6eb0fc4d86725623a4a6abf7de0a45efff6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173c6dca913f6bf2de763b12239823d247e590ffa0a0c9b873a68e6c437afcd32101bd4be6e7a6e94a3df292097b8ab4deb40f49dc2b1664400a182d4291b92aebf193d4667d924a21978ab30d4eba320c75ae64d3ee0aabd5b3bb9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7af3bd47666179fd15f43cab87e642f282da966900a4ec974dd207031e24a8a279e3a38dd948fc30ad128c26628655a1a1f4fbfa5455c91bef83c717bf2311671da8943cd052557dbdc22f2c13a07a05bf353bf771fb9e065e57f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13942648b601c6d5786c8a6d4cd61f0246e54edf868c0549400d3f17f60521574a607e5244db6cf2e5b2162ab0f5bb13a74b8cf1636114f0b420436c8dbf36ea4d30346b725a80bbba23a12b4ac3cf78669b448118b8f09d8505b16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1638c48db5010bf8fd4e7199c645fa9349e1f5dd1ecb08674a9829f8d473f8adcf7ff7b1ecb2cd155d1f1c6d872b946c6b78bf316f5c9754f7c2bb6ee0e8ecee3f5a8edf5d77b051a70656c70fa546db134819d51b1c74f2657c5ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6514ebc157beefd7e5bd9246ffb2d49426805fb48406212047f98332685479601347d453d46139df31627dccaa198c29d3825817c9aa9db8ab4b0554e73be41cfde0e9b797d2a765fe8fec46c4f157cc14bed0a375748bca9782a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e310860a60804992f9d59e7a9c9e91778ae981d4f60905836b2b7d5f07898c8ca1e482ef613b465fef5aba59269b3e0d3356df987a8ce79144dec1e5917cbd97b5b612d15a781ce1c4574891ce6f72c116747732090d8cdd7aaf0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b8915895ea2144ab3476d05349f62d0ec712825d35ab0897f036ed59c5a6eca33b723c873903f503dbdff98c162e62559dc1b4bc7d67f01f4100d56074ce57da079652a9a485cca62bf956d5cf539d8420bcc9ec51c645381f05b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f0b90e6da3241289713f7b4a152e83016c65d24c442abfb85ff9d0c5b7bd48be2c342db5568709422c6615af7502c4759211955fa63ba9def9dc7c55345f69eb72aa14a212cffa2a7cfaed85cfc8b1bbdb71a17694ec78c154a11;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb19190f13af960ee7f4e9b13b8ff613395649f320c2576ff661e831a635a864284c076a78daf729dbadf6b88b5cc418cbc1656fbf3d8bc8012e3ae6862d922e7e55b711defc28f264eab18bcd07207981c9c0c1df63a7b4aada548;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc3395f69379088123411d840f57d425f0dc5a47f7317dc00ed3c28601d859aab666d958ce33b6678c8fb311085f5c06f5c4db48e2a151966c9494cfb0da637e8c1555425f74e3c655d2ced17281caca249844557ed9f041a27b09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1841ba701f093e51061275ea74a38ef61d2773bffe60e2bd5bdbd45bdb12c31f3c45361f54eea0edffd36a944502712cab91bd163792448dbeaaa9fce9261866980d6ba5e4af8bc850f0a9fb8de66cb89a84f952113a213f7b88ce2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8bd537ef6b055d122ba1b030c867952a929e8e751346661374f49813ad9e43f7adc90218da89afe808ccac00e0b59075e6da7885ac49f5f89b77fdfaa102be7a40745c67cf73133ad2c42015673855020adc65a4ae0a8894fc13a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14508660556e9ab1deb128f80123c914584b507817601459a4fb7b2bbaf060b722f2b324ea6ce9e912ab7818f7b5415617b12b2d0445e7e132defe5145a100baa788d809985b294933a3e8e2dbb3a0522ced4adf35c18a401f8632b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b8a738396cb83ce726e1b0e686c0b00708675a4686b03f0a80465b20b58355b013add55a678afc95aff986a8284c8931369a0b8daefb56acb9fd468e9cd87f898cf72b0aa342f140dd29f6393894f2363dd76236c2dff61b9c22c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd31da1dcaa007bd77a99da5989dad3beb3f5e5c9453e0ad41fa90d6151076a2a990e446d1b6217b0ad55964be3128de66a9fe6248b587b184ef484bb3ee4bf6a08eae2a170ec4eaf029273e774856b946464418e6b707c999ac16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a367bee4dbb430ac0e4f7df6f0e72e97191667136cbe395eab4af88d6255fcaaf5c1975a997d71c37004603e72a7ec3e86a14653542591ff3d82fe50f8022607f67db46faaf2843d30ee6e3e498a956d9604cd758e67187ba646cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18400a4cf0a58b04c1633ac36299bf834cf47cf6a84b08095cc97e315f4c7ff993ceacd5006ab98997054d4e7bf46daed9759824a9e7f53b6d96912230743cc25973036136c29777ab42b9cdc4a167c8258a2934c29ffcb1630d96;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc80cea5b8a53893d9bf0c96568483da9dafd06cb5ffe5ab9d7ccd40a25412633827e11b3dcfabb48f45eb78fc0690832bb6a8f7435add02686e354d4cb7c2a5092a74ad571e5a4039c0953c14e86a6f690e861d7bb91564d14f0c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16af44211f780519ff687d2f31ea90cb85be77beaf0ce5fb38b0f388c35137871417b0ec2b2728e933d4a06f5989144af68eb8d521f109baf402292cf825906adedc660e36e037f9dcfd7f81af64fb0a7099110e47a5a85ba352cfd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10211322eca08834000f7b33b8bbd1df32fd5ff8cd85804ae37724f64fd299b854a494f343c0f94f93fe8222aab617827032a8c961a7939ab55fce8f87320e4708a463c450f745aa4bc338bc6fe3822f49381894b6415c37c1627b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1282d8d60389ff2489ba5fa182280a8ba7ef25dc87bbf8f161954f976dc0e53edb4a59a05401e28fcd30459fbdad18d20f00d234d2347931bd41cab37e5dfa90edd583c83100057acff9ffb9d9242102e2d9dc2feff0a1893b46dc4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b94e46f8eaec053a53639519bdf5ad3c6a65549641f273694ed9b5bb872f77b81545d57bfe447b12de8390aaa289800287fbb1dcb04ebee28f789837fad0b34827defe033951863a031b2c4dca6850ae03427ceff6392f8ef53714;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53808afcc033f5f2c659bf583066845b450f5aae9cd82aeac797f1d50663209723b0b1c18471d0c56fa56312f051c061fdfaffe83aa6172c37a1392d0d8b239076ff08a9f06383f8e45018a489ffb05ce202ffc3fe3b3e62b394cd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha97cfe56f396b537e3f34a1f283d6d96f6d8e2e04b4741a3bd6638cece6c9f78c4fe8c23d98328489088481829f131685ef24b533949ac904c5c163f3e0ca1f8587f954bd2f18c7483a7b9a72ee4c1ea696e80a16ae0aa6af690ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf1256fe1ce7c43d6261362eb7d6717405075a4fba1bf5be9c8054c1c6ccfd987a092f586d2d1bdc1edbfc742c698aa70c5283a51451c46e1d7f1645769cd8f1a98646eadfd3074ffcb5665cfb6f3f725abc1c9435c598671c17429;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc66253d34d05544b0c5d2db466ae028a19b067f250e4473b7d3513840824e5903947170d94a235f7d838d46524b0293fdc20ca4a100a9f2651ca9e384299106eded0c81d0b324c371aa3a30a5fe4d3a583cfedf0dfff7897fc7b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f07762eee6f3b8bcef3da3f8182cafcedce982bd1840bd801071dc38cf9ccf3958edfdefcf4e3b34a82758fdc8f273ab2954af567b24777e1f8ce2f52fae898158563af205242882b792d63406bb89a6ddfdcf375fe6f57fe5045;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ae3752cc3c7e9545ef909427fe5af1e0d5dce7615edba2532eca1c78de7da53703b28c5cac032623c51613c1ca99adbb697bcd901ad04774bf059ba06c56ba483c990e727fb42f0990f7900f005855bf64f1f3511a444e7ef5258;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1027bda790a2b3e4089bf3a1deacbd11873c6b97fcefe72db9a021759888666039153244dc790adcdbf46a32cb7fca260754398306175e6de91a73e95a19d68e5ebeccd36d87ff884c9ad39c2c4677d261600779e960f7d2ca5b7f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e1b9a5367ca77387113285412ed6598ff9f831e5dc4b7f09cfbb4001c8e9b20ca7d50df42acc159543ddc85c0a4808c443f809ba82dfaf4f240cedff1d68ee162ad68a22d8cf3f15d3be9deaf2b02bd5040731188d62b03c32899;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8796a53466435ec7b12ccff1d3ef302ca6065d8f4f8fffd7cec1667609cd3eef3785808887e4cf4172388ef388af8f079999ee168058bd08f2e33db7672c5e20a2614bfa8d848d329c0c09de282440a4fe0692fea90073299e37a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a8749cc078d6dd2654241bcd382121d560a5a31838ccc986cbd083c708d191d0023a9e181336d6b06273f7dcc38f7bc18c69ab0ffc1af090c2ba74a7c9167f0dec56fc46781081661e389491a22095bb43b440e624e8671f3ad0a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38f28a28a21b834031de229c2ab487b73f2e4186b6b0efb7a095e2b2a47a8f58e2c9b7b650abfbf95a16014f4fee7dd099fda8b9e985ef251a6eaecebae8f83377835b0469173302daca5b19bd3c8749c4deff7c699d1d317866b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f78c18c40a819921fc3e7f9f86088c857d488a6fd37288ccd66d90310b3cc1d3c10f854a02f5a34c554a3b8812a529fde7fa39d5ddecc1956a73f74cac64dfe2e237ec8941c4dc1ee28a46253873c11c0ba30fafb4bc0355f4d546;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158c74f5b7d50526a4933fbc9d861a281d0bf4b34ea4095e0a02d94e93dd21ac4c8e1f6688336fb264a8b6e2fc010366e5e61c9e0f8b35b0cf24bfac86a6d7eaa09fc8df9f3a68a6a0bd689864225bb696c01c54168f2b2e8f9600f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cac4fbd1072358d88dd62826724f63a6304d3a9f91863fe98b30ba0443a30f9bbc99aff99dd14ea0a18648dcf03bab8a51f9679b13a00279c05fa5a156a73a22816cdccdb5b9e18ee3fca93614a8b955f0202251c5b51906b91f1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0a8414d976795704b846fc757986561adccc104ffdd2338533acc09ce81350a8bd8ce5fcbeb8b00e7bac1144672ac1cdeafe3eff5b8bc2e4783fe673240390f26ae12fa7ca60549a8307e988cf37a1ee2926ecfaa1c1ef16ed255;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9fea521b834d5c2fbab6885a1f69d9cc72883b904e3b508c0213558d3ecf49427f9fca669e4f64c96833d5f80b23312640f5f17e089765876fc5cd056fc8114bf79b993f63ea38637dd9116a4966a618a84c47019d496fa843a55;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h181adc9a82665230f7ce567189a71b9832a2bf5bbd5d9eec20ec7a7c38602a9cf4b7e2e252ea5effbb46f39f9ca087e299bb8a0aa8f434e43897a9d73eb6db08c94020e254a2245ae1c62bc3b089aed76a8459501dfd93ffa87ccb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6c4bf8f86e9c271f637236bca040b3f9f46d4069cae907c2609fd424932c15a499d32bbd563d784522a39c66939a8b2c3c331b2d78b2847537f8f54cf67978dc5f5961d944cef699f245d328ee4b59ca59d7b0f26385f105b0c2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18bccb7ffd53203884c2145e3ab11d98457f061c5097774fae9ad2c25c4599e487d1c7edc99ad5f13b647aa2b22c8801078e25537dcc056cccb5fd2bb9eb63039c00b07a0840c3321b6be690a15d87ad9ab6a36ecdf2392acaef2f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8129cf301ae03ea84af4b62a3b2c51252555dfa473cadc2bd537943530f889b65095c5faade7e38c80ac6c1d8f28bcbb54690ad697f91b7a6775a8eb0f386347e5a24357546c195c0db503729e043dbe7be4ec311f463e90819d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b229ab7d84c9ea95d8d1238b5f2a88d486d991c128d046b9d09a7dd9c4542006a3224af815c4748fc986d6b25382a49df153d03fb40ba8d349b914ea1a35b1094db815c0192abaee3ab2d0f42cee956117971cb7ad7a9d84b2430;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c312390711893ac847a7695361c2f4857e1e595f8117e0bb8668008213c18eaae7fa2a18adc48408d17aaeb465888a889e3e65b67dd6804a71e8596a8868541b401d198b64fe6d178d14e458fef3e5c8ea4c244f05dda591a77485;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf5aaa689951ad418bb70204e4fcb4adcc2cd0a9cc91da63d50b7fe51a8a7f7deb068b56274654c880741295ecd99446539cef5ca4475229a272aafcbf559e22514ef39105ba8601d0ee8d8a3cd59f115c550021f22fe24d1119a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168ccd0e9e07ef7c12068352ae0730431a71c2bf91cf29553dbbf2546aa4f18102002e81f0df9a1cf351eb16223fc0fd1d5ab3afb1426654caa46f54cd5ae63e78711fa7b873c639327de160e6edc517f3ac092dbafc0326470075;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hac1fa56ef061d89dac87477e445b52d65b44e4bc160865913f8cd0ed53c0e4ecc6d0365a634cc73c839a192035a1502e513f159396070f7b94b5164a60fdeb75f5449f7d445b9db518aaea0611d0ad2165f79f2b0579b4b880e04c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11079537091dac6865e44752673b4a09cfdcf9b655e9c81e617eb070d19377acff74d5f896e73055793e286b5918fd0623bf1946ec97c82e8d26bddd8f39222de050bf3d2d8291ec19f121af8d9015150c7bc2fa1ee15d5527dcad9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f949d3300b4d0558d890ac7b2e225f7b19f130a943369a2b383096eca225d62c824f2439d91c0aa1bd34800e4427546f8c8cc72e531a57a4cda9cdd43f10122dbb49f26339c1c2955308939141f6f6fd3c42a322e60e616abfa6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd22226242d96f96867177db2d5c1fd2a7f6a7271cca2b69f554ee730107642c8583e5fd8409d822f90c7f661add953c032bb97e1f9ae5b85e09cfcd24d1323fe951bcda18f379fa99a61f398de7e7012796ce48b68ad528d3cc9f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13168e37a5bf55d963cbc7424f0ee93e1ae4fd7f541079fe713c8ad17259ea2131a835326be794cdde9690319786f82c6bd00f64375abcd3b66dcbcd03ff6474b7b3be9e44846d7628302646c6e83d8ebc1bc66b3425a399a530e98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7fefbf58ad38b93f7c19c0c23ee94d35c994256cd41ef00ced3f61a9ebb519763b8371654d395549a05e5865bfb1af45931d9f0d45063a8119aee101f971ba1400603e40b31f1dfec3cc23ca99130fa3efe42bd51414f0bd2b37d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c39e10c02680ed643148d1455a5ad4e36895cf7e1075062bacca3f93a0c25e73251fb66f6773a948897ba9a3a09341135deabde7c90ff02affd62c342b7a76ef8182318a98963c03089f8c95dd9fdc2e8481efc075ee6356ca10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c69d109c1ad0c714bb32cd3e43d2ae44f62a6956e778441e0ea1753d4f12881464156310ed11ed83fa9148ce515ec117ebe35e32a9be91328c028bec54bb98768b7c5edcd71b188410d4674a619f98fdef98b53def02bf2e1bd68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e0fc652c59f76c046f702796ea5c5a29d1acc9d647bb9879f079e5a17932a8959493001e178a0b79db0e062e9fb44f13b25c328fd90ff713973401bf5bdb16816b15666f6144dc09f8c1c482b3446a432021181e5b3d3f3d16b47;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfde3f830a36280357464f583eb03ca58cc0dadca407d9f551781225158193a9465c7ea19ff67a08774ac92fd4e754d6c1e366794d98155e1dfcf1f91f00ed38ea8c78765a7241319a6ea5f68e816ece8dc4687e5f1da4de191947;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cc9f778624516fa7dedddb9fbcf120c32084b7228adccd816ecc8f768301a3a57ece8a283069d49b60ca5df8a21170ebb556ec89799806879e824cea5b9ed67228e145ae619e68554c95ba90c3748683f65a0e21b4a62d546ed07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1327d2a63048a356e5298485fb427cfd77ed4bea67632c18d3687d159670576c548d47f6a4e05287393d8a80ce404e78c7f12344f4ef2a39f4263688f0b45c5ca8c4ddba78be86f039477ab207d8c6431192fae68dbb46a59b625a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18aaf9ed85fe192d7783b84e2a2a7ecb32c948d56c4c9a75a21c3edc68e72e12b1a05c10ecdd45d4681e24d4a9a7c1717a8b6f9407690f460ce82782aec9b1326c2e31986ee19e0ac650bf1ef342beec3f1cde35ddab65d8c17f96f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb98dedb7ee9b0107a1dba0f83f78e7551a500e0e84bd28bf27a510c13828c683d4b69c9d2400d3ff1df038e589cfb8e6269be20a3d70401913d8d3a297231721856f8139255e5ca217eb2ad4255cd40e8d457c926c22d042ae42;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bd5c4602c677390d222efd230040d8285d002fa0a25324774a898dc90c64a2550a66aa100a1c0d68037c20a66eb6852de1472579bdb1b837097f259373513a0811e1ec40392e3d480c301dffd539f350d64353846180dbe228d2c5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b15ea1d28730802b7666e1e992191e606923b42f3fb5333fbc427ff2e29d8120c25c9f6cd6632f44b978640e2cd03021501a822fe499434ea3ad737fda4f3762841361f9f969822ab37885f7890725129f5f781748034f61e9ba2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf10aca53c9855fb2fb0a64c8f1e1259891b16bcbc762fc78e0e73e72688697065dfe46bbd5219fed63dbb32eb64a1a76afc08ebe9eb066b13a984004faab2eb038cff980917c106c7171df6d85122c83b3d3bfbf8026573e400dee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0b16094201a8d152ae623a7d32924d7df97128a2a591f3a27bff10828bfc5f810000c6cae492453a52f8eeef2d0479fe9bb7248c469ae086e8c6eb80ec4d95e2c27f18d68ab97505a5ac816f21d3236a33411c2aad5c0fe118df1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a52ebdaab758606228ba99ee6e86e589c1b1115ef15a9d63399f0c5ae4d8cf6738510588e0bdbb90aa2f5c74d048adf4ac298bd0d607e2ce8127c8169229c3ec63c85bed12c825698be97b78dfe189c603d0a8f059d5e9d080f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1209849dae78f393196a6207a0213e49eef9c91f128012c117d7161185dc2d32bc1fb108dd833780bcaf5a3b54e145019854b7bb9890150d4c51acd845e68fe47a8e7c9c91a91cac434eb8ff2f860e07e7a5d7f645de2535a2a6804;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd6397d82cd252771e5220bab856ee1fa348766ba2c081e550e8cf058da7f88ca7dbe9b4b463d69ca81611e86ad709936c6e602de8ced703c06dbf600afe78bfc4ebade9ef6c345b53b4b072c4a8924ed21923c5ca278a879ee0ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b0320aa70a7f7c56c1dcd849ef235b1597666b75bc668023d81f9e93331ecb1a849d7f5bdc9b574262b7f49207f361f6251e93b6626e7abfd4fb9a3814855eba1e0dc3c3ddfe38edbd1ee88207989c9ec48063cdfccf779277e14;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70465413df4a6ac0c559e92d22d5d3c238717f3c10a779838bdca21349a7077d5e8982e4a43af8e6b3e12ed3b371ffab138d61f4582a055bcbb1f77129c08b882245bdfc8d508820763926455060be251af7858e3ec0e0a7d2297f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4247b7e338d22d8a8051ac435acf87d6d5ac9ab8a65a4b2d445a5a8508de49857e8ca9c2c29e4f06835a1433d5303965830c7b8717af8a747c7113d7c05d57eb1fd2ae170aa6f2f2c69b56561a92e15eafa90a0fce61c6f0229f2b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29437cf25529436144760d8319d4268810dceb932f2030c3dc1136b17ec32f4da207d693be08567b9e4700aef6f0821d95473e449e725137bfafcb43d2fa019bd40f9eec8ed45a4413bf29e58738472d3bc774a68829598e8c9842;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ff701b78f1c86371250de636b23a2ce005fecdb9f9ed4389d423f2bd5e02de3b67aac08afbfa7ce424108dd893298c7a1a2403a7dcd4abaacf245e12606f2e12885da816a7df2d45e33c1eb9b2813d9c513d79d1ed49501494a7c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfff3116f38ef2a95530fe6c5d8d050602847397d545b9116612d1f08baa8c3911a8de3f97702ffc5b13b18acf69523c63c538b43e8c151d69e743c580e92853a7e07c321dabfaef8241716f5d6f23f8887f48b0d56378f3f24f3ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16582bea239a7bdddabe0f5341e5c2c681b2eaedb0fd40cc8dd009f6c7107c883a527d785b25153a1e89360dfa5891558f436a29862723c014e64298a492a869de1c2b6bc570a3649afbe64ec80fdc0098e5f98c29fa3d67197e731;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b4494116e1f76b26fe27c1725d1762b5ab66f8f55ee201e973f3b95ce61c2ec46008eb0bc1bd4c014915cedfd661a14690977ea7862121e6d3703b5a6ca14cb472420826becfb22a9c10196ef59eb8ad2b466c9c4e7c78565c6c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2cdc0043a2ecf1fbd8f0a1b1343c078056e53a3e386e622087d9dfd2797fa1f152c216ea1c3dc399a4a31d6e2e853a61557ef9a92b1d6edac466e081302fe2e030680ee84d4a1a9719d4f4d769fb3cba997ec56f47531395d90bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1681bf08339087ff705a1aceb2fa8126e5949676d2e9eaca8b7b0340fe9e780be2fd3cd13bcdf69ebe0960c4db2aab66727113048396d9ca601455cab6c520d7381622bac17a7cbd1ce6b5c0ce539413f387569608a8d6e1af63758;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb3bfe977264628606c772927c43800af5d14b9d26066dfb586039a028b08977674baf3e445cc3368ced609a3e4ea03f29fff6c5261327e4f586a4d99354f7f66bbf06efa40b7f9c1d0f81ab4760ad8a662e28d4cc3874def63d120;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h124c9130cafc7b98a9d5ecdfe020f2e313abe7e0a3b6c1e452eebc80ab3e931c4f1ee0f3e7b502d61858367def7fa6a14c62e897e33f59e21e49abef5346b81bb28df4f9e9fb63b45eb414e4dd96aea40a5fcfcd68d0069324ce0d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hddc0c1aa8157be3c4ad6baa2df17f69034a183478bdd62abbbcedc88c3bba68bddbda71b882896468696f3456d993495d3fe0caab6d2e26d47036d2ac3a8044417515940bc2de8e47253b81490a728c20f55ed38211abc1943f1cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ec735e41313bd204b9e521153ff34e52920aefea3cf2ff37d8c1a848fb36f518ad18ad8bdd073cbce7019a6b1914a5392e2b0297f7ae4366c839b5b03e4f4002619a7cb177b3ff170aa5d5bb9408a1f6034551e43c5a92d8f7331;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb29cc9047ad1ff0fc8df77616ccba503c41355de8a47d57d33d08f8af3576d728e8e3ed1c060a4ab0119f178044f889560e77c585de7be87c92f7cd3beeabcf654c409f633ab2d92774ff6aad9df2c963640fccbb4370ae826bfc2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc63082f9e2914c8806d9f5e5e7770c1485d58014be9e37341368d242785368a359866c839cc2c52fb1d91ab5f4ec43c577df9c49153800ab200f81f3334c74986fb81f9e428d272474ddd5d4486a5f5f9aedaf678ac63be59ebe6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h388787a70c13e25c2532115c5bf67001b04a0df66b9cd3c212d81795caa9047fa3cace67a21623914d7c4c4ebe5640061d648713c689af99f905b7b20132e794022328ba4d49b3f1d482474f8df0462a56674b4e539d27dd86b196;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12df4e38bb5b581c59ef96110fb2ae4acd2c3a9d6037557694eedc95aeaf0ac52cb95416027a6b4f0c495a5e7e653f510334e7507c73029a5ddf0b6a2aadc3e3dfb867e7e5e308e94d7911d42407e21cb4548e5fc84d75512519223;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7cfb329de4b7827d04fd97e4e7072e8a4db97ee5dbc115f0cc094c42a2c9da9439cc844bb040579c0f758923b53b5e645904be9be5e5199d001cc13669019fc653b6e870bb1c178ca57669f642448f3df43b6457f9848119895825;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbeca62879c48cb44a5c5c28cad566ab92ab5762f4caf3d4192288c2972206bf9e2266cd52b1dac8c97c52515b567894d3351224212c21cffcf19914e576a408f003838835b88aad28e78415e29f931451290a2750234374f5f3a9f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1881dabc5943a937b0724df98d12e912dcc547d4a0512b591f87a3a31ae3e83d77819b8ef262fe10140e3bd5a2b90a5fe0799c59c622b369d7c33e1ff656e5c9dea368b1dcddf4b439690533f654879cdf0de528427b169e17e11bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aeac5beb718aa8d19e0c003ded4c6803547802e93590a01e0dc7e0bc0ac43dd7fccd1ee5fa3dc12126f091dd85de8b02d11f0c955fab131ee8049987aa915236ca792a48f0333985d1d7722b46f35651489df7714d7738c968ce02;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7174d420c2ff7f323a9b1ca47123fad67a90ce1959a5a8417af3818029ead64d26a1d266fcca457d68c9e131a459c27c32923325a569a4428ad933f6ddfbd6685f79b41dabcb4ed0ab8e0c4392de98927fbaea42e6f35557c526;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107d594f75ad00c8e2e51b05e9fac23ae61e0f3aab09177843baa6035b3bc9ef2e9b003a9a5e1a5e0829112087517b1c9020400470eaeeb70cab89eeca78630131a136c775a3601a5f7b7d77bff4dfddc2873237c13fcee6d2c6249;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36bb6a7876427e3ed112f6de738317fcff808f3e866ab2e9edcab50dfad6a90b001d6af7ae5a3e298ae14a679fc33d972ebc38746c019b65e468b1a1608f88de9a99697e8dc55f70a102cbe96a3f875d29bb1000b57d843a26d634;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b5ca2b0e0dbad09ff1baf826279a4d39e14586051204230e8ecb4b86c4dd718b7b0db95a59d09f987caf17c98e0d5114d677e19d17fae94f137273b726413bb4f47f113659972273f254195773b4f49d6da40f83263127238e247;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b620fca593be3adff5091fbac6e374267a916319ca9f963058a76eeb90d3578d81a0a558580bb17f312e48a417e8a72271d77a7a549babce342ad1cf07d35d6e23884fb575bc0b344210dbfbb4e9b09cdd27916afc90631dcdf108;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e200b318b82eb11ea001ebd121a953ec65e091998876029ca5dc0cbc9a95791d2bdcddd0c827025c989d52ffe18dfe34239fb1cfbbf0fa03c8c6ace435c885b4a7e31558efa498fb4fcddae5f541570c526aa907f6956f23d9bd1f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1080da0e6ce0811cf1f15fe4a0526fa954bf84e97f5220b72cb00ef5db6878ff76671b34d05c9ae5de1ca4bc0bc6f042a3ca67928621b90920df5f088212d75f937234a5135f89fc82c5a1581f5878d0d5466e35190631370875f4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e83c317c5f3aa03a076314f4efa48fb8ea584722eba7797f8fd5a8c89ca0eceecfbacc499fc646d1c03f5f86101d947cf5a7ea5e35cfb315b7863a89b017db6e2b557de0bce32d49e350a8e47126a4b55ed46858f363c6b9f8dff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182e8649bc703a0db459ac3e19fb29b9745c09ce9b71f7741fa20ae1cd6085684eb06c6b531a046cbc23773924c24f158939a1caed14cef3260287b49f86b77e5ec13a7441233f16d16ee6e62575b973fb1fc2576ab96d18fd6a82a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a392ce801089c181d6c78fbea74b3c652b0610cc56b8d5056b82daeaee35feece25b2cec8601258ba382e393806fb7463e2986f7b3c7d4fd8783fef499961acfd24261c0606c42a6bdcee319299817298a58d09a17e4b377bd981;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf66a79a36018240353a879653021027891b612dbb263705a6f4f7a96c62c0ebf048d36844cebc0b98ee83e1bc74b99b209b3b77c17ea268b1e798cddea37ad6415fbd19265f77631d4649bba9775ac6f288cf4fbb8285865b7c998;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e3ce6dadbccd3433a3da6d5fd50e6fc7470b876bfcdcb334921d58d5b4261c2531f0935bfd8e9ae826413e69bfe027cb664479cce3a6108330dabcc1e50a86104ccb4ee336b6ef3dcdab0a7e02df681c101f576ac46eebe700e17;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180d3996b654750f1a607e30647cd9c2b37194bcf0db85b17bee148fddc43c3758f738ed9303fa268ecda7506cb18c8c124cb764d371c75ac492a3c1c9a45ed3ffaefb6685a5a5e4ebca1f7d04cc8163e8fbe20a94658c4c20a2742;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef3c0d158162594f79f22fcd9de2e9e1cafc420b88dbde8f2ad3fafd3e54644836ead73bcb5ba4b6c7b3cfaa5d670277f42d46081825a97bc9749da086a75ea46aee5e0f5bf8adabe0964a7bf73f2705d4afe7d40d4e7b69bda482;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha58c5c7c4fca7332e45ad6a0072a74049b65294f0a601b97d0372f735a671ea147a36de87e5da0b48db0d1964ed6dac6f689d26eb072e3536d1753e52e5826c1aeccfd98152f27e41fc2c3f8366725202e10c4619c1c875932e4e2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6196bc41a05c5fdf1ad2217c89994a27db51634133bbb3160af4b57ca8f87f7b2ad845ce5a65805c940065162001eabdc852ee7087d9581a65cf0c719beecb1faf905d3e440d6591fbfed703e499117d01040ae3cf789f7bce6c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27ea07da4252b0d1b5248d32284e9575a928dfe819d6ce2bf68c98a4c5aed882fe5addee15082f2203a009144eef7251a3ddd25c789b7a381ccba588ad7301a0b61cd3f65857c7be4fcfbda0d66eef8097d94e82a137aa06fcba37;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7d431a04ad3edae9423e5b1520402181a6870be14e8a8bd63b0c551fe027bf10d70012a94ef7043ce0cad4fa7de56464da7b274428a1445f6117f64d04d7f72bd447c8c882f65b6ec8115406c741527da48e064ab21b53da7f7ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc3d05e0b642ce1dfd4240a0e3d9a8bb077e54016bf749cc1f27da300e12b0436e9fc1391b939963c703d8df95f0c4b95737abd69461e153f8972e01d85b95fe0e4d953e9ce47aa49ce77b38591d1845e5ac8c08a5dac9f1c409a33;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10151be73f5b34f5fae674d8fecc0ede522820f3b70fd0b106e38db11dd4186780b3acb44c444bfb01b3c3512cee74be28b1e2d9882412c4c0e0f092c22718e2d6e86d2b68b81d29ae1188e25b466c964081d1e2538860b8a0e82a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6629c53bf631cd949b9e8a98e71eb9782aea31d1554c6aebaeec761608535f8ae1eea9b4ec64fe70997f49146050323a35aa7d92986d42c3fc8f2953284da8cc314377e744ed07d151de77b6333254653bfc9337bced5c10880b75;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12834faf742acb75ee3fe764ea8c1174b66375c7c9eb058d0723bb022cf58e2e15c7ca0de304a258d2ee356cc7d9271406fb22965421e38b52b4625a4faf5bb525d52b8777da3968d1f5b782dd7c13d24975526978b2132c7b48020;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e0224496dbedbc207fe38317743ccba01e179e6364f290414faf9acdc630844dc9957420383053fd9d8a09f7b250ef65604544970d9309224249a840465bf7b597ae3fb30974103436f7a6bcdac912021dbf6ce595caa277ebaa7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf667a28bb4c946d56d1861b438e70b7ae681b56e5339022f94be770497aa5290167048121e72bae60d8a8d1941983fab7fc04e4dccde7c8f4965ede568b70762fc957c0a1cd9143da407c253c3402cd0053effd71ee5f9f6484eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef27d74c3d8d5110b23b861aa51c1c8d0154724010db53919723d8b2d7a55962820c2b01a2638ffa536cadcc4254d281af3b48a5426617f7b1759434be0d4a2e7495be4a604ae43c42cd6bfe2c99ae177d8afa1d278f91126c65ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf48f555ade2e385742282c8fe9995cd58e914d522e587638d18cbd502c917e2ef88c32dc95f663562f4676f40abb572dc2999c705f8656b964994aa5d49890b01f973ad146c5380927b9166fafe70e010e4ed79baa7c6a82d78d04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18813fbf3f18e3d771cb4c2ad8672e4072fd73980f2a07876d277948becc91e512a63a330066fc420cbc85073cbcba005da4deb09d73536e342c8b6b2e3c1582031efbed8ab21d431a5cca25849b926efc37af045fea85b1d20bb8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8482fd86648f3f17c1302c7c1496e619984000562b1b0a1a27a5e85d46b98a850bec074259d658522803e134ae43b79972a103b1ff68b4c4d0eed77e1f7a4662ac319f57dede7ddc2f1dfc5b4a8d8cc9815f881c4d2fa01f4abed5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9eed62f657a232ff1137100d150e6d5b7fca666df3e1788e68d74237f088936b62a2514d2e953d4c2a6380122d5c9d074636229d7b7d099951d20c129979b656e907b8258028211dda13267af19b6c7cba63c3ea1aa6b3006745a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26b6da4b5dd44c7650f14684868894a52413d9eb45a5d83054f81b06f77ce4cabe7abda6ca57606e09471af4a9e2a9c7452ab03b3a6be7e9d760932dea7dccdf9c7c43a9bc1f16d7c4dfd3424529b7b2d2a497865bafeee690849d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7613cb2f5b4ded47107859cf7dde1188aee1c033bb144c39317d002a0362ea44ed6c82510c8739e73010b2edd5ff60bf91f34c543569d6e87a53d0e601c638bde0bb5bf5aee7c0d64bf16511642fcc244180d77a0deda08ae4a2c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ebe730fbeb82dd3bdb53d66deae218698b76ca9eaf6c88814514716e5c11af8d50bf94525ba14b710498aced3bbb39edfe0e96ff7e075f77fb3c458735896876250afbfb6eb839dd2e97564522ee97c92ad5ee8c95421b74d960d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab9549f292e2c87c9a082a764cebb98107ea05393f9e95058021bc980b933121a12fed2c74ebe2a6be317977fe092153214594752b8631a177c8678ebf0acc259f0f4351d2b8d9ce393e9bd24c8b4bebe688b6e1a037932b4bf830;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b0644bac0b177d0d52f49ddcc351fdfc7ceeafc580224855813c1652bd5aef2562ada4d12588505ceab4253e608dc5634d25517dd25e073360467d00d0dedfce624b060cad3e30829a8f72432e6345ee6e699fbbd5bb5b5fab0f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d7aae49f2739280177633284e9c3c58419138cedb60df144fbb8e276e7564b6178c9eb7c97e8a9747922cef939a030aee01a835617e2eacc76265c14fde29aadb3b9784ecc1259277e85cec9681a198c6195ae5c92ff2c7c2f95b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h593661c44902c386908a89415bb963b4073d468bb6a9415ca46355c998e6b47e81ef45c94bf5547bb64673d00c9af8c9c9182ade718e359c64325135625996472edea368ea2616d63e32fb6720519bc6713c6fc52abd3a6b42642;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a4256c6ccbc283cc4da1adda105c78a5e645228aebf20f1318db25b2e5da27cbd6cef7a30d8a8778a39288e66629621d56a8f5bc8e51a5e744cd2409d0c4011e172bf3463722ee3cb867c30db628b6c2a1154b85b50bdd23c2e69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18731947b44a706a84df2288526f8fadf7213a7abdc7cd1be1187ffcda59be63860ee4a6203177146116f6716725b3888097f4ac11e9b7dfd2dce9fe6d97aa2c2aefa3587ce8ac54f42670afb1e663d3e5e69993385de51f096c906;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6f08150433a365a7603ab618d0d26a4752d11bd63c5e0b2c9d00989fa7452ef44b8446ea22765e4bf434f2373faf797644f1f2992dc9e17f59cbd3726cc07664676e6c54ef62717d2b11d23b75fead2111f67e555d4a7555821a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb936375a57269c4d2679da1216c4a7f60575177c1937b32d1f115087d910cbd64f4715b112810d463b4b67bd2ab3559a2c8e1521ebfb306088b224c9ee0ff1f8a27f8171b15796e74b21b0e86176d5919e11783173cea5a075e01f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h852daaddfb028a51cbf0266782019c6386f7562add37a582c29ed609f12f9d3f2e0a8e91a1db7a7699952448b43bc0af6a4db5fa52d967713c58e7da7f96b642ff456c6cbd8348b0adfc543045551ce7f5ba8930c347b7fe989959;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a592c57f9a0f65a7be9722cbd24969da110eb73e5fd2f6419180e568fcefd2cc05b293a231821889a3f830ca2d89eb6fa9ed66d581a812208449cab08e7176995ad93da20fe7655368ae1785c005d97e4908ebbecdba3bd3984cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fd316c482ba8725c8ac8e0e9488ff9e12b3bfedff41f7031ee5dd2bd04547ba320a8a747e47a35656812cda27458f294dab840da22c9598c3fb35b4bcb4f54628792272461cc19b5bee22377ab965d1ac8f527376975f294aa8d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43548e5ea90e03161f9a4dd9c2de7c627e4e480c64957dd628d40cbd1363c476d90926cbab3b33f7f4ce5fcf1c140ddefaaac0af42309831d269fa4fa5a74d5b78ce2980b835ad2c006c7bd129c5535d0a39850950176b0ce050b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h349c54a87407f4d3197bb1765868104e8c965e2d55479ec22dd8745e54cab5c14f96391340a702cb5258b21a66ba9da6c5e914a63872d6579fd059d45f8cf8c30ca8ae7e384ffb14f0ea83915c9d4c09563140c3d5023d5b08c215;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h52e4cd68aeef903dd55daf08f33f0399ffc147fd2ff9eee70d23ba8009f67ecc9e17d409ef37e416aca136d739d93024797d3af7a381b4c9be34aaac6c69c93fc0c424720ab2c81a0330c63c354ebbf211259974713c509a74efdf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3983c8bcb70273cbe5b11566426d8e7c9b5a09c01dacfb004cfd28a151a721ba4df6ae15133ba302022670faa3dfcc5cfb2843ab1fdb139bec775f5098f858af5bc9cb92af96104c02b6321fbc3e6d994d2f5c0a886b4726d4b029;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc7c3eba6de67851c32b0a6da64de23a7913deb9e2752abab62c7c6ff77e59718489c1689bb3e4e2d328eb2e335821054490cf0595330f0b4598fe61c8f6f4a65750eca412c863629c669180c474916012e2bbd0d20e2b317ee2c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43478c9844a46a442d20b0d6e5fd062bf363630202c2be7823eaadc9570e901ec6667931daacb7fd9dfe1aec352e6931458ca699e9622b6b0242e02b1465a028eb3afcb308f3528be853b85da7780bf7d51c8515a856a5e93eed88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0758224f4bfa21c7d3b0927711bad23e6e312aadd21331eba6c409a4540c15ee69c5fef221b3735368f8546925216c7be49a3d36f878f848df22a065bb894628972dd518f2ad2ed7a54ffaffbe4782c2e6b2ed2e9bef9076a1084;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67382b6ea3cfb42419eeb9610ff9df7302d9d4d2177b3cd28bf0c478b49521f1b8025d2628326e5cd5e1f8b0b94610304cf76266bc420afefec3741fc5df4f547d40aa27f6dcbe7f3e41eee755b1a9850cb62e1d3d6111c97fd5ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8492780a3f76e494e4f5477a323028338fe9a1e71edabf5fc34d73cb1d270cca8e67e8ea7128c767e59eee22e2372fd43e316fde7c1002bdfd08596f8faa9e640af63ec0643069f3976356769eef0af2ac93f1f539912621d840eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17d635a5c2c800d1f6d0a67b5fa0c296006ececb89c2ebab119eb2bbfb52d9041abf80275004b3b19f6d50478e34e10dc15addbe5ea11f25e11610e33b9cca813e1d3b45c92e7061baf5c7ff27d660ffa14c089e22675a904719c0e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha056b1c51446373a05564312af19a870da05fb5e06bbfc28fd8fd65d2b5dc2b79a9b91a9eb1ab3b7b2f31e267bab4b2a1b23876d66342214911611852f7d597f89b7326ac0659c998c6bd73f847109123040d85991fe6c3ad9c18c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cba00b8e2971044c137c54da5d7392b1205cd76d9fe954b6836f5e03e652aeff79c983c499e6204b22984089ae5777d3652c8fd08aae8e28ebdd82ba58476726be315240948215abce1ed4638bc7bc457dc79b5043bbae8236ae7f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h39a12a867e6f0c28d4d13d2d84e6fcd3059fab28be8767a702dadc1e351d2c3a48e1c398c2528e6160e3c09eb1bf07b71a9389724134aa82e749d4a9894b28191165ae3e96742ce3af5d11096a9e91efb59f65ae87abedb37fc03b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f62365877a629295b219dcd03131b861e442dfc599f446412a416a32fa9fd41a92cae528e0c476923ec1baab12a24a4023caa163ab8ef8176a4a553bbcf220486b23b8a68fe2041abab9b0c124de46d77bb9d637280afbbe944a9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18dd78bcc092c6362b5d176e6c0b361d9d92d09ca8229e8f56a7015046be0ca5a680c1ed1f95182e34188fa7160eba0f4db7db84349804972057903f4f4dd291b346a82044a4891beddd274b00918288b68dd1eca2c50b403837913;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h642e40c86791205f5aa7e3e8a3612a110d889aceb57ace8288b1e315f3c4cdeba0d2c600dba39d2f0095cef1881d656a03918ab93c511c1e9845dcb8df45a28247a17a0b7d22a2efbd99d6f8915cb948761db6ef7d192f693fa310;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e37a4e2de9a0a9168b7c613718d3e3ba71a710a3e88563263e148fbb378ecdf6eeab9b31de8faaefe744ed5ee8b2a19eccb591ad916980db91a62111ba6c8bdbc521c1b92e58aa742d61595208b18f8ffabb5350533820ba2fa5f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc35d9f844e0d7ed2433039f4ed6bae29c1efc8ca958e20281c788a8db836210bc41ed14aabf2bfd0d47d688a39b6a60f2ea471540b60213f5114ed156b773ca1f25f8b25ae05444f9a1b9c0a2598de05a20fb2a9964118a6c448d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86b8ec577a67e96ec19569ebecf48579b494f433f751b550d457e034e9a3b5ee0ca79a0c63462809a70bf75363a62d79c239896134c5ceea52d3844726e5876f9aa9e82bc02a18ea70883c6ee41f0c0fce31be4ea45efffba4b539;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h768c8b09693b269ec841ff00171e610822937eb753413b19c59a9a1fef974e116c1e7850ce53ec153983a97b939b6546488b280295a1f85f80b454319441127819da1c992ad1096789a08a4c7cba5a35a9597a400e23014d6d643e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13be207ab4c2e35f1e3eff2987336093299a2bb3f843004d763b1b08d5c326e5dd15b3218b9809ee2d1bf3f9f8123036a8f6d7da81b8fc5af18199db1a3fe0a0c81191833e57169a9e323a26a9a6206e10245e2338f6b8343196a58;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hadf0defd51c87cafc6888f2e9c043cf50958eb4260ecb7f5e7a08c1e5a40f4611468adf98b7a009bce574497fba03fc9cab79d6a52fb930bee68e4087f1aa050341a3abe154ac85471879c2354cd5ddb783937b94b7b76ea240bd9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8a1a3d460917a8569c1409776e2769c6a607a46da661a25655ae845a62f88e351262a865fdf6f1b664fca676daed0748b68a9d2e14308a980a6c0cc3006f7f639673c8571ec12c291355d40b8a1aac23abbd7e8955ad2c0f7396f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e1728ddb57795c6f28e7c6ddab952ab8bc65976079a8f68167c62553b5f8540b0f5826f6fb0a9e88c9cad504f9bf53041d9f632f8fe173bbe95fcc094d13d4d5b33ca5b14c9f29ced542ac788b9115f168e60508cdf838bbbe962;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185df9472bdbd720dbf65fff3ab6368c1793b2b7d3fc9ce69b04806c0e66f12eb4375bfddc1bb0352ec1d2333b5180e8c0362812ea7f58b4172553b58d5085d1c848dcd8f3f84ba05ae4e298923ab14ca568671bed4b678cb415436;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97431bcda2b5126f4c4183634512c3144e2361d415cecc101cf2ba00a6d39760b9535f93b96e19fb50b722bb1d9487ef8eb5e3a4d2725dc48499183302425d5cb0222c4e035b303c4b5286465eb0e7e9f880fe72bb014267fee5d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166e02607471a824e2de52a4bcbad0893578db2a80523aebf6bb0e3dafd254fbb0bb76cebf5e49eeecb30bb6455d6948191a98e8b34d5f1adacc05fe92e84e4c9b1a1ff1ec645fc130400c708a8036fb33e7051e2ae37754c7e84b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h45484f01108ef2d03960fa45c84740ffb0873907f927c4cb338ee5dec30f74d67f9a49d8c0baa624c5ba93dceef9e7ef494e233518033179217be114b9f65744bbbbf3550e78289f7a084bda5119eec50fff13a93b54b4682bd581;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a50e9b2556d8f314b51da8b3837b27e4b8f86391bd86836348113099725b8eb1123056a8e21d95defa58c8187286fae487d35530febf49bd70cbeec500099bf38a0d86788b0d82a1caf01e9b9b169b12ae28ca9f0ef80a5aeabc6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3dd2170cb4f568d525030b08162e9730ef0945ac56ad5b8d9607f21ed16ebd640e139be0b365e5a83365e204740c3f8039d49599af4507ed0c3292544b8c6831719d0722936408d78650cffc1905495358c8166b6af898d81f5f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h627dd9bedb49507b86f24a7a55594d813a5008e16cc64faac407ea09e9daa216efc181334b9f4ec489eab7d10d331d3d11e6b670b37da65006fd80445b105bd739891ded261a7aa6f40323d9ffca9a0594df3ddf1bb62dfe55e0fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h22abaf38ec42a0388a4643148c18d0d92f80fb4123ea9214285528f8d786e37a03bc1dcd074d7c9d17f595382da6c58fe99bf9d63ef3d7c47d4cb17c454537a68cea20744480534c9ed3b325ffeb5c1bebd6688cb45537f4b12a5f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf2392258fac15cfa90d7a0f67641d545ecbfeaf09c3dfaed74ff3efb37c4b94792bc8beec4a4d9bd54764e8798add530c53f03b2f41405bfa334aa5d8b2cf32383b7589f86bf729515f1938c641cef00dc85d295685ccd761e6d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70078d04296beefe34031635adf5a1b16ba98bb9b74d5a14fabb6f190349714810b4d33590c1ad7c00b5040fa8a7e45749e59d3a067504c9379c123ae973db36ebbe71104a2824ed8424fe0ad862a23396e4dd1d024dd735a163c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h199c2bf7455bdba887f3339cf1c21617f6059587c7bf6bca802f0b38f7df209d8afd450bae3cc46f7e50ee4e9ae20f469dbbaf211ee3d20461cc2ab358aed258f3b0b1b23f458aa5b4cf3f9684d9bafddcbf44cb559a13474e5beb2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h704c6a9cf98707de61451e0b53f01a6ea7eef562e45a6ab468bfffe12ff2bcafe175beb52e47f97e5a09308b2ff7b205ec576181597a5cb94803d7288df57e5c939fee31ace72e05c55f88939aaeee393863d553adb31be02a6146;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ae9b905399c76a671ea3f90e7ed3f13026ecdbaa880d1eba5b3a9ffc4908d70058783d808f6a204e9765196cac418549af9589c3962ab536d8f913a2bf3a61b9704d9eb0f30d76af8990896276257c4e048bfb19ba67b26dc8b8e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1865cc95867ed58d13d0ce8c27b32ee121e10b872cfec0134e4ee395ce5a7f4e08d586bdf524f9cdae3661a6767cdd807a07d8796fa319b487f280c5d99939ae2aedc35e529672401cbf5285c97a9fc31599313190738c0d0a808c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hadcb5590cfcfd0b9a3231cd85bc02f184640aa15239d69d44385ebae480488fd67ec739b2caebc3674a84edbf3429c2fdca60a5df099fcf58e251581c183be5d5be3c2cc4fdbf319ee552e2d1b6107fdb0a2c444c27350ac7eb755;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5f68a9b94d06aa11d8495bc7d93b809d5f43645fa865fa764df9d02eea1bb5298d9f1f5c2f80a630fc8b33e7babf08bf736c3cd2769f7d2bce09f246a57c23dac62850da74719176704ab4fe671a0ff1dbd4884d3a2fdc21ed37d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16918b4adb453a0b69c33fdba3c79d075da4b1b882428a4ba2cab67bf076c1f1ddef4f5b9073b831c20fe0ebe324b3166868987ffbd79fc076ac1c45ea90fc5e74b3152a02eceb3ec2be2364ce0180f9df4be74ad24e5c60bf62112;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107a0f08b250fa2ed96e6814d2b8afdcee2a6b2031e499b9b0194fc792bfd68137fba32b45649053468b57180756bc078098e6e1e32817b15dae0f9ce0dc0b7fc3bed6172fc67b899770127bddcdd33d3357d5d01f426ccc69bc687;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1845cc02a270a84811effe618e5852c2902802dcceb511e0f6b262f43a18904ba4a1d01dff6767421ac340095ec44a8cbe30b34ec14302b48f467e2ea5e4f3a2b9efa9a4c5281ebc6c020a18708fde9a58b5002c621e97456e55b6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2aa41b872061ee1655934695b4fd365ee86a6b1bd6c67b0c51d936367d024246406ca32863ecd552c8d3d42a380d862216eec29407cba21ff91799aabcc5a74e4535fd5a2d15b23cecb1ccc83b5f436eb080b563106c097fc4f59;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h139d6da095a614c486c1d0fba19dcdfb1f0742034bf2fd75cb0947dc8def604b5b42fe131696c51df1e5d91ee75bf335ac5016de25965030e244635e6c6b7b626e0dfa89c753ed20590d5c23d45385c8ebde727b409dc8cd8d29981;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h307fcda8297402caaf37b840d77eba7251d3809c48cecf41ddf3ebf58e99fc6c54e8e15fdbfdf8f580e605317365f22c310eba3853c5bf4f58e0c16fe0559f3bd706463af5aaa15f2c0fb4f3b2795d5b175d50cba3952a48a8883e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb92b6e41ffe7cc58206be8e4836c0b4081f4a40f363aee40b475a515827ad291e53857580109692b714c7c1d232bf1432e3f5a024fe809f72ab572814ce3457241262bedc50380d0ee4461f70db90c74815d40e02dd63fc00fcca3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7fd33002cdba73f41c4d3c33fd4513566c8cec0b66ea2750ff2a4a5322ab164d31ec79a0249a81246a878f2ce63db9f690f7748c0e16265aa033362146355e65155b031a8a9d965f9ddf870ec044b5cfdba1ebb122b12b9de9850;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb44db2d49efe594d45fe523688f8ef825c0ce27842c8cdf03b49713b69330fd7532e87ea809dda2133da117a22c7f6b1d30a23c0b057a2593facf9db2e98bab8a1ba171de651def42c74947b77a43a70cec0bebc8d425809436df4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1a3782de599bfb5c4420c0bbfeb3e657cb84a420d00730e3733a6b3e42f45be542bb7fc896abdca2aee31de169d3662e4024c77f6d46ae5afeed0c776275e1ee8f16915393199eaa172988857bb2f1011d40838acb63fa44e9d93;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11bf800d040d5231b44fde34fe7358213292f7175b84d3e6a9793cb24e92b407a5ffa00e701b0ac9210f54b5e2acd1e9d7d4c797ccfc666e7ad6a00ff243d3a65f0fc616d0a92c28005f23d7bf5bf95bf9beef34f72e1dd64513cd7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fde424e22359e638d06c907df2cb1747910cad8c95278f9413bb6b91f640b90c43467abafc43120b42b236bda10d4a7be81bd9f24dc3070a79e810b61aa7492b508faab2cfb4e544baa9aa8b191bd6730cd2c47f469bd86774b35e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c64ecb43d7bc43a6b572fb81b974ff662b5ada807f08a82e14129c4a025f0d18902678f22a283ca39099d918ab91e5619fa7f7f2b65aee1e302fcf59fa664e08a9d7df049ad7c98b6015777f73a5020358f738fcaa439db2d6ba9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3477194afde1573ef73db6c06f8e13e2ef4e21c682fbaa413808af0ce91fff74d39af6403996ce07bdd5db3d8edf2c511bf4c97348e7717979415629075ed8abdbeadf2e4154782b69b1dbfa94a939a46641482bdf9d74ecc61540;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h117855328457321cf7deaee841e3af7182568586b31f044a3fca02021d681e11e258765167f87a48e635f27ac5d6448fef471129a325291f5bfb7752eef144d844b30468ea10a315eccef4583aa0aab1c66c404917671ccdd60bac9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e896fa6e00eb385192f83f053c8c0b1b0330ea0784b5385c4486aa627382de0b9396cf2ece46a313d2e3995d372cf95701e1389cb6f1a234dd6f8e46a9b451e483568f93c3390a21713ce715560342dbd5129c90d2b48d89c1561d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbca9d59003815ba17e3d99718bfcc390abc38c35ae32f0b80a377144d4eb54e0e5c2864c5a1cdc9104917f6382722a785499fd7d57ee090083272ed89ae50839d71a0100454f96b044d62646435209455c80bc75f5bea871ff04f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a7c5d214f3f9aefa28cf689e4ade98bbaaf3e64ab4a7dc590628eace407698f9f4702679b123da0c2a68bbca2ed7682ac85edeff7d0eb7bde2a78496345b7a733484d5ae15b916955f3f800a1137d6261d202b07c3c8a002fa45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fdf96fc5ca73ef3b26c5a8faed472a3374660ee9bdcbb763918a5d15971f33e40fde416325ffb7dded113fbd3b42c1d5cb2d3e989c0d8195b5b61d3948de45cb5369e587ec316e6625bdf68e2a40c0904b7809d04d754b7eb250ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a9eb10f0ce69b464a5035ec701b85d9c2cc7813e8ce01bcd306310bcc45587e2e67ef274adeb42339422f87e7c36a0a76c582b037064a9589774230604ef06c3d28dfea0722636d9283292f67132671744b14fd51b1927d33ba12;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1519c97181e9dfbe9d816d7458f104d52f14710382c18afe6edf66674e68509b0de725fac9aabc44978826e99539368e9b23428ee5d0f4735d8adcabbd470b602998cb850963eea7777883096c45381bbb534eb8f454db846074e41;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3d45398ec8a8958199a5d1220c3641644fdee739cd0f8db7534ff1f10d003a5b969e0403f308906d73510db5e4d0155c2667ae28da73787a8f7edbb031de4129cdd2a40a8e39167a30fbdc2be4df0b35b73b3090a56824e9c4a6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2ec83ffbb367a357086953c28f5073613db334dffd62fbc923a12ac24127841aa169cdc2e35619548a86b2c727b9049536e6fc27dbd2014cc1ca4755529ffcdf3fc3ddad18d5ecf97bc42b108530875a14e2985cae2ee0a51887b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34065d37ad1c41d59be4027bdf159bfec64ef3fabfd5db6f8827dc8e9863cc2e7c336a2533763783df03332ea9f70e588702a789016851feb76c6b4ffc9cf24ffcec21cf420836004f8ea7326fd4afad0fc0d4760be5a03e0f372f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a0b170c4a3057708dd9ed98fd88a3671522cfe44f602b5d6467b1c7a5c69f50148315b8ffb3aa90cbb00faad8cb38697cede18549ecdb28a09dd01e78726212f855a7719fc8096d8109aa155c1531d0023c660cd999548da51e3f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e7bbff5111edb9cec65dc77e19eea4edfd72e43b9ba6c323a431c49340d69d9a205dae626d67bfc41064e6cbf1230e69f87cab904c9e1a8c83a8773a49f88d8a053527e4c426c4817ced27a87eb1d07543a4fddd64790b1ac86a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115c1697514303ba683e831b50aea700c66f3e413a91472449eccbe82d471326c4d2e87b91eccbef62797c2157099c1d13b40a6e46c35e4dd8ceda74b6e0e529737cb3adf5ff960950a1bb0f90bf5b0458d3d54cd7cfb881bfc8bb5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3c12eec797fbd4ebe2824e59fb3533a9ac64b3e2f1b606a9953ca7680ed3edb14148f402b8992cf70fb2a835c13304080fdcec57712687c3fa7d798ce58b59064c12f630cfad31b7fe7548343b1d902b345777cce06dd0622dda5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40dc8d0f5bf79a505b015bb4a9679167c24801a0dfc0fe6d3e95ef633f0c450e80c61a3419755803b6d6e6653c06ba6515378177d1231c22e3c60b69ef2d70d41f5eaade3c9d14e92805a8b85f8874b985dc0092d3645908532ab8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1916b718fe08875b99643a99b3ffddcef14f2393060894c7bbde255e400fe8b424baeff465911639c7be9a06bb2b03c55820a10cf6a524b088ad1a72b6607372063a57ecfaf95fd82755cb889cf9cce73e348926ceb95ebe5bc61;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h684392ca0e076c8fd8f7f48556a3b3d025531c41918c2250ea8ce5f6d273b09fe9eb17edd75440ccd53134d5e45c1c8a59de7887494d6bed0c443a1e0ae29de902b495059fb32314ddc6efe064f14d46a86a9fa9f86399e760565a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h74f7b02f4c108831d34bdc87957f25963ef1489f5a8cc7e3b2822ce0098e89c2e6b0098b868c8104e113fd524875cb2cc5d27f00aecf549a8101f44ce4890c4fa35066fab761a1bf5d4338597b5e5903482d662bd0b134b356b59c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf609b072ae982aa4d7f9c10c138757c7f9f89003189684ae66c9f55c46c5b8930eee8d5f2817c7a8f8d1a752960f013bff84706a019adf65fa79e1bd6e4170935bcd235ddddf10bd04de02a9279f697934b84dfb0649265030f2ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ded74c90622201b3b46aa30fa2b40ae7e203a30772a41c615af1b915fe04730f593cdc1e324caa4a33f632a907f7c81e0c51b6e079cc3dad1d3a45e49158b59d9d0767702905bc096334d76a6464a1b4bb3997086693d490889912;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d918e37f8563308415436658853a726b64ef036fd1663c61777a816a98942ee45f1b9d522cc79f627cf071390e9dd634d788e05b21d5f4ebaa2a691e86626e93db6ecff50fcb7a3ce87e31f26fea919ab1564b823bc76e5c83948;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1384b43181d90f28ff997cc7e4c5fea63fc75e98eb1297d5225175dd3bb4ac32c694d5c625bf3a1bb26f7f415d4b793fa4134c2600442730bf78e148ead1b49a3019fabf30b18723cbf023e2a718ab3b8aa5c7321dc5c76daef0e97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b53786d9c8e364144c2bbbcbdd5dee1d3fd62bba7882b944974b6e081f4b08511de2eea76987569921e86922477d8c86dc9a474b4d36b5e0a584f2ad0f7ec5265d701273b197b5f5783447464f9e8356ccf03c0dee26e2c493e31;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4165ed387245a2160182758f6b441a242ac843d579c3c7d6d60426cefef8b19073b853525ca3faa9f6861f795759b361ae1ab0599ea65b4be16c3ec99e368a8d0277f7aae24dce47de6e01fe34467df524bc58daa1334624242681;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152917bc80d15a41d54d2f0e3b3266fd3bf6cfdcbd5e686af27d51941e3cfc611356673f43a6681d4fd65c28bf36cd5e5504767289cf45b8b442db5ee9491d452e5f52433d0693718a73018ce6e846ef43307e168acdb4b00646271;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc59d237de35b4e9f4e428fc612f325278dcefafaf2bce94843f0d70848e643615d4e42ed074b954d42406bf64e8ef25f5d1b9528b1ca0d34242812ecc1d013af5ff0a0b4d8ab336768fb84c667696788bc7768e80712ccf3ed381;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a3d79d8c24928814a812e70dd82d86c6a38ab3e08625f4ab76a6ddc04213e4806af60d13bbbfe5597ffd593f037d5c4de524e024df00b54f43c9dcf0e1eada7a89e76fad26fd585137b041a1c451933efd3e66a5fe0f49b82d127;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14bc9e8d1cd5172e42dfac202a85f7a5779c12f23556ffd53e09c9f858ab7c7c755b18102652ff74bb12975216750287d08c873aa76d321acf2d942f2607670ae8bc283d74ec03760f55903e87d72ffe12207765e81090b6a50ecf4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30a553718061f900975d9cd1211aeb0f91f9e55ab4bbcb602e39ee931f9d37960b1dcc606fce4cc6385b7c44549c422ad943c761b5e7ca2f0f714dc4a24e53f35295e317dda1cb9dadce0a3e22a06fd33e4c6586a33ef3aee7ff25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e06c0f416d47189f460858f327f66ea5ed2d5a697a4086ded4381858cbba7998dfc3a632776fb155d3264209a2f4709e20aa31961f3519f1e5247e3d13b69d208f4218d3e46076aa5f9f0b61faf0e4d783ba35d14622034c87762a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105e210cd7ae04363a89415c318fa0ed5211d55f71baf6073762cd6fc00ee6f8907f5a6c4433faad192dbd610066466421efce357954ee4c0161fd9cc4feacc3e726f8e5ae9c4ac5d0cc1b8a7be4d58929af6e683235956e83091ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h766e5969fa53c585f9203ccc17991a4bab6433e44e93d1a93eaeb108aeabece48ed49a4c74dfc9b109a9793b415f99e1a75e3bc56be556e05c7a894aed97e91fb7e37639917cbdd0d934e31595b7c14042ae476cce8eaaa92cd728;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170865f57f373a483d0d517196b39bce3dad8fd8a6003c35c02b9f08b269350341990f2e5e8e01d9887f145534b28ad49fdc72d5dcfa42f62de2548c8b4f954a357af8e54097c1c4ca03ca80473431189a3844dac9633a2d1d9d2c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe91687318d535e6b8c7e2f2af67a88c41c882dc20178cac05d1ae647865a599ff2f29884d5c0621156e8a5b3f58281d5d26afab2d9743eb7a76f9dd0c42f31ef337ea9ce2ae732b508eae7a94c9d76716ecefcc0ff3bbff9b3431;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6122083d04bbc5c9ecce71f75a1d2e70e1a09f6abc0e9bcc4dba77ffedd103106390032c6bb482ff48735c35d23ae3e8bb10fc31c6a6b79072468632a48f4562dcee88dea8a0cca9d9f378f53635c363fa6e2c24cefd339d4859;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1532436ce8f30e7ac68446c73f7bbda12a4e9f9f332964910740abbed8606037e0bc3bee6a3f95085611c8452b8b9b2cf203f63692782e178ecc669d70d5d44424176efb2b74cf206381cf43991a5e2f866c1cbe2f199c5e305d817;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcbe78c8d5b51544fed39518fa69a2506678d9b74ee6fb073083b1e001e38c2b856b13d06902b7389a37669c800c73ecebe2591eaec346e4e4d682cd7dec0e2fedc773e41a0ce4de15b298e698eaece81de2bb5d5964820ca1d73de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb428f6ca8d4ae3b413138deba50bd0e15e563acadf52dc56295b9eccb5478777b8f0bfe175d1cbb8cd4e13e59a651efe8154475560ec27c170a8ec5aab60219fd67adc386b6eb356620ab999068e2e400d39c61e759c6802f3ddca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7b9badeb776945bb543375b1e036d69a0630709e904167b5dd8bd63b88d604d36aafbb4b8dbe3473686940d9d34e5a60eaa700fb9f22f48ed0b0e8481e9735acf6a5d3e5493917682dc035847b5e50a95859f319147676316b169;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf15b709e5d41803871e4f5709373b88f0863716234c2c6def24611575edcb39e3149b92f4f2b0f8c4b4a04bd95732d804105af997b5ba7db4b5faed266ae1306b22b167646114e7e359bbc724502f977cae37db3794ca1eaada1c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1091cb33480921cf20b05fc9244b6694bbb50b466e85004106a0bc4b7ba8459a50fcf08882a3aec711ebaaf979c729d53a72f5299724bf3c44373e61825a19c75b2a09c84d66a9f0aa32169e60e5123065bd7efbc9910686976d6d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8b1f97716e960ff805207ed64f76a1452287e8fefc9f29dfaf826673050f071cd309ec225dd362628feb44b9b5daea07adacb3c9b0299f8d065ab536616d037b5ea8fae85af1f3665137fae69069266adbfb47773fcaf4e5df919;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h312740a6b3825ee81bf38e116daa31ed76b4793aa8924a334e8d0449a754e1517f6782ec9c545529657ac7a129283a1c746e7c79bab9cc04e647a29ac17aeb4aa3e269ef18729213ca33f28f13550399a76c15dbbf986ecc336122;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcf25f27ffdae8fd9decd9db861756d90f4204f635455de624ec7b9dac2f519c5a343f8621d44536b72b217617529dd8d96b5cd54159e6187da4b18276e0b82e14fbd2b0e49e5e7c97e4788f0b2c4abe72f46fe7ce8b95f6979d57f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce84d0d8f5822aaed27074a05f16220c2509c8c1b926cdfe578a776c50cff100405515aebc942f8255fce3074d700d985c4e41e32533762a9ee2f4cec233efdefb9dc57677df62ea0a453b2230be917873f009170db662e0dd33c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec0fde6274699fe056bf630fe4608723eef18c032656f433358c674d50cf3ad81579b24943316310ca267e3c18bbbe69632c50fd4d9204491381971939140dc9806d6033111ef9a61630a43e0c9360af8437bd0b0e71ee30078a83;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f32cfa458233b4d23b2cbf392fe1461d712eb257600ba7457137102eabad8edd0cc2066dab900516bcef22d11f37d000b37eb3278bd55ae30593a87e505fa442f3806582d16babd050c6284fbc4f903cfa7acba896f4a3cb5c5ad7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11717e1dfd084578ef86efa8e2488312474e0325ecc1a2abf735330bfe3cd31cea5100d7e8c88e9b6196e3a892edf081ee814de01c8d3f8bdcdf012fe2bbb10df18a8de6514a3022e168c61b5d1d461701cd55a150c84721211ddd4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5fac308f9e39fe0b4853acb767675a2d5e1bd22d21d585af7def060275fd9b3f61aa43592211dbc3142c9f500ae2b1c92f913bb47938207b21ecea426e7c5cf7bcd07eb641082a9fb4ad1f58bb9de3b7dc8f834b580dde11d5319;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24621955071cb3612ee45adac5fb12431ed5b8752e5460dc39410369895ab5b00c8faaa7bfe7a38ace4d1330e7190f3589129f8b6676ce5d0bd7b69352797b2f458f791c790d72f2e77352307d4748299c8a3722053f870fc5c91d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffdf187de15e8d7ca8f86d6bb1dec9aad32d0404e982918dde1ad6e295e786697f53f5e52abbb70bc2d08afd11786bf0ed73a4c61ff23beb116f1ea9a7046d7c34e85e84d89a739a4886e546bbf43755ead6204445e3aeaef64d02;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86d172ebea6dfa32f061d2172c9c23d2aeabe3a47beb6cbd0e22314335d1072aca491b5812f2bf45df267747db92e6ac7a6bed7612d2c9da1cae1f6527100c2b35789d9ea6c12d4f61daacb72b4d42d4312559cf96a5ad36ddbcc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a06bb6a16a70409bb70f75aa4771562e81efbb0fbecd4011e61d1178cb896e8c70155e7f15e23ebfcdfebaa5db116d472a33eb467b4d06cee3c1e56794ecb9d793890426beebe718b1ecae8bdf5951d9fa661896d5ea122223e3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5827cae69079b8a68a689ffb1ebc8136a07e0035df84f3761076177520b5616a1f1ca2bc758854de21bbcd88d3862089d31bf1bc36eaa9a4e9264a6fffe6d340da84c63a83c896de8cec63602425d603e8dd4bab4f919704f826ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8f8abc7ea6205d7e9c0334593c14fcc32b13172770e1813424bad7cfe9645c8c5d5cca3588ab261fd8dd00caf3fab397cbd41abc3dedade9ddc10c8a6f039450e0ff86698ffb62144cf9a09e2ac6eace09cd1e2c36251c484f088;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h608351b383d46cd91ce8b4fe414a93858d35e69075a50b70dca1237f92c338cc4c80b78ce128e91749e34f38ef528840481ba3c50ee475c061efa315f68e0570390e24c668f2ab34aa5ecc5f889394beba06e494dda38673b27332;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ee0a32a4ea2057326981017cb190737d369a07f6565bc0b3c556e0d8489f2775f6f6d6bdb9eb2bf8d497897fd0940c4219efa31fdfc81d8a01d16eca2ed5adbd118478e9c98387de840aedf5cc1ffc2bd4797fe0ee183050baa2f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123c76cd5517d83f8c41ad695806f88af3c4d2fd8ce2da97b5392f051fa88a4319acb68d65cf4f64a517baa13c104a1ccbb686d04e9e62c098d0eb935ec8c9eebc2432e220cf593e6bfc571127199bdebd1db287c413bbd643455ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b6986e1c9e27710b391089e4587f88482c3b258d589eb77049705f68cba50089bd0224fb1a819ae30eff8067f4b608dd697f36b67c76aa203393f70dee05cf009c1c2d542769b7fc5cda8be9a82f17472ac814bc0b437289514e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14387aec8218b1ba5acc26f31b2ab8f8ca72f0ed8a7aa40926362f05386e2d4a7d7751fa203af8153f1004a2acaff403fc6c75cde1a1c3763b58d63ddfe9542fad5a7e016cf5ef632364d1ba44cc548265aa17484883d33d3f8a98e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbe761bc5f77d481d48bef96b6cc1dfdc550bfe85f6b9813d7259b6bb60e6ad5af49b883ab4a28eb887bbcceb349b745c4d2d6974ce5662bd45bae2bd0fe44ddab8708f6344600de834747faca8c665e53d7d7af9c53dd76842dc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd16128eeb032725c7fe450d2a73ae955a719a7a2de729cf0320c8db2251722512802654a6326357cb863cc455d05c7ccca4113cb87bc17cdb5c0b7da346565096feb2f60a060fc62b910810265a5ee202774ce3ccf99139883fdeb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha17e03fcd393a7d8cd8c7aa0ceed7c6bf60f802b3487d283877ef962fe5f45604b410f8e393233d389ba6b70bd14dd90e111e7231c6b8a1da750c19e52b19bfcf5bb2083c9c1c7d5a8825d677f67d2a83494c504e679a39ed46508;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h318fc69bb094ec360d5ac52439be6df2845593bc5ec0ef97d4347eabb3758a5d3284189cf8b517a828dfd2a824abfa49a175c31fe48fbf6110e013664b2debadc2aafda54dcbd7641832661d516a2143d6e72afeaff052a8967101;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137ee7a31eb14c81b86e0da8d4a809f2064e59aa08444744e78ad61e1b768746c2527942135513b5e8f0399dcca324f04708d3935365ab01b2b2918760e2c85c543771aed7c185de0687a43fc35878ee3de886477d317f5763109ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9c3abcaa1f42bd4646a4fb01a987392bed82cb176fb935cb7818653c7d8db0a74a470778c3ece44f4d838d2a296e06ad1abcef7c4cb39e64235f30c702e205400c855943eea321b3ad0e638a732e9d475287a53f1817f8fd45ae8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb18ff2976aaed1c5ada0e5e5be75ff55f2e6092dda7c94b48f6d8eca842b4d234ebf7f566d52a888036e1c6bf5dda98e7e82af25c0281cd3c452752973bf743f085aab8b2d1fddb5f700f809ab75bd7624b0326b4b5df7663099f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8753d9b33eae011f93fed01da4ae579d68b77e848b31ec4199887bce66f3c6eb3f7836232e1b8767ec1e6d3d167cd149e83e2feda313eb4e2e755c064817ede725f8129e4d3853cc6134f16c2fb25eb3bc1caf7f0b20d4f4359e46;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8e0ebd7a61ce0bf64cccef19514a858d1f9885cbf9555a6c574066f14755f4e3714d914e1146462ad99d22d10edb982016bd6d76e4b2d675d192b44bf8620be405e5a3a39688666861caec026fd25a36b95a707cf300c3f00765b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd3fb14b76501a602565a3b4e4c7a6c3ca5430c0df8e5905ed8282a0169c3a455fc1a9fede005800e0a041722fcf861203b3ebe0886685c7f90990f98b664c17801ec052277d761b9920a232b1e0ecb0dc465fa98770fb96fc490c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc568604995a23158e9e03e0920b74b25c8649e2107ac7f970d21f56f559ddd588a299531d7dbcb6a8892424120849a56a3c96470c8e77d66f98965eab5fc4d696cb8fa2c29bbd71a3a4c26a0e0dd5d88026d33cd8577cace9f01e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7161644febef8d60a7fc2b8db315b1da163fe26e1533ad6d4975d772fcb55dff12d4863fbcecdb5f7f578a176723a7c7f2647840afd54e36fafdca9d80afb4a4b0815e27574431f9205f814966f833b2bb9555bc3441449b668f45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1752f4b9a5a3dcd753b8b4a30d19ff5db6077f023ba4369913b45937059cf95e5597876c95963edb10b36ede34e9c36a078f4b17be4c99dbc4def66ae810475a971543e9ba92016383b52e1d64ddecd778e132068848680c1d01a39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c90117641230238a164830753107ebab536ce2940a6431ea4374a259de4436cfa30f5859e10e7f89462a784bd73fec60224ef275ccc65350868b4f163b47dafc57466718abf31bb6169e8075a964ac987b8f68c0d0b80bd027a631;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4d55fc7fa1c3d5bbb30afb8c6a0fc7557087d8d3cc7e453536cc6b616813fa4cebd1144d3d0a35eb0937af2e493b577a5a029f8cd5ca8f0bff496c45a34ba218ee5588db9ece79628af098d4d6d0cbe652a426ccae507ae1543b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f259737035a0cc1f975c781aaf3a561bc24edabb6083a58d1e02cb5fb8c220186ac4223c533f1779cb3be9c4762406a3a33fc5830dcb21a6832d97dca35c35cbeaa9a475262b53a8339ea328ada06b3e7bc5140ac7652753d21c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12aa61d9c0c18e5b02cc3d1c7b852d29185ab3f47495589a9d59277ee37d9c443cd05847025f716f38aa236f2b3613506aba75669066386de2293949035f11e0202b8574118c9e6587be1488cba3cafe35849ccfc5d501d954702bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b323b1bb536f1efc21d01a70a8be7f1bb350307a955599b1587562515e2b2552fb5673f148615c9d0f761f43180101859893e4805ee39acb3ea3196ba4467351102f9cb9f717ccb64e47063ba58a58249b05cbf69ee4a0c67ea208;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3742e7768cc3758991a73af3d3e83d34cbdcc7c8f98cbd6d3a59b004de2b51c8d9aa3c15f81a5f962b508f972bb54b9f223ae7abe1b06cc704a4c16e2451cf56503c0532b0ca68a0727d547a3d7047f5398348c9524ce2af29546;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18161b1a29840657de1c53d903a67105e89fd10600f9c234c9d96ff021beb2fa8c4bb8982ba2fb8254d0a66e2414f444f8de05cf3716f6b5cf821cd99927a40ebe982ce5a672797bacd4edd0d702566ccd14a826848e6701b15db5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a72a0800d252ca4c3f43170796e69012bdcfb6157c6a6f81a43b72b30690db373e47ddd837adb127044a4394c8e57fef23b323c20e32613f335490a71191a26c28e324574807ab173e1706e5fe3622a4753091aaec4da103dd0c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bcebdccbb2f9400f74d79124a81775a0730b2650db78510dfe987d654ec853dfdeb45ebd8d7ee4d75272ef432ab026ad65b74e1464a91338accc8a888e6b4e516b97db77e5b80c6ac0f13425c09512e0696dd138cec0e210817271;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha0301236c15eb9c348bcb4f235ee165737424fe76b8335c68375b6f49dfd1fc69997c2ee6739ab881d9b8030a5372bf9701f955e797f86e86a7ee591a07e99325eda1cd2fcbc3b7a58069ba7938ae2d6a8e0691cf534d8bba914fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6601868380a68cb7c50a8d38c7c5277f549b3cde2993e6309ebe84b44b0b551d7e3b99a09765f3b1eb11431115bbb417a92798172fff462223042a31382ad68d53d9c8216a529d87bf4dbc30feac8bf904a75155e50366128dcfe6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heacdd06cb93af7c8d9ded89af240bb08c688857dded43b5f44e2f4eb0d602d8d0981c1fe49e9834eeaaf1d91e335f79b2c629492b56aacfe6533c43bebc75a359fec1d63a22aaf7bb64e3286700c8b1d75ebd0d5542039688a073d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h321433942de12e452e04b4f750e9877c20e9953c6013f02c43fb233654306c8a96141732215826bcf6f87157401ca898caeebb1da06a21ed418abb92bbbd7cb72d66070c60436de5e335565b80609335c5a979307d28fe30b2bf13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb5854c07688b29d2a5b4b3e5372ee5056c4140d66d30d1189133553d54fc1ca9754aa405600cca07a14e187b7c293186998bb3e351207bf371dc7fe76c82126eb96261f831ad04349ce7f4c5b59bc5f5b424b6f25de4e09bc023fb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d30001a7d77ba5c0df1cbd36d9e18b4c79d8ba8b5eb8f71e214f79b9c6567c97837ea2e76aa25a4c8d07691546ca3798db611e53407de2852c1f6161dca41a620f264bbca9496d874c3b07b667c06c51c9e07e0c68b97b5227ef4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b493a0ea508f52953f3df89711e376dc4b4529b71daa4d9328ffa01a815d870182a0c48e4fc7cd2cc44c8fcdb22a26228911918b40ca45add11e7bf3c17279512980d94ea5bdea88a1442c2c4a1b9fd38de15caa061c8fdc05325f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0ab29bc50025f802e03d5350186268448b9a972ff9a772dd3d6a5ac77f902340aae73fb6e1307bf449f478c06e60a837991939a40b7e4286daa1e3601757722d2d37d4ff10c4ad88c0bbc977745ddc7af325acde92631be6a3230;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a09ed8abf7ed4191d1069145be97b2631f4d415f5fdbe064190ec8bbb38151f8cb6c57c34d5ed055a608f25e61390defdb6a04903f5e7bbb2a38198aa66a5e6ea0cd933059a551b846605e4e32f478fb8fb5f0f90787d48c73089;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h28d303328b9960ca59ca8e4aadd8db015091d7fda11c82f7f1a0d91618393f118bc8e44b10ee8a4f72ccd3e0a29a71294fbfbffc6116b92b878c3d9ee0a0ef2b6e3c9a00be8af91a11c3f70767642585e75a1ee83dff1f5136c10c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cbf485092af6f4b9e1b621644711df4fcae151111659babf9f939417724374df1d906c28fe8854e6524ef9f11ae9a02d3643106a962e348ac05016b2244fe24cb6aad7250e93b601895ec249bf963856bbca674e31e7b7bc1b8e6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heff53255d084c4784f3af64f83c3c467be1b4c12f887c2db49c785a47fc0c3152d8dc08c0ba565377123c0a8acbe2aad1f04e3b56d68ae7d0f8d00100102ead5a0a71d472392fb540903ae3fc11a65cb7b43456d8e902896bb8483;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aec7b87b3d523cb3b2a4b4035900130574134a209f7130d93a1cec68eb5755c5a64fb6a63066ad640961e2fb7634a7d384d06cb01052b07e03258bf14a0432354a4a514a69c6af69d34978bd4d33f1b4658df4e7f0f5aab1fc928e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f120083c0eff875f6954d69f8508d7afd4d0450e60cf5d52dec2a308eef9589e6a7879f8f014e2399c9a55c3484e60a9b8ac41bf46346b8a2ec8bba824830d1e6b0050f0eb234f5dc622f4b21c72a37166efea9de5c17102568df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1924270cebd30ea2fb683eebfc8c483cf4e633c707e7219c663048ef303b3728b056f989f760a564cffd195f66ba3e770c2efa22b6a166b5942a856b305e81a47576de2583912039b17aab10adeccedd48c7fd0708e5c1c6e4083;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6b37089a5cca74d2dab55ff4a392d431f228ea6233d8cadc82b30d938ff1dfb7b557e7b7e8bb2b1178511b6a951205e470129b20b17fc97ca3967b8bd2bc82bc1db5e94af33f4dde48a0f3aa22d1228f3ccab6c8c51f3b014558f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h198f27dc047dedfdafc3369d65cc1d316b058a35208bc8577cec32be187ea7c52cacca99e59d555f531f4c79f2734b7a0af284d61d1246c82745f976d3c738990ee34701c81d691b46410f4680d1299d5b92cae67c44e5cb8f3648e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd2ba33e078d807a92f7fcd5c8bc31965fe5b6f0b3ba2a3b5824589d12f68ccc0c97ea9b5a817029e76e1c2dbeaaab4ae83a0c4846de08081d9b01a4593a11667cde836aedf5a2f232e7a7eb0f067974460ac093b1d4f791763f4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79cdb2fcd47642503ba8490e44d4c57dc0a61d63cdd7a1ab1454130ffaf978abcca067c375dd3e748333e36e449b4f683344ac61892692d1b6b60f21bfa749f41bc8b17f260605c459b469fb733a1995ed3b89e841ebf0170e408b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h52e3cd8f2038fc2759e35a7eeddfd9bdbe704ecd5f2ff81b9dd7a37c7cc2404c293d8e0cbd35c343af9f22dcfecea0fc821626b2e90dc3134da294da132fa3013643567cfb8337e6ebf6dcd97ef7a3dcfb8844f7582d35b9c60365;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1debbf7e3bcdc462b63334e0b51780a5b0d0d120dfac9f209d0aa17581b13235eb3e08f4683907dea71bd2e773cded572f06f6d11127d6e6c815c2dc0aea533fbced4df7db90f7dc2d75168b267f79c863d716ea8a1122abaf02712;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4eaa0320050785d91f2d3e803c788ccf3f952178b6abab2935ed5fa971d52a08d1d8934414d5edbccd982422ac9a69174db1b27b9d35d4d6754c5749104bd1b8675cf77d226a6214bc3eb45808f80a2af6c662ad66fcb7b3553a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea1f0f9f7846eebe0961fd692a75dd353e91f9b45c14cb2c53d02c56d929367ba25b37d71e3783319e237217b936a48fa32c73c963b6f3d9229f7e13b642bafde5f51b2502fbd52331cbc7ab54f47754395d367ed5f14b3f06d26a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b7c613c453aab41c1ffbcafb9f02db855c55cca85a3fe94d5beab291f6b94a55facf2199c140d21b0c78102a116738f2d1930547c4af7e0343f852ee94fee8f65f91e97a5ab051707bfeec95c124fdb2a76ec12057cd8e4ff681c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc42919591add36f4e7edacac0baa3437766fa042913daf310f291b2f12f90396bcedf609d4a19729003bd1d6bbe04df6eb615b4035d36cd76e5a962dc0c427140f7b18e10e7d0a69caae6a3dbed2f46eaa239cfce9906a8938cf26;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a182bb8247790ffa4526019ecc26c7d41ad674b99779e6fc2c235f0e65ee62962a95fce89dc660d88e1ef0aa2c7c4e365bb7cbd3d641cf6f0991cb1471aa93adc40ca5bdd6ad2d16bb98e6dd543cedb028dc5ab559845a561abec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4becae95e2e246287cc47182ea8ec6e36a69a2a02655c2275b21425c537cdc39fd35dbd963324a21a48054e11220ad53840b06b33fa6b14e81dde46798e8e7d1132d2c894e99c0ff3dd42d8a85b0f1a4c5d9c41da9b14c723a127;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb8ad2dbf7b19505b707fcfc92011aad2fd3b2c711a63295c49e4601989bc346c386286470bf748ff2513809de2330bbb49257a5e941c37b93d1351eb068972bca4148d84878169bd1a3dd8e9a636c7532fe9208b879002e0cdae5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ca00ec9ad3d871d31d376cf9d51584ce99b9e18fe6cc3ddcb1566bca41c35a4c705cac4d0911ab59db58ab11cddee9aa43a05c45ba95d7e501b3594ed0adf71d9dac2d18c6ed9b397003848857476ab0659eb836f714096c1704d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e21489c69a380a1bc523b00499ec81384e7ed0fa9def34f2d496a3c83142fe387d14a1e6b4028012dc8f06a0d67bff05d3180354185dfef1c5895321712f3c4a579d130816790c9eafd393306857fd3ccbb2bc35c25201e7a8c390;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9800a3a4eeb79a31935b22c1f7b0ba990bb3c9af721a26ad97605d5628ff0bd777992494a3a4dfbfdf71afbd37794daf1724e42bcdb90fa794146060ccb781de9e70fbbbb8aedc6433f297501db9f249991cbb12feee99df8d93d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9c59b88c8eb41ba0e6c078bd9c485ac90e64d32b1a837b1cad71a2e2f23aa1aaa26fa7990d69402d66b92a67321cf1408835760fa38b2046b4e01112f82d528cd3acc05bfe2f76c9fa5cbd73c8dcb11a0fba67de531c2540ce623;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h599937baf2f1e2a0fdfed1a6ee05b56c42841336f41f5c77610fd9a9eb25a66da1d0b135c11ba7abefecbaaaf6d6f0fd374a82c2afd19975f75c142cca63ea604f6cfbf6882bc2bc9ff36e398fbe01807a776a79eea63c3185c43b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf140f912aff4532e5c4b938bf2dc01b6dd7403375c852e6ae9fd52d3885afaab911913543291c8c52baf4c4cac7fef1dc2b3c83259b796eb0ab75458afa3377a6fe75cad282443a4aa24003713c22bbf4a9010a0466a31b375ba9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd08b9b02037407dd2ebd23c37b1d640cc77008a255566367493e08ab48a8f85003f24d036abc28228ede1cada21c0d3638f7de89e47be2d18548972c676075c594ef6c19cb38eeb0c2d553281352437218a6e883b540f38fed395;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc343e93e7cb096fda014c509dd9f18109290fdf4e28456986b9dbccccf7226744ff6b7492722c5c0e1515ae25261d4e10cae93b0779e6dd712efed7e82dd8def818b15ee378a40d5e908c5686e9c4ab483846ca461f051a8c2563;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6e7a662e6219ee574f34853d842967774f8912cff4ec375856ae16f0bc88c45779e13a4e16cd7d2519cea90a2a65872ea369d2281e7507b3edb2dd1f08d723352efc9f6149a82d5a3abda16b48a2aa13381393039e0646dbba5af7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2dc0c826f9ce455a484a8046e7c090bce58c1811ac0e61103cb7cb343d98bde3e36e893592b47a2904201614f991798428b14af2783ee2a94e65ef53c0f5d254b868525f46887954d953ab273fa471eddd8b54e27a6cc40449cb64;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17433b9dcd8f99242f5bf8d267654b067e524a578e39dae295ac5ddf359210644feb30b70f4594348819f7226d377d793ac1cdb7c4d95369842b5c52a4ddf42ae63ceb551e5cfd7152e853cd4bf5c5814ec3c201cf05c9d0ba36451;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a82e4bedb3b1ba90cc642830cc921f00bfbafba113b7eb6a13d370e4ca4e237e7d1aba9ce07060851c9f2118e607812fdf586a6ea11561ba5ac0518d77e4f2b6f104299267e9ceb05b3bf54ce3556e855a51e3980fb4318a70483f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f50aab9cdc342f8065054d98a54a4ec245a267daa9c8395d2c8446c78f291b1b1af2af31b2307ba4abb9cf08c766360a2fdb0e39f06e09b3c4ddc6dad111aff977bdad1f44df362aa43b1846f4b6decb5c9d9a4fb61fd009b157d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1e0afc281abd70b72614cc0b18e02e2c84047387f549679e09ad40757c6c66a035f9fb81eb4bd895a26916a29b7bdf0b1793cab28326668143a362eb27465863eda641f1efaed7c6681e206fa1f089c106a85a02f70f0afa41284;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h774fcfd8025f499cd4589be1af8574ead41935de76229bfaa9e9b068dc6a50145cdf66e4ec1cc97829c1f56ab7414d9c5c585d8173ff1a4ff9d3676535b820d85518faa9854aa9c23ac71b74213f6697bca8f52ae6b3306bd3e973;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab0e75df96920598b9dd4a42f142629c3fdcad8279792c8e2d815492ded3ce690e6f001f43383b4eac5238ac79a0b61afd205ea73e792356742b7231e9762043db3fdf8c2c3e2afbcbab7bdec8f4c5801ef37ab532f2ad253a8fdd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d9768418d9bd6bf94a3ea4c0955db5be30f54b72504252f1a18806469529d34cd095631822826b2173c39aba570d52d360feba56b488d9108913190a3422176608217841f17df7a283c7a9b9714a0b34a92b7835c534a3b66847;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc3d795030447df1a5f0d891f2506435bad4a7b7a7baf602bd2e3c997b602642961cb391186b44da48575cbac9500d7b880146beb3aa1091281d3c3adec901763f9cd42c9906f8e78ee3c4614fa54204feff63d06822f71e03b77c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1164ebd52e188cf62354b412c3258f528fb28d75310990dc4124fe1a7621484c4fc33572302da6772b1fbc3ab21c4a55952c9ab5a12678e896d2a08eb1f8c858ca88b825b749ccdb4031d045420c92a7339b2550b6867eebb925366;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62fa40f5b413c0d388665abc430b25102f8becb4aade9475f3caec2473b89e43b993071fccf8ec2f30314a44be9ab7b76bb7fdd85b80ff0c32b335fe0c066e88befe6d15d2c5030316a40167bfc5865f2fee922f7f27abfd7b18d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bdb56ba65e1aa3af5bd673e113416a9c600e909423ae5855b74dab8a4f4fcabf20aa81924f4ff311b5a22e3e5e6294002df04706ae4fc1b13c70e9279113bcef9bdd0fadb757c68d76499416121a19fd540774ec7654cfd502fff5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40de57481d19e1cfabd9c020e5302323e002fde64eb5ae4a80f117425ad491c2e8dd9266a316a0ebc1ff177a5d4b38b38c5d132f89808caf63b616bb12f3da0d3a6bc8953dc0a27ded05e9548b2d1310f34863e678abf0f550d92;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc0793ea5f4cf5a10a7f5357999f8cc9085d2374078b022f5bebed32ffe5c780f5ddc416dda7116642186931289e74fecdd81b6b14705eba927b7a3d5a534fff983acd8075bbbcf3e08f81c4ce0cc97d006cc2e51ffaaa24558bcd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e9183d5c7e05d476c2b0dcb5e39dfe5f10f00a5e0d2ddb42a615cd9668af1e0b5ef9e4b0e541aec0fb406200fb3c85803e0b9e3b1088ebe315d9ffb7427392e24fffedc759794e0662e9fc7ec8e51bec72e7b3f4d3e875a458790;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h39571cfc7d5757ae873588cd42b862ae18b13a414daf4318aebc7734ed77cfaff61a9ad5bcea26cccaf3d6292a25ca1ddaaa85d021e27bb9d39bd4a5f43ccec74843ef50b608b73b8fbf1c3bf4e30458e478de9cf42f1748fa69b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1922eb80d4e27843a1b4df082a0c32131917e4c93e28120bf33f35d0602e7b07190af519f1d07de64e85d3758f24adc713604aa6dfb75e2cbba04288df4cab8fb39439eb4081ec917ef09ae8f96fb1816eafe6a176f871645caba20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1fd1e9a4bc93118e2e1bd9df58608f3f33fc33467fff4e12a62b816b6f54c0cf8444e529a6559d0dfc8629c3b1b0d84985f13d17ca111512415649146c327e16fa13d6218649e8b89fff14771e8cd18bdd89fc16f25382e2fcf98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e21921dfca0b3cf7544e7edf62aa61953ddda20d09a68698253c3e15d5d0607455f488849a8017e28988381c0fa4bc47b13c22deadf9480a7bf9a83d54b5acb32391e04e4de2fa6848327c8b7765d830190c3bcc2b628da9aa38d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h117981087e3ae18aa79bc69880b878f084bc3f1494b0b79b207ce201b1a1ab46f418609f1ff22f5bf46a1750ed499893b2e387a165d81ab5458db5ee66a1eec03bfc0bea9e35327be999290a77861f3682d6cf6d4aae4589f837afd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15edcbe5190a6ba8e6d9f3ecfcc9de562a4fa832c5176071bb1e647646553d5d58a245e06f6af906d2fb572d2e0d95e421b1e6a1979ca1bf850813a0cad5e4b37c49af1513f5de640c1d39c5abdf3f3aeb03c9c16d1288a440311ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16516e4bd7aa6d2cefa62fc6e46b9a11e1de7ff93d0607e797862ffdada83ab51c8d5a33782a9ecb0c394791239738475443bff3a4ae3323f1a79bbd53a4b790b013391ceb319114fc93b8076ad8202f65149d6e0be66b3ff082096;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ec2313d35e301aa5d8c39c34ccab252dfbf3423e0d3dcf80c76ce54e0bb1a7b20a28a5597da6b380c198686d6e50661c1f6cda60d619fdfdeb33bf48ec3b51354d6003364f82c56fe3cce15269e2cc7220c314a3e9237c5d31f77;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ea7fa3c7f16c42d86851f8541975991b6008202db01b24231a1e787b981197d02d76b2f5e90cc6162ec82a1420fdd5cc5c19a859e40e17605e91dfef2c5a502fccb28fd889b991e9506e5b46d69b050040d9d675f0467d797c116;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18fe8de1d9025535f9cfb890c8f93b3bce284e4fb33f6bed532059f7fdd4181128afe4b15bdbef6ed20039824d4c68fa5c6fd8fe0bda00e6df09a663d9a68ceef08804e86cdb1974a16b2bf5a59b4f6f4ab4af862f27017fcb33be6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ef2c213078c85145d64e43fabf64788246cb03081ef483f857925cba9ca11b6828ae3c9264aef5533807d45cbd05eeffd72b4cb77c0301e783326a6fd13b0c3380b6951e8929a975dc295e6c6b310a01bc556313aa13bb25c88fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1909ebd7b952237e91a003b7049e852849bff6bbe26b28fd78a1ff09d659e765c73ca42809f24d5dc26e278807aa2e8ef665618e70896a9bd8fb60673a9c4f2dfd9a75c2ca7bd89583bbc2c38d6c91fe803c43b278a48ee21c4b8d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7cfa6455bee57857483d27ddd20d315d3bffe22b390610e7602866d26f9fe6968fcd565cb47780a0e04ff6334f41d8053079244e974648df4292abb133c27c328f60fa47f1645d7ab501d55575ded32263862c708b613cbd8454;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9773106918dd6c7f5ae43072d995f3ea7d12858009044068d0e883acb5d2d9c56d91401cf6bc765e86a89b407e2370d0c8db618814eb1676ea94086f4e42f94198c407de169934e93bec7dde061c183a5614f9035e19a70ccd9696;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dfa81e98d3a80295fdbcf4e40014d7a118d3dfd31e4be45b0d752edc4204bd308ce23e3cb82e032bd9cefe49a6ab494aae3d5ff8a98971f282379894a917b4957fe899dbfe9a402070c90621e9b7a0a5fec7ba7f972f6b6f2e0d38;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he67aba99731c7c139979b95a50f0fbbaf7cff33c08c053ce09c01577e9920a7bf2e4a4229d63f6be0f3102840aeb026f1d96cb63b9cfcd331ff5832f7fe4a956f7fcedab6679ebcfae8e6ab1d33cfc36efd5de3e3088b2a29106b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5bf6e480529a6b8961ace9b9b473de49eae08a993c42996a3a8a7531f30c516a0ccaaafb39edabe76f5056257f0900d08c7a6c06e40335f41942681b936b1115a009be65ebc74dcc639737947cdba19fc491419e6a9c14017967;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8863cabc602734e1875f2638a7baae98132cc6bfca2a41de2e222ad6f3b8f78e6287b3e3c6e9e6e9beb997064317573000dbc56f7cdc75df798c89ee0f1b1517a2223a0f4cc86bf44e9ae36c2181ec02bb39ede91149212f854298;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefbde33db2cdf019607b0afd6641e452ee7d442b1da4c539acbb8cba6741c94350379e16e6741ae5d052dc10c760e25ecec741b2454bfa61138a4c1b46255285aa3bfd8593045509e5ffdcb1f790a6823e91677a3dcefc17ecb5ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16407d5ea2c71b5c256b2b6b44c54becf442e2b1a133421c19f862dd57a19c35df60b5ab2d1b5557276ad555f692328b333d43f1bdf733a56ef469f67a9adc35a23d2f1ec2b09e08346bf1a795d06aced73ec9c480f9fc5da13f17f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126794ef759e96dacae3c4dfdbc7c8ba02625df971a41c4aa7a1a3bf45b1191cc67f8d9fbad8530af666047e0e55bad723fc63ee5af120ab83794efd8bd5421470cb2ec6773d22be13ab555f2171282692abadb31a5dc6616806ee1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha3fe71b2cda1ce468152113f4bed02acf272f7675b35a886d38505dde25db15d707eef2b09b6c65848364b7c7f7918c2701a5b1c79433b3e3ce9b3f284ec4e032abddd13131c44aee09632c58b0aed1416ce45f6e1ae327742fc96;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc14ca3a239ecf5db594a0583f1ee305451528331ef3ce3010cc993440b403d79b504a09c2c4f55595c6d356f92e39309da4ad3bb8c11b614fe0d0b59e3fad0363024dc517c5b02858f8f6a35a0f58435155803dcf125808c84e3f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h138d5c9b49270046f4708d598308ca3bad0cd7f6d5bc48a107d5fee088314735a541eeceeed0c8ea6f571bd65b27237ea112f29e27cd41f08ca80a8c05723cd19489a873acf942a7ccb9d683827b5ba4c96f003faa59ec62781dda5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e2ce37abf8aca55dc9e77221d53e8894d3d387c2866fbc79a678a0fa97909217ec6571a4a0b4e8fddbf16dc1c4c1132879362a32fa4564ee3a17281c8ce17689e2e56e741d1669905e307e6cf591f73f79dec5ec1619656b581da;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14197c34962cad848b7c60c204413248e561708d6d9f5c4fa5c244d0ba54f45113a8af00349881461801920c52ffe351d95e918de998324b13aac6cd1bfa86a7e7bc8b6c946dc8024b0e6ccc494201959f279fc5a1f2476fb176810;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h740f007dc68a00e206da967778a366a42d91a6d4ddecf8ee9332d746321785461f3da807cb422f07caaaa556288bea3c1bc66ce7cb66471ac0b47776e413753112cd1ab444d9ed7b92e2a896e2d340a53d664789011eafd10e761b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2c50ab88484bbe096d2a19f68a958c1f74132bcac613264dd89675a16e43c6cfd4b1f8d72574deb4c342722bbd5cc411aba3225a16a6c386ba285cbb0d7fe78880dd55d77d3d7b3ccb510505c5fb9eb7c8157e3883257df4e4e0d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h162a54de8f760bfc24c5197c5cadc599beb13cd56ac9c001638e4e6bbc333c09124bb84cc258428371351003fcca31546c620cd67373368d82b609f85eef3c7a3a071cba7525ee7a3ec3832c4d90734d2f7a8ff473c984bbc32639e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdde02a51c62ee9267ac10a3028e840e9aa9e4c63cb3d5087e514b13e1951be97575a43e8b7795dd71ab03fe26629753bf8d29dce0b88b7bcc78d653dfddd676dcce154c6d0a4ab3d0bf436f7e42af3d538fe7bf78090a279f2e442;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13255e7950bbeccd6be24c6ab72e96647ae80c0895efdf5d64f6cb7548f94678fbfe1d5e1684ffd91feac62519adf147d4ea81374e89e12db706910bda24f673b7d834d2a28abddaad72a96a4bcf25df227c103418b146105961920;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14babf4cae8b5b435aa07dfcc56c6c21ccd561913c07164575eebc6d02ad0c38a166e4c61c4c5c8852c1313945ae4c9cf0a95eeb5c536a1e7404aaeb2755dccb7a050106f181fc29ef57d794536cc9d0a06b39d368623def1ee78ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h560dd208154ee910b934999dbab2ac3e2cf14def7e236d0e2ab12651a29abcd44cece56bfc1f72a3623edfebd71426ed5db2aead9481876df0dfb4890e2afed6d6161c4beef58f19cbe586b94aac1ac0f536be700f01fd09403874;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29cd8ac358359817fc3f3f2482e411b38eeadc9206a4c264776187d5776ce88557ae20277e6ef18bab4c1481736a8a74a0b78c205efd01fabf46cdaae76a7e39369e4818fcb16acfaa53ed5fea28eb076318725d2aa00d19189e15;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca9dd706599be69f6a7753261feb968b11bf38007ffa4d0043716237c03aa9d19c30540f3108d215a9db2a99769ac94052b095b36c52faa56ee365f1db319b7d6552821235e0e3701ed8555d5b9e26b951a4fe0d360a703031c7e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c2cec35e4ab033e741897d7a203bc2a50b437460b463e4e5d917f98dc544801c3e74ad16581ddfd4a677fb5e1456b664d90b5c596163a9123194d463af66a72dfe88b3873a3a52e4106118fec18e9c5d5eb82bcf57c78a935824dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6beed2998942244b85de663f9554abe58bd2c9a1f2087a8a8fc86d4ec8a47e733db0c1948f24287f47810576e7fedd3fd863afa48018657d0ad648cc6dcfa116bbc71ebb67e1faab46401fbf904b92ca49ae3258dba04ad0725a15;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3867cd6af5c04f73806b840f0f1c7718043df9ad2e896f3ba50f3722bdad72893003b0a792f76a75ea92dda7418da98d2e819df839008f9b8f8e27314201ded3eee94a263d0a590511a35a01d03e7bf1a9a3e4c91b6934164ea38b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d496b90d34a015c0ea7bfd209fe2d31b758e6342207511351f4caa47d4decaf054683671f59105bf866ed0cd822a63916c2c8eff6034904a5bc68565a29d3cc5fa4d50b7c3a46b54f8c38cad955b4644b7dbd8e19be2363b7f35f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ab18fc93eb631fc557aec9417eeb22ef2766271e0577d1cb54adb687e3a27888208a70ead82c53f146dccdb4b300bb14db10829847caa8ee3555edc227e7ecad35b3932a38f774006861219aa2c49d53856242868f06b7389417e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h865bcd7d26599ed562fc3539cdb5b0beac6d6869048dfe2863ff3d9aa2b314b5606432f8b756331cca80bb8cb8c7f79d7791c3dfc684354e61d20fd04a621b864346abce00ffdde8aa1f6345efbed2f8db104a5fb8712d5aab6d8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de223702e42308cc7f30477a7875fb27ad4519a1e22667b69bbd07d43eb83df1d88312efa56b9d61b93f55209aed733a2fa18a6d3dc1c5d27593a882bd1baf87c9ddda39b989ac3bfc2ce40736e6bfe290f54e15ae88923d718168;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ba6e6c4ce63a335c6b729a9b4607385063bc0ed6207d0f8222cf70c9e315b18e18c5fe2dfb4c4616bf2bf6ec43ce436765541e40f0f7b46354390ed0aef3e2096900ec4190342367acd00d6b09bad63d908bea8f45619f0c4aa2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he269436af7a248c74b516a93042e72e190fd7bc60d30b282dc300195c3e3307927a2d1e62749a18eb405c8038a91c454cbdadf97b7920fe5531cb75b3b9b572d94401768a22ca0acf92e6a37d3032d50336745c0309063fa4aa495;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb983350815f52988398a8e2d6d6fab5afc228c466d6f57251f0e19c0f9704c1ada2cf8d208961ccbd350852fd1e443a001c9f1f6819972e813059f67506b0e65bcb5daba15a7a92494985d56f4575cbcc20b385fb40ec692120c6d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13cdb8376d98117c8027c7baf69015092a02ed7d7d8122ba2310056e9066503317a4a7791da89e6465a6bb804c10716e4c70929c7229f29e6b57d8804c09f69824a1f7284fe4d3135845999944f6661af734f6a5be8f99663fc9e9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80716afd2305eaf09d3851c83c152d83d5dd7597a0a37dfe69f2ba5cc84ba0ca97eac97754f7f7722b742fa416e910e0b353b7e658588e8b83e413b6408ce6ef6e7efe43f7d9cfea486cebecbc1a788654983cbf013294296572be;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1caa513d93c549ee624f95e77768fa6c2294bf34f3048206b26bd2831e227314f1bfcb349cf735983d2250434c483e31ea1910bf9ed4ae3f8482c7f50d00c1352253e6fb737491cea5d1f01f7225623012ffe061227e93c4d4ad277;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85b2531be99e4abea2569deb36eebeb2462f35bc085157b8f1f0e40c5a65b669c610636dc2a8b4921357aadc187ebce1c40d730135efbe4467a8d6fa3e06b9bd81b9a1e175bd85401fda3d8156b7a6e99ac9f72a4e31ac4c1f6b03;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15cbeee67b484524f9c2a944038e523128fea065142e7a407761270a835ddaa6dcef57acfadd3a6e0d85a27676402f5ddcdccd728e07e60bf387bd3123a3ff74c18e81c19de9d8ce412e72807c44d5c1d380adeecb7171f25e26d15;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15241b719c783767d625651629d358a5f371e3a5675d896b57f3044bfd2b3ba38313ccf3ea7eebbe054ac1883e35858de43f8608bf8363dcdd68b7dde8b42ec6289bb6b81fed617021ef082c803d1fb3fd49aa264a949b0940990e4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd35ac47b0bca59439ceb883975edf749a7c8d8570b32d720dfc6b735dc1c91d45b93d41c68e3f5342105e7ac9070d52346a3f51000d5e57b7cabc15238c77ee01631550c56f75ba5856f206f262e69a667a79f802a7b68bbd7816;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197dbff0d032b26f4c7992b577542b753224843c1849ea82bc49a8873c8d578e8f2c1db220f942259a5fa9353a63dd7a2279606133c706938541fc0796b89610ec4b0c7796b75939541088d1125dead0f191b2e0def5abb398625b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6773efeefee7cba5ceacc5d03cfb5558271697786fb84f95ac9aa935b50cfc5925b01c2654f7568a4fca4ee7480306c6c359f5ca42212cb421e6be0e24391d6d806370e25120cc66927905dfcc004c1248baedfc9fc6656675d84;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93ae7580a634be5b937dbcb198f7e01f4cd01464917ba08588d651665513d53622b5ad6777af45b29f14c3b530aafab2ea1f7ba0b397084c1b987c2cbfc2e6988fc5ab470d3bcb0eb8960c243c98bc92ea78a82e11261e1d3645c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca503e58212c96ef9123e9a5eb559f28c2fe1aff8bf009f25e0dc09892cb582f684553f974c4ba730d947029a7cf52546bfee15bb89640726a100cff29053ec61779f201e83174ba035af5363bbd3422b7a929804de666f464b274;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95079194ca7f147ec343fa3b4a37b011bb079771fcc59c3ac6da7f70376a895508801056f45e30f1c7d5037cc4c7f417b071fddf168c866c0ec581eb761f86d09a1dde3bec81efc34edbaa198c6576639ea5483dde3929c2096373;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e9386d483a26939191b188e5dd00884ce392dcaee99306927f2dd680844082f790eba217961dc45f54b3ddbec1f82f6b6cc10052dc6017f584f7cba4330ba26bb843541a49067970c519643b72a2b625e5df6f17c30101aa003cc1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1146f625d485f129b06063a9af793bb1e3831d3235f6f55d51d513a60e0ca71ba7657d2aa2616eb69aa1078f5f1ce19f6c943102dffd04e162c10f799c1584821989763f6a96bd59323c33f33ca45492129a6ccd732ccac53deee3c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17be30ee5028ac8617e56cebd3e75b0ab95d32f0e0b01c78f9746adaa320e510cfa89d6f876ffd6d7ecb12b0b484b4884a492ef1d617b7f94bc34f76c2d2b7ace3b792ddf5c2a171c21f7337643671b7dfafcf70b2287c1c1f12dd0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7cd68cf0940db5fef2674cf2effea5880cece04fb91b4cef3fd94c01d7124c7bc53d9fa5fda0da304de03d59f04c96a11c1bc945355a58a2f92ef688437c6bc574ef6da5765e96489f3edef01b2fcb66dc2e3967b8309387c4e7af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115055bcb96c9c2c3e32acb49e266cf6b443291aa5fef2ba414f617fb3b61f4800368be654c6fb63d880b9995283687f5dac3554ce4177b702cbe46b9ad4cbfac9ff494e02fc578b5564e0cf4519a53d7489279986f44406c2bd2e1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7170027b09be28a2fc88b4f34366541d10d09dd3f2e45f18372d08fcacd8d0c50499bdf5188249b2c8458ae084d14140614e7d7758c1184cea9622dd65a5f7f46c43e76f9f0a38c9bd5c8616e469cd6ad1ee84e82aad9deb591bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33d4837b36f98f6af2fd1ddaea28177595cd233624162c7bb835599ced6541b1f3ae1fc44c1f050f51bca4f117b31cc4763b58922ad60f09404cde79bd03b66ea6b41131eaa58e62dfd656177dc01cfa112cef8d571630aed05042;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h108d9ca8a1ec86c7b41483f2adafd0a37b4383818449563810993c9ccfaa5c19e1d3a3c0469c14a94760ead3f8e016dd497941e5852d07bb1c0c87f5f4d875f99aadba62f7016b02ffe7e83eaff0c853cdb83b9f0445399095c8ce8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184587ae095791daf4d8a48a146af15f85301672129a42b92fd8e3e3a10d546817ddb14dc81f76781595c5aacab927db0b96ac0a6ceb927962b34130cac6489fec6d326973babc1275059af3ec6b30890468ca4d3cb0baf4047a382;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h691b322d162965bdcd18abd6a55958bf193dfeaff88565190c71ff23922508c9be7285377d1df32a1ac8599ab2915475c8528702056b7ffb1110a8d9dd0559241546c08aa3c4f031f04d6bf3db40ecbae8fd1a3b4f4c3dbbf89f2b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4aee5c119447f5de30f3e8ef26d71dd77031412a8594116380fdbd11cbe7e445057150f79812946813de059fea7d0002410146ee249c900f1718545066e2df0ff54826fc6f46a99a9b1504890b3f62d4dff24b4894cfc2ece8afb3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heca8303145cb43b8bfb8a4ba602ee3dd6f63bddf15455c2d4f1c7afe274f10ae3c8a8ada4c76feb699c14511f9e0bf4f80ad1b4b9aa38dadc8bae81875f57e5c700ec0b0ff4c37c21860bc66704db5a4c616e0b16e7e30a086fc1b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c14c710c33878c8470a538fe9d50209e7e7e78c5bd892d5ae57a0bec1af2041cdef112cbdfe2d42e58de6b74a5fd23c03f2f23c509e2204c9eea46160c42209fe3c0e4443ed6cfcf565bf899eccb7e33ca1ed2708470bbd80e41b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc6d3d80e2ebf5ddd3fa62c31e8d0dccf0d3b860f72c4450e2569afd1bffadb814146663854690b0386e55013ddbc64b2a78f66daf0bc298d38a069f637dd3982a2d708b8abd0e6a0c763cbb41471951752c0ade339dc03931d1fe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3526a932078a9c2581b7b8c1c62efb6e61ee797f059d8febc0b9549199724fc50099ada18baef2cec1d4d72554c6b6d6d55e952e9b52e634cbb99e0306174064a5903762453c45e0c5ad32a46f11a2bd93fda1939e529147cbf8ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a7c474b89fec39a2b18fb2507e4347a070bfde930374d46fd359eb66b5d5c869db844a4508ffee21ad85e49900305353117ea995397a43243ad4f23c6ea4e2e1de77c2b967ef2ec9898b88e8f6ee64f6aa39cb73e6c7b66ca9bd2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h175f9605da031a941082a02f91bf435f90a201d9ef0263924b2c5a2465360cb3b1395ae2e7d091265bb0136cbbb9f424f6bbd1dedef7a54135ee71bcb162240bd5eb229f3ef71174cb335f48146805ad41d915250f802a86d5c1d90;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a7624fd082c71bd806b039397d91b3d26cb344be6fc2f6bd200630a3be4b16bec8069b97dec5cc0d457ccdf12f6a5b90179ccf02fb954f17922ba4e28094a09d75ebcbc9e400b5849f23a0201797791bad0c97aaf60316d28a3765;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11624ad66b6dbefeccda012aab5fbea3cc649ae2366ad3b4517557eb699dfa95071a3dd07d7f0bb39242f897d905d058dd9ae8989576febcff8d3abcad7a43a845ace8f52a2dff2d1ac0adc2b18e24e51121e9aa1124745aff00ab2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec0353f9f06e01c2209d278ecd9679884a4b68a898ff8fea8028fae22cac3ec699cca2db35c513af575d48dbd384edd58203f55d29201f26715058d31fd7da9a5726ed0c89b9a73bf515bfc7ec4d3a9b9e7082e4c46d315e2597cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfced1173c0fe715b73b478f9826f48e3f068ab452b7aba688d835cb4d875c47339949115784ca4fb285fbc4ec84c613688fd54e60cff2860b9a8f085d6081efeeed46909daac5dfc7bc245fde72f9a3229e58fdc254b7b6f6c6417;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2c5ff448b370c81069fde916610e7f2057453052c916e9ad4d8c07662248a7a021ee89c4b5f4ca070a48f924165ea11e33701ae1c4c50634c33ed61df94b2ef531ea1a237cd3f810e7f1f561fa9563408a429bbd314db14dceac9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167908a79fee134c167b39a0f6de8b7f6fa4ccb89a23a8786becf03e28197f487a4b156017c34a32d37f12ab73d1478f748fa6440b17e6bf5f74ee43ff8c0bee5e7a498b006098ad6b53d6c8497af9bbd11c52237fa19e2a97b4832;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b4176f96bd01a67ea2c0dccd89222ded4c474f34a1bf322509acbf5b42798d6478b12511871a3a9f1149debe1ccd816cccbb270128a44ea0fe4a4420d588331035992c3b3813ccbb27b735cbbb5f7c09f358ba4a43f601bbeeea8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h581da7324c9d5b826dd26ea116f2a97579e5904ba2a68a359a0b8b0028475ec221b01ba4f908d3fa86e02178a83b779660b8fc80ca0296ac91e12cd6044580523a85863a7fc6ccfb9f59bff31eee154eba285466a31f86cd90155e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haadc9f95d0321e0c27510ba4897f41870493cedd1405bca7ae8d3084e59210bccc0cd304367df1018f14ed00d27ed62753f71e46bfc50c965656bc7b96aa8aca932f3c41140e0a2c7e8ed7dcfcd45c180d14bac5030e00badf7c27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heaf8b01c41479f9a32cab39cb6502eddcf84dab1873dc24c7d425ea96d5a570819ec57cef3168f2d35090c3a3b06b6ee85e432820dd76fe34b266cb9f27da4ed79289654414e80e5da91c30c2012850a3ede97c76dae861295e8e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97f60eefef1c5fa6499f4161e4a49521bdb175e73e9d27ab0a6851cfb7f9228aab1cbbdd6a0e86c1508a901661ace23105defa4cad862b570a64d9647f231107d08911770047d4c654b9b60e28b43931247496c7dc2cfa7ea98256;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f729ac0dac3e51743ef07a03e84e7eed14a6d367cb2f847cd4f243016595dcfa65756b1863e328836e64af1483b8bd76e80301b4f6045e5e1086a1798fc2d33f35e7ee1c41254109c8614a0514479b0e729a8a3f37ef2aa4121437;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd39f8acc045e3259d44584467063d4d66b1e9ad6ab0860d75fa9086a717dce5338066f89c73de47046aa58b3d90757591aa011c99497eb7f1c9927822480820bae91b33fab1ec684b7b8655ae5ab1925c1e3a255dea4d23bbcf4e4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c56d640a7bf89d8416ebf38380938f3e358ea43023ca7910b365f7261625e283afd4a117422691de57a67d75576e110636bd09f6358402bc78bef4a9135c4839be41dee332f97e3a506d7b1ab16d67d17dfdb733c5b0bd74d0006;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2c1093adc999d9c5c52470f3300d5439106d7852ff7b02949437d6ff1c631b9e00559437d52404d7a54abe182440fe6a83242adfafb2596b3c097736104b30222ad89d9024ac0725d505940648040c9bf3123b97baf6ebd3cd233;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18de58bcfd827cffda60c1c0f0aa4355fff477c6a9e45f8540375d3952c2c629be15e45e72251335721adff4677ec592dd5f1365285439e2fb998624a9fabb8d2f63737a2b02b8106e3b9834bd8c2e73a9c986c717b54710979e906;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h109f70b6bd854dfc5541b0ca56f7b9301ca0dbfaed430366a902c57726df12b006991101af9ec3a8e0bab0d86c7b8156b9ee38dcae7f22b3d938754635e02392fe730b953e735a9c7452a1afb2a037dcd2cbf606bd7263f60fb1b46;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58b6ac735b01c5a04497e07cb74ec191ea6fe19820e7032935b8a4e56d76b8bf972c28113cb06608ed6a7252bd53bd0b6c413fea7de3df9808b2d40e67e3136b0203a62469b61f8fecb2fdfcd9c85b7799d2a196d9a450cd003ebe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90e260d9ad7798dfd936638e28ef1648fac171822bbd56d9d1eec3ff56307592d08fe3525c20d381bacca15e9bbbc23290ec435066184e5daf5f7fbfb13985a2d2e36ad01e703560f801c1a146028731075db9bd7abb6f6fbd682e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f5e7b1436d8b41a1029c3fcd6b6471ebdf8e4bffe536f00b2bf5461b332f9f4d4c2e6536ef8dfb337fda221af7be2dacd9211ab7bee112f6d3369cff9e330f1851b9b7eb5bdaf29cf4ecfc5561c4cf9028330bb230b9a7f6b68a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d43e0b1293edff77691761c240082348b41c22c5a774b6b8564d6b163d49f3955f3548b3d5fe81233f1654d33574221fcf5f4559bc63514ac2e7f0c293cf479bde9664e36523f5593cce2de26eb1860d3c1fff12e65d9274b7de75;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h501a38ef039efcde4204385ea78c7db297a4386de838e6dbd002014155193cf555c54e1be35316a6ccfdcaf56b9faaacb6ea6b84e75021e97974f9efc65f71d2aad052e18ab2063487a3b38f3924e5b9b3fd20852d6fb6a8c13d82;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9ff60ff5d4711fc5f3d7e3adbd9c5a8c322b4bf16b4489e311cb4847e2fac807545108184c42a4d99e47aa0ee5ba07d5aa40609ae3c5a133877a60047c79cf240cee636858ce07f74802f947304b51d2cab5343b909cdb5fe2656;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18504cbf02e2c9dabdef28d71188c29b7f9c8830433d1142122e08d828774bffd0115f16c0d79aa1f2070ded794aff5e866f9f44313c3f39589ea09a8bf9cf3a20ef622318c6e7aaaac0442abc6045d06c25e8707fd135f47eb122e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147271345b722460421b745a6adbcc2ffbb11f67824e539702de2e10cce6428dc731b1eb0d2fe085cbab4c2a8275f859c77734f5c4cb3c6a6f4998927374f17b783bea858d5e8cd786ea04318e8103003fc1eda6f0d4b32b6d3cb3a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d55eb910dee7781b01b3ab9dfd01ccf98f58b420c10d8f24dd6bf737d017ef0b61c22e7aa2eaae00db30845b5960de546b52e636c67a0bbc35b1f4e34bdaf24698f9a605eac1ad3838080f16fb896f263fdf672181f407a280fe9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4913344e53ef5669ee408d28972a8607e2cd2a67f632a80c8b80d9ba299c22dc8bcbd60708ea8108ebabdb56218f175d0b4c3248cb902e9bd63b288bcf87065273d83a7592ff3de1e13b7df3bc36f32026a0db29ad5d936bf224f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e4591d362f98d03dfda6ce7c0bdbca5487aaf217b54fc0110db0736d96ee30bab7314d2684165bf6422f7964bf9a7342a1dda31d03930611eb70d2166166198c9b0d6e148889cb699e3202a0211450b52f1cca0b7bf7f83a322d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6149497a9c687c835ad1ef468d86b2dadd59c33a2cf2a215b5c28b8b4ec56df5f59be82690665c741ad070be9cf948196757ad52dc2491f6d1497912fb91ea71a8f8282d43a5e7f1454e2dc7a27a7fe68dd007e488ddd980c86d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123a12d2f80d9baf5cf882cc5297e4e63c2f81f88cf1b8021644582ddc0b20247a580fc0706c9791bab921c87265849d242a3ddb0081a1dbac3eea8af4215819331af745bae018a27424b21aea9a6ae0d2bc97afc57e49d5d00c1c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haeaa23b36f2bd5c50d60dc1c79f097960a48df42f7900ea13bac7d3988fe8a81c2a248bbbbc5b0c0a38d667903f90b94f773d8080a7b2500609e914b9accbdd49c8e7662ae7da37cef0f23947032eeb6596147525f00b8658e91e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd14b0d294fb94e11e38985943230f5ff65df06fb0f72b9feb040903abb19615e088efce2a7f2c136350da7bc37325feed0ffe46487ea9eaee04cc2a95991efea636966bc6696c90e96838662f6111ca3ba3827e3e65e20cc5640d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he2d45b18de71870fb5b25084252155aeebd4cbdce708eec793c1bf4319a73cc78b00dc41cdb0c507c0466d6fedd64e51ddb122e8d41abba5b8c87c0e4f1fe5807bcd87f14ead5ce88c83ff0d18f1ff47058754600cbc888a5bc4fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd876d1c077317c8245e8f000ae8bcdaea5c15729a9934d9ef3f00f664d8dcb64234af38f83cd32a41146c1bf0fa7ccdfc5df75049eef54c788c96c065b7dd5db62a18358c3415b656aae9a13cd53b5083547995b360fd26b7893e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff903e793752d6978085eabd9aaa5efc3bf54781654262e86c17d01dc7742bfb577aa14622c2339864486d07d127dd833e5320c557adfdbc1c9aca53bf9811eb630de4212ebe3e89acf333388840ec572ab5fc6857bab31432093e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd80c2e4eb802620b768d42ed861c97d852780e898b14f760519ea506d6a69d90260496412e56f7ff652d40f4ec14d1414e965a815cc9b642e8844398fb083efc4fb810f5460c941e68bd1e5ffe49df55e4d69a2cac3a5e300d9ab0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e9856d8651bf74692ce1e401ef96551bc8b848e6f8a192a4efccda03a029c60e7ee3a46cc14920f4bc2c6c63274da47a3f5f5a5fa835bc4f1e56bffc4226013b4117750b99ac12e5831aa5ea286783a2414fba25ea2bb4232107a7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h249b5e8547a4638481fd5a2aeabcbf3f9c4d36561db0e7c9fa0fa245b6185c7124c0a60f9d6184bd5bad9f77a80762f83cfc0ed353bd82a8a1fd4c55cf291cdd8e0262b5b0b59f29c244e4c42ebbf6e11abb12cdb27e7bec757cd3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f54ea7cf2a82625033e048224734606d5504fe8e95edaa335bdc3daed4e842d9c264b1c713cc467f983856b29c055ebd03b239b594bbe01acd43036cb17ba59504c3fac29172c8535457692dc8ca21bfdc99da0f3448e599fc6d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1937bc16465346317366848fd8dfd7f6d57686fb1d72b5efd3c4284e09c2dcb2764e4e78dde1af1484f2f3d43c88b6c8c0668525d45be22e1c053b8894eb1ef8c9d869517e640553e83746d9e12d860568b95c78c17971ca37fb05c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he3182ce547795e802be27e3fb8fe66ca459495a62401df2df0bbcf67794b8f943925c7f037da198d67d0f705813136ee633f3ca0ba10d9479b1f53456dc51b327af15fb89348e4e512c9f98056bb6bd655c7c7c4aebbe1805aee5f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h163af3e9a69a35e64ca3bce5f23c5ef4d42d437737a1b6a7edbab3cbce939fe8b3139723042840c5a268113536aa926cd7078a275102ec791c5be494a56539d70cdc7693c317024c3e5da1f18b4a6ecbfd11c417c7963c8fed04278;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4830af18f91480bf9ff1ad2e8a145299de6aa41372092b997c0c81dcdf1950d67b9c789de9b5655380686a3b02351c88b51778c14cc67daa1ca1946eff6d7ee2af1ad41f607ced3f611bd087f4337e301fd346d2ce69d84ea1fd0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb8629516b4f2cf39075684fc98b76ef7494b7c17b82a4ef9b6b2264234721d9172d6da9635cfcf482ec7dda6995a2c34efcb9c0ff2f59f5a58ea998198e16507fdff6795552c3b67fbe11b1c4726c3cc918c3e9c2e75c073dbe94;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3e39ca7e4dee965953885176981443d0d6d123e9a2656497bd5bc8786f6a0d9df2911191257e29874c09fe47c23e111c88b37b8f72959d4cfbe40a0d992714e5127b5030c895031659f66f5a8007297cbc4480181059e837ed4e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1df7c146e62f60e3250e57ad2a86a1aeed4ffbaaa2ae0384b59a173425096d50a5735dbc9c41424358db18a35fd3f75d49b0c0cd06bc80504b28ce468900044b22a8ee09e4e3164950c0e4f9e339eae1502a60dcd3ad2f40b9d643b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1196b33fcf424bc4af1fd27dab64cd2f461a4df712a3129062a8f471c6308e3c09c90086af8879650f18d320de2be6884aff02af92205e4afdf67303c1ba69518ec1254ce996b45b4d5df36b6562d8a40027bd2aca3b9c8ff11863d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d00df9347e1a22067d71d10b18bafd0334b90b48babde7da5842fc95fb26aa8e1a4a0d8b0b5c689933cd20dd3c48797c419957be0af0e07e60e61c634eca514255f3a9947dc4a8f8c0d4a18ac0dcf17971aace6676e4710d80ca6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8eaf54a3549d1cff33184ace4c028673c05231409685ef71ec3b8f7fd28a654b22582a3518634b76ce799d3727b9b2dc312d5036f263716b6f313a72ecd4f90e6c15b7fdc965efe42a49f88e25cce16e0f893c83d16c3c9a9b6d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b0fb16e6ce231050be9b899f056a9240db608f9ba3e893cad80cd0b3d344f030b9f5c63b149a0d673fa4f213193d808d23da1c1d54c971c52bdb8a39ffebadc35ae1888c26001533301e045b4323a727ecec6a1573a0abb34dee0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f2a8043ca6c355002e6771688584af312aeaba7544865df7335b1223fb4c143bb7774bcd49a2fd6fa465521c63b9450df4cde00a501414976e5c50648d2c2d60b093f41a4d365ec770f21a326aa442585e1e1326fb15775cefcf3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f74f974ebb99eb74dd19521b9da41825a7055ed391b9b3da19e4e53632760ef5e7e837b1dfa602b447b41507ac22ab878a4450db249ffd544ecbc5ceaeecc82057e52dad7ab3f6a9efb4ff236dae499e3ec9530b3cd152c918659;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9aad16a567c1fb2de387a9b4923792be84604ac0d3a696cba3255dc3ff335d404560122dfad2fe82858cf5b2250951cc97274bc7fd1a83184f13a0cc148f44162869071f6f051e64572465e33e5e362a281335d8165ece4ecef67c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h555060c1308e00c0d6ade59a1976f4cff286aeb1f5458099d2c68e668f1ea2c817c1d9289a66ba16437843733f9da964408b39868db6173953742ba7148b871af9680b1f3c5521287c66cba0b2e520faa82ea19fd2e34f3f8654ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1716a4a4cf883d4e7aa84e44617516f3ba1cd14dc29b6e9d84c08e47b7c25ebce3bd3bd742e72b6ccd0b6d3035abf27818e29a43d7b6ad76aecd7a2214a1e2a3c977a167a637286be8308ea9d1fea5299f8439266347eb75e206862;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167f9b0db288cc3723bd4ce2660f2bfdc6ef2a555553bb69b67ba3b3a50ca0011c49af3a42cd2956e780827d04c15b87740499f883796649079dbaca0b69fd272664b1bd787de386a27a1d27eea30953ce78c56f341617ec204e62;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha68bcb8de71abcb40db649aa4901f1abd5aa75f945ee65698ab3b4fa6782950b0fbc2db9a3103d3e629e072e39f348c906a803c6925f7a739ad79938115a06823576a191ac1352b25fa327a1c3eeb1fff8846d07af31e4c2c8d9d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1543e2c4038fb212161d57e108cfa5bf0d6e467688f4d136820c907b82bfe71d42ef11c4d63fe1184e616585ff08a3c006335c4262445e03aa065f20aed79b9dbf6fa9e3b1936e28daf6555f7085d55926dadc8b66da8facb89a784;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14177433380a4b6fd8ec49097df9de0ce71d37f5f184c7d7abc2b8562cc285cb4032baa1f19ab28cdcbc0f0a0d784087f7cb8677167ae47c11e8613c2191f0bbdde857b877ab51f1dd6e14640d66ef4e6e56e94acb87e975628ac78;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152db6dd6e783c6f64f8cb6259247ec3c8cb1d1f61443dd59ee82d1de144a1e62198db582d934aabfb6ae3b4e223af5970a579df38f8eafffe90512f263e7e5e8df9c679884b402d5d6e8f933ec353b0dd8237302cb0326e30360fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf83f125a406d4221f5aea7a53faf8f61de7b62655ed3e92a214b3683e7c256019d1a4161a458e074be46b380c6367c5e876dd710a2315b703f783282b13d9a995db4b45c90ba7787eca436a77ca90552595f847660dc1128d95bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d58c670860e1ffa8b0f85b91fc7e8adaf4be52752a7ac42c9249ca12ba3682d68925db8696f04f3e2ec3dcbb3e89cc813402b6511d0c38714f1a606e9adfb087326e6e6d720dcdc677aedbf42dea082fedb49cf6f18844cde03132;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h256188d4ef49333d5b5bec33228a613d169d49f28391a72160b901f9f84515443ff83aadcfd70fa052a4e62f67687b8c51bbe419987cbefde9c710e761264e1372075316071bdf696b648c07db38017c9a26fe4f65622c24acd31;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e45029a1fa0be388ad8833f79be8e7cdd6329891dca6d233c3cc29c2a81e08e16e0cc95abc070c47f8c4f534aa4bac368386bb9bf7f8936ccbcc0355354e4dd80d871ebf6b0daa9b68bc0f1fba346eed05faaec1c8f3961923464;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14bfa1efc573c7e3678c881c8ccc414a91caa67e7045dee411c89976d534a5897be986c9c244deffeb811d10a45bb5a09072a58d134dce01b73a8c972acef187ea1ca7d4ace484a6ab8917e1217b63d645786a55f6dc7bb3c54442c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e499dec5dd59b893d4508807491610f531c438c215c724aed3ab9147cdeb682840776258757c371f3c0e67973912fa0a8943b8b49429d8fa3df9167fbb71b3e87478bba20628378fe24314943a708f8d0b13df8675aaddb8e93788;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h674cddb379723775633410115719712a65570d4a81aedea2aed81194355444a5c5fdd68915c861ff7c57799c9e64e67ebb6f5bcfdbf4863513038d05d92ed5590dcdaa0a57b5845d018e3a8b44d19cd256a61b442927b5b5b21c0f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9fe3156a3e6ab1603821250794f3ab951cc0247ae9ef6f6c2d7fa7866385c9136e21d8a840efa4941ae0cd37f4e21c29e7c385e3f96d5f1aa7588a3624ff7249ef04c324dde92c4aae8ebbadb6a211d75451d46e41507c19fbb95;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113c413421c33435d988e9fad6cafefa21ee62be8bb113f2d94a491d1379676c8722eac948749c8c24434c6a46af7d28dd486826ed4d1c3f330af4e331bbf08ef3d9cd33ef34c293c31bfd5adfe8896912a58905850797da7f2b36b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c344be44e4d6f0f8e00c8e91737f02e3f35c092e1e8f74dd7a021644cae496f074797e8e19bce2fff1921a04433ecc99cc8b197f0704d9e7fd1a057833dd7eb962954b3d6dd802b9387145fb382522e9191438dd3adb679da85dd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h112f3d6539849d7b0be62b33a09b47bcb96cdd371a9b451ef2b9a3af6523aa380efd9fab22e68287c198624e5b2ac81824d9f2d3e7b12d0499cf89362932e45d459c4b228b9e51f6021f13f727114c5f27d3fd0872aaaae0850e551;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4a10b52d3e40ff2f3ddf9d723515db7eeddb4b42d9e38b28a066352f0fb48cef1f742880cba41f015293f0db31941ac5609bb9fcb7cac2a8b874976610a0da83c2e11ee0f1392b6b45ae6f8e91008a7fbfbbc57732a5516c3ca67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h385db4a65c8bd7762dbbd8319cadc815027491900869055a02eca839c92f29329ebef71ed78656849dbcc016bb10d833ad2e28a3fc2f67e12eb285b87e048169db8fd9c1e18cdaa0605900585dd797a0b94bc2a5c79f5c7581a2de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9db5a90518398b98d38a1a903f3ec43db73089085de3cfd1e6fd90e3609da92b3042d528adc2259485fbb079812f87f17f08c15110c8d17ee6983575e8165c1d8cc0a20acf51eefe66383a7181090e713887289d94c2b0a1b90519;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha0834dd64f1d0233ef5bc7dbe6ac04c24bb8e07f0c4b2e9ba2eed5ccdbc187f8a279b9baccac382e4c41984095d71f65979d6b0e8e7f63e5452ead85560c5c072c818ce1aa94d1314ddd2097444b2bf86812d44305b53cc369c10c;
        #1
        $finish();
    end
endmodule
