module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    compressor_CLA256_32 compressor_CLA256_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
        src12 <= 256'h0;
        src13 <= 256'h0;
        src14 <= 256'h0;
        src15 <= 256'h0;
        src16 <= 256'h0;
        src17 <= 256'h0;
        src18 <= 256'h0;
        src19 <= 256'h0;
        src20 <= 256'h0;
        src21 <= 256'h0;
        src22 <= 256'h0;
        src23 <= 256'h0;
        src24 <= 256'h0;
        src25 <= 256'h0;
        src26 <= 256'h0;
        src27 <= 256'h0;
        src28 <= 256'h0;
        src29 <= 256'h0;
        src30 <= 256'h0;
        src31 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA256_32(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    input [255:0]src12,
    input [255:0]src13,
    input [255:0]src14,
    input [255:0]src15,
    input [255:0]src16,
    input [255:0]src17,
    input [255:0]src18,
    input [255:0]src19,
    input [255:0]src20,
    input [255:0]src21,
    input [255:0]src22,
    input [255:0]src23,
    input [255:0]src24,
    input [255:0]src25,
    input [255:0]src26,
    input [255:0]src27,
    input [255:0]src28,
    input [255:0]src29,
    input [255:0]src30,
    input [255:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [0:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [0:0] comp_out38;
    wire [0:0] comp_out39;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], 1'h0, comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], 1'h0, comp_out2[1], comp_out1[1], 1'h0}),
        .dst({dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      input wire [255:0] src12,
      input wire [255:0] src13,
      input wire [255:0] src14,
      input wire [255:0] src15,
      input wire [255:0] src16,
      input wire [255:0] src17,
      input wire [255:0] src18,
      input wire [255:0] src19,
      input wire [255:0] src20,
      input wire [255:0] src21,
      input wire [255:0] src22,
      input wire [255:0] src23,
      input wire [255:0] src24,
      input wire [255:0] src25,
      input wire [255:0] src26,
      input wire [255:0] src27,
      input wire [255:0] src28,
      input wire [255:0] src29,
      input wire [255:0] src30,
      input wire [255:0] src31,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [0:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [0:0] dst38,
      output wire [0:0] dst39);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [255:0] stage0_12;
   wire [255:0] stage0_13;
   wire [255:0] stage0_14;
   wire [255:0] stage0_15;
   wire [255:0] stage0_16;
   wire [255:0] stage0_17;
   wire [255:0] stage0_18;
   wire [255:0] stage0_19;
   wire [255:0] stage0_20;
   wire [255:0] stage0_21;
   wire [255:0] stage0_22;
   wire [255:0] stage0_23;
   wire [255:0] stage0_24;
   wire [255:0] stage0_25;
   wire [255:0] stage0_26;
   wire [255:0] stage0_27;
   wire [255:0] stage0_28;
   wire [255:0] stage0_29;
   wire [255:0] stage0_30;
   wire [255:0] stage0_31;
   wire [49:0] stage1_0;
   wire [97:0] stage1_1;
   wire [91:0] stage1_2;
   wire [90:0] stage1_3;
   wire [148:0] stage1_4;
   wire [125:0] stage1_5;
   wire [95:0] stage1_6;
   wire [100:0] stage1_7;
   wire [119:0] stage1_8;
   wire [131:0] stage1_9;
   wire [96:0] stage1_10;
   wire [139:0] stage1_11;
   wire [197:0] stage1_12;
   wire [92:0] stage1_13;
   wire [113:0] stage1_14;
   wire [92:0] stage1_15;
   wire [95:0] stage1_16;
   wire [126:0] stage1_17;
   wire [150:0] stage1_18;
   wire [93:0] stage1_19;
   wire [115:0] stage1_20;
   wire [138:0] stage1_21;
   wire [93:0] stage1_22;
   wire [93:0] stage1_23;
   wire [253:0] stage1_24;
   wire [117:0] stage1_25;
   wire [236:0] stage1_26;
   wire [107:0] stage1_27;
   wire [101:0] stage1_28;
   wire [117:0] stage1_29;
   wire [96:0] stage1_30;
   wire [132:0] stage1_31;
   wire [73:0] stage1_32;
   wire [33:0] stage1_33;
   wire [23:0] stage2_0;
   wire [32:0] stage2_1;
   wire [34:0] stage2_2;
   wire [42:0] stage2_3;
   wire [73:0] stage2_4;
   wire [41:0] stage2_5;
   wire [52:0] stage2_6;
   wire [53:0] stage2_7;
   wire [55:0] stage2_8;
   wire [65:0] stage2_9;
   wire [48:0] stage2_10;
   wire [57:0] stage2_11;
   wire [74:0] stage2_12;
   wire [56:0] stage2_13;
   wire [89:0] stage2_14;
   wire [46:0] stage2_15;
   wire [40:0] stage2_16;
   wire [54:0] stage2_17;
   wire [90:0] stage2_18;
   wire [45:0] stage2_19;
   wire [125:0] stage2_20;
   wire [71:0] stage2_21;
   wire [46:0] stage2_22;
   wire [56:0] stage2_23;
   wire [63:0] stage2_24;
   wire [65:0] stage2_25;
   wire [67:0] stage2_26;
   wire [95:0] stage2_27;
   wire [71:0] stage2_28;
   wire [39:0] stage2_29;
   wire [44:0] stage2_30;
   wire [47:0] stage2_31;
   wire [43:0] stage2_32;
   wire [30:0] stage2_33;
   wire [16:0] stage2_34;
   wire [5:0] stage2_35;
   wire [5:0] stage3_0;
   wire [27:0] stage3_1;
   wire [24:0] stage3_2;
   wire [34:0] stage3_3;
   wire [35:0] stage3_4;
   wire [15:0] stage3_5;
   wire [19:0] stage3_6;
   wire [23:0] stage3_7;
   wire [26:0] stage3_8;
   wire [21:0] stage3_9;
   wire [18:0] stage3_10;
   wire [25:0] stage3_11;
   wire [31:0] stage3_12;
   wire [36:0] stage3_13;
   wire [25:0] stage3_14;
   wire [32:0] stage3_15;
   wire [26:0] stage3_16;
   wire [19:0] stage3_17;
   wire [37:0] stage3_18;
   wire [34:0] stage3_19;
   wire [36:0] stage3_20;
   wire [32:0] stage3_21;
   wire [34:0] stage3_22;
   wire [20:0] stage3_23;
   wire [23:0] stage3_24;
   wire [35:0] stage3_25;
   wire [23:0] stage3_26;
   wire [38:0] stage3_27;
   wire [44:0] stage3_28;
   wire [27:0] stage3_29;
   wire [17:0] stage3_30;
   wire [36:0] stage3_31;
   wire [19:0] stage3_32;
   wire [17:0] stage3_33;
   wire [9:0] stage3_34;
   wire [12:0] stage3_35;
   wire [2:0] stage3_36;
   wire [5:0] stage4_0;
   wire [12:0] stage4_1;
   wire [7:0] stage4_2;
   wire [11:0] stage4_3;
   wire [15:0] stage4_4;
   wire [11:0] stage4_5;
   wire [14:0] stage4_6;
   wire [14:0] stage4_7;
   wire [7:0] stage4_8;
   wire [9:0] stage4_9;
   wire [14:0] stage4_10;
   wire [10:0] stage4_11;
   wire [11:0] stage4_12;
   wire [20:0] stage4_13;
   wire [11:0] stage4_14;
   wire [16:0] stage4_15;
   wire [18:0] stage4_16;
   wire [7:0] stage4_17;
   wire [13:0] stage4_18;
   wire [13:0] stage4_19;
   wire [18:0] stage4_20;
   wire [11:0] stage4_21;
   wire [24:0] stage4_22;
   wire [10:0] stage4_23;
   wire [7:0] stage4_24;
   wire [11:0] stage4_25;
   wire [15:0] stage4_26;
   wire [16:0] stage4_27;
   wire [19:0] stage4_28;
   wire [23:0] stage4_29;
   wire [9:0] stage4_30;
   wire [16:0] stage4_31;
   wire [9:0] stage4_32;
   wire [8:0] stage4_33;
   wire [5:0] stage4_34;
   wire [11:0] stage4_35;
   wire [5:0] stage4_36;
   wire [0:0] stage4_37;
   wire [0:0] stage5_0;
   wire [3:0] stage5_1;
   wire [4:0] stage5_2;
   wire [2:0] stage5_3;
   wire [8:0] stage5_4;
   wire [5:0] stage5_5;
   wire [6:0] stage5_6;
   wire [6:0] stage5_7;
   wire [6:0] stage5_8;
   wire [12:0] stage5_9;
   wire [5:0] stage5_10;
   wire [6:0] stage5_11;
   wire [3:0] stage5_12;
   wire [7:0] stage5_13;
   wire [6:0] stage5_14;
   wire [8:0] stage5_15;
   wire [5:0] stage5_16;
   wire [7:0] stage5_17;
   wire [5:0] stage5_18;
   wire [6:0] stage5_19;
   wire [9:0] stage5_20;
   wire [5:0] stage5_21;
   wire [7:0] stage5_22;
   wire [6:0] stage5_23;
   wire [5:0] stage5_24;
   wire [2:0] stage5_25;
   wire [5:0] stage5_26;
   wire [7:0] stage5_27;
   wire [5:0] stage5_28;
   wire [6:0] stage5_29;
   wire [12:0] stage5_30;
   wire [5:0] stage5_31;
   wire [5:0] stage5_32;
   wire [5:0] stage5_33;
   wire [3:0] stage5_34;
   wire [7:0] stage5_35;
   wire [7:0] stage5_36;
   wire [1:0] stage5_37;
   wire [0:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [0:0] stage6_3;
   wire [3:0] stage6_4;
   wire [2:0] stage6_5;
   wire [2:0] stage6_6;
   wire [2:0] stage6_7;
   wire [4:0] stage6_8;
   wire [3:0] stage6_9;
   wire [5:0] stage6_10;
   wire [2:0] stage6_11;
   wire [5:0] stage6_12;
   wire [2:0] stage6_13;
   wire [3:0] stage6_14;
   wire [3:0] stage6_15;
   wire [1:0] stage6_16;
   wire [2:0] stage6_17;
   wire [4:0] stage6_18;
   wire [1:0] stage6_19;
   wire [5:0] stage6_20;
   wire [2:0] stage6_21;
   wire [5:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [2:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [2:0] stage6_28;
   wire [3:0] stage6_29;
   wire [5:0] stage6_30;
   wire [2:0] stage6_31;
   wire [2:0] stage6_32;
   wire [2:0] stage6_33;
   wire [2:0] stage6_34;
   wire [2:0] stage6_35;
   wire [3:0] stage6_36;
   wire [3:0] stage6_37;
   wire [0:0] stage6_38;
   wire [0:0] stage7_0;
   wire [1:0] stage7_1;
   wire [1:0] stage7_2;
   wire [0:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage7_24;
   wire [0:0] stage7_25;
   wire [1:0] stage7_26;
   wire [1:0] stage7_27;
   wire [1:0] stage7_28;
   wire [1:0] stage7_29;
   wire [1:0] stage7_30;
   wire [1:0] stage7_31;
   wire [1:0] stage7_32;
   wire [1:0] stage7_33;
   wire [1:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [0:0] stage7_38;
   wire [0:0] stage7_39;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;
   assign dst25 = stage7_25;
   assign dst26 = stage7_26;
   assign dst27 = stage7_27;
   assign dst28 = stage7_28;
   assign dst29 = stage7_29;
   assign dst30 = stage7_30;
   assign dst31 = stage7_31;
   assign dst32 = stage7_32;
   assign dst33 = stage7_33;
   assign dst34 = stage7_34;
   assign dst35 = stage7_35;
   assign dst36 = stage7_36;
   assign dst37 = stage7_37;
   assign dst38 = stage7_38;
   assign dst39 = stage7_39;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc135_4 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc135_4 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1406_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[7]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[8]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[3],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[4],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[5],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[6],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage1_4[7],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage1_4[8],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[9],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[10],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[11],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[12],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[13],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[14],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[15],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[16],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[17],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[18],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[19],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[20],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[21],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[22],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[23],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[24],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[25],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[26],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[27],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[28],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[29],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[30],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[31],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[32],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[33],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[34],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[35],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[36],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[37],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[38],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[39],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[40],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[41],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[42],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[43],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[44],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[5],stage1_4[45],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[6],stage1_4[46],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[7],stage1_4[47],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[8],stage1_4[48],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[9],stage1_4[49],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[10],stage1_4[50],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[11],stage1_4[51],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[12],stage1_4[52],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[13],stage1_4[53],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[14],stage1_4[54],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[15],stage1_4[55],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[16],stage1_4[56],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[17],stage1_4[57],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134]},
      {stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage1_5[18],stage1_4[58],stage1_3[61],stage1_2[61],stage1_1[61]}
   );
   gpc606_5 gpc62 (
      {stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140]},
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122]},
      {stage1_5[19],stage1_4[59],stage1_3[62],stage1_2[62],stage1_1[62]}
   );
   gpc606_5 gpc63 (
      {stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146]},
      {stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage1_5[20],stage1_4[60],stage1_3[63],stage1_2[63],stage1_1[63]}
   );
   gpc606_5 gpc64 (
      {stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152]},
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage1_5[21],stage1_4[61],stage1_3[64],stage1_2[64],stage1_1[64]}
   );
   gpc606_5 gpc65 (
      {stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158]},
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140]},
      {stage1_5[22],stage1_4[62],stage1_3[65],stage1_2[65],stage1_1[65]}
   );
   gpc606_5 gpc66 (
      {stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163], stage0_1[164]},
      {stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146]},
      {stage1_5[23],stage1_4[63],stage1_3[66],stage1_2[66],stage1_1[66]}
   );
   gpc606_5 gpc67 (
      {stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169], stage0_1[170]},
      {stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152]},
      {stage1_5[24],stage1_4[64],stage1_3[67],stage1_2[67],stage1_1[67]}
   );
   gpc606_5 gpc68 (
      {stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175], stage0_1[176]},
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage1_5[25],stage1_4[65],stage1_3[68],stage1_2[68],stage1_1[68]}
   );
   gpc606_5 gpc69 (
      {stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182]},
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage1_5[26],stage1_4[66],stage1_3[69],stage1_2[69],stage1_1[69]}
   );
   gpc606_5 gpc70 (
      {stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187], stage0_1[188]},
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170]},
      {stage1_5[27],stage1_4[67],stage1_3[70],stage1_2[70],stage1_1[70]}
   );
   gpc606_5 gpc71 (
      {stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193], stage0_1[194]},
      {stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage1_5[28],stage1_4[68],stage1_3[71],stage1_2[71],stage1_1[71]}
   );
   gpc606_5 gpc72 (
      {stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199], stage0_1[200]},
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182]},
      {stage1_5[29],stage1_4[69],stage1_3[72],stage1_2[72],stage1_1[72]}
   );
   gpc606_5 gpc73 (
      {stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205], stage0_1[206]},
      {stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage1_5[30],stage1_4[70],stage1_3[73],stage1_2[73],stage1_1[73]}
   );
   gpc606_5 gpc74 (
      {stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211], stage0_1[212]},
      {stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage1_5[31],stage1_4[71],stage1_3[74],stage1_2[74],stage1_1[74]}
   );
   gpc606_5 gpc75 (
      {stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217], stage0_1[218]},
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200]},
      {stage1_5[32],stage1_4[72],stage1_3[75],stage1_2[75],stage1_1[75]}
   );
   gpc606_5 gpc76 (
      {stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223], stage0_1[224]},
      {stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage1_5[33],stage1_4[73],stage1_3[76],stage1_2[76],stage1_1[76]}
   );
   gpc606_5 gpc77 (
      {stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229], stage0_1[230]},
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212]},
      {stage1_5[34],stage1_4[74],stage1_3[77],stage1_2[77],stage1_1[77]}
   );
   gpc606_5 gpc78 (
      {stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235], stage0_1[236]},
      {stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218]},
      {stage1_5[35],stage1_4[75],stage1_3[78],stage1_2[78],stage1_1[78]}
   );
   gpc606_5 gpc79 (
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[36],stage1_4[76],stage1_3[79],stage1_2[79]}
   );
   gpc606_5 gpc80 (
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[37],stage1_4[77],stage1_3[80],stage1_2[80]}
   );
   gpc623_5 gpc81 (
      {stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage0_3[219], stage0_3[220]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[38],stage1_4[78],stage1_3[81],stage1_2[81]}
   );
   gpc615_5 gpc82 (
      {stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225]},
      {stage0_4[18]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[3],stage1_5[39],stage1_4[79],stage1_3[82]}
   );
   gpc615_5 gpc83 (
      {stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230]},
      {stage0_4[19]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[4],stage1_5[40],stage1_4[80],stage1_3[83]}
   );
   gpc615_5 gpc84 (
      {stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235]},
      {stage0_4[20]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[5],stage1_5[41],stage1_4[81],stage1_3[84]}
   );
   gpc615_5 gpc85 (
      {stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240]},
      {stage0_4[21]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[6],stage1_5[42],stage1_4[82],stage1_3[85]}
   );
   gpc615_5 gpc86 (
      {stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245]},
      {stage0_4[22]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[7],stage1_5[43],stage1_4[83],stage1_3[86]}
   );
   gpc615_5 gpc87 (
      {stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250]},
      {stage0_4[23]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[8],stage1_5[44],stage1_4[84],stage1_3[87]}
   );
   gpc623_5 gpc88 (
      {stage0_3[251], stage0_3[252], stage0_3[253]},
      {stage0_4[24], stage0_4[25]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[9],stage1_5[45],stage1_4[85],stage1_3[88]}
   );
   gpc1163_5 gpc89 (
      {stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_6[0]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[7],stage1_6[10],stage1_5[46],stage1_4[86]}
   );
   gpc1163_5 gpc90 (
      {stage0_4[29], stage0_4[30], stage0_4[31]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[1]},
      {stage0_7[1]},
      {stage1_8[1],stage1_7[8],stage1_6[11],stage1_5[47],stage1_4[87]}
   );
   gpc1163_5 gpc91 (
      {stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_6[2]},
      {stage0_7[2]},
      {stage1_8[2],stage1_7[9],stage1_6[12],stage1_5[48],stage1_4[88]}
   );
   gpc1163_5 gpc92 (
      {stage0_4[35], stage0_4[36], stage0_4[37]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_6[3]},
      {stage0_7[3]},
      {stage1_8[3],stage1_7[10],stage1_6[13],stage1_5[49],stage1_4[89]}
   );
   gpc1163_5 gpc93 (
      {stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_6[4]},
      {stage0_7[4]},
      {stage1_8[4],stage1_7[11],stage1_6[14],stage1_5[50],stage1_4[90]}
   );
   gpc1163_5 gpc94 (
      {stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_6[5]},
      {stage0_7[5]},
      {stage1_8[5],stage1_7[12],stage1_6[15],stage1_5[51],stage1_4[91]}
   );
   gpc606_5 gpc95 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[6],stage1_7[13],stage1_6[16],stage1_5[52],stage1_4[92]}
   );
   gpc606_5 gpc96 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[7],stage1_7[14],stage1_6[17],stage1_5[53],stage1_4[93]}
   );
   gpc606_5 gpc97 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[8],stage1_7[15],stage1_6[18],stage1_5[54],stage1_4[94]}
   );
   gpc606_5 gpc98 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[9],stage1_7[16],stage1_6[19],stage1_5[55],stage1_4[95]}
   );
   gpc606_5 gpc99 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[10],stage1_7[17],stage1_6[20],stage1_5[56],stage1_4[96]}
   );
   gpc606_5 gpc100 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[11],stage1_7[18],stage1_6[21],stage1_5[57],stage1_4[97]}
   );
   gpc606_5 gpc101 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[12],stage1_7[19],stage1_6[22],stage1_5[58],stage1_4[98]}
   );
   gpc606_5 gpc102 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[13],stage1_7[20],stage1_6[23],stage1_5[59],stage1_4[99]}
   );
   gpc606_5 gpc103 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[14],stage1_7[21],stage1_6[24],stage1_5[60],stage1_4[100]}
   );
   gpc606_5 gpc104 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[15],stage1_7[22],stage1_6[25],stage1_5[61],stage1_4[101]}
   );
   gpc606_5 gpc105 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[16],stage1_7[23],stage1_6[26],stage1_5[62],stage1_4[102]}
   );
   gpc606_5 gpc106 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[17],stage1_7[24],stage1_6[27],stage1_5[63],stage1_4[103]}
   );
   gpc606_5 gpc107 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[18],stage1_7[25],stage1_6[28],stage1_5[64],stage1_4[104]}
   );
   gpc606_5 gpc108 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[19],stage1_7[26],stage1_6[29],stage1_5[65],stage1_4[105]}
   );
   gpc606_5 gpc109 (
      {stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[20],stage1_7[27],stage1_6[30],stage1_5[66],stage1_4[106]}
   );
   gpc606_5 gpc110 (
      {stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[21],stage1_7[28],stage1_6[31],stage1_5[67],stage1_4[107]}
   );
   gpc606_5 gpc111 (
      {stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[22],stage1_7[29],stage1_6[32],stage1_5[68],stage1_4[108]}
   );
   gpc606_5 gpc112 (
      {stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[23],stage1_7[30],stage1_6[33],stage1_5[69],stage1_4[109]}
   );
   gpc606_5 gpc113 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[24],stage1_7[31],stage1_6[34],stage1_5[70],stage1_4[110]}
   );
   gpc606_5 gpc114 (
      {stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[25],stage1_7[32],stage1_6[35],stage1_5[71],stage1_4[111]}
   );
   gpc606_5 gpc115 (
      {stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[26],stage1_7[33],stage1_6[36],stage1_5[72],stage1_4[112]}
   );
   gpc606_5 gpc116 (
      {stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[27],stage1_7[34],stage1_6[37],stage1_5[73],stage1_4[113]}
   );
   gpc606_5 gpc117 (
      {stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[28],stage1_7[35],stage1_6[38],stage1_5[74],stage1_4[114]}
   );
   gpc606_5 gpc118 (
      {stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[29],stage1_7[36],stage1_6[39],stage1_5[75],stage1_4[115]}
   );
   gpc606_5 gpc119 (
      {stage0_4[188], stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[30],stage1_7[37],stage1_6[40],stage1_5[76],stage1_4[116]}
   );
   gpc606_5 gpc120 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[31],stage1_7[38],stage1_6[41],stage1_5[77],stage1_4[117]}
   );
   gpc606_5 gpc121 (
      {stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[32],stage1_7[39],stage1_6[42],stage1_5[78],stage1_4[118]}
   );
   gpc606_5 gpc122 (
      {stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[33],stage1_7[40],stage1_6[43],stage1_5[79],stage1_4[119]}
   );
   gpc606_5 gpc123 (
      {stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[34],stage1_7[41],stage1_6[44],stage1_5[80],stage1_4[120]}
   );
   gpc606_5 gpc124 (
      {stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[35],stage1_7[42],stage1_6[45],stage1_5[81],stage1_4[121]}
   );
   gpc606_5 gpc125 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[36],stage1_7[43],stage1_6[46],stage1_5[82],stage1_4[122]}
   );
   gpc606_5 gpc126 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[0],stage1_8[37],stage1_7[44],stage1_6[47],stage1_5[83]}
   );
   gpc606_5 gpc127 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[1],stage1_8[38],stage1_7[45],stage1_6[48],stage1_5[84]}
   );
   gpc606_5 gpc128 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[2],stage1_8[39],stage1_7[46],stage1_6[49],stage1_5[85]}
   );
   gpc606_5 gpc129 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[3],stage1_8[40],stage1_7[47],stage1_6[50],stage1_5[86]}
   );
   gpc606_5 gpc130 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[4],stage1_8[41],stage1_7[48],stage1_6[51],stage1_5[87]}
   );
   gpc606_5 gpc131 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[5],stage1_8[42],stage1_7[49],stage1_6[52],stage1_5[88]}
   );
   gpc606_5 gpc132 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[6],stage1_8[43],stage1_7[50],stage1_6[53],stage1_5[89]}
   );
   gpc606_5 gpc133 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[7],stage1_8[44],stage1_7[51],stage1_6[54],stage1_5[90]}
   );
   gpc606_5 gpc134 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[8],stage1_8[45],stage1_7[52],stage1_6[55],stage1_5[91]}
   );
   gpc606_5 gpc135 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[9],stage1_8[46],stage1_7[53],stage1_6[56],stage1_5[92]}
   );
   gpc606_5 gpc136 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[10],stage1_8[47],stage1_7[54],stage1_6[57],stage1_5[93]}
   );
   gpc606_5 gpc137 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[11],stage1_8[48],stage1_7[55],stage1_6[58],stage1_5[94]}
   );
   gpc606_5 gpc138 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[12],stage1_8[49],stage1_7[56],stage1_6[59],stage1_5[95]}
   );
   gpc606_5 gpc139 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[13],stage1_8[50],stage1_7[57],stage1_6[60],stage1_5[96]}
   );
   gpc606_5 gpc140 (
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[14],stage1_8[51],stage1_7[58],stage1_6[61],stage1_5[97]}
   );
   gpc606_5 gpc141 (
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[15],stage1_8[52],stage1_7[59],stage1_6[62],stage1_5[98]}
   );
   gpc606_5 gpc142 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[16],stage1_8[53],stage1_7[60],stage1_6[63],stage1_5[99]}
   );
   gpc606_5 gpc143 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[17],stage1_8[54],stage1_7[61],stage1_6[64],stage1_5[100]}
   );
   gpc606_5 gpc144 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[18],stage1_8[55],stage1_7[62],stage1_6[65],stage1_5[101]}
   );
   gpc606_5 gpc145 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[19],stage1_8[56],stage1_7[63],stage1_6[66],stage1_5[102]}
   );
   gpc606_5 gpc146 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[20],stage1_8[57],stage1_7[64],stage1_6[67],stage1_5[103]}
   );
   gpc606_5 gpc147 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[21],stage1_8[58],stage1_7[65],stage1_6[68],stage1_5[104]}
   );
   gpc606_5 gpc148 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[22],stage1_8[59],stage1_7[66],stage1_6[69],stage1_5[105]}
   );
   gpc606_5 gpc149 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[23],stage1_8[60],stage1_7[67],stage1_6[70],stage1_5[106]}
   );
   gpc606_5 gpc150 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[24],stage1_8[61],stage1_7[68],stage1_6[71],stage1_5[107]}
   );
   gpc606_5 gpc151 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[25],stage1_8[62],stage1_7[69],stage1_6[72],stage1_5[108]}
   );
   gpc606_5 gpc152 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[26],stage1_8[63],stage1_7[70],stage1_6[73],stage1_5[109]}
   );
   gpc606_5 gpc153 (
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[27],stage1_8[64],stage1_7[71],stage1_6[74]}
   );
   gpc606_5 gpc154 (
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[28],stage1_8[65],stage1_7[72],stage1_6[75]}
   );
   gpc606_5 gpc155 (
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[29],stage1_8[66],stage1_7[73],stage1_6[76]}
   );
   gpc606_5 gpc156 (
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[30],stage1_8[67],stage1_7[74],stage1_6[77]}
   );
   gpc606_5 gpc157 (
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[31],stage1_8[68],stage1_7[75],stage1_6[78]}
   );
   gpc606_5 gpc158 (
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[32],stage1_8[69],stage1_7[76],stage1_6[79]}
   );
   gpc615_5 gpc159 (
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232]},
      {stage0_7[168]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[33],stage1_8[70],stage1_7[77],stage1_6[80]}
   );
   gpc615_5 gpc160 (
      {stage0_6[233], stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237]},
      {stage0_7[169]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[34],stage1_8[71],stage1_7[78],stage1_6[81]}
   );
   gpc615_5 gpc161 (
      {stage0_6[238], stage0_6[239], stage0_6[240], stage0_6[241], stage0_6[242]},
      {stage0_7[170]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[35],stage1_8[72],stage1_7[79],stage1_6[82]}
   );
   gpc615_5 gpc162 (
      {stage0_7[171], stage0_7[172], stage0_7[173], stage0_7[174], stage0_7[175]},
      {stage0_8[54]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[9],stage1_9[36],stage1_8[73],stage1_7[80]}
   );
   gpc615_5 gpc163 (
      {stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179], stage0_7[180]},
      {stage0_8[55]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[10],stage1_9[37],stage1_8[74],stage1_7[81]}
   );
   gpc615_5 gpc164 (
      {stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage0_8[56]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[11],stage1_9[38],stage1_8[75],stage1_7[82]}
   );
   gpc615_5 gpc165 (
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190]},
      {stage0_8[57]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[12],stage1_9[39],stage1_8[76],stage1_7[83]}
   );
   gpc615_5 gpc166 (
      {stage0_7[191], stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195]},
      {stage0_8[58]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[13],stage1_9[40],stage1_8[77],stage1_7[84]}
   );
   gpc615_5 gpc167 (
      {stage0_7[196], stage0_7[197], stage0_7[198], stage0_7[199], stage0_7[200]},
      {stage0_8[59]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[14],stage1_9[41],stage1_8[78],stage1_7[85]}
   );
   gpc615_5 gpc168 (
      {stage0_7[201], stage0_7[202], stage0_7[203], stage0_7[204], stage0_7[205]},
      {stage0_8[60]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[15],stage1_9[42],stage1_8[79],stage1_7[86]}
   );
   gpc615_5 gpc169 (
      {stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209], stage0_7[210]},
      {stage0_8[61]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[16],stage1_9[43],stage1_8[80],stage1_7[87]}
   );
   gpc615_5 gpc170 (
      {stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage0_8[62]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[17],stage1_9[44],stage1_8[81],stage1_7[88]}
   );
   gpc615_5 gpc171 (
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220]},
      {stage0_8[63]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[18],stage1_9[45],stage1_8[82],stage1_7[89]}
   );
   gpc615_5 gpc172 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[64]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[19],stage1_9[46],stage1_8[83],stage1_7[90]}
   );
   gpc615_5 gpc173 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[65]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[20],stage1_9[47],stage1_8[84],stage1_7[91]}
   );
   gpc615_5 gpc174 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[66]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[21],stage1_9[48],stage1_8[85],stage1_7[92]}
   );
   gpc615_5 gpc175 (
      {stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239], stage0_7[240]},
      {stage0_8[67]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[22],stage1_9[49],stage1_8[86],stage1_7[93]}
   );
   gpc615_5 gpc176 (
      {stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage0_8[68]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[23],stage1_9[50],stage1_8[87],stage1_7[94]}
   );
   gpc615_5 gpc177 (
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250]},
      {stage0_8[69]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[24],stage1_9[51],stage1_8[88],stage1_7[95]}
   );
   gpc606_5 gpc178 (
      {stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[16],stage1_10[25],stage1_9[52],stage1_8[89]}
   );
   gpc606_5 gpc179 (
      {stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[17],stage1_10[26],stage1_9[53],stage1_8[90]}
   );
   gpc606_5 gpc180 (
      {stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[18],stage1_10[27],stage1_9[54],stage1_8[91]}
   );
   gpc606_5 gpc181 (
      {stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[19],stage1_10[28],stage1_9[55],stage1_8[92]}
   );
   gpc606_5 gpc182 (
      {stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[20],stage1_10[29],stage1_9[56],stage1_8[93]}
   );
   gpc606_5 gpc183 (
      {stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[21],stage1_10[30],stage1_9[57],stage1_8[94]}
   );
   gpc606_5 gpc184 (
      {stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[22],stage1_10[31],stage1_9[58],stage1_8[95]}
   );
   gpc606_5 gpc185 (
      {stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[23],stage1_10[32],stage1_9[59],stage1_8[96]}
   );
   gpc606_5 gpc186 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[24],stage1_10[33],stage1_9[60],stage1_8[97]}
   );
   gpc606_5 gpc187 (
      {stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[25],stage1_10[34],stage1_9[61],stage1_8[98]}
   );
   gpc606_5 gpc188 (
      {stage0_8[130], stage0_8[131], stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[26],stage1_10[35],stage1_9[62],stage1_8[99]}
   );
   gpc606_5 gpc189 (
      {stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[27],stage1_10[36],stage1_9[63],stage1_8[100]}
   );
   gpc606_5 gpc190 (
      {stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[28],stage1_10[37],stage1_9[64],stage1_8[101]}
   );
   gpc606_5 gpc191 (
      {stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[29],stage1_10[38],stage1_9[65],stage1_8[102]}
   );
   gpc606_5 gpc192 (
      {stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[30],stage1_10[39],stage1_9[66],stage1_8[103]}
   );
   gpc606_5 gpc193 (
      {stage0_8[160], stage0_8[161], stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[31],stage1_10[40],stage1_9[67],stage1_8[104]}
   );
   gpc606_5 gpc194 (
      {stage0_8[166], stage0_8[167], stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[32],stage1_10[41],stage1_9[68],stage1_8[105]}
   );
   gpc606_5 gpc195 (
      {stage0_8[172], stage0_8[173], stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[33],stage1_10[42],stage1_9[69],stage1_8[106]}
   );
   gpc606_5 gpc196 (
      {stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[34],stage1_10[43],stage1_9[70],stage1_8[107]}
   );
   gpc606_5 gpc197 (
      {stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[35],stage1_10[44],stage1_9[71],stage1_8[108]}
   );
   gpc606_5 gpc198 (
      {stage0_8[190], stage0_8[191], stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[36],stage1_10[45],stage1_9[72],stage1_8[109]}
   );
   gpc606_5 gpc199 (
      {stage0_8[196], stage0_8[197], stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[37],stage1_10[46],stage1_9[73],stage1_8[110]}
   );
   gpc606_5 gpc200 (
      {stage0_8[202], stage0_8[203], stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[38],stage1_10[47],stage1_9[74],stage1_8[111]}
   );
   gpc606_5 gpc201 (
      {stage0_8[208], stage0_8[209], stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[39],stage1_10[48],stage1_9[75],stage1_8[112]}
   );
   gpc606_5 gpc202 (
      {stage0_8[214], stage0_8[215], stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[40],stage1_10[49],stage1_9[76],stage1_8[113]}
   );
   gpc606_5 gpc203 (
      {stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[41],stage1_10[50],stage1_9[77],stage1_8[114]}
   );
   gpc606_5 gpc204 (
      {stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[42],stage1_10[51],stage1_9[78],stage1_8[115]}
   );
   gpc606_5 gpc205 (
      {stage0_8[232], stage0_8[233], stage0_8[234], stage0_8[235], stage0_8[236], stage0_8[237]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[43],stage1_10[52],stage1_9[79],stage1_8[116]}
   );
   gpc606_5 gpc206 (
      {stage0_8[238], stage0_8[239], stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[44],stage1_10[53],stage1_9[80],stage1_8[117]}
   );
   gpc606_5 gpc207 (
      {stage0_8[244], stage0_8[245], stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[45],stage1_10[54],stage1_9[81],stage1_8[118]}
   );
   gpc606_5 gpc208 (
      {stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253], stage0_8[254], stage0_8[255]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[46],stage1_10[55],stage1_9[82],stage1_8[119]}
   );
   gpc606_5 gpc209 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[31],stage1_11[47],stage1_10[56],stage1_9[83]}
   );
   gpc606_5 gpc210 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[32],stage1_11[48],stage1_10[57],stage1_9[84]}
   );
   gpc606_5 gpc211 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[33],stage1_11[49],stage1_10[58],stage1_9[85]}
   );
   gpc606_5 gpc212 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[34],stage1_11[50],stage1_10[59],stage1_9[86]}
   );
   gpc606_5 gpc213 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[35],stage1_11[51],stage1_10[60],stage1_9[87]}
   );
   gpc606_5 gpc214 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[36],stage1_11[52],stage1_10[61],stage1_9[88]}
   );
   gpc606_5 gpc215 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[37],stage1_11[53],stage1_10[62],stage1_9[89]}
   );
   gpc606_5 gpc216 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[38],stage1_11[54],stage1_10[63],stage1_9[90]}
   );
   gpc606_5 gpc217 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[39],stage1_11[55],stage1_10[64],stage1_9[91]}
   );
   gpc606_5 gpc218 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[40],stage1_11[56],stage1_10[65],stage1_9[92]}
   );
   gpc606_5 gpc219 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[41],stage1_11[57],stage1_10[66],stage1_9[93]}
   );
   gpc606_5 gpc220 (
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[42],stage1_11[58],stage1_10[67],stage1_9[94]}
   );
   gpc606_5 gpc221 (
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[43],stage1_11[59],stage1_10[68],stage1_9[95]}
   );
   gpc606_5 gpc222 (
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[44],stage1_11[60],stage1_10[69],stage1_9[96]}
   );
   gpc606_5 gpc223 (
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[45],stage1_11[61],stage1_10[70],stage1_9[97]}
   );
   gpc606_5 gpc224 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[46],stage1_11[62],stage1_10[71],stage1_9[98]}
   );
   gpc606_5 gpc225 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[47],stage1_11[63],stage1_10[72],stage1_9[99]}
   );
   gpc606_5 gpc226 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[48],stage1_11[64],stage1_10[73],stage1_9[100]}
   );
   gpc606_5 gpc227 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[49],stage1_11[65],stage1_10[74],stage1_9[101]}
   );
   gpc615_5 gpc228 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214]},
      {stage0_10[186]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[50],stage1_11[66],stage1_10[75],stage1_9[102]}
   );
   gpc615_5 gpc229 (
      {stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219]},
      {stage0_10[187]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[51],stage1_11[67],stage1_10[76],stage1_9[103]}
   );
   gpc615_5 gpc230 (
      {stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224]},
      {stage0_10[188]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[52],stage1_11[68],stage1_10[77],stage1_9[104]}
   );
   gpc615_5 gpc231 (
      {stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229]},
      {stage0_10[189]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[53],stage1_11[69],stage1_10[78],stage1_9[105]}
   );
   gpc615_5 gpc232 (
      {stage0_10[190], stage0_10[191], stage0_10[192], stage0_10[193], stage0_10[194]},
      {stage0_11[138]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[23],stage1_12[54],stage1_11[70],stage1_10[79]}
   );
   gpc615_5 gpc233 (
      {stage0_10[195], stage0_10[196], stage0_10[197], stage0_10[198], stage0_10[199]},
      {stage0_11[139]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[24],stage1_12[55],stage1_11[71],stage1_10[80]}
   );
   gpc615_5 gpc234 (
      {stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203], stage0_10[204]},
      {stage0_11[140]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[25],stage1_12[56],stage1_11[72],stage1_10[81]}
   );
   gpc615_5 gpc235 (
      {stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage0_11[141]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[26],stage1_12[57],stage1_11[73],stage1_10[82]}
   );
   gpc615_5 gpc236 (
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214]},
      {stage0_11[142]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[27],stage1_12[58],stage1_11[74],stage1_10[83]}
   );
   gpc615_5 gpc237 (
      {stage0_10[215], stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219]},
      {stage0_11[143]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[28],stage1_12[59],stage1_11[75],stage1_10[84]}
   );
   gpc615_5 gpc238 (
      {stage0_10[220], stage0_10[221], stage0_10[222], stage0_10[223], stage0_10[224]},
      {stage0_11[144]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[29],stage1_12[60],stage1_11[76],stage1_10[85]}
   );
   gpc615_5 gpc239 (
      {stage0_10[225], stage0_10[226], stage0_10[227], stage0_10[228], stage0_10[229]},
      {stage0_11[145]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[30],stage1_12[61],stage1_11[77],stage1_10[86]}
   );
   gpc615_5 gpc240 (
      {stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233], stage0_10[234]},
      {stage0_11[146]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[31],stage1_12[62],stage1_11[78],stage1_10[87]}
   );
   gpc615_5 gpc241 (
      {stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage0_11[147]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[32],stage1_12[63],stage1_11[79],stage1_10[88]}
   );
   gpc615_5 gpc242 (
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244]},
      {stage0_11[148]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[33],stage1_12[64],stage1_11[80],stage1_10[89]}
   );
   gpc615_5 gpc243 (
      {stage0_10[245], stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249]},
      {stage0_11[149]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[34],stage1_12[65],stage1_11[81],stage1_10[90]}
   );
   gpc615_5 gpc244 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154]},
      {stage0_12[72]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[12],stage1_13[35],stage1_12[66],stage1_11[82]}
   );
   gpc615_5 gpc245 (
      {stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159]},
      {stage0_12[73]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[13],stage1_13[36],stage1_12[67],stage1_11[83]}
   );
   gpc615_5 gpc246 (
      {stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164]},
      {stage0_12[74]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[14],stage1_13[37],stage1_12[68],stage1_11[84]}
   );
   gpc615_5 gpc247 (
      {stage0_11[165], stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169]},
      {stage0_12[75]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[15],stage1_13[38],stage1_12[69],stage1_11[85]}
   );
   gpc615_5 gpc248 (
      {stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173], stage0_11[174]},
      {stage0_12[76]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[16],stage1_13[39],stage1_12[70],stage1_11[86]}
   );
   gpc615_5 gpc249 (
      {stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage0_12[77]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[17],stage1_13[40],stage1_12[71],stage1_11[87]}
   );
   gpc615_5 gpc250 (
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184]},
      {stage0_12[78]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[18],stage1_13[41],stage1_12[72],stage1_11[88]}
   );
   gpc615_5 gpc251 (
      {stage0_11[185], stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189]},
      {stage0_12[79]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[19],stage1_13[42],stage1_12[73],stage1_11[89]}
   );
   gpc615_5 gpc252 (
      {stage0_11[190], stage0_11[191], stage0_11[192], stage0_11[193], stage0_11[194]},
      {stage0_12[80]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[20],stage1_13[43],stage1_12[74],stage1_11[90]}
   );
   gpc615_5 gpc253 (
      {stage0_11[195], stage0_11[196], stage0_11[197], stage0_11[198], stage0_11[199]},
      {stage0_12[81]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[21],stage1_13[44],stage1_12[75],stage1_11[91]}
   );
   gpc615_5 gpc254 (
      {stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203], stage0_11[204]},
      {stage0_12[82]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[22],stage1_13[45],stage1_12[76],stage1_11[92]}
   );
   gpc615_5 gpc255 (
      {stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage0_12[83]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[23],stage1_13[46],stage1_12[77],stage1_11[93]}
   );
   gpc117_4 gpc256 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90]},
      {stage0_13[72]},
      {stage0_14[0]},
      {stage1_15[12],stage1_14[24],stage1_13[47],stage1_12[78]}
   );
   gpc606_5 gpc257 (
      {stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96]},
      {stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5], stage0_14[6]},
      {stage1_16[0],stage1_15[13],stage1_14[25],stage1_13[48],stage1_12[79]}
   );
   gpc606_5 gpc258 (
      {stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102]},
      {stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11], stage0_14[12]},
      {stage1_16[1],stage1_15[14],stage1_14[26],stage1_13[49],stage1_12[80]}
   );
   gpc615_5 gpc259 (
      {stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_13[73]},
      {stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17], stage0_14[18]},
      {stage1_16[2],stage1_15[15],stage1_14[27],stage1_13[50],stage1_12[81]}
   );
   gpc615_5 gpc260 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112]},
      {stage0_13[74]},
      {stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23], stage0_14[24]},
      {stage1_16[3],stage1_15[16],stage1_14[28],stage1_13[51],stage1_12[82]}
   );
   gpc615_5 gpc261 (
      {stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117]},
      {stage0_13[75]},
      {stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29], stage0_14[30]},
      {stage1_16[4],stage1_15[17],stage1_14[29],stage1_13[52],stage1_12[83]}
   );
   gpc615_5 gpc262 (
      {stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122]},
      {stage0_13[76]},
      {stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35], stage0_14[36]},
      {stage1_16[5],stage1_15[18],stage1_14[30],stage1_13[53],stage1_12[84]}
   );
   gpc615_5 gpc263 (
      {stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_13[77]},
      {stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41], stage0_14[42]},
      {stage1_16[6],stage1_15[19],stage1_14[31],stage1_13[54],stage1_12[85]}
   );
   gpc615_5 gpc264 (
      {stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132]},
      {stage0_13[78]},
      {stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47], stage0_14[48]},
      {stage1_16[7],stage1_15[20],stage1_14[32],stage1_13[55],stage1_12[86]}
   );
   gpc615_5 gpc265 (
      {stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_13[79]},
      {stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53], stage0_14[54]},
      {stage1_16[8],stage1_15[21],stage1_14[33],stage1_13[56],stage1_12[87]}
   );
   gpc615_5 gpc266 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142]},
      {stage0_13[80]},
      {stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59], stage0_14[60]},
      {stage1_16[9],stage1_15[22],stage1_14[34],stage1_13[57],stage1_12[88]}
   );
   gpc615_5 gpc267 (
      {stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147]},
      {stage0_13[81]},
      {stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65], stage0_14[66]},
      {stage1_16[10],stage1_15[23],stage1_14[35],stage1_13[58],stage1_12[89]}
   );
   gpc606_5 gpc268 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[11],stage1_15[24],stage1_14[36],stage1_13[59]}
   );
   gpc606_5 gpc269 (
      {stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[12],stage1_15[25],stage1_14[37],stage1_13[60]}
   );
   gpc606_5 gpc270 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[13],stage1_15[26],stage1_14[38],stage1_13[61]}
   );
   gpc606_5 gpc271 (
      {stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[14],stage1_15[27],stage1_14[39],stage1_13[62]}
   );
   gpc615_5 gpc272 (
      {stage0_13[106], stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110]},
      {stage0_14[67]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[15],stage1_15[28],stage1_14[40],stage1_13[63]}
   );
   gpc615_5 gpc273 (
      {stage0_13[111], stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115]},
      {stage0_14[68]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[16],stage1_15[29],stage1_14[41],stage1_13[64]}
   );
   gpc615_5 gpc274 (
      {stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119], stage0_13[120]},
      {stage0_14[69]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[17],stage1_15[30],stage1_14[42],stage1_13[65]}
   );
   gpc615_5 gpc275 (
      {stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_14[70]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[18],stage1_15[31],stage1_14[43],stage1_13[66]}
   );
   gpc615_5 gpc276 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130]},
      {stage0_14[71]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[19],stage1_15[32],stage1_14[44],stage1_13[67]}
   );
   gpc615_5 gpc277 (
      {stage0_13[131], stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135]},
      {stage0_14[72]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[20],stage1_15[33],stage1_14[45],stage1_13[68]}
   );
   gpc615_5 gpc278 (
      {stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139], stage0_13[140]},
      {stage0_14[73]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[21],stage1_15[34],stage1_14[46],stage1_13[69]}
   );
   gpc615_5 gpc279 (
      {stage0_13[141], stage0_13[142], stage0_13[143], stage0_13[144], stage0_13[145]},
      {stage0_14[74]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[22],stage1_15[35],stage1_14[47],stage1_13[70]}
   );
   gpc615_5 gpc280 (
      {stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149], stage0_13[150]},
      {stage0_14[75]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[23],stage1_15[36],stage1_14[48],stage1_13[71]}
   );
   gpc615_5 gpc281 (
      {stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_14[76]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[24],stage1_15[37],stage1_14[49],stage1_13[72]}
   );
   gpc615_5 gpc282 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160]},
      {stage0_14[77]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[25],stage1_15[38],stage1_14[50],stage1_13[73]}
   );
   gpc615_5 gpc283 (
      {stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165]},
      {stage0_14[78]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[26],stage1_15[39],stage1_14[51],stage1_13[74]}
   );
   gpc615_5 gpc284 (
      {stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170]},
      {stage0_14[79]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[27],stage1_15[40],stage1_14[52],stage1_13[75]}
   );
   gpc615_5 gpc285 (
      {stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175]},
      {stage0_14[80]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[28],stage1_15[41],stage1_14[53],stage1_13[76]}
   );
   gpc615_5 gpc286 (
      {stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180]},
      {stage0_14[81]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[29],stage1_15[42],stage1_14[54],stage1_13[77]}
   );
   gpc615_5 gpc287 (
      {stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185]},
      {stage0_14[82]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[30],stage1_15[43],stage1_14[55],stage1_13[78]}
   );
   gpc615_5 gpc288 (
      {stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190]},
      {stage0_14[83]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[31],stage1_15[44],stage1_14[56],stage1_13[79]}
   );
   gpc615_5 gpc289 (
      {stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195]},
      {stage0_14[84]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[32],stage1_15[45],stage1_14[57],stage1_13[80]}
   );
   gpc615_5 gpc290 (
      {stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200]},
      {stage0_14[85]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[33],stage1_15[46],stage1_14[58],stage1_13[81]}
   );
   gpc615_5 gpc291 (
      {stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205]},
      {stage0_14[86]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[34],stage1_15[47],stage1_14[59],stage1_13[82]}
   );
   gpc615_5 gpc292 (
      {stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210]},
      {stage0_14[87]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[35],stage1_15[48],stage1_14[60],stage1_13[83]}
   );
   gpc615_5 gpc293 (
      {stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage0_14[88]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[36],stage1_15[49],stage1_14[61],stage1_13[84]}
   );
   gpc615_5 gpc294 (
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220]},
      {stage0_14[89]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[37],stage1_15[50],stage1_14[62],stage1_13[85]}
   );
   gpc615_5 gpc295 (
      {stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225]},
      {stage0_14[90]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[38],stage1_15[51],stage1_14[63],stage1_13[86]}
   );
   gpc615_5 gpc296 (
      {stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_14[91]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[39],stage1_15[52],stage1_14[64],stage1_13[87]}
   );
   gpc615_5 gpc297 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_14[92]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[40],stage1_15[53],stage1_14[65],stage1_13[88]}
   );
   gpc615_5 gpc298 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240]},
      {stage0_14[93]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[41],stage1_15[54],stage1_14[66],stage1_13[89]}
   );
   gpc615_5 gpc299 (
      {stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_14[94]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[42],stage1_15[55],stage1_14[67],stage1_13[90]}
   );
   gpc615_5 gpc300 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250]},
      {stage0_14[95]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[43],stage1_15[56],stage1_14[68],stage1_13[91]}
   );
   gpc615_5 gpc301 (
      {stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255]},
      {stage0_14[96]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[44],stage1_15[57],stage1_14[69],stage1_13[92]}
   );
   gpc606_5 gpc302 (
      {stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101], stage0_14[102]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[34],stage1_16[45],stage1_15[58],stage1_14[70]}
   );
   gpc606_5 gpc303 (
      {stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107], stage0_14[108]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[35],stage1_16[46],stage1_15[59],stage1_14[71]}
   );
   gpc606_5 gpc304 (
      {stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113], stage0_14[114]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[36],stage1_16[47],stage1_15[60],stage1_14[72]}
   );
   gpc606_5 gpc305 (
      {stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119], stage0_14[120]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[37],stage1_16[48],stage1_15[61],stage1_14[73]}
   );
   gpc606_5 gpc306 (
      {stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125], stage0_14[126]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[38],stage1_16[49],stage1_15[62],stage1_14[74]}
   );
   gpc606_5 gpc307 (
      {stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[39],stage1_16[50],stage1_15[63],stage1_14[75]}
   );
   gpc606_5 gpc308 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[40],stage1_16[51],stage1_15[64],stage1_14[76]}
   );
   gpc606_5 gpc309 (
      {stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143], stage0_14[144]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[41],stage1_16[52],stage1_15[65],stage1_14[77]}
   );
   gpc606_5 gpc310 (
      {stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149], stage0_14[150]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[42],stage1_16[53],stage1_15[66],stage1_14[78]}
   );
   gpc606_5 gpc311 (
      {stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155], stage0_14[156]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[43],stage1_16[54],stage1_15[67],stage1_14[79]}
   );
   gpc606_5 gpc312 (
      {stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161], stage0_14[162]},
      {stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65]},
      {stage1_18[10],stage1_17[44],stage1_16[55],stage1_15[68],stage1_14[80]}
   );
   gpc606_5 gpc313 (
      {stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167], stage0_14[168]},
      {stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71]},
      {stage1_18[11],stage1_17[45],stage1_16[56],stage1_15[69],stage1_14[81]}
   );
   gpc606_5 gpc314 (
      {stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173], stage0_14[174]},
      {stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77]},
      {stage1_18[12],stage1_17[46],stage1_16[57],stage1_15[70],stage1_14[82]}
   );
   gpc606_5 gpc315 (
      {stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179], stage0_14[180]},
      {stage0_16[78], stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83]},
      {stage1_18[13],stage1_17[47],stage1_16[58],stage1_15[71],stage1_14[83]}
   );
   gpc606_5 gpc316 (
      {stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185], stage0_14[186]},
      {stage0_16[84], stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89]},
      {stage1_18[14],stage1_17[48],stage1_16[59],stage1_15[72],stage1_14[84]}
   );
   gpc606_5 gpc317 (
      {stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191], stage0_14[192]},
      {stage0_16[90], stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95]},
      {stage1_18[15],stage1_17[49],stage1_16[60],stage1_15[73],stage1_14[85]}
   );
   gpc606_5 gpc318 (
      {stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197], stage0_14[198]},
      {stage0_16[96], stage0_16[97], stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101]},
      {stage1_18[16],stage1_17[50],stage1_16[61],stage1_15[74],stage1_14[86]}
   );
   gpc606_5 gpc319 (
      {stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203], stage0_14[204]},
      {stage0_16[102], stage0_16[103], stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107]},
      {stage1_18[17],stage1_17[51],stage1_16[62],stage1_15[75],stage1_14[87]}
   );
   gpc606_5 gpc320 (
      {stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209], stage0_14[210]},
      {stage0_16[108], stage0_16[109], stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113]},
      {stage1_18[18],stage1_17[52],stage1_16[63],stage1_15[76],stage1_14[88]}
   );
   gpc606_5 gpc321 (
      {stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215], stage0_14[216]},
      {stage0_16[114], stage0_16[115], stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119]},
      {stage1_18[19],stage1_17[53],stage1_16[64],stage1_15[77],stage1_14[89]}
   );
   gpc606_5 gpc322 (
      {stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221], stage0_14[222]},
      {stage0_16[120], stage0_16[121], stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125]},
      {stage1_18[20],stage1_17[54],stage1_16[65],stage1_15[78],stage1_14[90]}
   );
   gpc606_5 gpc323 (
      {stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227], stage0_14[228]},
      {stage0_16[126], stage0_16[127], stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131]},
      {stage1_18[21],stage1_17[55],stage1_16[66],stage1_15[79],stage1_14[91]}
   );
   gpc606_5 gpc324 (
      {stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233], stage0_14[234]},
      {stage0_16[132], stage0_16[133], stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137]},
      {stage1_18[22],stage1_17[56],stage1_16[67],stage1_15[80],stage1_14[92]}
   );
   gpc615_5 gpc325 (
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208]},
      {stage0_16[138]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[23],stage1_17[57],stage1_16[68],stage1_15[81]}
   );
   gpc615_5 gpc326 (
      {stage0_15[209], stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213]},
      {stage0_16[139]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[24],stage1_17[58],stage1_16[69],stage1_15[82]}
   );
   gpc615_5 gpc327 (
      {stage0_15[214], stage0_15[215], stage0_15[216], stage0_15[217], stage0_15[218]},
      {stage0_16[140]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[25],stage1_17[59],stage1_16[70],stage1_15[83]}
   );
   gpc615_5 gpc328 (
      {stage0_15[219], stage0_15[220], stage0_15[221], stage0_15[222], stage0_15[223]},
      {stage0_16[141]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[26],stage1_17[60],stage1_16[71],stage1_15[84]}
   );
   gpc615_5 gpc329 (
      {stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227], stage0_15[228]},
      {stage0_16[142]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[27],stage1_17[61],stage1_16[72],stage1_15[85]}
   );
   gpc615_5 gpc330 (
      {stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage0_16[143]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[28],stage1_17[62],stage1_16[73],stage1_15[86]}
   );
   gpc615_5 gpc331 (
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238]},
      {stage0_16[144]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[29],stage1_17[63],stage1_16[74],stage1_15[87]}
   );
   gpc615_5 gpc332 (
      {stage0_15[239], stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243]},
      {stage0_16[145]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[30],stage1_17[64],stage1_16[75],stage1_15[88]}
   );
   gpc615_5 gpc333 (
      {stage0_15[244], stage0_15[245], stage0_15[246], stage0_15[247], stage0_15[248]},
      {stage0_16[146]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[31],stage1_17[65],stage1_16[76],stage1_15[89]}
   );
   gpc615_5 gpc334 (
      {stage0_15[249], stage0_15[250], stage0_15[251], stage0_15[252], stage0_15[253]},
      {stage0_16[147]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[32],stage1_17[66],stage1_16[77],stage1_15[90]}
   );
   gpc606_5 gpc335 (
      {stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151], stage0_16[152], stage0_16[153]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[10],stage1_18[33],stage1_17[67],stage1_16[78]}
   );
   gpc606_5 gpc336 (
      {stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157], stage0_16[158], stage0_16[159]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[11],stage1_18[34],stage1_17[68],stage1_16[79]}
   );
   gpc606_5 gpc337 (
      {stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163], stage0_16[164], stage0_16[165]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[12],stage1_18[35],stage1_17[69],stage1_16[80]}
   );
   gpc606_5 gpc338 (
      {stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169], stage0_16[170], stage0_16[171]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[13],stage1_18[36],stage1_17[70],stage1_16[81]}
   );
   gpc606_5 gpc339 (
      {stage0_16[172], stage0_16[173], stage0_16[174], stage0_16[175], stage0_16[176], stage0_16[177]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[14],stage1_18[37],stage1_17[71],stage1_16[82]}
   );
   gpc606_5 gpc340 (
      {stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181], stage0_16[182], stage0_16[183]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[15],stage1_18[38],stage1_17[72],stage1_16[83]}
   );
   gpc606_5 gpc341 (
      {stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187], stage0_16[188], stage0_16[189]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[16],stage1_18[39],stage1_17[73],stage1_16[84]}
   );
   gpc606_5 gpc342 (
      {stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193], stage0_16[194], stage0_16[195]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[17],stage1_18[40],stage1_17[74],stage1_16[85]}
   );
   gpc606_5 gpc343 (
      {stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199], stage0_16[200], stage0_16[201]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[18],stage1_18[41],stage1_17[75],stage1_16[86]}
   );
   gpc606_5 gpc344 (
      {stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205], stage0_16[206], stage0_16[207]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[19],stage1_18[42],stage1_17[76],stage1_16[87]}
   );
   gpc606_5 gpc345 (
      {stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211], stage0_16[212], stage0_16[213]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[20],stage1_18[43],stage1_17[77],stage1_16[88]}
   );
   gpc606_5 gpc346 (
      {stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217], stage0_16[218], stage0_16[219]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[21],stage1_18[44],stage1_17[78],stage1_16[89]}
   );
   gpc606_5 gpc347 (
      {stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223], stage0_16[224], stage0_16[225]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[22],stage1_18[45],stage1_17[79],stage1_16[90]}
   );
   gpc606_5 gpc348 (
      {stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229], stage0_16[230], stage0_16[231]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[23],stage1_18[46],stage1_17[80],stage1_16[91]}
   );
   gpc606_5 gpc349 (
      {stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235], stage0_16[236], stage0_16[237]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[24],stage1_18[47],stage1_17[81],stage1_16[92]}
   );
   gpc606_5 gpc350 (
      {stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241], stage0_16[242], stage0_16[243]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[25],stage1_18[48],stage1_17[82],stage1_16[93]}
   );
   gpc606_5 gpc351 (
      {stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247], stage0_16[248], stage0_16[249]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[26],stage1_18[49],stage1_17[83],stage1_16[94]}
   );
   gpc606_5 gpc352 (
      {stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253], stage0_16[254], stage0_16[255]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[27],stage1_18[50],stage1_17[84],stage1_16[95]}
   );
   gpc606_5 gpc353 (
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[18],stage1_19[28],stage1_18[51],stage1_17[85]}
   );
   gpc606_5 gpc354 (
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[19],stage1_19[29],stage1_18[52],stage1_17[86]}
   );
   gpc615_5 gpc355 (
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76]},
      {stage0_18[108]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[20],stage1_19[30],stage1_18[53],stage1_17[87]}
   );
   gpc615_5 gpc356 (
      {stage0_17[77], stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81]},
      {stage0_18[109]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[21],stage1_19[31],stage1_18[54],stage1_17[88]}
   );
   gpc615_5 gpc357 (
      {stage0_17[82], stage0_17[83], stage0_17[84], stage0_17[85], stage0_17[86]},
      {stage0_18[110]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[22],stage1_19[32],stage1_18[55],stage1_17[89]}
   );
   gpc615_5 gpc358 (
      {stage0_17[87], stage0_17[88], stage0_17[89], stage0_17[90], stage0_17[91]},
      {stage0_18[111]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[23],stage1_19[33],stage1_18[56],stage1_17[90]}
   );
   gpc615_5 gpc359 (
      {stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95], stage0_17[96]},
      {stage0_18[112]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[24],stage1_19[34],stage1_18[57],stage1_17[91]}
   );
   gpc615_5 gpc360 (
      {stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage0_18[113]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[25],stage1_19[35],stage1_18[58],stage1_17[92]}
   );
   gpc615_5 gpc361 (
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106]},
      {stage0_18[114]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[26],stage1_19[36],stage1_18[59],stage1_17[93]}
   );
   gpc615_5 gpc362 (
      {stage0_17[107], stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111]},
      {stage0_18[115]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[27],stage1_19[37],stage1_18[60],stage1_17[94]}
   );
   gpc615_5 gpc363 (
      {stage0_17[112], stage0_17[113], stage0_17[114], stage0_17[115], stage0_17[116]},
      {stage0_18[116]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[28],stage1_19[38],stage1_18[61],stage1_17[95]}
   );
   gpc615_5 gpc364 (
      {stage0_17[117], stage0_17[118], stage0_17[119], stage0_17[120], stage0_17[121]},
      {stage0_18[117]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[29],stage1_19[39],stage1_18[62],stage1_17[96]}
   );
   gpc615_5 gpc365 (
      {stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125], stage0_17[126]},
      {stage0_18[118]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[30],stage1_19[40],stage1_18[63],stage1_17[97]}
   );
   gpc615_5 gpc366 (
      {stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage0_18[119]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[31],stage1_19[41],stage1_18[64],stage1_17[98]}
   );
   gpc615_5 gpc367 (
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136]},
      {stage0_18[120]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[32],stage1_19[42],stage1_18[65],stage1_17[99]}
   );
   gpc615_5 gpc368 (
      {stage0_17[137], stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141]},
      {stage0_18[121]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[33],stage1_19[43],stage1_18[66],stage1_17[100]}
   );
   gpc615_5 gpc369 (
      {stage0_17[142], stage0_17[143], stage0_17[144], stage0_17[145], stage0_17[146]},
      {stage0_18[122]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[34],stage1_19[44],stage1_18[67],stage1_17[101]}
   );
   gpc615_5 gpc370 (
      {stage0_17[147], stage0_17[148], stage0_17[149], stage0_17[150], stage0_17[151]},
      {stage0_18[123]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[35],stage1_19[45],stage1_18[68],stage1_17[102]}
   );
   gpc615_5 gpc371 (
      {stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155], stage0_17[156]},
      {stage0_18[124]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[36],stage1_19[46],stage1_18[69],stage1_17[103]}
   );
   gpc615_5 gpc372 (
      {stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage0_18[125]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[37],stage1_19[47],stage1_18[70],stage1_17[104]}
   );
   gpc615_5 gpc373 (
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166]},
      {stage0_18[126]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[38],stage1_19[48],stage1_18[71],stage1_17[105]}
   );
   gpc615_5 gpc374 (
      {stage0_17[167], stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171]},
      {stage0_18[127]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[39],stage1_19[49],stage1_18[72],stage1_17[106]}
   );
   gpc615_5 gpc375 (
      {stage0_17[172], stage0_17[173], stage0_17[174], stage0_17[175], stage0_17[176]},
      {stage0_18[128]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[40],stage1_19[50],stage1_18[73],stage1_17[107]}
   );
   gpc615_5 gpc376 (
      {stage0_17[177], stage0_17[178], stage0_17[179], stage0_17[180], stage0_17[181]},
      {stage0_18[129]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[41],stage1_19[51],stage1_18[74],stage1_17[108]}
   );
   gpc615_5 gpc377 (
      {stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185], stage0_17[186]},
      {stage0_18[130]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[42],stage1_19[52],stage1_18[75],stage1_17[109]}
   );
   gpc615_5 gpc378 (
      {stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage0_18[131]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[43],stage1_19[53],stage1_18[76],stage1_17[110]}
   );
   gpc615_5 gpc379 (
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196]},
      {stage0_18[132]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[44],stage1_19[54],stage1_18[77],stage1_17[111]}
   );
   gpc615_5 gpc380 (
      {stage0_17[197], stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201]},
      {stage0_18[133]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[45],stage1_19[55],stage1_18[78],stage1_17[112]}
   );
   gpc615_5 gpc381 (
      {stage0_17[202], stage0_17[203], stage0_17[204], stage0_17[205], stage0_17[206]},
      {stage0_18[134]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[46],stage1_19[56],stage1_18[79],stage1_17[113]}
   );
   gpc615_5 gpc382 (
      {stage0_17[207], stage0_17[208], stage0_17[209], stage0_17[210], stage0_17[211]},
      {stage0_18[135]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[47],stage1_19[57],stage1_18[80],stage1_17[114]}
   );
   gpc615_5 gpc383 (
      {stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215], stage0_17[216]},
      {stage0_18[136]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[48],stage1_19[58],stage1_18[81],stage1_17[115]}
   );
   gpc615_5 gpc384 (
      {stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage0_18[137]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[49],stage1_19[59],stage1_18[82],stage1_17[116]}
   );
   gpc615_5 gpc385 (
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226]},
      {stage0_18[138]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[50],stage1_19[60],stage1_18[83],stage1_17[117]}
   );
   gpc615_5 gpc386 (
      {stage0_17[227], stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231]},
      {stage0_18[139]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[51],stage1_19[61],stage1_18[84],stage1_17[118]}
   );
   gpc615_5 gpc387 (
      {stage0_17[232], stage0_17[233], stage0_17[234], stage0_17[235], stage0_17[236]},
      {stage0_18[140]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[52],stage1_19[62],stage1_18[85],stage1_17[119]}
   );
   gpc615_5 gpc388 (
      {stage0_17[237], stage0_17[238], stage0_17[239], stage0_17[240], stage0_17[241]},
      {stage0_18[141]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[53],stage1_19[63],stage1_18[86],stage1_17[120]}
   );
   gpc615_5 gpc389 (
      {stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245], stage0_17[246]},
      {stage0_18[142]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[54],stage1_19[64],stage1_18[87],stage1_17[121]}
   );
   gpc615_5 gpc390 (
      {stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage0_18[143]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[55],stage1_19[65],stage1_18[88],stage1_17[122]}
   );
   gpc606_5 gpc391 (
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[38],stage1_20[56],stage1_19[66],stage1_18[89]}
   );
   gpc606_5 gpc392 (
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[39],stage1_20[57],stage1_19[67],stage1_18[90]}
   );
   gpc606_5 gpc393 (
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[40],stage1_20[58],stage1_19[68],stage1_18[91]}
   );
   gpc606_5 gpc394 (
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[41],stage1_20[59],stage1_19[69],stage1_18[92]}
   );
   gpc606_5 gpc395 (
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[42],stage1_20[60],stage1_19[70],stage1_18[93]}
   );
   gpc606_5 gpc396 (
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[43],stage1_20[61],stage1_19[71],stage1_18[94]}
   );
   gpc606_5 gpc397 (
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[44],stage1_20[62],stage1_19[72],stage1_18[95]}
   );
   gpc606_5 gpc398 (
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[45],stage1_20[63],stage1_19[73],stage1_18[96]}
   );
   gpc606_5 gpc399 (
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[46],stage1_20[64],stage1_19[74],stage1_18[97]}
   );
   gpc606_5 gpc400 (
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[47],stage1_20[65],stage1_19[75],stage1_18[98]}
   );
   gpc606_5 gpc401 (
      {stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231], stage0_19[232], stage0_19[233]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[10],stage1_21[48],stage1_20[66],stage1_19[76]}
   );
   gpc606_5 gpc402 (
      {stage0_19[234], stage0_19[235], stage0_19[236], stage0_19[237], stage0_19[238], stage0_19[239]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[11],stage1_21[49],stage1_20[67],stage1_19[77]}
   );
   gpc615_5 gpc403 (
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64]},
      {stage0_21[12]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[12],stage1_21[50],stage1_20[68]}
   );
   gpc615_5 gpc404 (
      {stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69]},
      {stage0_21[13]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[13],stage1_21[51],stage1_20[69]}
   );
   gpc615_5 gpc405 (
      {stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74]},
      {stage0_21[14]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[14],stage1_21[52],stage1_20[70]}
   );
   gpc615_5 gpc406 (
      {stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79]},
      {stage0_21[15]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[5],stage1_22[15],stage1_21[53],stage1_20[71]}
   );
   gpc615_5 gpc407 (
      {stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84]},
      {stage0_21[16]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[6],stage1_22[16],stage1_21[54],stage1_20[72]}
   );
   gpc615_5 gpc408 (
      {stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage0_21[17]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[7],stage1_22[17],stage1_21[55],stage1_20[73]}
   );
   gpc615_5 gpc409 (
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94]},
      {stage0_21[18]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[8],stage1_22[18],stage1_21[56],stage1_20[74]}
   );
   gpc615_5 gpc410 (
      {stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99]},
      {stage0_21[19]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[9],stage1_22[19],stage1_21[57],stage1_20[75]}
   );
   gpc615_5 gpc411 (
      {stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104]},
      {stage0_21[20]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[10],stage1_22[20],stage1_21[58],stage1_20[76]}
   );
   gpc615_5 gpc412 (
      {stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109]},
      {stage0_21[21]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[11],stage1_22[21],stage1_21[59],stage1_20[77]}
   );
   gpc615_5 gpc413 (
      {stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114]},
      {stage0_21[22]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[12],stage1_22[22],stage1_21[60],stage1_20[78]}
   );
   gpc615_5 gpc414 (
      {stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage0_21[23]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[13],stage1_22[23],stage1_21[61],stage1_20[79]}
   );
   gpc615_5 gpc415 (
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124]},
      {stage0_21[24]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[14],stage1_22[24],stage1_21[62],stage1_20[80]}
   );
   gpc615_5 gpc416 (
      {stage0_20[125], stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129]},
      {stage0_21[25]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[15],stage1_22[25],stage1_21[63],stage1_20[81]}
   );
   gpc615_5 gpc417 (
      {stage0_20[130], stage0_20[131], stage0_20[132], stage0_20[133], stage0_20[134]},
      {stage0_21[26]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[16],stage1_22[26],stage1_21[64],stage1_20[82]}
   );
   gpc615_5 gpc418 (
      {stage0_20[135], stage0_20[136], stage0_20[137], stage0_20[138], stage0_20[139]},
      {stage0_21[27]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[17],stage1_22[27],stage1_21[65],stage1_20[83]}
   );
   gpc615_5 gpc419 (
      {stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143], stage0_20[144]},
      {stage0_21[28]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[18],stage1_22[28],stage1_21[66],stage1_20[84]}
   );
   gpc615_5 gpc420 (
      {stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage0_21[29]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[19],stage1_22[29],stage1_21[67],stage1_20[85]}
   );
   gpc615_5 gpc421 (
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154]},
      {stage0_21[30]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[20],stage1_22[30],stage1_21[68],stage1_20[86]}
   );
   gpc615_5 gpc422 (
      {stage0_20[155], stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159]},
      {stage0_21[31]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[21],stage1_22[31],stage1_21[69],stage1_20[87]}
   );
   gpc615_5 gpc423 (
      {stage0_20[160], stage0_20[161], stage0_20[162], stage0_20[163], stage0_20[164]},
      {stage0_21[32]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[22],stage1_22[32],stage1_21[70],stage1_20[88]}
   );
   gpc615_5 gpc424 (
      {stage0_20[165], stage0_20[166], stage0_20[167], stage0_20[168], stage0_20[169]},
      {stage0_21[33]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[23],stage1_22[33],stage1_21[71],stage1_20[89]}
   );
   gpc615_5 gpc425 (
      {stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173], stage0_20[174]},
      {stage0_21[34]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[24],stage1_22[34],stage1_21[72],stage1_20[90]}
   );
   gpc615_5 gpc426 (
      {stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage0_21[35]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[25],stage1_22[35],stage1_21[73],stage1_20[91]}
   );
   gpc615_5 gpc427 (
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184]},
      {stage0_21[36]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[26],stage1_22[36],stage1_21[74],stage1_20[92]}
   );
   gpc615_5 gpc428 (
      {stage0_20[185], stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189]},
      {stage0_21[37]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[27],stage1_22[37],stage1_21[75],stage1_20[93]}
   );
   gpc615_5 gpc429 (
      {stage0_20[190], stage0_20[191], stage0_20[192], stage0_20[193], stage0_20[194]},
      {stage0_21[38]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[28],stage1_22[38],stage1_21[76],stage1_20[94]}
   );
   gpc615_5 gpc430 (
      {stage0_20[195], stage0_20[196], stage0_20[197], stage0_20[198], stage0_20[199]},
      {stage0_21[39]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[29],stage1_22[39],stage1_21[77],stage1_20[95]}
   );
   gpc615_5 gpc431 (
      {stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203], stage0_20[204]},
      {stage0_21[40]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[30],stage1_22[40],stage1_21[78],stage1_20[96]}
   );
   gpc615_5 gpc432 (
      {stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209]},
      {stage0_21[41]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[31],stage1_22[41],stage1_21[79],stage1_20[97]}
   );
   gpc615_5 gpc433 (
      {stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213], stage0_20[214]},
      {stage0_21[42]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[32],stage1_22[42],stage1_21[80],stage1_20[98]}
   );
   gpc615_5 gpc434 (
      {stage0_20[215], stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219]},
      {stage0_21[43]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[33],stage1_22[43],stage1_21[81],stage1_20[99]}
   );
   gpc615_5 gpc435 (
      {stage0_20[220], stage0_20[221], stage0_20[222], stage0_20[223], stage0_20[224]},
      {stage0_21[44]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[34],stage1_22[44],stage1_21[82],stage1_20[100]}
   );
   gpc615_5 gpc436 (
      {stage0_20[225], stage0_20[226], stage0_20[227], stage0_20[228], stage0_20[229]},
      {stage0_21[45]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[35],stage1_22[45],stage1_21[83],stage1_20[101]}
   );
   gpc615_5 gpc437 (
      {stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233], stage0_20[234]},
      {stage0_21[46]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[36],stage1_22[46],stage1_21[84],stage1_20[102]}
   );
   gpc615_5 gpc438 (
      {stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239]},
      {stage0_21[47]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[37],stage1_22[47],stage1_21[85],stage1_20[103]}
   );
   gpc615_5 gpc439 (
      {stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244]},
      {stage0_21[48]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[38],stage1_22[48],stage1_21[86],stage1_20[104]}
   );
   gpc606_5 gpc440 (
      {stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53], stage0_21[54]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[37],stage1_23[39],stage1_22[49],stage1_21[87]}
   );
   gpc606_5 gpc441 (
      {stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59], stage0_21[60]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[38],stage1_23[40],stage1_22[50],stage1_21[88]}
   );
   gpc606_5 gpc442 (
      {stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65], stage0_21[66]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[39],stage1_23[41],stage1_22[51],stage1_21[89]}
   );
   gpc606_5 gpc443 (
      {stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71], stage0_21[72]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[40],stage1_23[42],stage1_22[52],stage1_21[90]}
   );
   gpc606_5 gpc444 (
      {stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77], stage0_21[78]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[41],stage1_23[43],stage1_22[53],stage1_21[91]}
   );
   gpc606_5 gpc445 (
      {stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83], stage0_21[84]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[42],stage1_23[44],stage1_22[54],stage1_21[92]}
   );
   gpc606_5 gpc446 (
      {stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89], stage0_21[90]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[43],stage1_23[45],stage1_22[55],stage1_21[93]}
   );
   gpc606_5 gpc447 (
      {stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95], stage0_21[96]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[44],stage1_23[46],stage1_22[56],stage1_21[94]}
   );
   gpc606_5 gpc448 (
      {stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101], stage0_21[102]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[45],stage1_23[47],stage1_22[57],stage1_21[95]}
   );
   gpc606_5 gpc449 (
      {stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107], stage0_21[108]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[46],stage1_23[48],stage1_22[58],stage1_21[96]}
   );
   gpc606_5 gpc450 (
      {stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113], stage0_21[114]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[47],stage1_23[49],stage1_22[59],stage1_21[97]}
   );
   gpc606_5 gpc451 (
      {stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119], stage0_21[120]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[48],stage1_23[50],stage1_22[60],stage1_21[98]}
   );
   gpc606_5 gpc452 (
      {stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125], stage0_21[126]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[49],stage1_23[51],stage1_22[61],stage1_21[99]}
   );
   gpc606_5 gpc453 (
      {stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131], stage0_21[132]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[50],stage1_23[52],stage1_22[62],stage1_21[100]}
   );
   gpc606_5 gpc454 (
      {stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137], stage0_21[138]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[51],stage1_23[53],stage1_22[63],stage1_21[101]}
   );
   gpc606_5 gpc455 (
      {stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143], stage0_21[144]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[52],stage1_23[54],stage1_22[64],stage1_21[102]}
   );
   gpc606_5 gpc456 (
      {stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149], stage0_21[150]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[53],stage1_23[55],stage1_22[65],stage1_21[103]}
   );
   gpc606_5 gpc457 (
      {stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155], stage0_21[156]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[54],stage1_23[56],stage1_22[66],stage1_21[104]}
   );
   gpc606_5 gpc458 (
      {stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161], stage0_21[162]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[55],stage1_23[57],stage1_22[67],stage1_21[105]}
   );
   gpc606_5 gpc459 (
      {stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167], stage0_21[168]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[56],stage1_23[58],stage1_22[68],stage1_21[106]}
   );
   gpc606_5 gpc460 (
      {stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173], stage0_21[174]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[57],stage1_23[59],stage1_22[69],stage1_21[107]}
   );
   gpc606_5 gpc461 (
      {stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179], stage0_21[180]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[58],stage1_23[60],stage1_22[70],stage1_21[108]}
   );
   gpc606_5 gpc462 (
      {stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185], stage0_21[186]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[59],stage1_23[61],stage1_22[71],stage1_21[109]}
   );
   gpc606_5 gpc463 (
      {stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191], stage0_21[192]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[60],stage1_23[62],stage1_22[72],stage1_21[110]}
   );
   gpc606_5 gpc464 (
      {stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197], stage0_21[198]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[61],stage1_23[63],stage1_22[73],stage1_21[111]}
   );
   gpc606_5 gpc465 (
      {stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203], stage0_21[204]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[62],stage1_23[64],stage1_22[74],stage1_21[112]}
   );
   gpc606_5 gpc466 (
      {stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209], stage0_21[210]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[63],stage1_23[65],stage1_22[75],stage1_21[113]}
   );
   gpc606_5 gpc467 (
      {stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215], stage0_21[216]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[64],stage1_23[66],stage1_22[76],stage1_21[114]}
   );
   gpc606_5 gpc468 (
      {stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221], stage0_21[222]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[65],stage1_23[67],stage1_22[77],stage1_21[115]}
   );
   gpc606_5 gpc469 (
      {stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227], stage0_21[228]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[66],stage1_23[68],stage1_22[78],stage1_21[116]}
   );
   gpc606_5 gpc470 (
      {stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233], stage0_21[234]},
      {stage0_23[180], stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage1_25[30],stage1_24[67],stage1_23[69],stage1_22[79],stage1_21[117]}
   );
   gpc606_5 gpc471 (
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[31],stage1_24[68],stage1_23[70],stage1_22[80]}
   );
   gpc606_5 gpc472 (
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[32],stage1_24[69],stage1_23[71],stage1_22[81]}
   );
   gpc606_5 gpc473 (
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[33],stage1_24[70],stage1_23[72],stage1_22[82]}
   );
   gpc606_5 gpc474 (
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[34],stage1_24[71],stage1_23[73],stage1_22[83]}
   );
   gpc606_5 gpc475 (
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190], stage0_23[191]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[4],stage1_25[35],stage1_24[72],stage1_23[74]}
   );
   gpc606_5 gpc476 (
      {stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196], stage0_23[197]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[5],stage1_25[36],stage1_24[73],stage1_23[75]}
   );
   gpc606_5 gpc477 (
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202], stage0_23[203]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[6],stage1_25[37],stage1_24[74],stage1_23[76]}
   );
   gpc606_5 gpc478 (
      {stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[7],stage1_25[38],stage1_24[75],stage1_23[77]}
   );
   gpc606_5 gpc479 (
      {stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[8],stage1_25[39],stage1_24[76],stage1_23[78]}
   );
   gpc606_5 gpc480 (
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[9],stage1_25[40],stage1_24[77],stage1_23[79]}
   );
   gpc606_5 gpc481 (
      {stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[10],stage1_25[41],stage1_24[78],stage1_23[80]}
   );
   gpc606_5 gpc482 (
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232], stage0_23[233]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[11],stage1_25[42],stage1_24[79],stage1_23[81]}
   );
   gpc606_5 gpc483 (
      {stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238], stage0_23[239]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[12],stage1_25[43],stage1_24[80],stage1_23[82]}
   );
   gpc606_5 gpc484 (
      {stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244], stage0_23[245]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[13],stage1_25[44],stage1_24[81],stage1_23[83]}
   );
   gpc606_5 gpc485 (
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[10],stage1_26[14],stage1_25[45],stage1_24[82]}
   );
   gpc606_5 gpc486 (
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[11],stage1_26[15],stage1_25[46],stage1_24[83]}
   );
   gpc606_5 gpc487 (
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[12],stage1_26[16],stage1_25[47],stage1_24[84]}
   );
   gpc606_5 gpc488 (
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[13],stage1_26[17],stage1_25[48],stage1_24[85]}
   );
   gpc606_5 gpc489 (
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[14],stage1_26[18],stage1_25[49],stage1_24[86]}
   );
   gpc606_5 gpc490 (
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[15],stage1_26[19],stage1_25[50],stage1_24[87]}
   );
   gpc606_5 gpc491 (
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[16],stage1_26[20],stage1_25[51],stage1_24[88]}
   );
   gpc606_5 gpc492 (
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[17],stage1_26[21],stage1_25[52],stage1_24[89]}
   );
   gpc606_5 gpc493 (
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[18],stage1_26[22],stage1_25[53],stage1_24[90]}
   );
   gpc606_5 gpc494 (
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[19],stage1_26[23],stage1_25[54],stage1_24[91]}
   );
   gpc606_5 gpc495 (
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[20],stage1_26[24],stage1_25[55],stage1_24[92]}
   );
   gpc606_5 gpc496 (
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[21],stage1_26[25],stage1_25[56],stage1_24[93]}
   );
   gpc606_5 gpc497 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[12],stage1_27[22],stage1_26[26],stage1_25[57]}
   );
   gpc606_5 gpc498 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[13],stage1_27[23],stage1_26[27],stage1_25[58]}
   );
   gpc606_5 gpc499 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[14],stage1_27[24],stage1_26[28],stage1_25[59]}
   );
   gpc606_5 gpc500 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[15],stage1_27[25],stage1_26[29],stage1_25[60]}
   );
   gpc606_5 gpc501 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[16],stage1_27[26],stage1_26[30],stage1_25[61]}
   );
   gpc606_5 gpc502 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[17],stage1_27[27],stage1_26[31],stage1_25[62]}
   );
   gpc606_5 gpc503 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[18],stage1_27[28],stage1_26[32],stage1_25[63]}
   );
   gpc606_5 gpc504 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[19],stage1_27[29],stage1_26[33],stage1_25[64]}
   );
   gpc606_5 gpc505 (
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[20],stage1_27[30],stage1_26[34],stage1_25[65]}
   );
   gpc606_5 gpc506 (
      {stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[21],stage1_27[31],stage1_26[35],stage1_25[66]}
   );
   gpc606_5 gpc507 (
      {stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[22],stage1_27[32],stage1_26[36],stage1_25[67]}
   );
   gpc606_5 gpc508 (
      {stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[23],stage1_27[33],stage1_26[37],stage1_25[68]}
   );
   gpc606_5 gpc509 (
      {stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[24],stage1_27[34],stage1_26[38],stage1_25[69]}
   );
   gpc606_5 gpc510 (
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[25],stage1_27[35],stage1_26[39],stage1_25[70]}
   );
   gpc606_5 gpc511 (
      {stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[26],stage1_27[36],stage1_26[40],stage1_25[71]}
   );
   gpc606_5 gpc512 (
      {stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[27],stage1_27[37],stage1_26[41],stage1_25[72]}
   );
   gpc606_5 gpc513 (
      {stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[28],stage1_27[38],stage1_26[42],stage1_25[73]}
   );
   gpc606_5 gpc514 (
      {stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[29],stage1_27[39],stage1_26[43],stage1_25[74]}
   );
   gpc606_5 gpc515 (
      {stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[30],stage1_27[40],stage1_26[44],stage1_25[75]}
   );
   gpc606_5 gpc516 (
      {stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[31],stage1_27[41],stage1_26[45],stage1_25[76]}
   );
   gpc606_5 gpc517 (
      {stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[32],stage1_27[42],stage1_26[46],stage1_25[77]}
   );
   gpc606_5 gpc518 (
      {stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[33],stage1_27[43],stage1_26[47],stage1_25[78]}
   );
   gpc606_5 gpc519 (
      {stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[34],stage1_27[44],stage1_26[48],stage1_25[79]}
   );
   gpc606_5 gpc520 (
      {stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[35],stage1_27[45],stage1_26[49],stage1_25[80]}
   );
   gpc606_5 gpc521 (
      {stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[36],stage1_27[46],stage1_26[50],stage1_25[81]}
   );
   gpc606_5 gpc522 (
      {stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[37],stage1_27[47],stage1_26[51],stage1_25[82]}
   );
   gpc606_5 gpc523 (
      {stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[38],stage1_27[48],stage1_26[52],stage1_25[83]}
   );
   gpc606_5 gpc524 (
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[0],stage1_29[27],stage1_28[39],stage1_27[49]}
   );
   gpc606_5 gpc525 (
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[1],stage1_29[28],stage1_28[40],stage1_27[50]}
   );
   gpc606_5 gpc526 (
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[2],stage1_29[29],stage1_28[41],stage1_27[51]}
   );
   gpc606_5 gpc527 (
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[3],stage1_29[30],stage1_28[42],stage1_27[52]}
   );
   gpc606_5 gpc528 (
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[4],stage1_29[31],stage1_28[43],stage1_27[53]}
   );
   gpc606_5 gpc529 (
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[5],stage1_29[32],stage1_28[44],stage1_27[54]}
   );
   gpc606_5 gpc530 (
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[6],stage1_29[33],stage1_28[45],stage1_27[55]}
   );
   gpc606_5 gpc531 (
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[7],stage1_30[7],stage1_29[34],stage1_28[46]}
   );
   gpc606_5 gpc532 (
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[8],stage1_30[8],stage1_29[35],stage1_28[47]}
   );
   gpc606_5 gpc533 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[9],stage1_30[9],stage1_29[36],stage1_28[48]}
   );
   gpc606_5 gpc534 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[10],stage1_30[10],stage1_29[37],stage1_28[49]}
   );
   gpc606_5 gpc535 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[11],stage1_30[11],stage1_29[38],stage1_28[50]}
   );
   gpc606_5 gpc536 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[12],stage1_30[12],stage1_29[39],stage1_28[51]}
   );
   gpc606_5 gpc537 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[13],stage1_30[13],stage1_29[40],stage1_28[52]}
   );
   gpc606_5 gpc538 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[14],stage1_30[14],stage1_29[41],stage1_28[53]}
   );
   gpc606_5 gpc539 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[15],stage1_30[15],stage1_29[42],stage1_28[54]}
   );
   gpc606_5 gpc540 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[16],stage1_30[16],stage1_29[43],stage1_28[55]}
   );
   gpc606_5 gpc541 (
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[17],stage1_30[17],stage1_29[44],stage1_28[56]}
   );
   gpc606_5 gpc542 (
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[18],stage1_30[18],stage1_29[45],stage1_28[57]}
   );
   gpc606_5 gpc543 (
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[19],stage1_30[19],stage1_29[46],stage1_28[58]}
   );
   gpc606_5 gpc544 (
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[20],stage1_30[20],stage1_29[47],stage1_28[59]}
   );
   gpc606_5 gpc545 (
      {stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[21],stage1_30[21],stage1_29[48],stage1_28[60]}
   );
   gpc606_5 gpc546 (
      {stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[22],stage1_30[22],stage1_29[49],stage1_28[61]}
   );
   gpc606_5 gpc547 (
      {stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[23],stage1_30[23],stage1_29[50],stage1_28[62]}
   );
   gpc606_5 gpc548 (
      {stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[24],stage1_30[24],stage1_29[51],stage1_28[63]}
   );
   gpc606_5 gpc549 (
      {stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[25],stage1_30[25],stage1_29[52],stage1_28[64]}
   );
   gpc606_5 gpc550 (
      {stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[26],stage1_30[26],stage1_29[53],stage1_28[65]}
   );
   gpc606_5 gpc551 (
      {stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[27],stage1_30[27],stage1_29[54],stage1_28[66]}
   );
   gpc606_5 gpc552 (
      {stage0_28[126], stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[28],stage1_30[28],stage1_29[55],stage1_28[67]}
   );
   gpc606_5 gpc553 (
      {stage0_28[132], stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[29],stage1_30[29],stage1_29[56],stage1_28[68]}
   );
   gpc606_5 gpc554 (
      {stage0_28[138], stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[30],stage1_30[30],stage1_29[57],stage1_28[69]}
   );
   gpc606_5 gpc555 (
      {stage0_28[144], stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[31],stage1_30[31],stage1_29[58],stage1_28[70]}
   );
   gpc606_5 gpc556 (
      {stage0_28[150], stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[32],stage1_30[32],stage1_29[59],stage1_28[71]}
   );
   gpc606_5 gpc557 (
      {stage0_28[156], stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[33],stage1_30[33],stage1_29[60],stage1_28[72]}
   );
   gpc606_5 gpc558 (
      {stage0_28[162], stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[34],stage1_30[34],stage1_29[61],stage1_28[73]}
   );
   gpc606_5 gpc559 (
      {stage0_28[168], stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[35],stage1_30[35],stage1_29[62],stage1_28[74]}
   );
   gpc606_5 gpc560 (
      {stage0_28[174], stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[36],stage1_30[36],stage1_29[63],stage1_28[75]}
   );
   gpc606_5 gpc561 (
      {stage0_28[180], stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[37],stage1_30[37],stage1_29[64],stage1_28[76]}
   );
   gpc606_5 gpc562 (
      {stage0_28[186], stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[38],stage1_30[38],stage1_29[65],stage1_28[77]}
   );
   gpc606_5 gpc563 (
      {stage0_28[192], stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[39],stage1_30[39],stage1_29[66],stage1_28[78]}
   );
   gpc606_5 gpc564 (
      {stage0_28[198], stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[40],stage1_30[40],stage1_29[67],stage1_28[79]}
   );
   gpc606_5 gpc565 (
      {stage0_28[204], stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[41],stage1_30[41],stage1_29[68],stage1_28[80]}
   );
   gpc606_5 gpc566 (
      {stage0_28[210], stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[42],stage1_30[42],stage1_29[69],stage1_28[81]}
   );
   gpc606_5 gpc567 (
      {stage0_28[216], stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[43],stage1_30[43],stage1_29[70],stage1_28[82]}
   );
   gpc606_5 gpc568 (
      {stage0_28[222], stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[44],stage1_30[44],stage1_29[71],stage1_28[83]}
   );
   gpc606_5 gpc569 (
      {stage0_28[228], stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[45],stage1_30[45],stage1_29[72],stage1_28[84]}
   );
   gpc606_5 gpc570 (
      {stage0_28[234], stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[46],stage1_30[46],stage1_29[73],stage1_28[85]}
   );
   gpc606_5 gpc571 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[40],stage1_31[47],stage1_30[47],stage1_29[74]}
   );
   gpc606_5 gpc572 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[41],stage1_31[48],stage1_30[48],stage1_29[75]}
   );
   gpc606_5 gpc573 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[42],stage1_31[49],stage1_30[49],stage1_29[76]}
   );
   gpc606_5 gpc574 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[43],stage1_31[50],stage1_30[50],stage1_29[77]}
   );
   gpc606_5 gpc575 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[44],stage1_31[51],stage1_30[51],stage1_29[78]}
   );
   gpc606_5 gpc576 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[45],stage1_31[52],stage1_30[52],stage1_29[79]}
   );
   gpc606_5 gpc577 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[46],stage1_31[53],stage1_30[53],stage1_29[80]}
   );
   gpc606_5 gpc578 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[47],stage1_31[54],stage1_30[54],stage1_29[81]}
   );
   gpc606_5 gpc579 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[48],stage1_31[55],stage1_30[55],stage1_29[82]}
   );
   gpc606_5 gpc580 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[49],stage1_31[56],stage1_30[56],stage1_29[83]}
   );
   gpc606_5 gpc581 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[50],stage1_31[57],stage1_30[57],stage1_29[84]}
   );
   gpc606_5 gpc582 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[51],stage1_31[58],stage1_30[58],stage1_29[85]}
   );
   gpc606_5 gpc583 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[52],stage1_31[59],stage1_30[59],stage1_29[86]}
   );
   gpc606_5 gpc584 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[53],stage1_31[60],stage1_30[60],stage1_29[87]}
   );
   gpc606_5 gpc585 (
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[54],stage1_31[61],stage1_30[61],stage1_29[88]}
   );
   gpc606_5 gpc586 (
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[55],stage1_31[62],stage1_30[62],stage1_29[89]}
   );
   gpc606_5 gpc587 (
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[56],stage1_31[63],stage1_30[63],stage1_29[90]}
   );
   gpc606_5 gpc588 (
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[57],stage1_31[64],stage1_30[64],stage1_29[91]}
   );
   gpc606_5 gpc589 (
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[58],stage1_31[65],stage1_30[65],stage1_29[92]}
   );
   gpc606_5 gpc590 (
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[59],stage1_31[66],stage1_30[66],stage1_29[93]}
   );
   gpc606_5 gpc591 (
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[60],stage1_31[67],stage1_30[67],stage1_29[94]}
   );
   gpc606_5 gpc592 (
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[61],stage1_31[68],stage1_30[68],stage1_29[95]}
   );
   gpc606_5 gpc593 (
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[62],stage1_31[69],stage1_30[69],stage1_29[96]}
   );
   gpc606_5 gpc594 (
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[63],stage1_31[70],stage1_30[70],stage1_29[97]}
   );
   gpc606_5 gpc595 (
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[64],stage1_31[71],stage1_30[71],stage1_29[98]}
   );
   gpc606_5 gpc596 (
      {stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[65],stage1_31[72],stage1_30[72],stage1_29[99]}
   );
   gpc606_5 gpc597 (
      {stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[66],stage1_31[73],stage1_30[73],stage1_29[100]}
   );
   gpc606_5 gpc598 (
      {stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[67],stage1_31[74],stage1_30[74],stage1_29[101]}
   );
   gpc606_5 gpc599 (
      {stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[68],stage1_31[75],stage1_30[75],stage1_29[102]}
   );
   gpc606_5 gpc600 (
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[69],stage1_31[76],stage1_30[76],stage1_29[103]}
   );
   gpc606_5 gpc601 (
      {stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[70],stage1_31[77],stage1_30[77],stage1_29[104]}
   );
   gpc606_5 gpc602 (
      {stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[71],stage1_31[78],stage1_30[78],stage1_29[105]}
   );
   gpc606_5 gpc603 (
      {stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[72],stage1_31[79],stage1_30[79],stage1_29[106]}
   );
   gpc606_5 gpc604 (
      {stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[73],stage1_31[80],stage1_30[80],stage1_29[107]}
   );
   gpc1_1 gpc605 (
      {stage0_0[249]},
      {stage1_0[43]}
   );
   gpc1_1 gpc606 (
      {stage0_0[250]},
      {stage1_0[44]}
   );
   gpc1_1 gpc607 (
      {stage0_0[251]},
      {stage1_0[45]}
   );
   gpc1_1 gpc608 (
      {stage0_0[252]},
      {stage1_0[46]}
   );
   gpc1_1 gpc609 (
      {stage0_0[253]},
      {stage1_0[47]}
   );
   gpc1_1 gpc610 (
      {stage0_0[254]},
      {stage1_0[48]}
   );
   gpc1_1 gpc611 (
      {stage0_0[255]},
      {stage1_0[49]}
   );
   gpc1_1 gpc612 (
      {stage0_1[237]},
      {stage1_1[79]}
   );
   gpc1_1 gpc613 (
      {stage0_1[238]},
      {stage1_1[80]}
   );
   gpc1_1 gpc614 (
      {stage0_1[239]},
      {stage1_1[81]}
   );
   gpc1_1 gpc615 (
      {stage0_1[240]},
      {stage1_1[82]}
   );
   gpc1_1 gpc616 (
      {stage0_1[241]},
      {stage1_1[83]}
   );
   gpc1_1 gpc617 (
      {stage0_1[242]},
      {stage1_1[84]}
   );
   gpc1_1 gpc618 (
      {stage0_1[243]},
      {stage1_1[85]}
   );
   gpc1_1 gpc619 (
      {stage0_1[244]},
      {stage1_1[86]}
   );
   gpc1_1 gpc620 (
      {stage0_1[245]},
      {stage1_1[87]}
   );
   gpc1_1 gpc621 (
      {stage0_1[246]},
      {stage1_1[88]}
   );
   gpc1_1 gpc622 (
      {stage0_1[247]},
      {stage1_1[89]}
   );
   gpc1_1 gpc623 (
      {stage0_1[248]},
      {stage1_1[90]}
   );
   gpc1_1 gpc624 (
      {stage0_1[249]},
      {stage1_1[91]}
   );
   gpc1_1 gpc625 (
      {stage0_1[250]},
      {stage1_1[92]}
   );
   gpc1_1 gpc626 (
      {stage0_1[251]},
      {stage1_1[93]}
   );
   gpc1_1 gpc627 (
      {stage0_1[252]},
      {stage1_1[94]}
   );
   gpc1_1 gpc628 (
      {stage0_1[253]},
      {stage1_1[95]}
   );
   gpc1_1 gpc629 (
      {stage0_1[254]},
      {stage1_1[96]}
   );
   gpc1_1 gpc630 (
      {stage0_1[255]},
      {stage1_1[97]}
   );
   gpc1_1 gpc631 (
      {stage0_2[246]},
      {stage1_2[82]}
   );
   gpc1_1 gpc632 (
      {stage0_2[247]},
      {stage1_2[83]}
   );
   gpc1_1 gpc633 (
      {stage0_2[248]},
      {stage1_2[84]}
   );
   gpc1_1 gpc634 (
      {stage0_2[249]},
      {stage1_2[85]}
   );
   gpc1_1 gpc635 (
      {stage0_2[250]},
      {stage1_2[86]}
   );
   gpc1_1 gpc636 (
      {stage0_2[251]},
      {stage1_2[87]}
   );
   gpc1_1 gpc637 (
      {stage0_2[252]},
      {stage1_2[88]}
   );
   gpc1_1 gpc638 (
      {stage0_2[253]},
      {stage1_2[89]}
   );
   gpc1_1 gpc639 (
      {stage0_2[254]},
      {stage1_2[90]}
   );
   gpc1_1 gpc640 (
      {stage0_2[255]},
      {stage1_2[91]}
   );
   gpc1_1 gpc641 (
      {stage0_3[254]},
      {stage1_3[89]}
   );
   gpc1_1 gpc642 (
      {stage0_3[255]},
      {stage1_3[90]}
   );
   gpc1_1 gpc643 (
      {stage0_4[230]},
      {stage1_4[123]}
   );
   gpc1_1 gpc644 (
      {stage0_4[231]},
      {stage1_4[124]}
   );
   gpc1_1 gpc645 (
      {stage0_4[232]},
      {stage1_4[125]}
   );
   gpc1_1 gpc646 (
      {stage0_4[233]},
      {stage1_4[126]}
   );
   gpc1_1 gpc647 (
      {stage0_4[234]},
      {stage1_4[127]}
   );
   gpc1_1 gpc648 (
      {stage0_4[235]},
      {stage1_4[128]}
   );
   gpc1_1 gpc649 (
      {stage0_4[236]},
      {stage1_4[129]}
   );
   gpc1_1 gpc650 (
      {stage0_4[237]},
      {stage1_4[130]}
   );
   gpc1_1 gpc651 (
      {stage0_4[238]},
      {stage1_4[131]}
   );
   gpc1_1 gpc652 (
      {stage0_4[239]},
      {stage1_4[132]}
   );
   gpc1_1 gpc653 (
      {stage0_4[240]},
      {stage1_4[133]}
   );
   gpc1_1 gpc654 (
      {stage0_4[241]},
      {stage1_4[134]}
   );
   gpc1_1 gpc655 (
      {stage0_4[242]},
      {stage1_4[135]}
   );
   gpc1_1 gpc656 (
      {stage0_4[243]},
      {stage1_4[136]}
   );
   gpc1_1 gpc657 (
      {stage0_4[244]},
      {stage1_4[137]}
   );
   gpc1_1 gpc658 (
      {stage0_4[245]},
      {stage1_4[138]}
   );
   gpc1_1 gpc659 (
      {stage0_4[246]},
      {stage1_4[139]}
   );
   gpc1_1 gpc660 (
      {stage0_4[247]},
      {stage1_4[140]}
   );
   gpc1_1 gpc661 (
      {stage0_4[248]},
      {stage1_4[141]}
   );
   gpc1_1 gpc662 (
      {stage0_4[249]},
      {stage1_4[142]}
   );
   gpc1_1 gpc663 (
      {stage0_4[250]},
      {stage1_4[143]}
   );
   gpc1_1 gpc664 (
      {stage0_4[251]},
      {stage1_4[144]}
   );
   gpc1_1 gpc665 (
      {stage0_4[252]},
      {stage1_4[145]}
   );
   gpc1_1 gpc666 (
      {stage0_4[253]},
      {stage1_4[146]}
   );
   gpc1_1 gpc667 (
      {stage0_4[254]},
      {stage1_4[147]}
   );
   gpc1_1 gpc668 (
      {stage0_4[255]},
      {stage1_4[148]}
   );
   gpc1_1 gpc669 (
      {stage0_5[240]},
      {stage1_5[110]}
   );
   gpc1_1 gpc670 (
      {stage0_5[241]},
      {stage1_5[111]}
   );
   gpc1_1 gpc671 (
      {stage0_5[242]},
      {stage1_5[112]}
   );
   gpc1_1 gpc672 (
      {stage0_5[243]},
      {stage1_5[113]}
   );
   gpc1_1 gpc673 (
      {stage0_5[244]},
      {stage1_5[114]}
   );
   gpc1_1 gpc674 (
      {stage0_5[245]},
      {stage1_5[115]}
   );
   gpc1_1 gpc675 (
      {stage0_5[246]},
      {stage1_5[116]}
   );
   gpc1_1 gpc676 (
      {stage0_5[247]},
      {stage1_5[117]}
   );
   gpc1_1 gpc677 (
      {stage0_5[248]},
      {stage1_5[118]}
   );
   gpc1_1 gpc678 (
      {stage0_5[249]},
      {stage1_5[119]}
   );
   gpc1_1 gpc679 (
      {stage0_5[250]},
      {stage1_5[120]}
   );
   gpc1_1 gpc680 (
      {stage0_5[251]},
      {stage1_5[121]}
   );
   gpc1_1 gpc681 (
      {stage0_5[252]},
      {stage1_5[122]}
   );
   gpc1_1 gpc682 (
      {stage0_5[253]},
      {stage1_5[123]}
   );
   gpc1_1 gpc683 (
      {stage0_5[254]},
      {stage1_5[124]}
   );
   gpc1_1 gpc684 (
      {stage0_5[255]},
      {stage1_5[125]}
   );
   gpc1_1 gpc685 (
      {stage0_6[243]},
      {stage1_6[83]}
   );
   gpc1_1 gpc686 (
      {stage0_6[244]},
      {stage1_6[84]}
   );
   gpc1_1 gpc687 (
      {stage0_6[245]},
      {stage1_6[85]}
   );
   gpc1_1 gpc688 (
      {stage0_6[246]},
      {stage1_6[86]}
   );
   gpc1_1 gpc689 (
      {stage0_6[247]},
      {stage1_6[87]}
   );
   gpc1_1 gpc690 (
      {stage0_6[248]},
      {stage1_6[88]}
   );
   gpc1_1 gpc691 (
      {stage0_6[249]},
      {stage1_6[89]}
   );
   gpc1_1 gpc692 (
      {stage0_6[250]},
      {stage1_6[90]}
   );
   gpc1_1 gpc693 (
      {stage0_6[251]},
      {stage1_6[91]}
   );
   gpc1_1 gpc694 (
      {stage0_6[252]},
      {stage1_6[92]}
   );
   gpc1_1 gpc695 (
      {stage0_6[253]},
      {stage1_6[93]}
   );
   gpc1_1 gpc696 (
      {stage0_6[254]},
      {stage1_6[94]}
   );
   gpc1_1 gpc697 (
      {stage0_6[255]},
      {stage1_6[95]}
   );
   gpc1_1 gpc698 (
      {stage0_7[251]},
      {stage1_7[96]}
   );
   gpc1_1 gpc699 (
      {stage0_7[252]},
      {stage1_7[97]}
   );
   gpc1_1 gpc700 (
      {stage0_7[253]},
      {stage1_7[98]}
   );
   gpc1_1 gpc701 (
      {stage0_7[254]},
      {stage1_7[99]}
   );
   gpc1_1 gpc702 (
      {stage0_7[255]},
      {stage1_7[100]}
   );
   gpc1_1 gpc703 (
      {stage0_9[230]},
      {stage1_9[106]}
   );
   gpc1_1 gpc704 (
      {stage0_9[231]},
      {stage1_9[107]}
   );
   gpc1_1 gpc705 (
      {stage0_9[232]},
      {stage1_9[108]}
   );
   gpc1_1 gpc706 (
      {stage0_9[233]},
      {stage1_9[109]}
   );
   gpc1_1 gpc707 (
      {stage0_9[234]},
      {stage1_9[110]}
   );
   gpc1_1 gpc708 (
      {stage0_9[235]},
      {stage1_9[111]}
   );
   gpc1_1 gpc709 (
      {stage0_9[236]},
      {stage1_9[112]}
   );
   gpc1_1 gpc710 (
      {stage0_9[237]},
      {stage1_9[113]}
   );
   gpc1_1 gpc711 (
      {stage0_9[238]},
      {stage1_9[114]}
   );
   gpc1_1 gpc712 (
      {stage0_9[239]},
      {stage1_9[115]}
   );
   gpc1_1 gpc713 (
      {stage0_9[240]},
      {stage1_9[116]}
   );
   gpc1_1 gpc714 (
      {stage0_9[241]},
      {stage1_9[117]}
   );
   gpc1_1 gpc715 (
      {stage0_9[242]},
      {stage1_9[118]}
   );
   gpc1_1 gpc716 (
      {stage0_9[243]},
      {stage1_9[119]}
   );
   gpc1_1 gpc717 (
      {stage0_9[244]},
      {stage1_9[120]}
   );
   gpc1_1 gpc718 (
      {stage0_9[245]},
      {stage1_9[121]}
   );
   gpc1_1 gpc719 (
      {stage0_9[246]},
      {stage1_9[122]}
   );
   gpc1_1 gpc720 (
      {stage0_9[247]},
      {stage1_9[123]}
   );
   gpc1_1 gpc721 (
      {stage0_9[248]},
      {stage1_9[124]}
   );
   gpc1_1 gpc722 (
      {stage0_9[249]},
      {stage1_9[125]}
   );
   gpc1_1 gpc723 (
      {stage0_9[250]},
      {stage1_9[126]}
   );
   gpc1_1 gpc724 (
      {stage0_9[251]},
      {stage1_9[127]}
   );
   gpc1_1 gpc725 (
      {stage0_9[252]},
      {stage1_9[128]}
   );
   gpc1_1 gpc726 (
      {stage0_9[253]},
      {stage1_9[129]}
   );
   gpc1_1 gpc727 (
      {stage0_9[254]},
      {stage1_9[130]}
   );
   gpc1_1 gpc728 (
      {stage0_9[255]},
      {stage1_9[131]}
   );
   gpc1_1 gpc729 (
      {stage0_10[250]},
      {stage1_10[91]}
   );
   gpc1_1 gpc730 (
      {stage0_10[251]},
      {stage1_10[92]}
   );
   gpc1_1 gpc731 (
      {stage0_10[252]},
      {stage1_10[93]}
   );
   gpc1_1 gpc732 (
      {stage0_10[253]},
      {stage1_10[94]}
   );
   gpc1_1 gpc733 (
      {stage0_10[254]},
      {stage1_10[95]}
   );
   gpc1_1 gpc734 (
      {stage0_10[255]},
      {stage1_10[96]}
   );
   gpc1_1 gpc735 (
      {stage0_11[210]},
      {stage1_11[94]}
   );
   gpc1_1 gpc736 (
      {stage0_11[211]},
      {stage1_11[95]}
   );
   gpc1_1 gpc737 (
      {stage0_11[212]},
      {stage1_11[96]}
   );
   gpc1_1 gpc738 (
      {stage0_11[213]},
      {stage1_11[97]}
   );
   gpc1_1 gpc739 (
      {stage0_11[214]},
      {stage1_11[98]}
   );
   gpc1_1 gpc740 (
      {stage0_11[215]},
      {stage1_11[99]}
   );
   gpc1_1 gpc741 (
      {stage0_11[216]},
      {stage1_11[100]}
   );
   gpc1_1 gpc742 (
      {stage0_11[217]},
      {stage1_11[101]}
   );
   gpc1_1 gpc743 (
      {stage0_11[218]},
      {stage1_11[102]}
   );
   gpc1_1 gpc744 (
      {stage0_11[219]},
      {stage1_11[103]}
   );
   gpc1_1 gpc745 (
      {stage0_11[220]},
      {stage1_11[104]}
   );
   gpc1_1 gpc746 (
      {stage0_11[221]},
      {stage1_11[105]}
   );
   gpc1_1 gpc747 (
      {stage0_11[222]},
      {stage1_11[106]}
   );
   gpc1_1 gpc748 (
      {stage0_11[223]},
      {stage1_11[107]}
   );
   gpc1_1 gpc749 (
      {stage0_11[224]},
      {stage1_11[108]}
   );
   gpc1_1 gpc750 (
      {stage0_11[225]},
      {stage1_11[109]}
   );
   gpc1_1 gpc751 (
      {stage0_11[226]},
      {stage1_11[110]}
   );
   gpc1_1 gpc752 (
      {stage0_11[227]},
      {stage1_11[111]}
   );
   gpc1_1 gpc753 (
      {stage0_11[228]},
      {stage1_11[112]}
   );
   gpc1_1 gpc754 (
      {stage0_11[229]},
      {stage1_11[113]}
   );
   gpc1_1 gpc755 (
      {stage0_11[230]},
      {stage1_11[114]}
   );
   gpc1_1 gpc756 (
      {stage0_11[231]},
      {stage1_11[115]}
   );
   gpc1_1 gpc757 (
      {stage0_11[232]},
      {stage1_11[116]}
   );
   gpc1_1 gpc758 (
      {stage0_11[233]},
      {stage1_11[117]}
   );
   gpc1_1 gpc759 (
      {stage0_11[234]},
      {stage1_11[118]}
   );
   gpc1_1 gpc760 (
      {stage0_11[235]},
      {stage1_11[119]}
   );
   gpc1_1 gpc761 (
      {stage0_11[236]},
      {stage1_11[120]}
   );
   gpc1_1 gpc762 (
      {stage0_11[237]},
      {stage1_11[121]}
   );
   gpc1_1 gpc763 (
      {stage0_11[238]},
      {stage1_11[122]}
   );
   gpc1_1 gpc764 (
      {stage0_11[239]},
      {stage1_11[123]}
   );
   gpc1_1 gpc765 (
      {stage0_11[240]},
      {stage1_11[124]}
   );
   gpc1_1 gpc766 (
      {stage0_11[241]},
      {stage1_11[125]}
   );
   gpc1_1 gpc767 (
      {stage0_11[242]},
      {stage1_11[126]}
   );
   gpc1_1 gpc768 (
      {stage0_11[243]},
      {stage1_11[127]}
   );
   gpc1_1 gpc769 (
      {stage0_11[244]},
      {stage1_11[128]}
   );
   gpc1_1 gpc770 (
      {stage0_11[245]},
      {stage1_11[129]}
   );
   gpc1_1 gpc771 (
      {stage0_11[246]},
      {stage1_11[130]}
   );
   gpc1_1 gpc772 (
      {stage0_11[247]},
      {stage1_11[131]}
   );
   gpc1_1 gpc773 (
      {stage0_11[248]},
      {stage1_11[132]}
   );
   gpc1_1 gpc774 (
      {stage0_11[249]},
      {stage1_11[133]}
   );
   gpc1_1 gpc775 (
      {stage0_11[250]},
      {stage1_11[134]}
   );
   gpc1_1 gpc776 (
      {stage0_11[251]},
      {stage1_11[135]}
   );
   gpc1_1 gpc777 (
      {stage0_11[252]},
      {stage1_11[136]}
   );
   gpc1_1 gpc778 (
      {stage0_11[253]},
      {stage1_11[137]}
   );
   gpc1_1 gpc779 (
      {stage0_11[254]},
      {stage1_11[138]}
   );
   gpc1_1 gpc780 (
      {stage0_11[255]},
      {stage1_11[139]}
   );
   gpc1_1 gpc781 (
      {stage0_12[148]},
      {stage1_12[90]}
   );
   gpc1_1 gpc782 (
      {stage0_12[149]},
      {stage1_12[91]}
   );
   gpc1_1 gpc783 (
      {stage0_12[150]},
      {stage1_12[92]}
   );
   gpc1_1 gpc784 (
      {stage0_12[151]},
      {stage1_12[93]}
   );
   gpc1_1 gpc785 (
      {stage0_12[152]},
      {stage1_12[94]}
   );
   gpc1_1 gpc786 (
      {stage0_12[153]},
      {stage1_12[95]}
   );
   gpc1_1 gpc787 (
      {stage0_12[154]},
      {stage1_12[96]}
   );
   gpc1_1 gpc788 (
      {stage0_12[155]},
      {stage1_12[97]}
   );
   gpc1_1 gpc789 (
      {stage0_12[156]},
      {stage1_12[98]}
   );
   gpc1_1 gpc790 (
      {stage0_12[157]},
      {stage1_12[99]}
   );
   gpc1_1 gpc791 (
      {stage0_12[158]},
      {stage1_12[100]}
   );
   gpc1_1 gpc792 (
      {stage0_12[159]},
      {stage1_12[101]}
   );
   gpc1_1 gpc793 (
      {stage0_12[160]},
      {stage1_12[102]}
   );
   gpc1_1 gpc794 (
      {stage0_12[161]},
      {stage1_12[103]}
   );
   gpc1_1 gpc795 (
      {stage0_12[162]},
      {stage1_12[104]}
   );
   gpc1_1 gpc796 (
      {stage0_12[163]},
      {stage1_12[105]}
   );
   gpc1_1 gpc797 (
      {stage0_12[164]},
      {stage1_12[106]}
   );
   gpc1_1 gpc798 (
      {stage0_12[165]},
      {stage1_12[107]}
   );
   gpc1_1 gpc799 (
      {stage0_12[166]},
      {stage1_12[108]}
   );
   gpc1_1 gpc800 (
      {stage0_12[167]},
      {stage1_12[109]}
   );
   gpc1_1 gpc801 (
      {stage0_12[168]},
      {stage1_12[110]}
   );
   gpc1_1 gpc802 (
      {stage0_12[169]},
      {stage1_12[111]}
   );
   gpc1_1 gpc803 (
      {stage0_12[170]},
      {stage1_12[112]}
   );
   gpc1_1 gpc804 (
      {stage0_12[171]},
      {stage1_12[113]}
   );
   gpc1_1 gpc805 (
      {stage0_12[172]},
      {stage1_12[114]}
   );
   gpc1_1 gpc806 (
      {stage0_12[173]},
      {stage1_12[115]}
   );
   gpc1_1 gpc807 (
      {stage0_12[174]},
      {stage1_12[116]}
   );
   gpc1_1 gpc808 (
      {stage0_12[175]},
      {stage1_12[117]}
   );
   gpc1_1 gpc809 (
      {stage0_12[176]},
      {stage1_12[118]}
   );
   gpc1_1 gpc810 (
      {stage0_12[177]},
      {stage1_12[119]}
   );
   gpc1_1 gpc811 (
      {stage0_12[178]},
      {stage1_12[120]}
   );
   gpc1_1 gpc812 (
      {stage0_12[179]},
      {stage1_12[121]}
   );
   gpc1_1 gpc813 (
      {stage0_12[180]},
      {stage1_12[122]}
   );
   gpc1_1 gpc814 (
      {stage0_12[181]},
      {stage1_12[123]}
   );
   gpc1_1 gpc815 (
      {stage0_12[182]},
      {stage1_12[124]}
   );
   gpc1_1 gpc816 (
      {stage0_12[183]},
      {stage1_12[125]}
   );
   gpc1_1 gpc817 (
      {stage0_12[184]},
      {stage1_12[126]}
   );
   gpc1_1 gpc818 (
      {stage0_12[185]},
      {stage1_12[127]}
   );
   gpc1_1 gpc819 (
      {stage0_12[186]},
      {stage1_12[128]}
   );
   gpc1_1 gpc820 (
      {stage0_12[187]},
      {stage1_12[129]}
   );
   gpc1_1 gpc821 (
      {stage0_12[188]},
      {stage1_12[130]}
   );
   gpc1_1 gpc822 (
      {stage0_12[189]},
      {stage1_12[131]}
   );
   gpc1_1 gpc823 (
      {stage0_12[190]},
      {stage1_12[132]}
   );
   gpc1_1 gpc824 (
      {stage0_12[191]},
      {stage1_12[133]}
   );
   gpc1_1 gpc825 (
      {stage0_12[192]},
      {stage1_12[134]}
   );
   gpc1_1 gpc826 (
      {stage0_12[193]},
      {stage1_12[135]}
   );
   gpc1_1 gpc827 (
      {stage0_12[194]},
      {stage1_12[136]}
   );
   gpc1_1 gpc828 (
      {stage0_12[195]},
      {stage1_12[137]}
   );
   gpc1_1 gpc829 (
      {stage0_12[196]},
      {stage1_12[138]}
   );
   gpc1_1 gpc830 (
      {stage0_12[197]},
      {stage1_12[139]}
   );
   gpc1_1 gpc831 (
      {stage0_12[198]},
      {stage1_12[140]}
   );
   gpc1_1 gpc832 (
      {stage0_12[199]},
      {stage1_12[141]}
   );
   gpc1_1 gpc833 (
      {stage0_12[200]},
      {stage1_12[142]}
   );
   gpc1_1 gpc834 (
      {stage0_12[201]},
      {stage1_12[143]}
   );
   gpc1_1 gpc835 (
      {stage0_12[202]},
      {stage1_12[144]}
   );
   gpc1_1 gpc836 (
      {stage0_12[203]},
      {stage1_12[145]}
   );
   gpc1_1 gpc837 (
      {stage0_12[204]},
      {stage1_12[146]}
   );
   gpc1_1 gpc838 (
      {stage0_12[205]},
      {stage1_12[147]}
   );
   gpc1_1 gpc839 (
      {stage0_12[206]},
      {stage1_12[148]}
   );
   gpc1_1 gpc840 (
      {stage0_12[207]},
      {stage1_12[149]}
   );
   gpc1_1 gpc841 (
      {stage0_12[208]},
      {stage1_12[150]}
   );
   gpc1_1 gpc842 (
      {stage0_12[209]},
      {stage1_12[151]}
   );
   gpc1_1 gpc843 (
      {stage0_12[210]},
      {stage1_12[152]}
   );
   gpc1_1 gpc844 (
      {stage0_12[211]},
      {stage1_12[153]}
   );
   gpc1_1 gpc845 (
      {stage0_12[212]},
      {stage1_12[154]}
   );
   gpc1_1 gpc846 (
      {stage0_12[213]},
      {stage1_12[155]}
   );
   gpc1_1 gpc847 (
      {stage0_12[214]},
      {stage1_12[156]}
   );
   gpc1_1 gpc848 (
      {stage0_12[215]},
      {stage1_12[157]}
   );
   gpc1_1 gpc849 (
      {stage0_12[216]},
      {stage1_12[158]}
   );
   gpc1_1 gpc850 (
      {stage0_12[217]},
      {stage1_12[159]}
   );
   gpc1_1 gpc851 (
      {stage0_12[218]},
      {stage1_12[160]}
   );
   gpc1_1 gpc852 (
      {stage0_12[219]},
      {stage1_12[161]}
   );
   gpc1_1 gpc853 (
      {stage0_12[220]},
      {stage1_12[162]}
   );
   gpc1_1 gpc854 (
      {stage0_12[221]},
      {stage1_12[163]}
   );
   gpc1_1 gpc855 (
      {stage0_12[222]},
      {stage1_12[164]}
   );
   gpc1_1 gpc856 (
      {stage0_12[223]},
      {stage1_12[165]}
   );
   gpc1_1 gpc857 (
      {stage0_12[224]},
      {stage1_12[166]}
   );
   gpc1_1 gpc858 (
      {stage0_12[225]},
      {stage1_12[167]}
   );
   gpc1_1 gpc859 (
      {stage0_12[226]},
      {stage1_12[168]}
   );
   gpc1_1 gpc860 (
      {stage0_12[227]},
      {stage1_12[169]}
   );
   gpc1_1 gpc861 (
      {stage0_12[228]},
      {stage1_12[170]}
   );
   gpc1_1 gpc862 (
      {stage0_12[229]},
      {stage1_12[171]}
   );
   gpc1_1 gpc863 (
      {stage0_12[230]},
      {stage1_12[172]}
   );
   gpc1_1 gpc864 (
      {stage0_12[231]},
      {stage1_12[173]}
   );
   gpc1_1 gpc865 (
      {stage0_12[232]},
      {stage1_12[174]}
   );
   gpc1_1 gpc866 (
      {stage0_12[233]},
      {stage1_12[175]}
   );
   gpc1_1 gpc867 (
      {stage0_12[234]},
      {stage1_12[176]}
   );
   gpc1_1 gpc868 (
      {stage0_12[235]},
      {stage1_12[177]}
   );
   gpc1_1 gpc869 (
      {stage0_12[236]},
      {stage1_12[178]}
   );
   gpc1_1 gpc870 (
      {stage0_12[237]},
      {stage1_12[179]}
   );
   gpc1_1 gpc871 (
      {stage0_12[238]},
      {stage1_12[180]}
   );
   gpc1_1 gpc872 (
      {stage0_12[239]},
      {stage1_12[181]}
   );
   gpc1_1 gpc873 (
      {stage0_12[240]},
      {stage1_12[182]}
   );
   gpc1_1 gpc874 (
      {stage0_12[241]},
      {stage1_12[183]}
   );
   gpc1_1 gpc875 (
      {stage0_12[242]},
      {stage1_12[184]}
   );
   gpc1_1 gpc876 (
      {stage0_12[243]},
      {stage1_12[185]}
   );
   gpc1_1 gpc877 (
      {stage0_12[244]},
      {stage1_12[186]}
   );
   gpc1_1 gpc878 (
      {stage0_12[245]},
      {stage1_12[187]}
   );
   gpc1_1 gpc879 (
      {stage0_12[246]},
      {stage1_12[188]}
   );
   gpc1_1 gpc880 (
      {stage0_12[247]},
      {stage1_12[189]}
   );
   gpc1_1 gpc881 (
      {stage0_12[248]},
      {stage1_12[190]}
   );
   gpc1_1 gpc882 (
      {stage0_12[249]},
      {stage1_12[191]}
   );
   gpc1_1 gpc883 (
      {stage0_12[250]},
      {stage1_12[192]}
   );
   gpc1_1 gpc884 (
      {stage0_12[251]},
      {stage1_12[193]}
   );
   gpc1_1 gpc885 (
      {stage0_12[252]},
      {stage1_12[194]}
   );
   gpc1_1 gpc886 (
      {stage0_12[253]},
      {stage1_12[195]}
   );
   gpc1_1 gpc887 (
      {stage0_12[254]},
      {stage1_12[196]}
   );
   gpc1_1 gpc888 (
      {stage0_12[255]},
      {stage1_12[197]}
   );
   gpc1_1 gpc889 (
      {stage0_14[235]},
      {stage1_14[93]}
   );
   gpc1_1 gpc890 (
      {stage0_14[236]},
      {stage1_14[94]}
   );
   gpc1_1 gpc891 (
      {stage0_14[237]},
      {stage1_14[95]}
   );
   gpc1_1 gpc892 (
      {stage0_14[238]},
      {stage1_14[96]}
   );
   gpc1_1 gpc893 (
      {stage0_14[239]},
      {stage1_14[97]}
   );
   gpc1_1 gpc894 (
      {stage0_14[240]},
      {stage1_14[98]}
   );
   gpc1_1 gpc895 (
      {stage0_14[241]},
      {stage1_14[99]}
   );
   gpc1_1 gpc896 (
      {stage0_14[242]},
      {stage1_14[100]}
   );
   gpc1_1 gpc897 (
      {stage0_14[243]},
      {stage1_14[101]}
   );
   gpc1_1 gpc898 (
      {stage0_14[244]},
      {stage1_14[102]}
   );
   gpc1_1 gpc899 (
      {stage0_14[245]},
      {stage1_14[103]}
   );
   gpc1_1 gpc900 (
      {stage0_14[246]},
      {stage1_14[104]}
   );
   gpc1_1 gpc901 (
      {stage0_14[247]},
      {stage1_14[105]}
   );
   gpc1_1 gpc902 (
      {stage0_14[248]},
      {stage1_14[106]}
   );
   gpc1_1 gpc903 (
      {stage0_14[249]},
      {stage1_14[107]}
   );
   gpc1_1 gpc904 (
      {stage0_14[250]},
      {stage1_14[108]}
   );
   gpc1_1 gpc905 (
      {stage0_14[251]},
      {stage1_14[109]}
   );
   gpc1_1 gpc906 (
      {stage0_14[252]},
      {stage1_14[110]}
   );
   gpc1_1 gpc907 (
      {stage0_14[253]},
      {stage1_14[111]}
   );
   gpc1_1 gpc908 (
      {stage0_14[254]},
      {stage1_14[112]}
   );
   gpc1_1 gpc909 (
      {stage0_14[255]},
      {stage1_14[113]}
   );
   gpc1_1 gpc910 (
      {stage0_15[254]},
      {stage1_15[91]}
   );
   gpc1_1 gpc911 (
      {stage0_15[255]},
      {stage1_15[92]}
   );
   gpc1_1 gpc912 (
      {stage0_17[252]},
      {stage1_17[123]}
   );
   gpc1_1 gpc913 (
      {stage0_17[253]},
      {stage1_17[124]}
   );
   gpc1_1 gpc914 (
      {stage0_17[254]},
      {stage1_17[125]}
   );
   gpc1_1 gpc915 (
      {stage0_17[255]},
      {stage1_17[126]}
   );
   gpc1_1 gpc916 (
      {stage0_18[204]},
      {stage1_18[99]}
   );
   gpc1_1 gpc917 (
      {stage0_18[205]},
      {stage1_18[100]}
   );
   gpc1_1 gpc918 (
      {stage0_18[206]},
      {stage1_18[101]}
   );
   gpc1_1 gpc919 (
      {stage0_18[207]},
      {stage1_18[102]}
   );
   gpc1_1 gpc920 (
      {stage0_18[208]},
      {stage1_18[103]}
   );
   gpc1_1 gpc921 (
      {stage0_18[209]},
      {stage1_18[104]}
   );
   gpc1_1 gpc922 (
      {stage0_18[210]},
      {stage1_18[105]}
   );
   gpc1_1 gpc923 (
      {stage0_18[211]},
      {stage1_18[106]}
   );
   gpc1_1 gpc924 (
      {stage0_18[212]},
      {stage1_18[107]}
   );
   gpc1_1 gpc925 (
      {stage0_18[213]},
      {stage1_18[108]}
   );
   gpc1_1 gpc926 (
      {stage0_18[214]},
      {stage1_18[109]}
   );
   gpc1_1 gpc927 (
      {stage0_18[215]},
      {stage1_18[110]}
   );
   gpc1_1 gpc928 (
      {stage0_18[216]},
      {stage1_18[111]}
   );
   gpc1_1 gpc929 (
      {stage0_18[217]},
      {stage1_18[112]}
   );
   gpc1_1 gpc930 (
      {stage0_18[218]},
      {stage1_18[113]}
   );
   gpc1_1 gpc931 (
      {stage0_18[219]},
      {stage1_18[114]}
   );
   gpc1_1 gpc932 (
      {stage0_18[220]},
      {stage1_18[115]}
   );
   gpc1_1 gpc933 (
      {stage0_18[221]},
      {stage1_18[116]}
   );
   gpc1_1 gpc934 (
      {stage0_18[222]},
      {stage1_18[117]}
   );
   gpc1_1 gpc935 (
      {stage0_18[223]},
      {stage1_18[118]}
   );
   gpc1_1 gpc936 (
      {stage0_18[224]},
      {stage1_18[119]}
   );
   gpc1_1 gpc937 (
      {stage0_18[225]},
      {stage1_18[120]}
   );
   gpc1_1 gpc938 (
      {stage0_18[226]},
      {stage1_18[121]}
   );
   gpc1_1 gpc939 (
      {stage0_18[227]},
      {stage1_18[122]}
   );
   gpc1_1 gpc940 (
      {stage0_18[228]},
      {stage1_18[123]}
   );
   gpc1_1 gpc941 (
      {stage0_18[229]},
      {stage1_18[124]}
   );
   gpc1_1 gpc942 (
      {stage0_18[230]},
      {stage1_18[125]}
   );
   gpc1_1 gpc943 (
      {stage0_18[231]},
      {stage1_18[126]}
   );
   gpc1_1 gpc944 (
      {stage0_18[232]},
      {stage1_18[127]}
   );
   gpc1_1 gpc945 (
      {stage0_18[233]},
      {stage1_18[128]}
   );
   gpc1_1 gpc946 (
      {stage0_18[234]},
      {stage1_18[129]}
   );
   gpc1_1 gpc947 (
      {stage0_18[235]},
      {stage1_18[130]}
   );
   gpc1_1 gpc948 (
      {stage0_18[236]},
      {stage1_18[131]}
   );
   gpc1_1 gpc949 (
      {stage0_18[237]},
      {stage1_18[132]}
   );
   gpc1_1 gpc950 (
      {stage0_18[238]},
      {stage1_18[133]}
   );
   gpc1_1 gpc951 (
      {stage0_18[239]},
      {stage1_18[134]}
   );
   gpc1_1 gpc952 (
      {stage0_18[240]},
      {stage1_18[135]}
   );
   gpc1_1 gpc953 (
      {stage0_18[241]},
      {stage1_18[136]}
   );
   gpc1_1 gpc954 (
      {stage0_18[242]},
      {stage1_18[137]}
   );
   gpc1_1 gpc955 (
      {stage0_18[243]},
      {stage1_18[138]}
   );
   gpc1_1 gpc956 (
      {stage0_18[244]},
      {stage1_18[139]}
   );
   gpc1_1 gpc957 (
      {stage0_18[245]},
      {stage1_18[140]}
   );
   gpc1_1 gpc958 (
      {stage0_18[246]},
      {stage1_18[141]}
   );
   gpc1_1 gpc959 (
      {stage0_18[247]},
      {stage1_18[142]}
   );
   gpc1_1 gpc960 (
      {stage0_18[248]},
      {stage1_18[143]}
   );
   gpc1_1 gpc961 (
      {stage0_18[249]},
      {stage1_18[144]}
   );
   gpc1_1 gpc962 (
      {stage0_18[250]},
      {stage1_18[145]}
   );
   gpc1_1 gpc963 (
      {stage0_18[251]},
      {stage1_18[146]}
   );
   gpc1_1 gpc964 (
      {stage0_18[252]},
      {stage1_18[147]}
   );
   gpc1_1 gpc965 (
      {stage0_18[253]},
      {stage1_18[148]}
   );
   gpc1_1 gpc966 (
      {stage0_18[254]},
      {stage1_18[149]}
   );
   gpc1_1 gpc967 (
      {stage0_18[255]},
      {stage1_18[150]}
   );
   gpc1_1 gpc968 (
      {stage0_19[240]},
      {stage1_19[78]}
   );
   gpc1_1 gpc969 (
      {stage0_19[241]},
      {stage1_19[79]}
   );
   gpc1_1 gpc970 (
      {stage0_19[242]},
      {stage1_19[80]}
   );
   gpc1_1 gpc971 (
      {stage0_19[243]},
      {stage1_19[81]}
   );
   gpc1_1 gpc972 (
      {stage0_19[244]},
      {stage1_19[82]}
   );
   gpc1_1 gpc973 (
      {stage0_19[245]},
      {stage1_19[83]}
   );
   gpc1_1 gpc974 (
      {stage0_19[246]},
      {stage1_19[84]}
   );
   gpc1_1 gpc975 (
      {stage0_19[247]},
      {stage1_19[85]}
   );
   gpc1_1 gpc976 (
      {stage0_19[248]},
      {stage1_19[86]}
   );
   gpc1_1 gpc977 (
      {stage0_19[249]},
      {stage1_19[87]}
   );
   gpc1_1 gpc978 (
      {stage0_19[250]},
      {stage1_19[88]}
   );
   gpc1_1 gpc979 (
      {stage0_19[251]},
      {stage1_19[89]}
   );
   gpc1_1 gpc980 (
      {stage0_19[252]},
      {stage1_19[90]}
   );
   gpc1_1 gpc981 (
      {stage0_19[253]},
      {stage1_19[91]}
   );
   gpc1_1 gpc982 (
      {stage0_19[254]},
      {stage1_19[92]}
   );
   gpc1_1 gpc983 (
      {stage0_19[255]},
      {stage1_19[93]}
   );
   gpc1_1 gpc984 (
      {stage0_20[245]},
      {stage1_20[105]}
   );
   gpc1_1 gpc985 (
      {stage0_20[246]},
      {stage1_20[106]}
   );
   gpc1_1 gpc986 (
      {stage0_20[247]},
      {stage1_20[107]}
   );
   gpc1_1 gpc987 (
      {stage0_20[248]},
      {stage1_20[108]}
   );
   gpc1_1 gpc988 (
      {stage0_20[249]},
      {stage1_20[109]}
   );
   gpc1_1 gpc989 (
      {stage0_20[250]},
      {stage1_20[110]}
   );
   gpc1_1 gpc990 (
      {stage0_20[251]},
      {stage1_20[111]}
   );
   gpc1_1 gpc991 (
      {stage0_20[252]},
      {stage1_20[112]}
   );
   gpc1_1 gpc992 (
      {stage0_20[253]},
      {stage1_20[113]}
   );
   gpc1_1 gpc993 (
      {stage0_20[254]},
      {stage1_20[114]}
   );
   gpc1_1 gpc994 (
      {stage0_20[255]},
      {stage1_20[115]}
   );
   gpc1_1 gpc995 (
      {stage0_21[235]},
      {stage1_21[118]}
   );
   gpc1_1 gpc996 (
      {stage0_21[236]},
      {stage1_21[119]}
   );
   gpc1_1 gpc997 (
      {stage0_21[237]},
      {stage1_21[120]}
   );
   gpc1_1 gpc998 (
      {stage0_21[238]},
      {stage1_21[121]}
   );
   gpc1_1 gpc999 (
      {stage0_21[239]},
      {stage1_21[122]}
   );
   gpc1_1 gpc1000 (
      {stage0_21[240]},
      {stage1_21[123]}
   );
   gpc1_1 gpc1001 (
      {stage0_21[241]},
      {stage1_21[124]}
   );
   gpc1_1 gpc1002 (
      {stage0_21[242]},
      {stage1_21[125]}
   );
   gpc1_1 gpc1003 (
      {stage0_21[243]},
      {stage1_21[126]}
   );
   gpc1_1 gpc1004 (
      {stage0_21[244]},
      {stage1_21[127]}
   );
   gpc1_1 gpc1005 (
      {stage0_21[245]},
      {stage1_21[128]}
   );
   gpc1_1 gpc1006 (
      {stage0_21[246]},
      {stage1_21[129]}
   );
   gpc1_1 gpc1007 (
      {stage0_21[247]},
      {stage1_21[130]}
   );
   gpc1_1 gpc1008 (
      {stage0_21[248]},
      {stage1_21[131]}
   );
   gpc1_1 gpc1009 (
      {stage0_21[249]},
      {stage1_21[132]}
   );
   gpc1_1 gpc1010 (
      {stage0_21[250]},
      {stage1_21[133]}
   );
   gpc1_1 gpc1011 (
      {stage0_21[251]},
      {stage1_21[134]}
   );
   gpc1_1 gpc1012 (
      {stage0_21[252]},
      {stage1_21[135]}
   );
   gpc1_1 gpc1013 (
      {stage0_21[253]},
      {stage1_21[136]}
   );
   gpc1_1 gpc1014 (
      {stage0_21[254]},
      {stage1_21[137]}
   );
   gpc1_1 gpc1015 (
      {stage0_21[255]},
      {stage1_21[138]}
   );
   gpc1_1 gpc1016 (
      {stage0_22[246]},
      {stage1_22[84]}
   );
   gpc1_1 gpc1017 (
      {stage0_22[247]},
      {stage1_22[85]}
   );
   gpc1_1 gpc1018 (
      {stage0_22[248]},
      {stage1_22[86]}
   );
   gpc1_1 gpc1019 (
      {stage0_22[249]},
      {stage1_22[87]}
   );
   gpc1_1 gpc1020 (
      {stage0_22[250]},
      {stage1_22[88]}
   );
   gpc1_1 gpc1021 (
      {stage0_22[251]},
      {stage1_22[89]}
   );
   gpc1_1 gpc1022 (
      {stage0_22[252]},
      {stage1_22[90]}
   );
   gpc1_1 gpc1023 (
      {stage0_22[253]},
      {stage1_22[91]}
   );
   gpc1_1 gpc1024 (
      {stage0_22[254]},
      {stage1_22[92]}
   );
   gpc1_1 gpc1025 (
      {stage0_22[255]},
      {stage1_22[93]}
   );
   gpc1_1 gpc1026 (
      {stage0_23[246]},
      {stage1_23[84]}
   );
   gpc1_1 gpc1027 (
      {stage0_23[247]},
      {stage1_23[85]}
   );
   gpc1_1 gpc1028 (
      {stage0_23[248]},
      {stage1_23[86]}
   );
   gpc1_1 gpc1029 (
      {stage0_23[249]},
      {stage1_23[87]}
   );
   gpc1_1 gpc1030 (
      {stage0_23[250]},
      {stage1_23[88]}
   );
   gpc1_1 gpc1031 (
      {stage0_23[251]},
      {stage1_23[89]}
   );
   gpc1_1 gpc1032 (
      {stage0_23[252]},
      {stage1_23[90]}
   );
   gpc1_1 gpc1033 (
      {stage0_23[253]},
      {stage1_23[91]}
   );
   gpc1_1 gpc1034 (
      {stage0_23[254]},
      {stage1_23[92]}
   );
   gpc1_1 gpc1035 (
      {stage0_23[255]},
      {stage1_23[93]}
   );
   gpc1_1 gpc1036 (
      {stage0_24[96]},
      {stage1_24[94]}
   );
   gpc1_1 gpc1037 (
      {stage0_24[97]},
      {stage1_24[95]}
   );
   gpc1_1 gpc1038 (
      {stage0_24[98]},
      {stage1_24[96]}
   );
   gpc1_1 gpc1039 (
      {stage0_24[99]},
      {stage1_24[97]}
   );
   gpc1_1 gpc1040 (
      {stage0_24[100]},
      {stage1_24[98]}
   );
   gpc1_1 gpc1041 (
      {stage0_24[101]},
      {stage1_24[99]}
   );
   gpc1_1 gpc1042 (
      {stage0_24[102]},
      {stage1_24[100]}
   );
   gpc1_1 gpc1043 (
      {stage0_24[103]},
      {stage1_24[101]}
   );
   gpc1_1 gpc1044 (
      {stage0_24[104]},
      {stage1_24[102]}
   );
   gpc1_1 gpc1045 (
      {stage0_24[105]},
      {stage1_24[103]}
   );
   gpc1_1 gpc1046 (
      {stage0_24[106]},
      {stage1_24[104]}
   );
   gpc1_1 gpc1047 (
      {stage0_24[107]},
      {stage1_24[105]}
   );
   gpc1_1 gpc1048 (
      {stage0_24[108]},
      {stage1_24[106]}
   );
   gpc1_1 gpc1049 (
      {stage0_24[109]},
      {stage1_24[107]}
   );
   gpc1_1 gpc1050 (
      {stage0_24[110]},
      {stage1_24[108]}
   );
   gpc1_1 gpc1051 (
      {stage0_24[111]},
      {stage1_24[109]}
   );
   gpc1_1 gpc1052 (
      {stage0_24[112]},
      {stage1_24[110]}
   );
   gpc1_1 gpc1053 (
      {stage0_24[113]},
      {stage1_24[111]}
   );
   gpc1_1 gpc1054 (
      {stage0_24[114]},
      {stage1_24[112]}
   );
   gpc1_1 gpc1055 (
      {stage0_24[115]},
      {stage1_24[113]}
   );
   gpc1_1 gpc1056 (
      {stage0_24[116]},
      {stage1_24[114]}
   );
   gpc1_1 gpc1057 (
      {stage0_24[117]},
      {stage1_24[115]}
   );
   gpc1_1 gpc1058 (
      {stage0_24[118]},
      {stage1_24[116]}
   );
   gpc1_1 gpc1059 (
      {stage0_24[119]},
      {stage1_24[117]}
   );
   gpc1_1 gpc1060 (
      {stage0_24[120]},
      {stage1_24[118]}
   );
   gpc1_1 gpc1061 (
      {stage0_24[121]},
      {stage1_24[119]}
   );
   gpc1_1 gpc1062 (
      {stage0_24[122]},
      {stage1_24[120]}
   );
   gpc1_1 gpc1063 (
      {stage0_24[123]},
      {stage1_24[121]}
   );
   gpc1_1 gpc1064 (
      {stage0_24[124]},
      {stage1_24[122]}
   );
   gpc1_1 gpc1065 (
      {stage0_24[125]},
      {stage1_24[123]}
   );
   gpc1_1 gpc1066 (
      {stage0_24[126]},
      {stage1_24[124]}
   );
   gpc1_1 gpc1067 (
      {stage0_24[127]},
      {stage1_24[125]}
   );
   gpc1_1 gpc1068 (
      {stage0_24[128]},
      {stage1_24[126]}
   );
   gpc1_1 gpc1069 (
      {stage0_24[129]},
      {stage1_24[127]}
   );
   gpc1_1 gpc1070 (
      {stage0_24[130]},
      {stage1_24[128]}
   );
   gpc1_1 gpc1071 (
      {stage0_24[131]},
      {stage1_24[129]}
   );
   gpc1_1 gpc1072 (
      {stage0_24[132]},
      {stage1_24[130]}
   );
   gpc1_1 gpc1073 (
      {stage0_24[133]},
      {stage1_24[131]}
   );
   gpc1_1 gpc1074 (
      {stage0_24[134]},
      {stage1_24[132]}
   );
   gpc1_1 gpc1075 (
      {stage0_24[135]},
      {stage1_24[133]}
   );
   gpc1_1 gpc1076 (
      {stage0_24[136]},
      {stage1_24[134]}
   );
   gpc1_1 gpc1077 (
      {stage0_24[137]},
      {stage1_24[135]}
   );
   gpc1_1 gpc1078 (
      {stage0_24[138]},
      {stage1_24[136]}
   );
   gpc1_1 gpc1079 (
      {stage0_24[139]},
      {stage1_24[137]}
   );
   gpc1_1 gpc1080 (
      {stage0_24[140]},
      {stage1_24[138]}
   );
   gpc1_1 gpc1081 (
      {stage0_24[141]},
      {stage1_24[139]}
   );
   gpc1_1 gpc1082 (
      {stage0_24[142]},
      {stage1_24[140]}
   );
   gpc1_1 gpc1083 (
      {stage0_24[143]},
      {stage1_24[141]}
   );
   gpc1_1 gpc1084 (
      {stage0_24[144]},
      {stage1_24[142]}
   );
   gpc1_1 gpc1085 (
      {stage0_24[145]},
      {stage1_24[143]}
   );
   gpc1_1 gpc1086 (
      {stage0_24[146]},
      {stage1_24[144]}
   );
   gpc1_1 gpc1087 (
      {stage0_24[147]},
      {stage1_24[145]}
   );
   gpc1_1 gpc1088 (
      {stage0_24[148]},
      {stage1_24[146]}
   );
   gpc1_1 gpc1089 (
      {stage0_24[149]},
      {stage1_24[147]}
   );
   gpc1_1 gpc1090 (
      {stage0_24[150]},
      {stage1_24[148]}
   );
   gpc1_1 gpc1091 (
      {stage0_24[151]},
      {stage1_24[149]}
   );
   gpc1_1 gpc1092 (
      {stage0_24[152]},
      {stage1_24[150]}
   );
   gpc1_1 gpc1093 (
      {stage0_24[153]},
      {stage1_24[151]}
   );
   gpc1_1 gpc1094 (
      {stage0_24[154]},
      {stage1_24[152]}
   );
   gpc1_1 gpc1095 (
      {stage0_24[155]},
      {stage1_24[153]}
   );
   gpc1_1 gpc1096 (
      {stage0_24[156]},
      {stage1_24[154]}
   );
   gpc1_1 gpc1097 (
      {stage0_24[157]},
      {stage1_24[155]}
   );
   gpc1_1 gpc1098 (
      {stage0_24[158]},
      {stage1_24[156]}
   );
   gpc1_1 gpc1099 (
      {stage0_24[159]},
      {stage1_24[157]}
   );
   gpc1_1 gpc1100 (
      {stage0_24[160]},
      {stage1_24[158]}
   );
   gpc1_1 gpc1101 (
      {stage0_24[161]},
      {stage1_24[159]}
   );
   gpc1_1 gpc1102 (
      {stage0_24[162]},
      {stage1_24[160]}
   );
   gpc1_1 gpc1103 (
      {stage0_24[163]},
      {stage1_24[161]}
   );
   gpc1_1 gpc1104 (
      {stage0_24[164]},
      {stage1_24[162]}
   );
   gpc1_1 gpc1105 (
      {stage0_24[165]},
      {stage1_24[163]}
   );
   gpc1_1 gpc1106 (
      {stage0_24[166]},
      {stage1_24[164]}
   );
   gpc1_1 gpc1107 (
      {stage0_24[167]},
      {stage1_24[165]}
   );
   gpc1_1 gpc1108 (
      {stage0_24[168]},
      {stage1_24[166]}
   );
   gpc1_1 gpc1109 (
      {stage0_24[169]},
      {stage1_24[167]}
   );
   gpc1_1 gpc1110 (
      {stage0_24[170]},
      {stage1_24[168]}
   );
   gpc1_1 gpc1111 (
      {stage0_24[171]},
      {stage1_24[169]}
   );
   gpc1_1 gpc1112 (
      {stage0_24[172]},
      {stage1_24[170]}
   );
   gpc1_1 gpc1113 (
      {stage0_24[173]},
      {stage1_24[171]}
   );
   gpc1_1 gpc1114 (
      {stage0_24[174]},
      {stage1_24[172]}
   );
   gpc1_1 gpc1115 (
      {stage0_24[175]},
      {stage1_24[173]}
   );
   gpc1_1 gpc1116 (
      {stage0_24[176]},
      {stage1_24[174]}
   );
   gpc1_1 gpc1117 (
      {stage0_24[177]},
      {stage1_24[175]}
   );
   gpc1_1 gpc1118 (
      {stage0_24[178]},
      {stage1_24[176]}
   );
   gpc1_1 gpc1119 (
      {stage0_24[179]},
      {stage1_24[177]}
   );
   gpc1_1 gpc1120 (
      {stage0_24[180]},
      {stage1_24[178]}
   );
   gpc1_1 gpc1121 (
      {stage0_24[181]},
      {stage1_24[179]}
   );
   gpc1_1 gpc1122 (
      {stage0_24[182]},
      {stage1_24[180]}
   );
   gpc1_1 gpc1123 (
      {stage0_24[183]},
      {stage1_24[181]}
   );
   gpc1_1 gpc1124 (
      {stage0_24[184]},
      {stage1_24[182]}
   );
   gpc1_1 gpc1125 (
      {stage0_24[185]},
      {stage1_24[183]}
   );
   gpc1_1 gpc1126 (
      {stage0_24[186]},
      {stage1_24[184]}
   );
   gpc1_1 gpc1127 (
      {stage0_24[187]},
      {stage1_24[185]}
   );
   gpc1_1 gpc1128 (
      {stage0_24[188]},
      {stage1_24[186]}
   );
   gpc1_1 gpc1129 (
      {stage0_24[189]},
      {stage1_24[187]}
   );
   gpc1_1 gpc1130 (
      {stage0_24[190]},
      {stage1_24[188]}
   );
   gpc1_1 gpc1131 (
      {stage0_24[191]},
      {stage1_24[189]}
   );
   gpc1_1 gpc1132 (
      {stage0_24[192]},
      {stage1_24[190]}
   );
   gpc1_1 gpc1133 (
      {stage0_24[193]},
      {stage1_24[191]}
   );
   gpc1_1 gpc1134 (
      {stage0_24[194]},
      {stage1_24[192]}
   );
   gpc1_1 gpc1135 (
      {stage0_24[195]},
      {stage1_24[193]}
   );
   gpc1_1 gpc1136 (
      {stage0_24[196]},
      {stage1_24[194]}
   );
   gpc1_1 gpc1137 (
      {stage0_24[197]},
      {stage1_24[195]}
   );
   gpc1_1 gpc1138 (
      {stage0_24[198]},
      {stage1_24[196]}
   );
   gpc1_1 gpc1139 (
      {stage0_24[199]},
      {stage1_24[197]}
   );
   gpc1_1 gpc1140 (
      {stage0_24[200]},
      {stage1_24[198]}
   );
   gpc1_1 gpc1141 (
      {stage0_24[201]},
      {stage1_24[199]}
   );
   gpc1_1 gpc1142 (
      {stage0_24[202]},
      {stage1_24[200]}
   );
   gpc1_1 gpc1143 (
      {stage0_24[203]},
      {stage1_24[201]}
   );
   gpc1_1 gpc1144 (
      {stage0_24[204]},
      {stage1_24[202]}
   );
   gpc1_1 gpc1145 (
      {stage0_24[205]},
      {stage1_24[203]}
   );
   gpc1_1 gpc1146 (
      {stage0_24[206]},
      {stage1_24[204]}
   );
   gpc1_1 gpc1147 (
      {stage0_24[207]},
      {stage1_24[205]}
   );
   gpc1_1 gpc1148 (
      {stage0_24[208]},
      {stage1_24[206]}
   );
   gpc1_1 gpc1149 (
      {stage0_24[209]},
      {stage1_24[207]}
   );
   gpc1_1 gpc1150 (
      {stage0_24[210]},
      {stage1_24[208]}
   );
   gpc1_1 gpc1151 (
      {stage0_24[211]},
      {stage1_24[209]}
   );
   gpc1_1 gpc1152 (
      {stage0_24[212]},
      {stage1_24[210]}
   );
   gpc1_1 gpc1153 (
      {stage0_24[213]},
      {stage1_24[211]}
   );
   gpc1_1 gpc1154 (
      {stage0_24[214]},
      {stage1_24[212]}
   );
   gpc1_1 gpc1155 (
      {stage0_24[215]},
      {stage1_24[213]}
   );
   gpc1_1 gpc1156 (
      {stage0_24[216]},
      {stage1_24[214]}
   );
   gpc1_1 gpc1157 (
      {stage0_24[217]},
      {stage1_24[215]}
   );
   gpc1_1 gpc1158 (
      {stage0_24[218]},
      {stage1_24[216]}
   );
   gpc1_1 gpc1159 (
      {stage0_24[219]},
      {stage1_24[217]}
   );
   gpc1_1 gpc1160 (
      {stage0_24[220]},
      {stage1_24[218]}
   );
   gpc1_1 gpc1161 (
      {stage0_24[221]},
      {stage1_24[219]}
   );
   gpc1_1 gpc1162 (
      {stage0_24[222]},
      {stage1_24[220]}
   );
   gpc1_1 gpc1163 (
      {stage0_24[223]},
      {stage1_24[221]}
   );
   gpc1_1 gpc1164 (
      {stage0_24[224]},
      {stage1_24[222]}
   );
   gpc1_1 gpc1165 (
      {stage0_24[225]},
      {stage1_24[223]}
   );
   gpc1_1 gpc1166 (
      {stage0_24[226]},
      {stage1_24[224]}
   );
   gpc1_1 gpc1167 (
      {stage0_24[227]},
      {stage1_24[225]}
   );
   gpc1_1 gpc1168 (
      {stage0_24[228]},
      {stage1_24[226]}
   );
   gpc1_1 gpc1169 (
      {stage0_24[229]},
      {stage1_24[227]}
   );
   gpc1_1 gpc1170 (
      {stage0_24[230]},
      {stage1_24[228]}
   );
   gpc1_1 gpc1171 (
      {stage0_24[231]},
      {stage1_24[229]}
   );
   gpc1_1 gpc1172 (
      {stage0_24[232]},
      {stage1_24[230]}
   );
   gpc1_1 gpc1173 (
      {stage0_24[233]},
      {stage1_24[231]}
   );
   gpc1_1 gpc1174 (
      {stage0_24[234]},
      {stage1_24[232]}
   );
   gpc1_1 gpc1175 (
      {stage0_24[235]},
      {stage1_24[233]}
   );
   gpc1_1 gpc1176 (
      {stage0_24[236]},
      {stage1_24[234]}
   );
   gpc1_1 gpc1177 (
      {stage0_24[237]},
      {stage1_24[235]}
   );
   gpc1_1 gpc1178 (
      {stage0_24[238]},
      {stage1_24[236]}
   );
   gpc1_1 gpc1179 (
      {stage0_24[239]},
      {stage1_24[237]}
   );
   gpc1_1 gpc1180 (
      {stage0_24[240]},
      {stage1_24[238]}
   );
   gpc1_1 gpc1181 (
      {stage0_24[241]},
      {stage1_24[239]}
   );
   gpc1_1 gpc1182 (
      {stage0_24[242]},
      {stage1_24[240]}
   );
   gpc1_1 gpc1183 (
      {stage0_24[243]},
      {stage1_24[241]}
   );
   gpc1_1 gpc1184 (
      {stage0_24[244]},
      {stage1_24[242]}
   );
   gpc1_1 gpc1185 (
      {stage0_24[245]},
      {stage1_24[243]}
   );
   gpc1_1 gpc1186 (
      {stage0_24[246]},
      {stage1_24[244]}
   );
   gpc1_1 gpc1187 (
      {stage0_24[247]},
      {stage1_24[245]}
   );
   gpc1_1 gpc1188 (
      {stage0_24[248]},
      {stage1_24[246]}
   );
   gpc1_1 gpc1189 (
      {stage0_24[249]},
      {stage1_24[247]}
   );
   gpc1_1 gpc1190 (
      {stage0_24[250]},
      {stage1_24[248]}
   );
   gpc1_1 gpc1191 (
      {stage0_24[251]},
      {stage1_24[249]}
   );
   gpc1_1 gpc1192 (
      {stage0_24[252]},
      {stage1_24[250]}
   );
   gpc1_1 gpc1193 (
      {stage0_24[253]},
      {stage1_24[251]}
   );
   gpc1_1 gpc1194 (
      {stage0_24[254]},
      {stage1_24[252]}
   );
   gpc1_1 gpc1195 (
      {stage0_24[255]},
      {stage1_24[253]}
   );
   gpc1_1 gpc1196 (
      {stage0_25[222]},
      {stage1_25[84]}
   );
   gpc1_1 gpc1197 (
      {stage0_25[223]},
      {stage1_25[85]}
   );
   gpc1_1 gpc1198 (
      {stage0_25[224]},
      {stage1_25[86]}
   );
   gpc1_1 gpc1199 (
      {stage0_25[225]},
      {stage1_25[87]}
   );
   gpc1_1 gpc1200 (
      {stage0_25[226]},
      {stage1_25[88]}
   );
   gpc1_1 gpc1201 (
      {stage0_25[227]},
      {stage1_25[89]}
   );
   gpc1_1 gpc1202 (
      {stage0_25[228]},
      {stage1_25[90]}
   );
   gpc1_1 gpc1203 (
      {stage0_25[229]},
      {stage1_25[91]}
   );
   gpc1_1 gpc1204 (
      {stage0_25[230]},
      {stage1_25[92]}
   );
   gpc1_1 gpc1205 (
      {stage0_25[231]},
      {stage1_25[93]}
   );
   gpc1_1 gpc1206 (
      {stage0_25[232]},
      {stage1_25[94]}
   );
   gpc1_1 gpc1207 (
      {stage0_25[233]},
      {stage1_25[95]}
   );
   gpc1_1 gpc1208 (
      {stage0_25[234]},
      {stage1_25[96]}
   );
   gpc1_1 gpc1209 (
      {stage0_25[235]},
      {stage1_25[97]}
   );
   gpc1_1 gpc1210 (
      {stage0_25[236]},
      {stage1_25[98]}
   );
   gpc1_1 gpc1211 (
      {stage0_25[237]},
      {stage1_25[99]}
   );
   gpc1_1 gpc1212 (
      {stage0_25[238]},
      {stage1_25[100]}
   );
   gpc1_1 gpc1213 (
      {stage0_25[239]},
      {stage1_25[101]}
   );
   gpc1_1 gpc1214 (
      {stage0_25[240]},
      {stage1_25[102]}
   );
   gpc1_1 gpc1215 (
      {stage0_25[241]},
      {stage1_25[103]}
   );
   gpc1_1 gpc1216 (
      {stage0_25[242]},
      {stage1_25[104]}
   );
   gpc1_1 gpc1217 (
      {stage0_25[243]},
      {stage1_25[105]}
   );
   gpc1_1 gpc1218 (
      {stage0_25[244]},
      {stage1_25[106]}
   );
   gpc1_1 gpc1219 (
      {stage0_25[245]},
      {stage1_25[107]}
   );
   gpc1_1 gpc1220 (
      {stage0_25[246]},
      {stage1_25[108]}
   );
   gpc1_1 gpc1221 (
      {stage0_25[247]},
      {stage1_25[109]}
   );
   gpc1_1 gpc1222 (
      {stage0_25[248]},
      {stage1_25[110]}
   );
   gpc1_1 gpc1223 (
      {stage0_25[249]},
      {stage1_25[111]}
   );
   gpc1_1 gpc1224 (
      {stage0_25[250]},
      {stage1_25[112]}
   );
   gpc1_1 gpc1225 (
      {stage0_25[251]},
      {stage1_25[113]}
   );
   gpc1_1 gpc1226 (
      {stage0_25[252]},
      {stage1_25[114]}
   );
   gpc1_1 gpc1227 (
      {stage0_25[253]},
      {stage1_25[115]}
   );
   gpc1_1 gpc1228 (
      {stage0_25[254]},
      {stage1_25[116]}
   );
   gpc1_1 gpc1229 (
      {stage0_25[255]},
      {stage1_25[117]}
   );
   gpc1_1 gpc1230 (
      {stage0_26[72]},
      {stage1_26[53]}
   );
   gpc1_1 gpc1231 (
      {stage0_26[73]},
      {stage1_26[54]}
   );
   gpc1_1 gpc1232 (
      {stage0_26[74]},
      {stage1_26[55]}
   );
   gpc1_1 gpc1233 (
      {stage0_26[75]},
      {stage1_26[56]}
   );
   gpc1_1 gpc1234 (
      {stage0_26[76]},
      {stage1_26[57]}
   );
   gpc1_1 gpc1235 (
      {stage0_26[77]},
      {stage1_26[58]}
   );
   gpc1_1 gpc1236 (
      {stage0_26[78]},
      {stage1_26[59]}
   );
   gpc1_1 gpc1237 (
      {stage0_26[79]},
      {stage1_26[60]}
   );
   gpc1_1 gpc1238 (
      {stage0_26[80]},
      {stage1_26[61]}
   );
   gpc1_1 gpc1239 (
      {stage0_26[81]},
      {stage1_26[62]}
   );
   gpc1_1 gpc1240 (
      {stage0_26[82]},
      {stage1_26[63]}
   );
   gpc1_1 gpc1241 (
      {stage0_26[83]},
      {stage1_26[64]}
   );
   gpc1_1 gpc1242 (
      {stage0_26[84]},
      {stage1_26[65]}
   );
   gpc1_1 gpc1243 (
      {stage0_26[85]},
      {stage1_26[66]}
   );
   gpc1_1 gpc1244 (
      {stage0_26[86]},
      {stage1_26[67]}
   );
   gpc1_1 gpc1245 (
      {stage0_26[87]},
      {stage1_26[68]}
   );
   gpc1_1 gpc1246 (
      {stage0_26[88]},
      {stage1_26[69]}
   );
   gpc1_1 gpc1247 (
      {stage0_26[89]},
      {stage1_26[70]}
   );
   gpc1_1 gpc1248 (
      {stage0_26[90]},
      {stage1_26[71]}
   );
   gpc1_1 gpc1249 (
      {stage0_26[91]},
      {stage1_26[72]}
   );
   gpc1_1 gpc1250 (
      {stage0_26[92]},
      {stage1_26[73]}
   );
   gpc1_1 gpc1251 (
      {stage0_26[93]},
      {stage1_26[74]}
   );
   gpc1_1 gpc1252 (
      {stage0_26[94]},
      {stage1_26[75]}
   );
   gpc1_1 gpc1253 (
      {stage0_26[95]},
      {stage1_26[76]}
   );
   gpc1_1 gpc1254 (
      {stage0_26[96]},
      {stage1_26[77]}
   );
   gpc1_1 gpc1255 (
      {stage0_26[97]},
      {stage1_26[78]}
   );
   gpc1_1 gpc1256 (
      {stage0_26[98]},
      {stage1_26[79]}
   );
   gpc1_1 gpc1257 (
      {stage0_26[99]},
      {stage1_26[80]}
   );
   gpc1_1 gpc1258 (
      {stage0_26[100]},
      {stage1_26[81]}
   );
   gpc1_1 gpc1259 (
      {stage0_26[101]},
      {stage1_26[82]}
   );
   gpc1_1 gpc1260 (
      {stage0_26[102]},
      {stage1_26[83]}
   );
   gpc1_1 gpc1261 (
      {stage0_26[103]},
      {stage1_26[84]}
   );
   gpc1_1 gpc1262 (
      {stage0_26[104]},
      {stage1_26[85]}
   );
   gpc1_1 gpc1263 (
      {stage0_26[105]},
      {stage1_26[86]}
   );
   gpc1_1 gpc1264 (
      {stage0_26[106]},
      {stage1_26[87]}
   );
   gpc1_1 gpc1265 (
      {stage0_26[107]},
      {stage1_26[88]}
   );
   gpc1_1 gpc1266 (
      {stage0_26[108]},
      {stage1_26[89]}
   );
   gpc1_1 gpc1267 (
      {stage0_26[109]},
      {stage1_26[90]}
   );
   gpc1_1 gpc1268 (
      {stage0_26[110]},
      {stage1_26[91]}
   );
   gpc1_1 gpc1269 (
      {stage0_26[111]},
      {stage1_26[92]}
   );
   gpc1_1 gpc1270 (
      {stage0_26[112]},
      {stage1_26[93]}
   );
   gpc1_1 gpc1271 (
      {stage0_26[113]},
      {stage1_26[94]}
   );
   gpc1_1 gpc1272 (
      {stage0_26[114]},
      {stage1_26[95]}
   );
   gpc1_1 gpc1273 (
      {stage0_26[115]},
      {stage1_26[96]}
   );
   gpc1_1 gpc1274 (
      {stage0_26[116]},
      {stage1_26[97]}
   );
   gpc1_1 gpc1275 (
      {stage0_26[117]},
      {stage1_26[98]}
   );
   gpc1_1 gpc1276 (
      {stage0_26[118]},
      {stage1_26[99]}
   );
   gpc1_1 gpc1277 (
      {stage0_26[119]},
      {stage1_26[100]}
   );
   gpc1_1 gpc1278 (
      {stage0_26[120]},
      {stage1_26[101]}
   );
   gpc1_1 gpc1279 (
      {stage0_26[121]},
      {stage1_26[102]}
   );
   gpc1_1 gpc1280 (
      {stage0_26[122]},
      {stage1_26[103]}
   );
   gpc1_1 gpc1281 (
      {stage0_26[123]},
      {stage1_26[104]}
   );
   gpc1_1 gpc1282 (
      {stage0_26[124]},
      {stage1_26[105]}
   );
   gpc1_1 gpc1283 (
      {stage0_26[125]},
      {stage1_26[106]}
   );
   gpc1_1 gpc1284 (
      {stage0_26[126]},
      {stage1_26[107]}
   );
   gpc1_1 gpc1285 (
      {stage0_26[127]},
      {stage1_26[108]}
   );
   gpc1_1 gpc1286 (
      {stage0_26[128]},
      {stage1_26[109]}
   );
   gpc1_1 gpc1287 (
      {stage0_26[129]},
      {stage1_26[110]}
   );
   gpc1_1 gpc1288 (
      {stage0_26[130]},
      {stage1_26[111]}
   );
   gpc1_1 gpc1289 (
      {stage0_26[131]},
      {stage1_26[112]}
   );
   gpc1_1 gpc1290 (
      {stage0_26[132]},
      {stage1_26[113]}
   );
   gpc1_1 gpc1291 (
      {stage0_26[133]},
      {stage1_26[114]}
   );
   gpc1_1 gpc1292 (
      {stage0_26[134]},
      {stage1_26[115]}
   );
   gpc1_1 gpc1293 (
      {stage0_26[135]},
      {stage1_26[116]}
   );
   gpc1_1 gpc1294 (
      {stage0_26[136]},
      {stage1_26[117]}
   );
   gpc1_1 gpc1295 (
      {stage0_26[137]},
      {stage1_26[118]}
   );
   gpc1_1 gpc1296 (
      {stage0_26[138]},
      {stage1_26[119]}
   );
   gpc1_1 gpc1297 (
      {stage0_26[139]},
      {stage1_26[120]}
   );
   gpc1_1 gpc1298 (
      {stage0_26[140]},
      {stage1_26[121]}
   );
   gpc1_1 gpc1299 (
      {stage0_26[141]},
      {stage1_26[122]}
   );
   gpc1_1 gpc1300 (
      {stage0_26[142]},
      {stage1_26[123]}
   );
   gpc1_1 gpc1301 (
      {stage0_26[143]},
      {stage1_26[124]}
   );
   gpc1_1 gpc1302 (
      {stage0_26[144]},
      {stage1_26[125]}
   );
   gpc1_1 gpc1303 (
      {stage0_26[145]},
      {stage1_26[126]}
   );
   gpc1_1 gpc1304 (
      {stage0_26[146]},
      {stage1_26[127]}
   );
   gpc1_1 gpc1305 (
      {stage0_26[147]},
      {stage1_26[128]}
   );
   gpc1_1 gpc1306 (
      {stage0_26[148]},
      {stage1_26[129]}
   );
   gpc1_1 gpc1307 (
      {stage0_26[149]},
      {stage1_26[130]}
   );
   gpc1_1 gpc1308 (
      {stage0_26[150]},
      {stage1_26[131]}
   );
   gpc1_1 gpc1309 (
      {stage0_26[151]},
      {stage1_26[132]}
   );
   gpc1_1 gpc1310 (
      {stage0_26[152]},
      {stage1_26[133]}
   );
   gpc1_1 gpc1311 (
      {stage0_26[153]},
      {stage1_26[134]}
   );
   gpc1_1 gpc1312 (
      {stage0_26[154]},
      {stage1_26[135]}
   );
   gpc1_1 gpc1313 (
      {stage0_26[155]},
      {stage1_26[136]}
   );
   gpc1_1 gpc1314 (
      {stage0_26[156]},
      {stage1_26[137]}
   );
   gpc1_1 gpc1315 (
      {stage0_26[157]},
      {stage1_26[138]}
   );
   gpc1_1 gpc1316 (
      {stage0_26[158]},
      {stage1_26[139]}
   );
   gpc1_1 gpc1317 (
      {stage0_26[159]},
      {stage1_26[140]}
   );
   gpc1_1 gpc1318 (
      {stage0_26[160]},
      {stage1_26[141]}
   );
   gpc1_1 gpc1319 (
      {stage0_26[161]},
      {stage1_26[142]}
   );
   gpc1_1 gpc1320 (
      {stage0_26[162]},
      {stage1_26[143]}
   );
   gpc1_1 gpc1321 (
      {stage0_26[163]},
      {stage1_26[144]}
   );
   gpc1_1 gpc1322 (
      {stage0_26[164]},
      {stage1_26[145]}
   );
   gpc1_1 gpc1323 (
      {stage0_26[165]},
      {stage1_26[146]}
   );
   gpc1_1 gpc1324 (
      {stage0_26[166]},
      {stage1_26[147]}
   );
   gpc1_1 gpc1325 (
      {stage0_26[167]},
      {stage1_26[148]}
   );
   gpc1_1 gpc1326 (
      {stage0_26[168]},
      {stage1_26[149]}
   );
   gpc1_1 gpc1327 (
      {stage0_26[169]},
      {stage1_26[150]}
   );
   gpc1_1 gpc1328 (
      {stage0_26[170]},
      {stage1_26[151]}
   );
   gpc1_1 gpc1329 (
      {stage0_26[171]},
      {stage1_26[152]}
   );
   gpc1_1 gpc1330 (
      {stage0_26[172]},
      {stage1_26[153]}
   );
   gpc1_1 gpc1331 (
      {stage0_26[173]},
      {stage1_26[154]}
   );
   gpc1_1 gpc1332 (
      {stage0_26[174]},
      {stage1_26[155]}
   );
   gpc1_1 gpc1333 (
      {stage0_26[175]},
      {stage1_26[156]}
   );
   gpc1_1 gpc1334 (
      {stage0_26[176]},
      {stage1_26[157]}
   );
   gpc1_1 gpc1335 (
      {stage0_26[177]},
      {stage1_26[158]}
   );
   gpc1_1 gpc1336 (
      {stage0_26[178]},
      {stage1_26[159]}
   );
   gpc1_1 gpc1337 (
      {stage0_26[179]},
      {stage1_26[160]}
   );
   gpc1_1 gpc1338 (
      {stage0_26[180]},
      {stage1_26[161]}
   );
   gpc1_1 gpc1339 (
      {stage0_26[181]},
      {stage1_26[162]}
   );
   gpc1_1 gpc1340 (
      {stage0_26[182]},
      {stage1_26[163]}
   );
   gpc1_1 gpc1341 (
      {stage0_26[183]},
      {stage1_26[164]}
   );
   gpc1_1 gpc1342 (
      {stage0_26[184]},
      {stage1_26[165]}
   );
   gpc1_1 gpc1343 (
      {stage0_26[185]},
      {stage1_26[166]}
   );
   gpc1_1 gpc1344 (
      {stage0_26[186]},
      {stage1_26[167]}
   );
   gpc1_1 gpc1345 (
      {stage0_26[187]},
      {stage1_26[168]}
   );
   gpc1_1 gpc1346 (
      {stage0_26[188]},
      {stage1_26[169]}
   );
   gpc1_1 gpc1347 (
      {stage0_26[189]},
      {stage1_26[170]}
   );
   gpc1_1 gpc1348 (
      {stage0_26[190]},
      {stage1_26[171]}
   );
   gpc1_1 gpc1349 (
      {stage0_26[191]},
      {stage1_26[172]}
   );
   gpc1_1 gpc1350 (
      {stage0_26[192]},
      {stage1_26[173]}
   );
   gpc1_1 gpc1351 (
      {stage0_26[193]},
      {stage1_26[174]}
   );
   gpc1_1 gpc1352 (
      {stage0_26[194]},
      {stage1_26[175]}
   );
   gpc1_1 gpc1353 (
      {stage0_26[195]},
      {stage1_26[176]}
   );
   gpc1_1 gpc1354 (
      {stage0_26[196]},
      {stage1_26[177]}
   );
   gpc1_1 gpc1355 (
      {stage0_26[197]},
      {stage1_26[178]}
   );
   gpc1_1 gpc1356 (
      {stage0_26[198]},
      {stage1_26[179]}
   );
   gpc1_1 gpc1357 (
      {stage0_26[199]},
      {stage1_26[180]}
   );
   gpc1_1 gpc1358 (
      {stage0_26[200]},
      {stage1_26[181]}
   );
   gpc1_1 gpc1359 (
      {stage0_26[201]},
      {stage1_26[182]}
   );
   gpc1_1 gpc1360 (
      {stage0_26[202]},
      {stage1_26[183]}
   );
   gpc1_1 gpc1361 (
      {stage0_26[203]},
      {stage1_26[184]}
   );
   gpc1_1 gpc1362 (
      {stage0_26[204]},
      {stage1_26[185]}
   );
   gpc1_1 gpc1363 (
      {stage0_26[205]},
      {stage1_26[186]}
   );
   gpc1_1 gpc1364 (
      {stage0_26[206]},
      {stage1_26[187]}
   );
   gpc1_1 gpc1365 (
      {stage0_26[207]},
      {stage1_26[188]}
   );
   gpc1_1 gpc1366 (
      {stage0_26[208]},
      {stage1_26[189]}
   );
   gpc1_1 gpc1367 (
      {stage0_26[209]},
      {stage1_26[190]}
   );
   gpc1_1 gpc1368 (
      {stage0_26[210]},
      {stage1_26[191]}
   );
   gpc1_1 gpc1369 (
      {stage0_26[211]},
      {stage1_26[192]}
   );
   gpc1_1 gpc1370 (
      {stage0_26[212]},
      {stage1_26[193]}
   );
   gpc1_1 gpc1371 (
      {stage0_26[213]},
      {stage1_26[194]}
   );
   gpc1_1 gpc1372 (
      {stage0_26[214]},
      {stage1_26[195]}
   );
   gpc1_1 gpc1373 (
      {stage0_26[215]},
      {stage1_26[196]}
   );
   gpc1_1 gpc1374 (
      {stage0_26[216]},
      {stage1_26[197]}
   );
   gpc1_1 gpc1375 (
      {stage0_26[217]},
      {stage1_26[198]}
   );
   gpc1_1 gpc1376 (
      {stage0_26[218]},
      {stage1_26[199]}
   );
   gpc1_1 gpc1377 (
      {stage0_26[219]},
      {stage1_26[200]}
   );
   gpc1_1 gpc1378 (
      {stage0_26[220]},
      {stage1_26[201]}
   );
   gpc1_1 gpc1379 (
      {stage0_26[221]},
      {stage1_26[202]}
   );
   gpc1_1 gpc1380 (
      {stage0_26[222]},
      {stage1_26[203]}
   );
   gpc1_1 gpc1381 (
      {stage0_26[223]},
      {stage1_26[204]}
   );
   gpc1_1 gpc1382 (
      {stage0_26[224]},
      {stage1_26[205]}
   );
   gpc1_1 gpc1383 (
      {stage0_26[225]},
      {stage1_26[206]}
   );
   gpc1_1 gpc1384 (
      {stage0_26[226]},
      {stage1_26[207]}
   );
   gpc1_1 gpc1385 (
      {stage0_26[227]},
      {stage1_26[208]}
   );
   gpc1_1 gpc1386 (
      {stage0_26[228]},
      {stage1_26[209]}
   );
   gpc1_1 gpc1387 (
      {stage0_26[229]},
      {stage1_26[210]}
   );
   gpc1_1 gpc1388 (
      {stage0_26[230]},
      {stage1_26[211]}
   );
   gpc1_1 gpc1389 (
      {stage0_26[231]},
      {stage1_26[212]}
   );
   gpc1_1 gpc1390 (
      {stage0_26[232]},
      {stage1_26[213]}
   );
   gpc1_1 gpc1391 (
      {stage0_26[233]},
      {stage1_26[214]}
   );
   gpc1_1 gpc1392 (
      {stage0_26[234]},
      {stage1_26[215]}
   );
   gpc1_1 gpc1393 (
      {stage0_26[235]},
      {stage1_26[216]}
   );
   gpc1_1 gpc1394 (
      {stage0_26[236]},
      {stage1_26[217]}
   );
   gpc1_1 gpc1395 (
      {stage0_26[237]},
      {stage1_26[218]}
   );
   gpc1_1 gpc1396 (
      {stage0_26[238]},
      {stage1_26[219]}
   );
   gpc1_1 gpc1397 (
      {stage0_26[239]},
      {stage1_26[220]}
   );
   gpc1_1 gpc1398 (
      {stage0_26[240]},
      {stage1_26[221]}
   );
   gpc1_1 gpc1399 (
      {stage0_26[241]},
      {stage1_26[222]}
   );
   gpc1_1 gpc1400 (
      {stage0_26[242]},
      {stage1_26[223]}
   );
   gpc1_1 gpc1401 (
      {stage0_26[243]},
      {stage1_26[224]}
   );
   gpc1_1 gpc1402 (
      {stage0_26[244]},
      {stage1_26[225]}
   );
   gpc1_1 gpc1403 (
      {stage0_26[245]},
      {stage1_26[226]}
   );
   gpc1_1 gpc1404 (
      {stage0_26[246]},
      {stage1_26[227]}
   );
   gpc1_1 gpc1405 (
      {stage0_26[247]},
      {stage1_26[228]}
   );
   gpc1_1 gpc1406 (
      {stage0_26[248]},
      {stage1_26[229]}
   );
   gpc1_1 gpc1407 (
      {stage0_26[249]},
      {stage1_26[230]}
   );
   gpc1_1 gpc1408 (
      {stage0_26[250]},
      {stage1_26[231]}
   );
   gpc1_1 gpc1409 (
      {stage0_26[251]},
      {stage1_26[232]}
   );
   gpc1_1 gpc1410 (
      {stage0_26[252]},
      {stage1_26[233]}
   );
   gpc1_1 gpc1411 (
      {stage0_26[253]},
      {stage1_26[234]}
   );
   gpc1_1 gpc1412 (
      {stage0_26[254]},
      {stage1_26[235]}
   );
   gpc1_1 gpc1413 (
      {stage0_26[255]},
      {stage1_26[236]}
   );
   gpc1_1 gpc1414 (
      {stage0_27[204]},
      {stage1_27[56]}
   );
   gpc1_1 gpc1415 (
      {stage0_27[205]},
      {stage1_27[57]}
   );
   gpc1_1 gpc1416 (
      {stage0_27[206]},
      {stage1_27[58]}
   );
   gpc1_1 gpc1417 (
      {stage0_27[207]},
      {stage1_27[59]}
   );
   gpc1_1 gpc1418 (
      {stage0_27[208]},
      {stage1_27[60]}
   );
   gpc1_1 gpc1419 (
      {stage0_27[209]},
      {stage1_27[61]}
   );
   gpc1_1 gpc1420 (
      {stage0_27[210]},
      {stage1_27[62]}
   );
   gpc1_1 gpc1421 (
      {stage0_27[211]},
      {stage1_27[63]}
   );
   gpc1_1 gpc1422 (
      {stage0_27[212]},
      {stage1_27[64]}
   );
   gpc1_1 gpc1423 (
      {stage0_27[213]},
      {stage1_27[65]}
   );
   gpc1_1 gpc1424 (
      {stage0_27[214]},
      {stage1_27[66]}
   );
   gpc1_1 gpc1425 (
      {stage0_27[215]},
      {stage1_27[67]}
   );
   gpc1_1 gpc1426 (
      {stage0_27[216]},
      {stage1_27[68]}
   );
   gpc1_1 gpc1427 (
      {stage0_27[217]},
      {stage1_27[69]}
   );
   gpc1_1 gpc1428 (
      {stage0_27[218]},
      {stage1_27[70]}
   );
   gpc1_1 gpc1429 (
      {stage0_27[219]},
      {stage1_27[71]}
   );
   gpc1_1 gpc1430 (
      {stage0_27[220]},
      {stage1_27[72]}
   );
   gpc1_1 gpc1431 (
      {stage0_27[221]},
      {stage1_27[73]}
   );
   gpc1_1 gpc1432 (
      {stage0_27[222]},
      {stage1_27[74]}
   );
   gpc1_1 gpc1433 (
      {stage0_27[223]},
      {stage1_27[75]}
   );
   gpc1_1 gpc1434 (
      {stage0_27[224]},
      {stage1_27[76]}
   );
   gpc1_1 gpc1435 (
      {stage0_27[225]},
      {stage1_27[77]}
   );
   gpc1_1 gpc1436 (
      {stage0_27[226]},
      {stage1_27[78]}
   );
   gpc1_1 gpc1437 (
      {stage0_27[227]},
      {stage1_27[79]}
   );
   gpc1_1 gpc1438 (
      {stage0_27[228]},
      {stage1_27[80]}
   );
   gpc1_1 gpc1439 (
      {stage0_27[229]},
      {stage1_27[81]}
   );
   gpc1_1 gpc1440 (
      {stage0_27[230]},
      {stage1_27[82]}
   );
   gpc1_1 gpc1441 (
      {stage0_27[231]},
      {stage1_27[83]}
   );
   gpc1_1 gpc1442 (
      {stage0_27[232]},
      {stage1_27[84]}
   );
   gpc1_1 gpc1443 (
      {stage0_27[233]},
      {stage1_27[85]}
   );
   gpc1_1 gpc1444 (
      {stage0_27[234]},
      {stage1_27[86]}
   );
   gpc1_1 gpc1445 (
      {stage0_27[235]},
      {stage1_27[87]}
   );
   gpc1_1 gpc1446 (
      {stage0_27[236]},
      {stage1_27[88]}
   );
   gpc1_1 gpc1447 (
      {stage0_27[237]},
      {stage1_27[89]}
   );
   gpc1_1 gpc1448 (
      {stage0_27[238]},
      {stage1_27[90]}
   );
   gpc1_1 gpc1449 (
      {stage0_27[239]},
      {stage1_27[91]}
   );
   gpc1_1 gpc1450 (
      {stage0_27[240]},
      {stage1_27[92]}
   );
   gpc1_1 gpc1451 (
      {stage0_27[241]},
      {stage1_27[93]}
   );
   gpc1_1 gpc1452 (
      {stage0_27[242]},
      {stage1_27[94]}
   );
   gpc1_1 gpc1453 (
      {stage0_27[243]},
      {stage1_27[95]}
   );
   gpc1_1 gpc1454 (
      {stage0_27[244]},
      {stage1_27[96]}
   );
   gpc1_1 gpc1455 (
      {stage0_27[245]},
      {stage1_27[97]}
   );
   gpc1_1 gpc1456 (
      {stage0_27[246]},
      {stage1_27[98]}
   );
   gpc1_1 gpc1457 (
      {stage0_27[247]},
      {stage1_27[99]}
   );
   gpc1_1 gpc1458 (
      {stage0_27[248]},
      {stage1_27[100]}
   );
   gpc1_1 gpc1459 (
      {stage0_27[249]},
      {stage1_27[101]}
   );
   gpc1_1 gpc1460 (
      {stage0_27[250]},
      {stage1_27[102]}
   );
   gpc1_1 gpc1461 (
      {stage0_27[251]},
      {stage1_27[103]}
   );
   gpc1_1 gpc1462 (
      {stage0_27[252]},
      {stage1_27[104]}
   );
   gpc1_1 gpc1463 (
      {stage0_27[253]},
      {stage1_27[105]}
   );
   gpc1_1 gpc1464 (
      {stage0_27[254]},
      {stage1_27[106]}
   );
   gpc1_1 gpc1465 (
      {stage0_27[255]},
      {stage1_27[107]}
   );
   gpc1_1 gpc1466 (
      {stage0_28[240]},
      {stage1_28[86]}
   );
   gpc1_1 gpc1467 (
      {stage0_28[241]},
      {stage1_28[87]}
   );
   gpc1_1 gpc1468 (
      {stage0_28[242]},
      {stage1_28[88]}
   );
   gpc1_1 gpc1469 (
      {stage0_28[243]},
      {stage1_28[89]}
   );
   gpc1_1 gpc1470 (
      {stage0_28[244]},
      {stage1_28[90]}
   );
   gpc1_1 gpc1471 (
      {stage0_28[245]},
      {stage1_28[91]}
   );
   gpc1_1 gpc1472 (
      {stage0_28[246]},
      {stage1_28[92]}
   );
   gpc1_1 gpc1473 (
      {stage0_28[247]},
      {stage1_28[93]}
   );
   gpc1_1 gpc1474 (
      {stage0_28[248]},
      {stage1_28[94]}
   );
   gpc1_1 gpc1475 (
      {stage0_28[249]},
      {stage1_28[95]}
   );
   gpc1_1 gpc1476 (
      {stage0_28[250]},
      {stage1_28[96]}
   );
   gpc1_1 gpc1477 (
      {stage0_28[251]},
      {stage1_28[97]}
   );
   gpc1_1 gpc1478 (
      {stage0_28[252]},
      {stage1_28[98]}
   );
   gpc1_1 gpc1479 (
      {stage0_28[253]},
      {stage1_28[99]}
   );
   gpc1_1 gpc1480 (
      {stage0_28[254]},
      {stage1_28[100]}
   );
   gpc1_1 gpc1481 (
      {stage0_28[255]},
      {stage1_28[101]}
   );
   gpc1_1 gpc1482 (
      {stage0_29[246]},
      {stage1_29[108]}
   );
   gpc1_1 gpc1483 (
      {stage0_29[247]},
      {stage1_29[109]}
   );
   gpc1_1 gpc1484 (
      {stage0_29[248]},
      {stage1_29[110]}
   );
   gpc1_1 gpc1485 (
      {stage0_29[249]},
      {stage1_29[111]}
   );
   gpc1_1 gpc1486 (
      {stage0_29[250]},
      {stage1_29[112]}
   );
   gpc1_1 gpc1487 (
      {stage0_29[251]},
      {stage1_29[113]}
   );
   gpc1_1 gpc1488 (
      {stage0_29[252]},
      {stage1_29[114]}
   );
   gpc1_1 gpc1489 (
      {stage0_29[253]},
      {stage1_29[115]}
   );
   gpc1_1 gpc1490 (
      {stage0_29[254]},
      {stage1_29[116]}
   );
   gpc1_1 gpc1491 (
      {stage0_29[255]},
      {stage1_29[117]}
   );
   gpc1_1 gpc1492 (
      {stage0_30[240]},
      {stage1_30[81]}
   );
   gpc1_1 gpc1493 (
      {stage0_30[241]},
      {stage1_30[82]}
   );
   gpc1_1 gpc1494 (
      {stage0_30[242]},
      {stage1_30[83]}
   );
   gpc1_1 gpc1495 (
      {stage0_30[243]},
      {stage1_30[84]}
   );
   gpc1_1 gpc1496 (
      {stage0_30[244]},
      {stage1_30[85]}
   );
   gpc1_1 gpc1497 (
      {stage0_30[245]},
      {stage1_30[86]}
   );
   gpc1_1 gpc1498 (
      {stage0_30[246]},
      {stage1_30[87]}
   );
   gpc1_1 gpc1499 (
      {stage0_30[247]},
      {stage1_30[88]}
   );
   gpc1_1 gpc1500 (
      {stage0_30[248]},
      {stage1_30[89]}
   );
   gpc1_1 gpc1501 (
      {stage0_30[249]},
      {stage1_30[90]}
   );
   gpc1_1 gpc1502 (
      {stage0_30[250]},
      {stage1_30[91]}
   );
   gpc1_1 gpc1503 (
      {stage0_30[251]},
      {stage1_30[92]}
   );
   gpc1_1 gpc1504 (
      {stage0_30[252]},
      {stage1_30[93]}
   );
   gpc1_1 gpc1505 (
      {stage0_30[253]},
      {stage1_30[94]}
   );
   gpc1_1 gpc1506 (
      {stage0_30[254]},
      {stage1_30[95]}
   );
   gpc1_1 gpc1507 (
      {stage0_30[255]},
      {stage1_30[96]}
   );
   gpc1_1 gpc1508 (
      {stage0_31[204]},
      {stage1_31[81]}
   );
   gpc1_1 gpc1509 (
      {stage0_31[205]},
      {stage1_31[82]}
   );
   gpc1_1 gpc1510 (
      {stage0_31[206]},
      {stage1_31[83]}
   );
   gpc1_1 gpc1511 (
      {stage0_31[207]},
      {stage1_31[84]}
   );
   gpc1_1 gpc1512 (
      {stage0_31[208]},
      {stage1_31[85]}
   );
   gpc1_1 gpc1513 (
      {stage0_31[209]},
      {stage1_31[86]}
   );
   gpc1_1 gpc1514 (
      {stage0_31[210]},
      {stage1_31[87]}
   );
   gpc1_1 gpc1515 (
      {stage0_31[211]},
      {stage1_31[88]}
   );
   gpc1_1 gpc1516 (
      {stage0_31[212]},
      {stage1_31[89]}
   );
   gpc1_1 gpc1517 (
      {stage0_31[213]},
      {stage1_31[90]}
   );
   gpc1_1 gpc1518 (
      {stage0_31[214]},
      {stage1_31[91]}
   );
   gpc1_1 gpc1519 (
      {stage0_31[215]},
      {stage1_31[92]}
   );
   gpc1_1 gpc1520 (
      {stage0_31[216]},
      {stage1_31[93]}
   );
   gpc1_1 gpc1521 (
      {stage0_31[217]},
      {stage1_31[94]}
   );
   gpc1_1 gpc1522 (
      {stage0_31[218]},
      {stage1_31[95]}
   );
   gpc1_1 gpc1523 (
      {stage0_31[219]},
      {stage1_31[96]}
   );
   gpc1_1 gpc1524 (
      {stage0_31[220]},
      {stage1_31[97]}
   );
   gpc1_1 gpc1525 (
      {stage0_31[221]},
      {stage1_31[98]}
   );
   gpc1_1 gpc1526 (
      {stage0_31[222]},
      {stage1_31[99]}
   );
   gpc1_1 gpc1527 (
      {stage0_31[223]},
      {stage1_31[100]}
   );
   gpc1_1 gpc1528 (
      {stage0_31[224]},
      {stage1_31[101]}
   );
   gpc1_1 gpc1529 (
      {stage0_31[225]},
      {stage1_31[102]}
   );
   gpc1_1 gpc1530 (
      {stage0_31[226]},
      {stage1_31[103]}
   );
   gpc1_1 gpc1531 (
      {stage0_31[227]},
      {stage1_31[104]}
   );
   gpc1_1 gpc1532 (
      {stage0_31[228]},
      {stage1_31[105]}
   );
   gpc1_1 gpc1533 (
      {stage0_31[229]},
      {stage1_31[106]}
   );
   gpc1_1 gpc1534 (
      {stage0_31[230]},
      {stage1_31[107]}
   );
   gpc1_1 gpc1535 (
      {stage0_31[231]},
      {stage1_31[108]}
   );
   gpc1_1 gpc1536 (
      {stage0_31[232]},
      {stage1_31[109]}
   );
   gpc1_1 gpc1537 (
      {stage0_31[233]},
      {stage1_31[110]}
   );
   gpc1_1 gpc1538 (
      {stage0_31[234]},
      {stage1_31[111]}
   );
   gpc1_1 gpc1539 (
      {stage0_31[235]},
      {stage1_31[112]}
   );
   gpc1_1 gpc1540 (
      {stage0_31[236]},
      {stage1_31[113]}
   );
   gpc1_1 gpc1541 (
      {stage0_31[237]},
      {stage1_31[114]}
   );
   gpc1_1 gpc1542 (
      {stage0_31[238]},
      {stage1_31[115]}
   );
   gpc1_1 gpc1543 (
      {stage0_31[239]},
      {stage1_31[116]}
   );
   gpc1_1 gpc1544 (
      {stage0_31[240]},
      {stage1_31[117]}
   );
   gpc1_1 gpc1545 (
      {stage0_31[241]},
      {stage1_31[118]}
   );
   gpc1_1 gpc1546 (
      {stage0_31[242]},
      {stage1_31[119]}
   );
   gpc1_1 gpc1547 (
      {stage0_31[243]},
      {stage1_31[120]}
   );
   gpc1_1 gpc1548 (
      {stage0_31[244]},
      {stage1_31[121]}
   );
   gpc1_1 gpc1549 (
      {stage0_31[245]},
      {stage1_31[122]}
   );
   gpc1_1 gpc1550 (
      {stage0_31[246]},
      {stage1_31[123]}
   );
   gpc1_1 gpc1551 (
      {stage0_31[247]},
      {stage1_31[124]}
   );
   gpc1_1 gpc1552 (
      {stage0_31[248]},
      {stage1_31[125]}
   );
   gpc1_1 gpc1553 (
      {stage0_31[249]},
      {stage1_31[126]}
   );
   gpc1_1 gpc1554 (
      {stage0_31[250]},
      {stage1_31[127]}
   );
   gpc1_1 gpc1555 (
      {stage0_31[251]},
      {stage1_31[128]}
   );
   gpc1_1 gpc1556 (
      {stage0_31[252]},
      {stage1_31[129]}
   );
   gpc1_1 gpc1557 (
      {stage0_31[253]},
      {stage1_31[130]}
   );
   gpc1_1 gpc1558 (
      {stage0_31[254]},
      {stage1_31[131]}
   );
   gpc1_1 gpc1559 (
      {stage0_31[255]},
      {stage1_31[132]}
   );
   gpc1163_5 gpc1560 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc1561 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc1562 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc1563 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc1564 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc1565 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc1566 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc1567 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc1568 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc1569 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc1570 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc1571 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1163_5 gpc1572 (
      {stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_2[12]},
      {stage1_3[12]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc1573 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc1574 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_3[13]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc1575 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28]},
      {stage1_3[14]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[15],stage2_3[15],stage2_2[15]}
   );
   gpc615_5 gpc1576 (
      {stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage1_3[15]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[16],stage2_3[16],stage2_2[16]}
   );
   gpc615_5 gpc1577 (
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38]},
      {stage1_3[16]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[17],stage2_3[17],stage2_2[17]}
   );
   gpc615_5 gpc1578 (
      {stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43]},
      {stage1_3[17]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[18],stage2_3[18],stage2_2[18]}
   );
   gpc615_5 gpc1579 (
      {stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48]},
      {stage1_3[18]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[19],stage2_3[19],stage2_2[19]}
   );
   gpc615_5 gpc1580 (
      {stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage1_3[19]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[20],stage2_3[20],stage2_2[20]}
   );
   gpc615_5 gpc1581 (
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58]},
      {stage1_3[20]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[8],stage2_4[21],stage2_3[21],stage2_2[21]}
   );
   gpc615_5 gpc1582 (
      {stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage1_3[21]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[9],stage2_4[22],stage2_3[22],stage2_2[22]}
   );
   gpc615_5 gpc1583 (
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68]},
      {stage1_3[22]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[10],stage2_4[23],stage2_3[23],stage2_2[23]}
   );
   gpc615_5 gpc1584 (
      {stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73]},
      {stage1_3[23]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[11],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc615_5 gpc1585 (
      {stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77], stage1_2[78]},
      {stage1_3[24]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[12],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc615_5 gpc1586 (
      {stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83]},
      {stage1_3[25]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[13],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc606_5 gpc1587 (
      {stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[14],stage2_5[14],stage2_4[27],stage2_3[27]}
   );
   gpc615_5 gpc1588 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[84]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[15],stage2_5[15],stage2_4[28],stage2_3[28]}
   );
   gpc615_5 gpc1589 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[85]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[16],stage2_5[16],stage2_4[29],stage2_3[29]}
   );
   gpc615_5 gpc1590 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[86]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[17],stage2_5[17],stage2_4[30],stage2_3[30]}
   );
   gpc615_5 gpc1591 (
      {stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage1_4[87]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[18],stage2_5[18],stage2_4[31],stage2_3[31]}
   );
   gpc615_5 gpc1592 (
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56]},
      {stage1_4[88]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[19],stage2_5[19],stage2_4[32],stage2_3[32]}
   );
   gpc615_5 gpc1593 (
      {stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage1_4[89]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[20],stage2_5[20],stage2_4[33],stage2_3[33]}
   );
   gpc615_5 gpc1594 (
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66]},
      {stage1_4[90]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[21],stage2_5[21],stage2_4[34],stage2_3[34]}
   );
   gpc615_5 gpc1595 (
      {stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage1_4[91]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[22],stage2_5[22],stage2_4[35],stage2_3[35]}
   );
   gpc615_5 gpc1596 (
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_4[92]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[23],stage2_5[23],stage2_4[36],stage2_3[36]}
   );
   gpc615_5 gpc1597 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage1_4[93]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[24],stage2_5[24],stage2_4[37],stage2_3[37]}
   );
   gpc615_5 gpc1598 (
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86]},
      {stage1_4[94]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[25],stage2_5[25],stage2_4[38],stage2_3[38]}
   );
   gpc207_4 gpc1599 (
      {stage1_4[95], stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage1_6[0], stage1_6[1]},
      {stage2_7[12],stage2_6[26],stage2_5[26],stage2_4[39]}
   );
   gpc606_5 gpc1600 (
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[13],stage2_6[27],stage2_5[27],stage2_4[40]}
   );
   gpc615_5 gpc1601 (
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112]},
      {stage1_5[72]},
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage2_8[1],stage2_7[14],stage2_6[28],stage2_5[28],stage2_4[41]}
   );
   gpc615_5 gpc1602 (
      {stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117]},
      {stage1_5[73]},
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18], stage1_6[19]},
      {stage2_8[2],stage2_7[15],stage2_6[29],stage2_5[29],stage2_4[42]}
   );
   gpc606_5 gpc1603 (
      {stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[3],stage2_7[16],stage2_6[30],stage2_5[30]}
   );
   gpc606_5 gpc1604 (
      {stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[4],stage2_7[17],stage2_6[31],stage2_5[31]}
   );
   gpc606_5 gpc1605 (
      {stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[5],stage2_7[18],stage2_6[32],stage2_5[32]}
   );
   gpc606_5 gpc1606 (
      {stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[6],stage2_7[19],stage2_6[33],stage2_5[33]}
   );
   gpc606_5 gpc1607 (
      {stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[7],stage2_7[20],stage2_6[34],stage2_5[34]}
   );
   gpc606_5 gpc1608 (
      {stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[8],stage2_7[21],stage2_6[35],stage2_5[35]}
   );
   gpc606_5 gpc1609 (
      {stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[9],stage2_7[22],stage2_6[36],stage2_5[36]}
   );
   gpc606_5 gpc1610 (
      {stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[10],stage2_7[23],stage2_6[37],stage2_5[37]}
   );
   gpc606_5 gpc1611 (
      {stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[8],stage2_8[11],stage2_7[24],stage2_6[38]}
   );
   gpc615_5 gpc1612 (
      {stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage1_7[48]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[9],stage2_8[12],stage2_7[25],stage2_6[39]}
   );
   gpc615_5 gpc1613 (
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_7[49]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[10],stage2_8[13],stage2_7[26],stage2_6[40]}
   );
   gpc615_5 gpc1614 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40]},
      {stage1_7[50]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[11],stage2_8[14],stage2_7[27],stage2_6[41]}
   );
   gpc615_5 gpc1615 (
      {stage1_6[41], stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45]},
      {stage1_7[51]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[12],stage2_8[15],stage2_7[28],stage2_6[42]}
   );
   gpc615_5 gpc1616 (
      {stage1_6[46], stage1_6[47], stage1_6[48], stage1_6[49], stage1_6[50]},
      {stage1_7[52]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[13],stage2_8[16],stage2_7[29],stage2_6[43]}
   );
   gpc615_5 gpc1617 (
      {stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55]},
      {stage1_7[53]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[14],stage2_8[17],stage2_7[30],stage2_6[44]}
   );
   gpc615_5 gpc1618 (
      {stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage1_7[54]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[15],stage2_8[18],stage2_7[31],stage2_6[45]}
   );
   gpc615_5 gpc1619 (
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage1_7[55]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[16],stage2_8[19],stage2_7[32],stage2_6[46]}
   );
   gpc615_5 gpc1620 (
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70]},
      {stage1_7[56]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[17],stage2_8[20],stage2_7[33],stage2_6[47]}
   );
   gpc615_5 gpc1621 (
      {stage1_6[71], stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75]},
      {stage1_7[57]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[18],stage2_8[21],stage2_7[34],stage2_6[48]}
   );
   gpc615_5 gpc1622 (
      {stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80]},
      {stage1_7[58]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[19],stage2_8[22],stage2_7[35],stage2_6[49]}
   );
   gpc615_5 gpc1623 (
      {stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85]},
      {stage1_7[59]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[20],stage2_8[23],stage2_7[36],stage2_6[50]}
   );
   gpc615_5 gpc1624 (
      {stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage1_7[60]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[21],stage2_8[24],stage2_7[37],stage2_6[51]}
   );
   gpc615_5 gpc1625 (
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_7[61]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[22],stage2_8[25],stage2_7[38],stage2_6[52]}
   );
   gpc615_5 gpc1626 (
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage1_8[90]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[15],stage2_9[23],stage2_8[26],stage2_7[39]}
   );
   gpc615_5 gpc1627 (
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage1_8[91]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[16],stage2_9[24],stage2_8[27],stage2_7[40]}
   );
   gpc615_5 gpc1628 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[92]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[17],stage2_9[25],stage2_8[28],stage2_7[41]}
   );
   gpc615_5 gpc1629 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[93]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[18],stage2_9[26],stage2_8[29],stage2_7[42]}
   );
   gpc615_5 gpc1630 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[94]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[19],stage2_9[27],stage2_8[30],stage2_7[43]}
   );
   gpc615_5 gpc1631 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage1_8[95]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[20],stage2_9[28],stage2_8[31],stage2_7[44]}
   );
   gpc606_5 gpc1632 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[6],stage2_10[21],stage2_9[29]}
   );
   gpc606_5 gpc1633 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[1],stage2_11[7],stage2_10[22],stage2_9[30]}
   );
   gpc606_5 gpc1634 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[2],stage2_11[8],stage2_10[23],stage2_9[31]}
   );
   gpc606_5 gpc1635 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[3],stage2_11[9],stage2_10[24],stage2_9[32]}
   );
   gpc606_5 gpc1636 (
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[4],stage2_11[10],stage2_10[25],stage2_9[33]}
   );
   gpc606_5 gpc1637 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[5],stage2_11[11],stage2_10[26],stage2_9[34]}
   );
   gpc606_5 gpc1638 (
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[6],stage2_11[12],stage2_10[27],stage2_9[35]}
   );
   gpc606_5 gpc1639 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[7],stage2_11[13],stage2_10[28],stage2_9[36]}
   );
   gpc606_5 gpc1640 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[8],stage2_11[14],stage2_10[29],stage2_9[37]}
   );
   gpc606_5 gpc1641 (
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[9],stage2_11[15],stage2_10[30],stage2_9[38]}
   );
   gpc606_5 gpc1642 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[10],stage2_11[16],stage2_10[31],stage2_9[39]}
   );
   gpc615_5 gpc1643 (
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106]},
      {stage1_10[0]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[11],stage2_11[17],stage2_10[32],stage2_9[40]}
   );
   gpc606_5 gpc1644 (
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[12],stage2_12[12],stage2_11[18],stage2_10[33]}
   );
   gpc606_5 gpc1645 (
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[13],stage2_12[13],stage2_11[19],stage2_10[34]}
   );
   gpc606_5 gpc1646 (
      {stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[14],stage2_12[14],stage2_11[20],stage2_10[35]}
   );
   gpc606_5 gpc1647 (
      {stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[15],stage2_12[15],stage2_11[21],stage2_10[36]}
   );
   gpc606_5 gpc1648 (
      {stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[16],stage2_12[16],stage2_11[22],stage2_10[37]}
   );
   gpc606_5 gpc1649 (
      {stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[17],stage2_12[17],stage2_11[23],stage2_10[38]}
   );
   gpc606_5 gpc1650 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[18],stage2_12[18],stage2_11[24],stage2_10[39]}
   );
   gpc606_5 gpc1651 (
      {stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[19],stage2_12[19],stage2_11[25],stage2_10[40]}
   );
   gpc606_5 gpc1652 (
      {stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[20],stage2_12[20],stage2_11[26],stage2_10[41]}
   );
   gpc606_5 gpc1653 (
      {stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[21],stage2_12[21],stage2_11[27],stage2_10[42]}
   );
   gpc606_5 gpc1654 (
      {stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[22],stage2_12[22],stage2_11[28],stage2_10[43]}
   );
   gpc606_5 gpc1655 (
      {stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[23],stage2_12[23],stage2_11[29],stage2_10[44]}
   );
   gpc606_5 gpc1656 (
      {stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[24],stage2_12[24],stage2_11[30],stage2_10[45]}
   );
   gpc606_5 gpc1657 (
      {stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83], stage1_10[84]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[25],stage2_12[25],stage2_11[31],stage2_10[46]}
   );
   gpc606_5 gpc1658 (
      {stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[26],stage2_12[26],stage2_11[32],stage2_10[47]}
   );
   gpc606_5 gpc1659 (
      {stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage2_14[15],stage2_13[27],stage2_12[27],stage2_11[33],stage2_10[48]}
   );
   gpc615_5 gpc1660 (
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76]},
      {stage1_12[96]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[16],stage2_13[28],stage2_12[28],stage2_11[34]}
   );
   gpc615_5 gpc1661 (
      {stage1_11[77], stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81]},
      {stage1_12[97]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[17],stage2_13[29],stage2_12[29],stage2_11[35]}
   );
   gpc615_5 gpc1662 (
      {stage1_11[82], stage1_11[83], stage1_11[84], stage1_11[85], stage1_11[86]},
      {stage1_12[98]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[18],stage2_13[30],stage2_12[30],stage2_11[36]}
   );
   gpc615_5 gpc1663 (
      {stage1_11[87], stage1_11[88], stage1_11[89], stage1_11[90], stage1_11[91]},
      {stage1_12[99]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[19],stage2_13[31],stage2_12[31],stage2_11[37]}
   );
   gpc615_5 gpc1664 (
      {stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95], stage1_11[96]},
      {stage1_12[100]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[20],stage2_13[32],stage2_12[32],stage2_11[38]}
   );
   gpc615_5 gpc1665 (
      {stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage1_12[101]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[21],stage2_13[33],stage2_12[33],stage2_11[39]}
   );
   gpc615_5 gpc1666 (
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106]},
      {stage1_12[102]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[22],stage2_13[34],stage2_12[34],stage2_11[40]}
   );
   gpc615_5 gpc1667 (
      {stage1_11[107], stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111]},
      {stage1_12[103]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[23],stage2_13[35],stage2_12[35],stage2_11[41]}
   );
   gpc615_5 gpc1668 (
      {stage1_11[112], stage1_11[113], stage1_11[114], stage1_11[115], stage1_11[116]},
      {stage1_12[104]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[24],stage2_13[36],stage2_12[36],stage2_11[42]}
   );
   gpc615_5 gpc1669 (
      {stage1_11[117], stage1_11[118], stage1_11[119], stage1_11[120], stage1_11[121]},
      {stage1_12[105]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[25],stage2_13[37],stage2_12[37],stage2_11[43]}
   );
   gpc615_5 gpc1670 (
      {stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125], stage1_11[126]},
      {stage1_12[106]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[26],stage2_13[38],stage2_12[38],stage2_11[44]}
   );
   gpc606_5 gpc1671 (
      {stage1_12[107], stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[11],stage2_14[27],stage2_13[39],stage2_12[39]}
   );
   gpc606_5 gpc1672 (
      {stage1_12[113], stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[12],stage2_14[28],stage2_13[40],stage2_12[40]}
   );
   gpc606_5 gpc1673 (
      {stage1_12[119], stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[13],stage2_14[29],stage2_13[41],stage2_12[41]}
   );
   gpc606_5 gpc1674 (
      {stage1_12[125], stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[14],stage2_14[30],stage2_13[42],stage2_12[42]}
   );
   gpc606_5 gpc1675 (
      {stage1_12[131], stage1_12[132], stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[15],stage2_14[31],stage2_13[43],stage2_12[43]}
   );
   gpc606_5 gpc1676 (
      {stage1_12[137], stage1_12[138], stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[16],stage2_14[32],stage2_13[44],stage2_12[44]}
   );
   gpc606_5 gpc1677 (
      {stage1_12[143], stage1_12[144], stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[17],stage2_14[33],stage2_13[45],stage2_12[45]}
   );
   gpc606_5 gpc1678 (
      {stage1_12[149], stage1_12[150], stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[18],stage2_14[34],stage2_13[46],stage2_12[46]}
   );
   gpc606_5 gpc1679 (
      {stage1_12[155], stage1_12[156], stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[19],stage2_14[35],stage2_13[47],stage2_12[47]}
   );
   gpc606_5 gpc1680 (
      {stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164], stage1_12[165], stage1_12[166]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[20],stage2_14[36],stage2_13[48],stage2_12[48]}
   );
   gpc606_5 gpc1681 (
      {stage1_12[167], stage1_12[168], stage1_12[169], stage1_12[170], stage1_12[171], stage1_12[172]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[21],stage2_14[37],stage2_13[49],stage2_12[49]}
   );
   gpc606_5 gpc1682 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[11],stage2_15[22],stage2_14[38],stage2_13[50]}
   );
   gpc606_5 gpc1683 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[12],stage2_15[23],stage2_14[39],stage2_13[51]}
   );
   gpc606_5 gpc1684 (
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[13],stage2_15[24],stage2_14[40],stage2_13[52]}
   );
   gpc606_5 gpc1685 (
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[14],stage2_15[25],stage2_14[41],stage2_13[53]}
   );
   gpc615_5 gpc1686 (
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[0],stage2_17[4],stage2_16[15],stage2_15[26]}
   );
   gpc615_5 gpc1687 (
      {stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33]},
      {stage1_16[1]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[1],stage2_17[5],stage2_16[16],stage2_15[27]}
   );
   gpc615_5 gpc1688 (
      {stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37], stage1_15[38]},
      {stage1_16[2]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[2],stage2_17[6],stage2_16[17],stage2_15[28]}
   );
   gpc615_5 gpc1689 (
      {stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage1_16[3]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[3],stage2_17[7],stage2_16[18],stage2_15[29]}
   );
   gpc615_5 gpc1690 (
      {stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48]},
      {stage1_16[4]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[4],stage2_17[8],stage2_16[19],stage2_15[30]}
   );
   gpc615_5 gpc1691 (
      {stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage1_16[5]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[5],stage2_17[9],stage2_16[20],stage2_15[31]}
   );
   gpc615_5 gpc1692 (
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58]},
      {stage1_16[6]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[6],stage2_17[10],stage2_16[21],stage2_15[32]}
   );
   gpc615_5 gpc1693 (
      {stage1_15[59], stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63]},
      {stage1_16[7]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[7],stage2_17[11],stage2_16[22],stage2_15[33]}
   );
   gpc615_5 gpc1694 (
      {stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67], stage1_15[68]},
      {stage1_16[8]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[8],stage2_17[12],stage2_16[23],stage2_15[34]}
   );
   gpc615_5 gpc1695 (
      {stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72], stage1_15[73]},
      {stage1_16[9]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[9],stage2_17[13],stage2_16[24],stage2_15[35]}
   );
   gpc615_5 gpc1696 (
      {stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77], stage1_15[78]},
      {stage1_16[10]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[10],stage2_17[14],stage2_16[25],stage2_15[36]}
   );
   gpc615_5 gpc1697 (
      {stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage1_16[11]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[11],stage2_17[15],stage2_16[26],stage2_15[37]}
   );
   gpc606_5 gpc1698 (
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[12],stage2_18[12],stage2_17[16],stage2_16[27]}
   );
   gpc606_5 gpc1699 (
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[13],stage2_18[13],stage2_17[17],stage2_16[28]}
   );
   gpc606_5 gpc1700 (
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[14],stage2_18[14],stage2_17[18],stage2_16[29]}
   );
   gpc606_5 gpc1701 (
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[15],stage2_18[15],stage2_17[19],stage2_16[30]}
   );
   gpc606_5 gpc1702 (
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[16],stage2_18[16],stage2_17[20],stage2_16[31]}
   );
   gpc606_5 gpc1703 (
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[17],stage2_18[17],stage2_17[21],stage2_16[32]}
   );
   gpc606_5 gpc1704 (
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[18],stage2_18[18],stage2_17[22],stage2_16[33]}
   );
   gpc606_5 gpc1705 (
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[19],stage2_18[19],stage2_17[23],stage2_16[34]}
   );
   gpc606_5 gpc1706 (
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage2_20[8],stage2_19[20],stage2_18[20],stage2_17[24],stage2_16[35]}
   );
   gpc606_5 gpc1707 (
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage2_20[9],stage2_19[21],stage2_18[21],stage2_17[25],stage2_16[36]}
   );
   gpc606_5 gpc1708 (
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage2_20[10],stage2_19[22],stage2_18[22],stage2_17[26],stage2_16[37]}
   );
   gpc606_5 gpc1709 (
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage2_20[11],stage2_19[23],stage2_18[23],stage2_17[27],stage2_16[38]}
   );
   gpc606_5 gpc1710 (
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage2_20[12],stage2_19[24],stage2_18[24],stage2_17[28],stage2_16[39]}
   );
   gpc606_5 gpc1711 (
      {stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95]},
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage2_20[13],stage2_19[25],stage2_18[25],stage2_17[29],stage2_16[40]}
   );
   gpc606_5 gpc1712 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[14],stage2_19[26],stage2_18[26],stage2_17[30]}
   );
   gpc606_5 gpc1713 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[15],stage2_19[27],stage2_18[27],stage2_17[31]}
   );
   gpc606_5 gpc1714 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[16],stage2_19[28],stage2_18[28],stage2_17[32]}
   );
   gpc606_5 gpc1715 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[17],stage2_19[29],stage2_18[29],stage2_17[33]}
   );
   gpc606_5 gpc1716 (
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[18],stage2_19[30],stage2_18[30],stage2_17[34]}
   );
   gpc606_5 gpc1717 (
      {stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105], stage1_17[106], stage1_17[107]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[19],stage2_19[31],stage2_18[31],stage2_17[35]}
   );
   gpc615_5 gpc1718 (
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88]},
      {stage1_19[36]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[6],stage2_20[20],stage2_19[32],stage2_18[32]}
   );
   gpc615_5 gpc1719 (
      {stage1_18[89], stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93]},
      {stage1_19[37]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[7],stage2_20[21],stage2_19[33],stage2_18[33]}
   );
   gpc615_5 gpc1720 (
      {stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41], stage1_19[42]},
      {stage1_20[12]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[2],stage2_21[8],stage2_20[22],stage2_19[34]}
   );
   gpc615_5 gpc1721 (
      {stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage1_20[13]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[3],stage2_21[9],stage2_20[23],stage2_19[35]}
   );
   gpc615_5 gpc1722 (
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52]},
      {stage1_20[14]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[4],stage2_21[10],stage2_20[24],stage2_19[36]}
   );
   gpc615_5 gpc1723 (
      {stage1_19[53], stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57]},
      {stage1_20[15]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[5],stage2_21[11],stage2_20[25],stage2_19[37]}
   );
   gpc615_5 gpc1724 (
      {stage1_19[58], stage1_19[59], stage1_19[60], stage1_19[61], stage1_19[62]},
      {stage1_20[16]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[6],stage2_21[12],stage2_20[26],stage2_19[38]}
   );
   gpc615_5 gpc1725 (
      {stage1_19[63], stage1_19[64], stage1_19[65], stage1_19[66], stage1_19[67]},
      {stage1_20[17]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[7],stage2_21[13],stage2_20[27],stage2_19[39]}
   );
   gpc615_5 gpc1726 (
      {stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71], stage1_19[72]},
      {stage1_20[18]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[8],stage2_21[14],stage2_20[28],stage2_19[40]}
   );
   gpc615_5 gpc1727 (
      {stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage1_20[19]},
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage2_23[7],stage2_22[9],stage2_21[15],stage2_20[29],stage2_19[41]}
   );
   gpc615_5 gpc1728 (
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82]},
      {stage1_20[20]},
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage2_23[8],stage2_22[10],stage2_21[16],stage2_20[30],stage2_19[42]}
   );
   gpc615_5 gpc1729 (
      {stage1_19[83], stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87]},
      {stage1_20[21]},
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage2_23[9],stage2_22[11],stage2_21[17],stage2_20[31],stage2_19[43]}
   );
   gpc615_5 gpc1730 (
      {stage1_19[88], stage1_19[89], stage1_19[90], stage1_19[91], stage1_19[92]},
      {stage1_20[22]},
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage2_23[10],stage2_22[12],stage2_21[18],stage2_20[32],stage2_19[44]}
   );
   gpc606_5 gpc1731 (
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[0],stage2_23[11],stage2_22[13],stage2_21[19]}
   );
   gpc606_5 gpc1732 (
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[1],stage2_23[12],stage2_22[14],stage2_21[20]}
   );
   gpc606_5 gpc1733 (
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[2],stage2_23[13],stage2_22[15],stage2_21[21]}
   );
   gpc606_5 gpc1734 (
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[3],stage2_23[14],stage2_22[16],stage2_21[22]}
   );
   gpc606_5 gpc1735 (
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[4],stage2_23[15],stage2_22[17]}
   );
   gpc606_5 gpc1736 (
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[5],stage2_24[5],stage2_23[16],stage2_22[18]}
   );
   gpc606_5 gpc1737 (
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[6],stage2_24[6],stage2_23[17],stage2_22[19]}
   );
   gpc606_5 gpc1738 (
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[7],stage2_24[7],stage2_23[18],stage2_22[20]}
   );
   gpc606_5 gpc1739 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[8],stage2_24[8],stage2_23[19],stage2_22[21]}
   );
   gpc606_5 gpc1740 (
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[9],stage2_24[9],stage2_23[20],stage2_22[22]}
   );
   gpc606_5 gpc1741 (
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[10],stage2_24[10],stage2_23[21],stage2_22[23]}
   );
   gpc606_5 gpc1742 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[11],stage2_24[11],stage2_23[22],stage2_22[24]}
   );
   gpc606_5 gpc1743 (
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[12],stage2_24[12],stage2_23[23],stage2_22[25]}
   );
   gpc606_5 gpc1744 (
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[13],stage2_24[13],stage2_23[24],stage2_22[26]}
   );
   gpc606_5 gpc1745 (
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[14],stage2_24[14],stage2_23[25],stage2_22[27]}
   );
   gpc606_5 gpc1746 (
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[15],stage2_24[15],stage2_23[26],stage2_22[28]}
   );
   gpc615_5 gpc1747 (
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76]},
      {stage1_23[24]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[16],stage2_24[16],stage2_23[27],stage2_22[29]}
   );
   gpc606_5 gpc1748 (
      {stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29], stage1_23[30]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[13],stage2_25[17],stage2_24[17],stage2_23[28]}
   );
   gpc606_5 gpc1749 (
      {stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35], stage1_23[36]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[14],stage2_25[18],stage2_24[18],stage2_23[29]}
   );
   gpc606_5 gpc1750 (
      {stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41], stage1_23[42]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[15],stage2_25[19],stage2_24[19],stage2_23[30]}
   );
   gpc606_5 gpc1751 (
      {stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47], stage1_23[48]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[16],stage2_25[20],stage2_24[20],stage2_23[31]}
   );
   gpc606_5 gpc1752 (
      {stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53], stage1_23[54]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[17],stage2_25[21],stage2_24[21],stage2_23[32]}
   );
   gpc606_5 gpc1753 (
      {stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59], stage1_23[60]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[18],stage2_25[22],stage2_24[22],stage2_23[33]}
   );
   gpc606_5 gpc1754 (
      {stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65], stage1_23[66]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[19],stage2_25[23],stage2_24[23],stage2_23[34]}
   );
   gpc606_5 gpc1755 (
      {stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71], stage1_23[72]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[20],stage2_25[24],stage2_24[24],stage2_23[35]}
   );
   gpc606_5 gpc1756 (
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[8],stage2_26[21],stage2_25[25],stage2_24[25]}
   );
   gpc615_5 gpc1757 (
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88]},
      {stage1_25[48]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[9],stage2_26[22],stage2_25[26],stage2_24[26]}
   );
   gpc615_5 gpc1758 (
      {stage1_24[89], stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93]},
      {stage1_25[49]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[10],stage2_26[23],stage2_25[27],stage2_24[27]}
   );
   gpc615_5 gpc1759 (
      {stage1_24[94], stage1_24[95], stage1_24[96], stage1_24[97], stage1_24[98]},
      {stage1_25[50]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[11],stage2_26[24],stage2_25[28],stage2_24[28]}
   );
   gpc615_5 gpc1760 (
      {stage1_24[99], stage1_24[100], stage1_24[101], stage1_24[102], stage1_24[103]},
      {stage1_25[51]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[12],stage2_26[25],stage2_25[29],stage2_24[29]}
   );
   gpc615_5 gpc1761 (
      {stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107], stage1_24[108]},
      {stage1_25[52]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[13],stage2_26[26],stage2_25[30],stage2_24[30]}
   );
   gpc615_5 gpc1762 (
      {stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage1_25[53]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[14],stage2_26[27],stage2_25[31],stage2_24[31]}
   );
   gpc615_5 gpc1763 (
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118]},
      {stage1_25[54]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[15],stage2_26[28],stage2_25[32],stage2_24[32]}
   );
   gpc615_5 gpc1764 (
      {stage1_24[119], stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123]},
      {stage1_25[55]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[16],stage2_26[29],stage2_25[33],stage2_24[33]}
   );
   gpc615_5 gpc1765 (
      {stage1_24[124], stage1_24[125], stage1_24[126], stage1_24[127], stage1_24[128]},
      {stage1_25[56]},
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage2_28[9],stage2_27[17],stage2_26[30],stage2_25[34],stage2_24[34]}
   );
   gpc615_5 gpc1766 (
      {stage1_24[129], stage1_24[130], stage1_24[131], stage1_24[132], stage1_24[133]},
      {stage1_25[57]},
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage2_28[10],stage2_27[18],stage2_26[31],stage2_25[35],stage2_24[35]}
   );
   gpc615_5 gpc1767 (
      {stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137], stage1_24[138]},
      {stage1_25[58]},
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70], stage1_26[71]},
      {stage2_28[11],stage2_27[19],stage2_26[32],stage2_25[36],stage2_24[36]}
   );
   gpc615_5 gpc1768 (
      {stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143]},
      {stage1_25[59]},
      {stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77]},
      {stage2_28[12],stage2_27[20],stage2_26[33],stage2_25[37],stage2_24[37]}
   );
   gpc615_5 gpc1769 (
      {stage1_24[144], stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148]},
      {stage1_25[60]},
      {stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83]},
      {stage2_28[13],stage2_27[21],stage2_26[34],stage2_25[38],stage2_24[38]}
   );
   gpc615_5 gpc1770 (
      {stage1_24[149], stage1_24[150], stage1_24[151], stage1_24[152], stage1_24[153]},
      {stage1_25[61]},
      {stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage2_28[14],stage2_27[22],stage2_26[35],stage2_25[39],stage2_24[39]}
   );
   gpc615_5 gpc1771 (
      {stage1_24[154], stage1_24[155], stage1_24[156], stage1_24[157], stage1_24[158]},
      {stage1_25[62]},
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage2_28[15],stage2_27[23],stage2_26[36],stage2_25[40],stage2_24[40]}
   );
   gpc615_5 gpc1772 (
      {stage1_24[159], stage1_24[160], stage1_24[161], stage1_24[162], stage1_24[163]},
      {stage1_25[63]},
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100], stage1_26[101]},
      {stage2_28[16],stage2_27[24],stage2_26[37],stage2_25[41],stage2_24[41]}
   );
   gpc615_5 gpc1773 (
      {stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167], stage1_24[168]},
      {stage1_25[64]},
      {stage1_26[102], stage1_26[103], stage1_26[104], stage1_26[105], stage1_26[106], stage1_26[107]},
      {stage2_28[17],stage2_27[25],stage2_26[38],stage2_25[42],stage2_24[42]}
   );
   gpc615_5 gpc1774 (
      {stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage1_25[65]},
      {stage1_26[108], stage1_26[109], stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113]},
      {stage2_28[18],stage2_27[26],stage2_26[39],stage2_25[43],stage2_24[43]}
   );
   gpc615_5 gpc1775 (
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178]},
      {stage1_25[66]},
      {stage1_26[114], stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119]},
      {stage2_28[19],stage2_27[27],stage2_26[40],stage2_25[44],stage2_24[44]}
   );
   gpc615_5 gpc1776 (
      {stage1_24[179], stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183]},
      {stage1_25[67]},
      {stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage2_28[20],stage2_27[28],stage2_26[41],stage2_25[45],stage2_24[45]}
   );
   gpc615_5 gpc1777 (
      {stage1_24[184], stage1_24[185], stage1_24[186], stage1_24[187], stage1_24[188]},
      {stage1_25[68]},
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130], stage1_26[131]},
      {stage2_28[21],stage2_27[29],stage2_26[42],stage2_25[46],stage2_24[46]}
   );
   gpc615_5 gpc1778 (
      {stage1_24[189], stage1_24[190], stage1_24[191], stage1_24[192], stage1_24[193]},
      {stage1_25[69]},
      {stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135], stage1_26[136], stage1_26[137]},
      {stage2_28[22],stage2_27[30],stage2_26[43],stage2_25[47],stage2_24[47]}
   );
   gpc615_5 gpc1779 (
      {stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197], stage1_24[198]},
      {stage1_25[70]},
      {stage1_26[138], stage1_26[139], stage1_26[140], stage1_26[141], stage1_26[142], stage1_26[143]},
      {stage2_28[23],stage2_27[31],stage2_26[44],stage2_25[48],stage2_24[48]}
   );
   gpc615_5 gpc1780 (
      {stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203]},
      {stage1_25[71]},
      {stage1_26[144], stage1_26[145], stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149]},
      {stage2_28[24],stage2_27[32],stage2_26[45],stage2_25[49],stage2_24[49]}
   );
   gpc615_5 gpc1781 (
      {stage1_24[204], stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208]},
      {stage1_25[72]},
      {stage1_26[150], stage1_26[151], stage1_26[152], stage1_26[153], stage1_26[154], stage1_26[155]},
      {stage2_28[25],stage2_27[33],stage2_26[46],stage2_25[50],stage2_24[50]}
   );
   gpc615_5 gpc1782 (
      {stage1_24[209], stage1_24[210], stage1_24[211], stage1_24[212], stage1_24[213]},
      {stage1_25[73]},
      {stage1_26[156], stage1_26[157], stage1_26[158], stage1_26[159], stage1_26[160], stage1_26[161]},
      {stage2_28[26],stage2_27[34],stage2_26[47],stage2_25[51],stage2_24[51]}
   );
   gpc615_5 gpc1783 (
      {stage1_24[214], stage1_24[215], stage1_24[216], stage1_24[217], stage1_24[218]},
      {stage1_25[74]},
      {stage1_26[162], stage1_26[163], stage1_26[164], stage1_26[165], stage1_26[166], stage1_26[167]},
      {stage2_28[27],stage2_27[35],stage2_26[48],stage2_25[52],stage2_24[52]}
   );
   gpc615_5 gpc1784 (
      {stage1_24[219], stage1_24[220], stage1_24[221], stage1_24[222], stage1_24[223]},
      {stage1_25[75]},
      {stage1_26[168], stage1_26[169], stage1_26[170], stage1_26[171], stage1_26[172], stage1_26[173]},
      {stage2_28[28],stage2_27[36],stage2_26[49],stage2_25[53],stage2_24[53]}
   );
   gpc615_5 gpc1785 (
      {stage1_24[224], stage1_24[225], stage1_24[226], stage1_24[227], stage1_24[228]},
      {stage1_25[76]},
      {stage1_26[174], stage1_26[175], stage1_26[176], stage1_26[177], stage1_26[178], stage1_26[179]},
      {stage2_28[29],stage2_27[37],stage2_26[50],stage2_25[54],stage2_24[54]}
   );
   gpc615_5 gpc1786 (
      {stage1_24[229], stage1_24[230], stage1_24[231], stage1_24[232], stage1_24[233]},
      {stage1_25[77]},
      {stage1_26[180], stage1_26[181], stage1_26[182], stage1_26[183], stage1_26[184], stage1_26[185]},
      {stage2_28[30],stage2_27[38],stage2_26[51],stage2_25[55],stage2_24[55]}
   );
   gpc615_5 gpc1787 (
      {stage1_24[234], stage1_24[235], stage1_24[236], stage1_24[237], stage1_24[238]},
      {stage1_25[78]},
      {stage1_26[186], stage1_26[187], stage1_26[188], stage1_26[189], stage1_26[190], stage1_26[191]},
      {stage2_28[31],stage2_27[39],stage2_26[52],stage2_25[56],stage2_24[56]}
   );
   gpc615_5 gpc1788 (
      {stage1_24[239], stage1_24[240], stage1_24[241], stage1_24[242], stage1_24[243]},
      {stage1_25[79]},
      {stage1_26[192], stage1_26[193], stage1_26[194], stage1_26[195], stage1_26[196], stage1_26[197]},
      {stage2_28[32],stage2_27[40],stage2_26[53],stage2_25[57],stage2_24[57]}
   );
   gpc615_5 gpc1789 (
      {stage1_24[244], stage1_24[245], stage1_24[246], stage1_24[247], stage1_24[248]},
      {stage1_25[80]},
      {stage1_26[198], stage1_26[199], stage1_26[200], stage1_26[201], stage1_26[202], stage1_26[203]},
      {stage2_28[33],stage2_27[41],stage2_26[54],stage2_25[58],stage2_24[58]}
   );
   gpc606_5 gpc1790 (
      {stage1_25[81], stage1_25[82], stage1_25[83], stage1_25[84], stage1_25[85], stage1_25[86]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[34],stage2_27[42],stage2_26[55],stage2_25[59]}
   );
   gpc606_5 gpc1791 (
      {stage1_25[87], stage1_25[88], stage1_25[89], stage1_25[90], stage1_25[91], stage1_25[92]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[35],stage2_27[43],stage2_26[56],stage2_25[60]}
   );
   gpc606_5 gpc1792 (
      {stage1_25[93], stage1_25[94], stage1_25[95], stage1_25[96], stage1_25[97], stage1_25[98]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[36],stage2_27[44],stage2_26[57],stage2_25[61]}
   );
   gpc606_5 gpc1793 (
      {stage1_25[99], stage1_25[100], stage1_25[101], stage1_25[102], stage1_25[103], stage1_25[104]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[37],stage2_27[45],stage2_26[58],stage2_25[62]}
   );
   gpc606_5 gpc1794 (
      {stage1_25[105], stage1_25[106], stage1_25[107], stage1_25[108], stage1_25[109], stage1_25[110]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[38],stage2_27[46],stage2_26[59],stage2_25[63]}
   );
   gpc606_5 gpc1795 (
      {stage1_25[111], stage1_25[112], stage1_25[113], stage1_25[114], stage1_25[115], stage1_25[116]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[39],stage2_27[47],stage2_26[60],stage2_25[64]}
   );
   gpc615_5 gpc1796 (
      {stage1_26[204], stage1_26[205], stage1_26[206], stage1_26[207], stage1_26[208]},
      {stage1_27[36]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[6],stage2_28[40],stage2_27[48],stage2_26[61]}
   );
   gpc615_5 gpc1797 (
      {stage1_26[209], stage1_26[210], stage1_26[211], stage1_26[212], stage1_26[213]},
      {stage1_27[37]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[7],stage2_28[41],stage2_27[49],stage2_26[62]}
   );
   gpc615_5 gpc1798 (
      {stage1_26[214], stage1_26[215], stage1_26[216], stage1_26[217], stage1_26[218]},
      {stage1_27[38]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[8],stage2_28[42],stage2_27[50],stage2_26[63]}
   );
   gpc615_5 gpc1799 (
      {stage1_26[219], stage1_26[220], stage1_26[221], stage1_26[222], stage1_26[223]},
      {stage1_27[39]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[9],stage2_28[43],stage2_27[51],stage2_26[64]}
   );
   gpc615_5 gpc1800 (
      {stage1_26[224], stage1_26[225], stage1_26[226], stage1_26[227], stage1_26[228]},
      {stage1_27[40]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[10],stage2_28[44],stage2_27[52],stage2_26[65]}
   );
   gpc615_5 gpc1801 (
      {stage1_26[229], stage1_26[230], stage1_26[231], stage1_26[232], stage1_26[233]},
      {stage1_27[41]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[11],stage2_28[45],stage2_27[53],stage2_26[66]}
   );
   gpc615_5 gpc1802 (
      {stage1_26[234], stage1_26[235], stage1_26[236], 1'b0, 1'b0},
      {stage1_27[42]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[12],stage2_28[46],stage2_27[54],stage2_26[67]}
   );
   gpc615_5 gpc1803 (
      {stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage1_28[42]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[7],stage2_29[13],stage2_28[47],stage2_27[55]}
   );
   gpc615_5 gpc1804 (
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_28[43]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[8],stage2_29[14],stage2_28[48],stage2_27[56]}
   );
   gpc615_5 gpc1805 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[44]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[9],stage2_29[15],stage2_28[49],stage2_27[57]}
   );
   gpc615_5 gpc1806 (
      {stage1_27[58], stage1_27[59], stage1_27[60], stage1_27[61], stage1_27[62]},
      {stage1_28[45]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[10],stage2_29[16],stage2_28[50],stage2_27[58]}
   );
   gpc615_5 gpc1807 (
      {stage1_27[63], stage1_27[64], stage1_27[65], stage1_27[66], stage1_27[67]},
      {stage1_28[46]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[11],stage2_29[17],stage2_28[51],stage2_27[59]}
   );
   gpc615_5 gpc1808 (
      {stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71], stage1_27[72]},
      {stage1_28[47]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[12],stage2_29[18],stage2_28[52],stage2_27[60]}
   );
   gpc606_5 gpc1809 (
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[6],stage2_30[13],stage2_29[19],stage2_28[53]}
   );
   gpc606_5 gpc1810 (
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[7],stage2_30[14],stage2_29[20],stage2_28[54]}
   );
   gpc606_5 gpc1811 (
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[8],stage2_30[15],stage2_29[21],stage2_28[55]}
   );
   gpc606_5 gpc1812 (
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[9],stage2_30[16],stage2_29[22],stage2_28[56]}
   );
   gpc606_5 gpc1813 (
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[10],stage2_30[17],stage2_29[23],stage2_28[57]}
   );
   gpc606_5 gpc1814 (
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[11],stage2_30[18],stage2_29[24],stage2_28[58]}
   );
   gpc606_5 gpc1815 (
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[12],stage2_30[19],stage2_29[25],stage2_28[59]}
   );
   gpc606_5 gpc1816 (
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[7],stage2_31[13],stage2_30[20],stage2_29[26]}
   );
   gpc606_5 gpc1817 (
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[8],stage2_31[14],stage2_30[21],stage2_29[27]}
   );
   gpc606_5 gpc1818 (
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[9],stage2_31[15],stage2_30[22],stage2_29[28]}
   );
   gpc606_5 gpc1819 (
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[10],stage2_31[16],stage2_30[23],stage2_29[29]}
   );
   gpc606_5 gpc1820 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[11],stage2_31[17],stage2_30[24],stage2_29[30]}
   );
   gpc606_5 gpc1821 (
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[12],stage2_31[18],stage2_30[25],stage2_29[31]}
   );
   gpc606_5 gpc1822 (
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[13],stage2_31[19],stage2_30[26],stage2_29[32]}
   );
   gpc606_5 gpc1823 (
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[14],stage2_31[20],stage2_30[27],stage2_29[33]}
   );
   gpc606_5 gpc1824 (
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[15],stage2_31[21],stage2_30[28],stage2_29[34]}
   );
   gpc606_5 gpc1825 (
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[16],stage2_31[22],stage2_30[29],stage2_29[35]}
   );
   gpc606_5 gpc1826 (
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage2_33[10],stage2_32[17],stage2_31[23],stage2_30[30],stage2_29[36]}
   );
   gpc606_5 gpc1827 (
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69], stage1_31[70], stage1_31[71]},
      {stage2_33[11],stage2_32[18],stage2_31[24],stage2_30[31],stage2_29[37]}
   );
   gpc606_5 gpc1828 (
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage1_31[72], stage1_31[73], stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77]},
      {stage2_33[12],stage2_32[19],stage2_31[25],stage2_30[32],stage2_29[38]}
   );
   gpc606_5 gpc1829 (
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], 1'b0, 1'b0},
      {stage1_31[78], stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage2_33[13],stage2_32[20],stage2_31[26],stage2_30[33],stage2_29[39]}
   );
   gpc615_5 gpc1830 (
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46]},
      {stage1_31[84]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[14],stage2_32[21],stage2_31[27],stage2_30[34]}
   );
   gpc615_5 gpc1831 (
      {stage1_30[47], stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51]},
      {stage1_31[85]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[15],stage2_32[22],stage2_31[28],stage2_30[35]}
   );
   gpc615_5 gpc1832 (
      {stage1_30[52], stage1_30[53], stage1_30[54], stage1_30[55], stage1_30[56]},
      {stage1_31[86]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[16],stage2_32[23],stage2_31[29],stage2_30[36]}
   );
   gpc615_5 gpc1833 (
      {stage1_30[57], stage1_30[58], stage1_30[59], stage1_30[60], stage1_30[61]},
      {stage1_31[87]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[17],stage2_32[24],stage2_31[30],stage2_30[37]}
   );
   gpc615_5 gpc1834 (
      {stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65], stage1_30[66]},
      {stage1_31[88]},
      {stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28], stage1_32[29]},
      {stage2_34[4],stage2_33[18],stage2_32[25],stage2_31[31],stage2_30[38]}
   );
   gpc615_5 gpc1835 (
      {stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_31[89]},
      {stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34], stage1_32[35]},
      {stage2_34[5],stage2_33[19],stage2_32[26],stage2_31[32],stage2_30[39]}
   );
   gpc615_5 gpc1836 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76]},
      {stage1_31[90]},
      {stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41]},
      {stage2_34[6],stage2_33[20],stage2_32[27],stage2_31[33],stage2_30[40]}
   );
   gpc615_5 gpc1837 (
      {stage1_30[77], stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81]},
      {stage1_31[91]},
      {stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47]},
      {stage2_34[7],stage2_33[21],stage2_32[28],stage2_31[34],stage2_30[41]}
   );
   gpc615_5 gpc1838 (
      {stage1_30[82], stage1_30[83], stage1_30[84], stage1_30[85], stage1_30[86]},
      {stage1_31[92]},
      {stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53]},
      {stage2_34[8],stage2_33[22],stage2_32[29],stage2_31[35],stage2_30[42]}
   );
   gpc615_5 gpc1839 (
      {stage1_30[87], stage1_30[88], stage1_30[89], stage1_30[90], stage1_30[91]},
      {stage1_31[93]},
      {stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59]},
      {stage2_34[9],stage2_33[23],stage2_32[30],stage2_31[36],stage2_30[43]}
   );
   gpc615_5 gpc1840 (
      {stage1_30[92], stage1_30[93], stage1_30[94], stage1_30[95], stage1_30[96]},
      {stage1_31[94]},
      {stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65]},
      {stage2_34[10],stage2_33[24],stage2_32[31],stage2_31[37],stage2_30[44]}
   );
   gpc606_5 gpc1841 (
      {stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99], stage1_31[100]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[11],stage2_33[25],stage2_32[32],stage2_31[38]}
   );
   gpc606_5 gpc1842 (
      {stage1_31[101], stage1_31[102], stage1_31[103], stage1_31[104], stage1_31[105], stage1_31[106]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[12],stage2_33[26],stage2_32[33],stage2_31[39]}
   );
   gpc606_5 gpc1843 (
      {stage1_31[107], stage1_31[108], stage1_31[109], stage1_31[110], stage1_31[111], stage1_31[112]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[13],stage2_33[27],stage2_32[34],stage2_31[40]}
   );
   gpc606_5 gpc1844 (
      {stage1_31[113], stage1_31[114], stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[14],stage2_33[28],stage2_32[35],stage2_31[41]}
   );
   gpc615_5 gpc1845 (
      {stage1_31[119], stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123]},
      {stage1_32[66]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[15],stage2_33[29],stage2_32[36],stage2_31[42]}
   );
   gpc615_5 gpc1846 (
      {stage1_31[124], stage1_31[125], stage1_31[126], stage1_31[127], stage1_31[128]},
      {stage1_32[67]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], 1'b0, 1'b0},
      {stage2_35[5],stage2_34[16],stage2_33[30],stage2_32[37],stage2_31[43]}
   );
   gpc1_1 gpc1847 (
      {stage1_0[39]},
      {stage2_0[13]}
   );
   gpc1_1 gpc1848 (
      {stage1_0[40]},
      {stage2_0[14]}
   );
   gpc1_1 gpc1849 (
      {stage1_0[41]},
      {stage2_0[15]}
   );
   gpc1_1 gpc1850 (
      {stage1_0[42]},
      {stage2_0[16]}
   );
   gpc1_1 gpc1851 (
      {stage1_0[43]},
      {stage2_0[17]}
   );
   gpc1_1 gpc1852 (
      {stage1_0[44]},
      {stage2_0[18]}
   );
   gpc1_1 gpc1853 (
      {stage1_0[45]},
      {stage2_0[19]}
   );
   gpc1_1 gpc1854 (
      {stage1_0[46]},
      {stage2_0[20]}
   );
   gpc1_1 gpc1855 (
      {stage1_0[47]},
      {stage2_0[21]}
   );
   gpc1_1 gpc1856 (
      {stage1_0[48]},
      {stage2_0[22]}
   );
   gpc1_1 gpc1857 (
      {stage1_0[49]},
      {stage2_0[23]}
   );
   gpc1_1 gpc1858 (
      {stage1_1[78]},
      {stage2_1[13]}
   );
   gpc1_1 gpc1859 (
      {stage1_1[79]},
      {stage2_1[14]}
   );
   gpc1_1 gpc1860 (
      {stage1_1[80]},
      {stage2_1[15]}
   );
   gpc1_1 gpc1861 (
      {stage1_1[81]},
      {stage2_1[16]}
   );
   gpc1_1 gpc1862 (
      {stage1_1[82]},
      {stage2_1[17]}
   );
   gpc1_1 gpc1863 (
      {stage1_1[83]},
      {stage2_1[18]}
   );
   gpc1_1 gpc1864 (
      {stage1_1[84]},
      {stage2_1[19]}
   );
   gpc1_1 gpc1865 (
      {stage1_1[85]},
      {stage2_1[20]}
   );
   gpc1_1 gpc1866 (
      {stage1_1[86]},
      {stage2_1[21]}
   );
   gpc1_1 gpc1867 (
      {stage1_1[87]},
      {stage2_1[22]}
   );
   gpc1_1 gpc1868 (
      {stage1_1[88]},
      {stage2_1[23]}
   );
   gpc1_1 gpc1869 (
      {stage1_1[89]},
      {stage2_1[24]}
   );
   gpc1_1 gpc1870 (
      {stage1_1[90]},
      {stage2_1[25]}
   );
   gpc1_1 gpc1871 (
      {stage1_1[91]},
      {stage2_1[26]}
   );
   gpc1_1 gpc1872 (
      {stage1_1[92]},
      {stage2_1[27]}
   );
   gpc1_1 gpc1873 (
      {stage1_1[93]},
      {stage2_1[28]}
   );
   gpc1_1 gpc1874 (
      {stage1_1[94]},
      {stage2_1[29]}
   );
   gpc1_1 gpc1875 (
      {stage1_1[95]},
      {stage2_1[30]}
   );
   gpc1_1 gpc1876 (
      {stage1_1[96]},
      {stage2_1[31]}
   );
   gpc1_1 gpc1877 (
      {stage1_1[97]},
      {stage2_1[32]}
   );
   gpc1_1 gpc1878 (
      {stage1_2[84]},
      {stage2_2[27]}
   );
   gpc1_1 gpc1879 (
      {stage1_2[85]},
      {stage2_2[28]}
   );
   gpc1_1 gpc1880 (
      {stage1_2[86]},
      {stage2_2[29]}
   );
   gpc1_1 gpc1881 (
      {stage1_2[87]},
      {stage2_2[30]}
   );
   gpc1_1 gpc1882 (
      {stage1_2[88]},
      {stage2_2[31]}
   );
   gpc1_1 gpc1883 (
      {stage1_2[89]},
      {stage2_2[32]}
   );
   gpc1_1 gpc1884 (
      {stage1_2[90]},
      {stage2_2[33]}
   );
   gpc1_1 gpc1885 (
      {stage1_2[91]},
      {stage2_2[34]}
   );
   gpc1_1 gpc1886 (
      {stage1_3[87]},
      {stage2_3[39]}
   );
   gpc1_1 gpc1887 (
      {stage1_3[88]},
      {stage2_3[40]}
   );
   gpc1_1 gpc1888 (
      {stage1_3[89]},
      {stage2_3[41]}
   );
   gpc1_1 gpc1889 (
      {stage1_3[90]},
      {stage2_3[42]}
   );
   gpc1_1 gpc1890 (
      {stage1_4[118]},
      {stage2_4[43]}
   );
   gpc1_1 gpc1891 (
      {stage1_4[119]},
      {stage2_4[44]}
   );
   gpc1_1 gpc1892 (
      {stage1_4[120]},
      {stage2_4[45]}
   );
   gpc1_1 gpc1893 (
      {stage1_4[121]},
      {stage2_4[46]}
   );
   gpc1_1 gpc1894 (
      {stage1_4[122]},
      {stage2_4[47]}
   );
   gpc1_1 gpc1895 (
      {stage1_4[123]},
      {stage2_4[48]}
   );
   gpc1_1 gpc1896 (
      {stage1_4[124]},
      {stage2_4[49]}
   );
   gpc1_1 gpc1897 (
      {stage1_4[125]},
      {stage2_4[50]}
   );
   gpc1_1 gpc1898 (
      {stage1_4[126]},
      {stage2_4[51]}
   );
   gpc1_1 gpc1899 (
      {stage1_4[127]},
      {stage2_4[52]}
   );
   gpc1_1 gpc1900 (
      {stage1_4[128]},
      {stage2_4[53]}
   );
   gpc1_1 gpc1901 (
      {stage1_4[129]},
      {stage2_4[54]}
   );
   gpc1_1 gpc1902 (
      {stage1_4[130]},
      {stage2_4[55]}
   );
   gpc1_1 gpc1903 (
      {stage1_4[131]},
      {stage2_4[56]}
   );
   gpc1_1 gpc1904 (
      {stage1_4[132]},
      {stage2_4[57]}
   );
   gpc1_1 gpc1905 (
      {stage1_4[133]},
      {stage2_4[58]}
   );
   gpc1_1 gpc1906 (
      {stage1_4[134]},
      {stage2_4[59]}
   );
   gpc1_1 gpc1907 (
      {stage1_4[135]},
      {stage2_4[60]}
   );
   gpc1_1 gpc1908 (
      {stage1_4[136]},
      {stage2_4[61]}
   );
   gpc1_1 gpc1909 (
      {stage1_4[137]},
      {stage2_4[62]}
   );
   gpc1_1 gpc1910 (
      {stage1_4[138]},
      {stage2_4[63]}
   );
   gpc1_1 gpc1911 (
      {stage1_4[139]},
      {stage2_4[64]}
   );
   gpc1_1 gpc1912 (
      {stage1_4[140]},
      {stage2_4[65]}
   );
   gpc1_1 gpc1913 (
      {stage1_4[141]},
      {stage2_4[66]}
   );
   gpc1_1 gpc1914 (
      {stage1_4[142]},
      {stage2_4[67]}
   );
   gpc1_1 gpc1915 (
      {stage1_4[143]},
      {stage2_4[68]}
   );
   gpc1_1 gpc1916 (
      {stage1_4[144]},
      {stage2_4[69]}
   );
   gpc1_1 gpc1917 (
      {stage1_4[145]},
      {stage2_4[70]}
   );
   gpc1_1 gpc1918 (
      {stage1_4[146]},
      {stage2_4[71]}
   );
   gpc1_1 gpc1919 (
      {stage1_4[147]},
      {stage2_4[72]}
   );
   gpc1_1 gpc1920 (
      {stage1_4[148]},
      {stage2_4[73]}
   );
   gpc1_1 gpc1921 (
      {stage1_5[122]},
      {stage2_5[38]}
   );
   gpc1_1 gpc1922 (
      {stage1_5[123]},
      {stage2_5[39]}
   );
   gpc1_1 gpc1923 (
      {stage1_5[124]},
      {stage2_5[40]}
   );
   gpc1_1 gpc1924 (
      {stage1_5[125]},
      {stage2_5[41]}
   );
   gpc1_1 gpc1925 (
      {stage1_7[92]},
      {stage2_7[45]}
   );
   gpc1_1 gpc1926 (
      {stage1_7[93]},
      {stage2_7[46]}
   );
   gpc1_1 gpc1927 (
      {stage1_7[94]},
      {stage2_7[47]}
   );
   gpc1_1 gpc1928 (
      {stage1_7[95]},
      {stage2_7[48]}
   );
   gpc1_1 gpc1929 (
      {stage1_7[96]},
      {stage2_7[49]}
   );
   gpc1_1 gpc1930 (
      {stage1_7[97]},
      {stage2_7[50]}
   );
   gpc1_1 gpc1931 (
      {stage1_7[98]},
      {stage2_7[51]}
   );
   gpc1_1 gpc1932 (
      {stage1_7[99]},
      {stage2_7[52]}
   );
   gpc1_1 gpc1933 (
      {stage1_7[100]},
      {stage2_7[53]}
   );
   gpc1_1 gpc1934 (
      {stage1_8[96]},
      {stage2_8[32]}
   );
   gpc1_1 gpc1935 (
      {stage1_8[97]},
      {stage2_8[33]}
   );
   gpc1_1 gpc1936 (
      {stage1_8[98]},
      {stage2_8[34]}
   );
   gpc1_1 gpc1937 (
      {stage1_8[99]},
      {stage2_8[35]}
   );
   gpc1_1 gpc1938 (
      {stage1_8[100]},
      {stage2_8[36]}
   );
   gpc1_1 gpc1939 (
      {stage1_8[101]},
      {stage2_8[37]}
   );
   gpc1_1 gpc1940 (
      {stage1_8[102]},
      {stage2_8[38]}
   );
   gpc1_1 gpc1941 (
      {stage1_8[103]},
      {stage2_8[39]}
   );
   gpc1_1 gpc1942 (
      {stage1_8[104]},
      {stage2_8[40]}
   );
   gpc1_1 gpc1943 (
      {stage1_8[105]},
      {stage2_8[41]}
   );
   gpc1_1 gpc1944 (
      {stage1_8[106]},
      {stage2_8[42]}
   );
   gpc1_1 gpc1945 (
      {stage1_8[107]},
      {stage2_8[43]}
   );
   gpc1_1 gpc1946 (
      {stage1_8[108]},
      {stage2_8[44]}
   );
   gpc1_1 gpc1947 (
      {stage1_8[109]},
      {stage2_8[45]}
   );
   gpc1_1 gpc1948 (
      {stage1_8[110]},
      {stage2_8[46]}
   );
   gpc1_1 gpc1949 (
      {stage1_8[111]},
      {stage2_8[47]}
   );
   gpc1_1 gpc1950 (
      {stage1_8[112]},
      {stage2_8[48]}
   );
   gpc1_1 gpc1951 (
      {stage1_8[113]},
      {stage2_8[49]}
   );
   gpc1_1 gpc1952 (
      {stage1_8[114]},
      {stage2_8[50]}
   );
   gpc1_1 gpc1953 (
      {stage1_8[115]},
      {stage2_8[51]}
   );
   gpc1_1 gpc1954 (
      {stage1_8[116]},
      {stage2_8[52]}
   );
   gpc1_1 gpc1955 (
      {stage1_8[117]},
      {stage2_8[53]}
   );
   gpc1_1 gpc1956 (
      {stage1_8[118]},
      {stage2_8[54]}
   );
   gpc1_1 gpc1957 (
      {stage1_8[119]},
      {stage2_8[55]}
   );
   gpc1_1 gpc1958 (
      {stage1_9[107]},
      {stage2_9[41]}
   );
   gpc1_1 gpc1959 (
      {stage1_9[108]},
      {stage2_9[42]}
   );
   gpc1_1 gpc1960 (
      {stage1_9[109]},
      {stage2_9[43]}
   );
   gpc1_1 gpc1961 (
      {stage1_9[110]},
      {stage2_9[44]}
   );
   gpc1_1 gpc1962 (
      {stage1_9[111]},
      {stage2_9[45]}
   );
   gpc1_1 gpc1963 (
      {stage1_9[112]},
      {stage2_9[46]}
   );
   gpc1_1 gpc1964 (
      {stage1_9[113]},
      {stage2_9[47]}
   );
   gpc1_1 gpc1965 (
      {stage1_9[114]},
      {stage2_9[48]}
   );
   gpc1_1 gpc1966 (
      {stage1_9[115]},
      {stage2_9[49]}
   );
   gpc1_1 gpc1967 (
      {stage1_9[116]},
      {stage2_9[50]}
   );
   gpc1_1 gpc1968 (
      {stage1_9[117]},
      {stage2_9[51]}
   );
   gpc1_1 gpc1969 (
      {stage1_9[118]},
      {stage2_9[52]}
   );
   gpc1_1 gpc1970 (
      {stage1_9[119]},
      {stage2_9[53]}
   );
   gpc1_1 gpc1971 (
      {stage1_9[120]},
      {stage2_9[54]}
   );
   gpc1_1 gpc1972 (
      {stage1_9[121]},
      {stage2_9[55]}
   );
   gpc1_1 gpc1973 (
      {stage1_9[122]},
      {stage2_9[56]}
   );
   gpc1_1 gpc1974 (
      {stage1_9[123]},
      {stage2_9[57]}
   );
   gpc1_1 gpc1975 (
      {stage1_9[124]},
      {stage2_9[58]}
   );
   gpc1_1 gpc1976 (
      {stage1_9[125]},
      {stage2_9[59]}
   );
   gpc1_1 gpc1977 (
      {stage1_9[126]},
      {stage2_9[60]}
   );
   gpc1_1 gpc1978 (
      {stage1_9[127]},
      {stage2_9[61]}
   );
   gpc1_1 gpc1979 (
      {stage1_9[128]},
      {stage2_9[62]}
   );
   gpc1_1 gpc1980 (
      {stage1_9[129]},
      {stage2_9[63]}
   );
   gpc1_1 gpc1981 (
      {stage1_9[130]},
      {stage2_9[64]}
   );
   gpc1_1 gpc1982 (
      {stage1_9[131]},
      {stage2_9[65]}
   );
   gpc1_1 gpc1983 (
      {stage1_11[127]},
      {stage2_11[45]}
   );
   gpc1_1 gpc1984 (
      {stage1_11[128]},
      {stage2_11[46]}
   );
   gpc1_1 gpc1985 (
      {stage1_11[129]},
      {stage2_11[47]}
   );
   gpc1_1 gpc1986 (
      {stage1_11[130]},
      {stage2_11[48]}
   );
   gpc1_1 gpc1987 (
      {stage1_11[131]},
      {stage2_11[49]}
   );
   gpc1_1 gpc1988 (
      {stage1_11[132]},
      {stage2_11[50]}
   );
   gpc1_1 gpc1989 (
      {stage1_11[133]},
      {stage2_11[51]}
   );
   gpc1_1 gpc1990 (
      {stage1_11[134]},
      {stage2_11[52]}
   );
   gpc1_1 gpc1991 (
      {stage1_11[135]},
      {stage2_11[53]}
   );
   gpc1_1 gpc1992 (
      {stage1_11[136]},
      {stage2_11[54]}
   );
   gpc1_1 gpc1993 (
      {stage1_11[137]},
      {stage2_11[55]}
   );
   gpc1_1 gpc1994 (
      {stage1_11[138]},
      {stage2_11[56]}
   );
   gpc1_1 gpc1995 (
      {stage1_11[139]},
      {stage2_11[57]}
   );
   gpc1_1 gpc1996 (
      {stage1_12[173]},
      {stage2_12[50]}
   );
   gpc1_1 gpc1997 (
      {stage1_12[174]},
      {stage2_12[51]}
   );
   gpc1_1 gpc1998 (
      {stage1_12[175]},
      {stage2_12[52]}
   );
   gpc1_1 gpc1999 (
      {stage1_12[176]},
      {stage2_12[53]}
   );
   gpc1_1 gpc2000 (
      {stage1_12[177]},
      {stage2_12[54]}
   );
   gpc1_1 gpc2001 (
      {stage1_12[178]},
      {stage2_12[55]}
   );
   gpc1_1 gpc2002 (
      {stage1_12[179]},
      {stage2_12[56]}
   );
   gpc1_1 gpc2003 (
      {stage1_12[180]},
      {stage2_12[57]}
   );
   gpc1_1 gpc2004 (
      {stage1_12[181]},
      {stage2_12[58]}
   );
   gpc1_1 gpc2005 (
      {stage1_12[182]},
      {stage2_12[59]}
   );
   gpc1_1 gpc2006 (
      {stage1_12[183]},
      {stage2_12[60]}
   );
   gpc1_1 gpc2007 (
      {stage1_12[184]},
      {stage2_12[61]}
   );
   gpc1_1 gpc2008 (
      {stage1_12[185]},
      {stage2_12[62]}
   );
   gpc1_1 gpc2009 (
      {stage1_12[186]},
      {stage2_12[63]}
   );
   gpc1_1 gpc2010 (
      {stage1_12[187]},
      {stage2_12[64]}
   );
   gpc1_1 gpc2011 (
      {stage1_12[188]},
      {stage2_12[65]}
   );
   gpc1_1 gpc2012 (
      {stage1_12[189]},
      {stage2_12[66]}
   );
   gpc1_1 gpc2013 (
      {stage1_12[190]},
      {stage2_12[67]}
   );
   gpc1_1 gpc2014 (
      {stage1_12[191]},
      {stage2_12[68]}
   );
   gpc1_1 gpc2015 (
      {stage1_12[192]},
      {stage2_12[69]}
   );
   gpc1_1 gpc2016 (
      {stage1_12[193]},
      {stage2_12[70]}
   );
   gpc1_1 gpc2017 (
      {stage1_12[194]},
      {stage2_12[71]}
   );
   gpc1_1 gpc2018 (
      {stage1_12[195]},
      {stage2_12[72]}
   );
   gpc1_1 gpc2019 (
      {stage1_12[196]},
      {stage2_12[73]}
   );
   gpc1_1 gpc2020 (
      {stage1_12[197]},
      {stage2_12[74]}
   );
   gpc1_1 gpc2021 (
      {stage1_13[90]},
      {stage2_13[54]}
   );
   gpc1_1 gpc2022 (
      {stage1_13[91]},
      {stage2_13[55]}
   );
   gpc1_1 gpc2023 (
      {stage1_13[92]},
      {stage2_13[56]}
   );
   gpc1_1 gpc2024 (
      {stage1_14[66]},
      {stage2_14[42]}
   );
   gpc1_1 gpc2025 (
      {stage1_14[67]},
      {stage2_14[43]}
   );
   gpc1_1 gpc2026 (
      {stage1_14[68]},
      {stage2_14[44]}
   );
   gpc1_1 gpc2027 (
      {stage1_14[69]},
      {stage2_14[45]}
   );
   gpc1_1 gpc2028 (
      {stage1_14[70]},
      {stage2_14[46]}
   );
   gpc1_1 gpc2029 (
      {stage1_14[71]},
      {stage2_14[47]}
   );
   gpc1_1 gpc2030 (
      {stage1_14[72]},
      {stage2_14[48]}
   );
   gpc1_1 gpc2031 (
      {stage1_14[73]},
      {stage2_14[49]}
   );
   gpc1_1 gpc2032 (
      {stage1_14[74]},
      {stage2_14[50]}
   );
   gpc1_1 gpc2033 (
      {stage1_14[75]},
      {stage2_14[51]}
   );
   gpc1_1 gpc2034 (
      {stage1_14[76]},
      {stage2_14[52]}
   );
   gpc1_1 gpc2035 (
      {stage1_14[77]},
      {stage2_14[53]}
   );
   gpc1_1 gpc2036 (
      {stage1_14[78]},
      {stage2_14[54]}
   );
   gpc1_1 gpc2037 (
      {stage1_14[79]},
      {stage2_14[55]}
   );
   gpc1_1 gpc2038 (
      {stage1_14[80]},
      {stage2_14[56]}
   );
   gpc1_1 gpc2039 (
      {stage1_14[81]},
      {stage2_14[57]}
   );
   gpc1_1 gpc2040 (
      {stage1_14[82]},
      {stage2_14[58]}
   );
   gpc1_1 gpc2041 (
      {stage1_14[83]},
      {stage2_14[59]}
   );
   gpc1_1 gpc2042 (
      {stage1_14[84]},
      {stage2_14[60]}
   );
   gpc1_1 gpc2043 (
      {stage1_14[85]},
      {stage2_14[61]}
   );
   gpc1_1 gpc2044 (
      {stage1_14[86]},
      {stage2_14[62]}
   );
   gpc1_1 gpc2045 (
      {stage1_14[87]},
      {stage2_14[63]}
   );
   gpc1_1 gpc2046 (
      {stage1_14[88]},
      {stage2_14[64]}
   );
   gpc1_1 gpc2047 (
      {stage1_14[89]},
      {stage2_14[65]}
   );
   gpc1_1 gpc2048 (
      {stage1_14[90]},
      {stage2_14[66]}
   );
   gpc1_1 gpc2049 (
      {stage1_14[91]},
      {stage2_14[67]}
   );
   gpc1_1 gpc2050 (
      {stage1_14[92]},
      {stage2_14[68]}
   );
   gpc1_1 gpc2051 (
      {stage1_14[93]},
      {stage2_14[69]}
   );
   gpc1_1 gpc2052 (
      {stage1_14[94]},
      {stage2_14[70]}
   );
   gpc1_1 gpc2053 (
      {stage1_14[95]},
      {stage2_14[71]}
   );
   gpc1_1 gpc2054 (
      {stage1_14[96]},
      {stage2_14[72]}
   );
   gpc1_1 gpc2055 (
      {stage1_14[97]},
      {stage2_14[73]}
   );
   gpc1_1 gpc2056 (
      {stage1_14[98]},
      {stage2_14[74]}
   );
   gpc1_1 gpc2057 (
      {stage1_14[99]},
      {stage2_14[75]}
   );
   gpc1_1 gpc2058 (
      {stage1_14[100]},
      {stage2_14[76]}
   );
   gpc1_1 gpc2059 (
      {stage1_14[101]},
      {stage2_14[77]}
   );
   gpc1_1 gpc2060 (
      {stage1_14[102]},
      {stage2_14[78]}
   );
   gpc1_1 gpc2061 (
      {stage1_14[103]},
      {stage2_14[79]}
   );
   gpc1_1 gpc2062 (
      {stage1_14[104]},
      {stage2_14[80]}
   );
   gpc1_1 gpc2063 (
      {stage1_14[105]},
      {stage2_14[81]}
   );
   gpc1_1 gpc2064 (
      {stage1_14[106]},
      {stage2_14[82]}
   );
   gpc1_1 gpc2065 (
      {stage1_14[107]},
      {stage2_14[83]}
   );
   gpc1_1 gpc2066 (
      {stage1_14[108]},
      {stage2_14[84]}
   );
   gpc1_1 gpc2067 (
      {stage1_14[109]},
      {stage2_14[85]}
   );
   gpc1_1 gpc2068 (
      {stage1_14[110]},
      {stage2_14[86]}
   );
   gpc1_1 gpc2069 (
      {stage1_14[111]},
      {stage2_14[87]}
   );
   gpc1_1 gpc2070 (
      {stage1_14[112]},
      {stage2_14[88]}
   );
   gpc1_1 gpc2071 (
      {stage1_14[113]},
      {stage2_14[89]}
   );
   gpc1_1 gpc2072 (
      {stage1_15[84]},
      {stage2_15[38]}
   );
   gpc1_1 gpc2073 (
      {stage1_15[85]},
      {stage2_15[39]}
   );
   gpc1_1 gpc2074 (
      {stage1_15[86]},
      {stage2_15[40]}
   );
   gpc1_1 gpc2075 (
      {stage1_15[87]},
      {stage2_15[41]}
   );
   gpc1_1 gpc2076 (
      {stage1_15[88]},
      {stage2_15[42]}
   );
   gpc1_1 gpc2077 (
      {stage1_15[89]},
      {stage2_15[43]}
   );
   gpc1_1 gpc2078 (
      {stage1_15[90]},
      {stage2_15[44]}
   );
   gpc1_1 gpc2079 (
      {stage1_15[91]},
      {stage2_15[45]}
   );
   gpc1_1 gpc2080 (
      {stage1_15[92]},
      {stage2_15[46]}
   );
   gpc1_1 gpc2081 (
      {stage1_17[108]},
      {stage2_17[36]}
   );
   gpc1_1 gpc2082 (
      {stage1_17[109]},
      {stage2_17[37]}
   );
   gpc1_1 gpc2083 (
      {stage1_17[110]},
      {stage2_17[38]}
   );
   gpc1_1 gpc2084 (
      {stage1_17[111]},
      {stage2_17[39]}
   );
   gpc1_1 gpc2085 (
      {stage1_17[112]},
      {stage2_17[40]}
   );
   gpc1_1 gpc2086 (
      {stage1_17[113]},
      {stage2_17[41]}
   );
   gpc1_1 gpc2087 (
      {stage1_17[114]},
      {stage2_17[42]}
   );
   gpc1_1 gpc2088 (
      {stage1_17[115]},
      {stage2_17[43]}
   );
   gpc1_1 gpc2089 (
      {stage1_17[116]},
      {stage2_17[44]}
   );
   gpc1_1 gpc2090 (
      {stage1_17[117]},
      {stage2_17[45]}
   );
   gpc1_1 gpc2091 (
      {stage1_17[118]},
      {stage2_17[46]}
   );
   gpc1_1 gpc2092 (
      {stage1_17[119]},
      {stage2_17[47]}
   );
   gpc1_1 gpc2093 (
      {stage1_17[120]},
      {stage2_17[48]}
   );
   gpc1_1 gpc2094 (
      {stage1_17[121]},
      {stage2_17[49]}
   );
   gpc1_1 gpc2095 (
      {stage1_17[122]},
      {stage2_17[50]}
   );
   gpc1_1 gpc2096 (
      {stage1_17[123]},
      {stage2_17[51]}
   );
   gpc1_1 gpc2097 (
      {stage1_17[124]},
      {stage2_17[52]}
   );
   gpc1_1 gpc2098 (
      {stage1_17[125]},
      {stage2_17[53]}
   );
   gpc1_1 gpc2099 (
      {stage1_17[126]},
      {stage2_17[54]}
   );
   gpc1_1 gpc2100 (
      {stage1_18[94]},
      {stage2_18[34]}
   );
   gpc1_1 gpc2101 (
      {stage1_18[95]},
      {stage2_18[35]}
   );
   gpc1_1 gpc2102 (
      {stage1_18[96]},
      {stage2_18[36]}
   );
   gpc1_1 gpc2103 (
      {stage1_18[97]},
      {stage2_18[37]}
   );
   gpc1_1 gpc2104 (
      {stage1_18[98]},
      {stage2_18[38]}
   );
   gpc1_1 gpc2105 (
      {stage1_18[99]},
      {stage2_18[39]}
   );
   gpc1_1 gpc2106 (
      {stage1_18[100]},
      {stage2_18[40]}
   );
   gpc1_1 gpc2107 (
      {stage1_18[101]},
      {stage2_18[41]}
   );
   gpc1_1 gpc2108 (
      {stage1_18[102]},
      {stage2_18[42]}
   );
   gpc1_1 gpc2109 (
      {stage1_18[103]},
      {stage2_18[43]}
   );
   gpc1_1 gpc2110 (
      {stage1_18[104]},
      {stage2_18[44]}
   );
   gpc1_1 gpc2111 (
      {stage1_18[105]},
      {stage2_18[45]}
   );
   gpc1_1 gpc2112 (
      {stage1_18[106]},
      {stage2_18[46]}
   );
   gpc1_1 gpc2113 (
      {stage1_18[107]},
      {stage2_18[47]}
   );
   gpc1_1 gpc2114 (
      {stage1_18[108]},
      {stage2_18[48]}
   );
   gpc1_1 gpc2115 (
      {stage1_18[109]},
      {stage2_18[49]}
   );
   gpc1_1 gpc2116 (
      {stage1_18[110]},
      {stage2_18[50]}
   );
   gpc1_1 gpc2117 (
      {stage1_18[111]},
      {stage2_18[51]}
   );
   gpc1_1 gpc2118 (
      {stage1_18[112]},
      {stage2_18[52]}
   );
   gpc1_1 gpc2119 (
      {stage1_18[113]},
      {stage2_18[53]}
   );
   gpc1_1 gpc2120 (
      {stage1_18[114]},
      {stage2_18[54]}
   );
   gpc1_1 gpc2121 (
      {stage1_18[115]},
      {stage2_18[55]}
   );
   gpc1_1 gpc2122 (
      {stage1_18[116]},
      {stage2_18[56]}
   );
   gpc1_1 gpc2123 (
      {stage1_18[117]},
      {stage2_18[57]}
   );
   gpc1_1 gpc2124 (
      {stage1_18[118]},
      {stage2_18[58]}
   );
   gpc1_1 gpc2125 (
      {stage1_18[119]},
      {stage2_18[59]}
   );
   gpc1_1 gpc2126 (
      {stage1_18[120]},
      {stage2_18[60]}
   );
   gpc1_1 gpc2127 (
      {stage1_18[121]},
      {stage2_18[61]}
   );
   gpc1_1 gpc2128 (
      {stage1_18[122]},
      {stage2_18[62]}
   );
   gpc1_1 gpc2129 (
      {stage1_18[123]},
      {stage2_18[63]}
   );
   gpc1_1 gpc2130 (
      {stage1_18[124]},
      {stage2_18[64]}
   );
   gpc1_1 gpc2131 (
      {stage1_18[125]},
      {stage2_18[65]}
   );
   gpc1_1 gpc2132 (
      {stage1_18[126]},
      {stage2_18[66]}
   );
   gpc1_1 gpc2133 (
      {stage1_18[127]},
      {stage2_18[67]}
   );
   gpc1_1 gpc2134 (
      {stage1_18[128]},
      {stage2_18[68]}
   );
   gpc1_1 gpc2135 (
      {stage1_18[129]},
      {stage2_18[69]}
   );
   gpc1_1 gpc2136 (
      {stage1_18[130]},
      {stage2_18[70]}
   );
   gpc1_1 gpc2137 (
      {stage1_18[131]},
      {stage2_18[71]}
   );
   gpc1_1 gpc2138 (
      {stage1_18[132]},
      {stage2_18[72]}
   );
   gpc1_1 gpc2139 (
      {stage1_18[133]},
      {stage2_18[73]}
   );
   gpc1_1 gpc2140 (
      {stage1_18[134]},
      {stage2_18[74]}
   );
   gpc1_1 gpc2141 (
      {stage1_18[135]},
      {stage2_18[75]}
   );
   gpc1_1 gpc2142 (
      {stage1_18[136]},
      {stage2_18[76]}
   );
   gpc1_1 gpc2143 (
      {stage1_18[137]},
      {stage2_18[77]}
   );
   gpc1_1 gpc2144 (
      {stage1_18[138]},
      {stage2_18[78]}
   );
   gpc1_1 gpc2145 (
      {stage1_18[139]},
      {stage2_18[79]}
   );
   gpc1_1 gpc2146 (
      {stage1_18[140]},
      {stage2_18[80]}
   );
   gpc1_1 gpc2147 (
      {stage1_18[141]},
      {stage2_18[81]}
   );
   gpc1_1 gpc2148 (
      {stage1_18[142]},
      {stage2_18[82]}
   );
   gpc1_1 gpc2149 (
      {stage1_18[143]},
      {stage2_18[83]}
   );
   gpc1_1 gpc2150 (
      {stage1_18[144]},
      {stage2_18[84]}
   );
   gpc1_1 gpc2151 (
      {stage1_18[145]},
      {stage2_18[85]}
   );
   gpc1_1 gpc2152 (
      {stage1_18[146]},
      {stage2_18[86]}
   );
   gpc1_1 gpc2153 (
      {stage1_18[147]},
      {stage2_18[87]}
   );
   gpc1_1 gpc2154 (
      {stage1_18[148]},
      {stage2_18[88]}
   );
   gpc1_1 gpc2155 (
      {stage1_18[149]},
      {stage2_18[89]}
   );
   gpc1_1 gpc2156 (
      {stage1_18[150]},
      {stage2_18[90]}
   );
   gpc1_1 gpc2157 (
      {stage1_19[93]},
      {stage2_19[45]}
   );
   gpc1_1 gpc2158 (
      {stage1_20[23]},
      {stage2_20[33]}
   );
   gpc1_1 gpc2159 (
      {stage1_20[24]},
      {stage2_20[34]}
   );
   gpc1_1 gpc2160 (
      {stage1_20[25]},
      {stage2_20[35]}
   );
   gpc1_1 gpc2161 (
      {stage1_20[26]},
      {stage2_20[36]}
   );
   gpc1_1 gpc2162 (
      {stage1_20[27]},
      {stage2_20[37]}
   );
   gpc1_1 gpc2163 (
      {stage1_20[28]},
      {stage2_20[38]}
   );
   gpc1_1 gpc2164 (
      {stage1_20[29]},
      {stage2_20[39]}
   );
   gpc1_1 gpc2165 (
      {stage1_20[30]},
      {stage2_20[40]}
   );
   gpc1_1 gpc2166 (
      {stage1_20[31]},
      {stage2_20[41]}
   );
   gpc1_1 gpc2167 (
      {stage1_20[32]},
      {stage2_20[42]}
   );
   gpc1_1 gpc2168 (
      {stage1_20[33]},
      {stage2_20[43]}
   );
   gpc1_1 gpc2169 (
      {stage1_20[34]},
      {stage2_20[44]}
   );
   gpc1_1 gpc2170 (
      {stage1_20[35]},
      {stage2_20[45]}
   );
   gpc1_1 gpc2171 (
      {stage1_20[36]},
      {stage2_20[46]}
   );
   gpc1_1 gpc2172 (
      {stage1_20[37]},
      {stage2_20[47]}
   );
   gpc1_1 gpc2173 (
      {stage1_20[38]},
      {stage2_20[48]}
   );
   gpc1_1 gpc2174 (
      {stage1_20[39]},
      {stage2_20[49]}
   );
   gpc1_1 gpc2175 (
      {stage1_20[40]},
      {stage2_20[50]}
   );
   gpc1_1 gpc2176 (
      {stage1_20[41]},
      {stage2_20[51]}
   );
   gpc1_1 gpc2177 (
      {stage1_20[42]},
      {stage2_20[52]}
   );
   gpc1_1 gpc2178 (
      {stage1_20[43]},
      {stage2_20[53]}
   );
   gpc1_1 gpc2179 (
      {stage1_20[44]},
      {stage2_20[54]}
   );
   gpc1_1 gpc2180 (
      {stage1_20[45]},
      {stage2_20[55]}
   );
   gpc1_1 gpc2181 (
      {stage1_20[46]},
      {stage2_20[56]}
   );
   gpc1_1 gpc2182 (
      {stage1_20[47]},
      {stage2_20[57]}
   );
   gpc1_1 gpc2183 (
      {stage1_20[48]},
      {stage2_20[58]}
   );
   gpc1_1 gpc2184 (
      {stage1_20[49]},
      {stage2_20[59]}
   );
   gpc1_1 gpc2185 (
      {stage1_20[50]},
      {stage2_20[60]}
   );
   gpc1_1 gpc2186 (
      {stage1_20[51]},
      {stage2_20[61]}
   );
   gpc1_1 gpc2187 (
      {stage1_20[52]},
      {stage2_20[62]}
   );
   gpc1_1 gpc2188 (
      {stage1_20[53]},
      {stage2_20[63]}
   );
   gpc1_1 gpc2189 (
      {stage1_20[54]},
      {stage2_20[64]}
   );
   gpc1_1 gpc2190 (
      {stage1_20[55]},
      {stage2_20[65]}
   );
   gpc1_1 gpc2191 (
      {stage1_20[56]},
      {stage2_20[66]}
   );
   gpc1_1 gpc2192 (
      {stage1_20[57]},
      {stage2_20[67]}
   );
   gpc1_1 gpc2193 (
      {stage1_20[58]},
      {stage2_20[68]}
   );
   gpc1_1 gpc2194 (
      {stage1_20[59]},
      {stage2_20[69]}
   );
   gpc1_1 gpc2195 (
      {stage1_20[60]},
      {stage2_20[70]}
   );
   gpc1_1 gpc2196 (
      {stage1_20[61]},
      {stage2_20[71]}
   );
   gpc1_1 gpc2197 (
      {stage1_20[62]},
      {stage2_20[72]}
   );
   gpc1_1 gpc2198 (
      {stage1_20[63]},
      {stage2_20[73]}
   );
   gpc1_1 gpc2199 (
      {stage1_20[64]},
      {stage2_20[74]}
   );
   gpc1_1 gpc2200 (
      {stage1_20[65]},
      {stage2_20[75]}
   );
   gpc1_1 gpc2201 (
      {stage1_20[66]},
      {stage2_20[76]}
   );
   gpc1_1 gpc2202 (
      {stage1_20[67]},
      {stage2_20[77]}
   );
   gpc1_1 gpc2203 (
      {stage1_20[68]},
      {stage2_20[78]}
   );
   gpc1_1 gpc2204 (
      {stage1_20[69]},
      {stage2_20[79]}
   );
   gpc1_1 gpc2205 (
      {stage1_20[70]},
      {stage2_20[80]}
   );
   gpc1_1 gpc2206 (
      {stage1_20[71]},
      {stage2_20[81]}
   );
   gpc1_1 gpc2207 (
      {stage1_20[72]},
      {stage2_20[82]}
   );
   gpc1_1 gpc2208 (
      {stage1_20[73]},
      {stage2_20[83]}
   );
   gpc1_1 gpc2209 (
      {stage1_20[74]},
      {stage2_20[84]}
   );
   gpc1_1 gpc2210 (
      {stage1_20[75]},
      {stage2_20[85]}
   );
   gpc1_1 gpc2211 (
      {stage1_20[76]},
      {stage2_20[86]}
   );
   gpc1_1 gpc2212 (
      {stage1_20[77]},
      {stage2_20[87]}
   );
   gpc1_1 gpc2213 (
      {stage1_20[78]},
      {stage2_20[88]}
   );
   gpc1_1 gpc2214 (
      {stage1_20[79]},
      {stage2_20[89]}
   );
   gpc1_1 gpc2215 (
      {stage1_20[80]},
      {stage2_20[90]}
   );
   gpc1_1 gpc2216 (
      {stage1_20[81]},
      {stage2_20[91]}
   );
   gpc1_1 gpc2217 (
      {stage1_20[82]},
      {stage2_20[92]}
   );
   gpc1_1 gpc2218 (
      {stage1_20[83]},
      {stage2_20[93]}
   );
   gpc1_1 gpc2219 (
      {stage1_20[84]},
      {stage2_20[94]}
   );
   gpc1_1 gpc2220 (
      {stage1_20[85]},
      {stage2_20[95]}
   );
   gpc1_1 gpc2221 (
      {stage1_20[86]},
      {stage2_20[96]}
   );
   gpc1_1 gpc2222 (
      {stage1_20[87]},
      {stage2_20[97]}
   );
   gpc1_1 gpc2223 (
      {stage1_20[88]},
      {stage2_20[98]}
   );
   gpc1_1 gpc2224 (
      {stage1_20[89]},
      {stage2_20[99]}
   );
   gpc1_1 gpc2225 (
      {stage1_20[90]},
      {stage2_20[100]}
   );
   gpc1_1 gpc2226 (
      {stage1_20[91]},
      {stage2_20[101]}
   );
   gpc1_1 gpc2227 (
      {stage1_20[92]},
      {stage2_20[102]}
   );
   gpc1_1 gpc2228 (
      {stage1_20[93]},
      {stage2_20[103]}
   );
   gpc1_1 gpc2229 (
      {stage1_20[94]},
      {stage2_20[104]}
   );
   gpc1_1 gpc2230 (
      {stage1_20[95]},
      {stage2_20[105]}
   );
   gpc1_1 gpc2231 (
      {stage1_20[96]},
      {stage2_20[106]}
   );
   gpc1_1 gpc2232 (
      {stage1_20[97]},
      {stage2_20[107]}
   );
   gpc1_1 gpc2233 (
      {stage1_20[98]},
      {stage2_20[108]}
   );
   gpc1_1 gpc2234 (
      {stage1_20[99]},
      {stage2_20[109]}
   );
   gpc1_1 gpc2235 (
      {stage1_20[100]},
      {stage2_20[110]}
   );
   gpc1_1 gpc2236 (
      {stage1_20[101]},
      {stage2_20[111]}
   );
   gpc1_1 gpc2237 (
      {stage1_20[102]},
      {stage2_20[112]}
   );
   gpc1_1 gpc2238 (
      {stage1_20[103]},
      {stage2_20[113]}
   );
   gpc1_1 gpc2239 (
      {stage1_20[104]},
      {stage2_20[114]}
   );
   gpc1_1 gpc2240 (
      {stage1_20[105]},
      {stage2_20[115]}
   );
   gpc1_1 gpc2241 (
      {stage1_20[106]},
      {stage2_20[116]}
   );
   gpc1_1 gpc2242 (
      {stage1_20[107]},
      {stage2_20[117]}
   );
   gpc1_1 gpc2243 (
      {stage1_20[108]},
      {stage2_20[118]}
   );
   gpc1_1 gpc2244 (
      {stage1_20[109]},
      {stage2_20[119]}
   );
   gpc1_1 gpc2245 (
      {stage1_20[110]},
      {stage2_20[120]}
   );
   gpc1_1 gpc2246 (
      {stage1_20[111]},
      {stage2_20[121]}
   );
   gpc1_1 gpc2247 (
      {stage1_20[112]},
      {stage2_20[122]}
   );
   gpc1_1 gpc2248 (
      {stage1_20[113]},
      {stage2_20[123]}
   );
   gpc1_1 gpc2249 (
      {stage1_20[114]},
      {stage2_20[124]}
   );
   gpc1_1 gpc2250 (
      {stage1_20[115]},
      {stage2_20[125]}
   );
   gpc1_1 gpc2251 (
      {stage1_21[90]},
      {stage2_21[23]}
   );
   gpc1_1 gpc2252 (
      {stage1_21[91]},
      {stage2_21[24]}
   );
   gpc1_1 gpc2253 (
      {stage1_21[92]},
      {stage2_21[25]}
   );
   gpc1_1 gpc2254 (
      {stage1_21[93]},
      {stage2_21[26]}
   );
   gpc1_1 gpc2255 (
      {stage1_21[94]},
      {stage2_21[27]}
   );
   gpc1_1 gpc2256 (
      {stage1_21[95]},
      {stage2_21[28]}
   );
   gpc1_1 gpc2257 (
      {stage1_21[96]},
      {stage2_21[29]}
   );
   gpc1_1 gpc2258 (
      {stage1_21[97]},
      {stage2_21[30]}
   );
   gpc1_1 gpc2259 (
      {stage1_21[98]},
      {stage2_21[31]}
   );
   gpc1_1 gpc2260 (
      {stage1_21[99]},
      {stage2_21[32]}
   );
   gpc1_1 gpc2261 (
      {stage1_21[100]},
      {stage2_21[33]}
   );
   gpc1_1 gpc2262 (
      {stage1_21[101]},
      {stage2_21[34]}
   );
   gpc1_1 gpc2263 (
      {stage1_21[102]},
      {stage2_21[35]}
   );
   gpc1_1 gpc2264 (
      {stage1_21[103]},
      {stage2_21[36]}
   );
   gpc1_1 gpc2265 (
      {stage1_21[104]},
      {stage2_21[37]}
   );
   gpc1_1 gpc2266 (
      {stage1_21[105]},
      {stage2_21[38]}
   );
   gpc1_1 gpc2267 (
      {stage1_21[106]},
      {stage2_21[39]}
   );
   gpc1_1 gpc2268 (
      {stage1_21[107]},
      {stage2_21[40]}
   );
   gpc1_1 gpc2269 (
      {stage1_21[108]},
      {stage2_21[41]}
   );
   gpc1_1 gpc2270 (
      {stage1_21[109]},
      {stage2_21[42]}
   );
   gpc1_1 gpc2271 (
      {stage1_21[110]},
      {stage2_21[43]}
   );
   gpc1_1 gpc2272 (
      {stage1_21[111]},
      {stage2_21[44]}
   );
   gpc1_1 gpc2273 (
      {stage1_21[112]},
      {stage2_21[45]}
   );
   gpc1_1 gpc2274 (
      {stage1_21[113]},
      {stage2_21[46]}
   );
   gpc1_1 gpc2275 (
      {stage1_21[114]},
      {stage2_21[47]}
   );
   gpc1_1 gpc2276 (
      {stage1_21[115]},
      {stage2_21[48]}
   );
   gpc1_1 gpc2277 (
      {stage1_21[116]},
      {stage2_21[49]}
   );
   gpc1_1 gpc2278 (
      {stage1_21[117]},
      {stage2_21[50]}
   );
   gpc1_1 gpc2279 (
      {stage1_21[118]},
      {stage2_21[51]}
   );
   gpc1_1 gpc2280 (
      {stage1_21[119]},
      {stage2_21[52]}
   );
   gpc1_1 gpc2281 (
      {stage1_21[120]},
      {stage2_21[53]}
   );
   gpc1_1 gpc2282 (
      {stage1_21[121]},
      {stage2_21[54]}
   );
   gpc1_1 gpc2283 (
      {stage1_21[122]},
      {stage2_21[55]}
   );
   gpc1_1 gpc2284 (
      {stage1_21[123]},
      {stage2_21[56]}
   );
   gpc1_1 gpc2285 (
      {stage1_21[124]},
      {stage2_21[57]}
   );
   gpc1_1 gpc2286 (
      {stage1_21[125]},
      {stage2_21[58]}
   );
   gpc1_1 gpc2287 (
      {stage1_21[126]},
      {stage2_21[59]}
   );
   gpc1_1 gpc2288 (
      {stage1_21[127]},
      {stage2_21[60]}
   );
   gpc1_1 gpc2289 (
      {stage1_21[128]},
      {stage2_21[61]}
   );
   gpc1_1 gpc2290 (
      {stage1_21[129]},
      {stage2_21[62]}
   );
   gpc1_1 gpc2291 (
      {stage1_21[130]},
      {stage2_21[63]}
   );
   gpc1_1 gpc2292 (
      {stage1_21[131]},
      {stage2_21[64]}
   );
   gpc1_1 gpc2293 (
      {stage1_21[132]},
      {stage2_21[65]}
   );
   gpc1_1 gpc2294 (
      {stage1_21[133]},
      {stage2_21[66]}
   );
   gpc1_1 gpc2295 (
      {stage1_21[134]},
      {stage2_21[67]}
   );
   gpc1_1 gpc2296 (
      {stage1_21[135]},
      {stage2_21[68]}
   );
   gpc1_1 gpc2297 (
      {stage1_21[136]},
      {stage2_21[69]}
   );
   gpc1_1 gpc2298 (
      {stage1_21[137]},
      {stage2_21[70]}
   );
   gpc1_1 gpc2299 (
      {stage1_21[138]},
      {stage2_21[71]}
   );
   gpc1_1 gpc2300 (
      {stage1_22[77]},
      {stage2_22[30]}
   );
   gpc1_1 gpc2301 (
      {stage1_22[78]},
      {stage2_22[31]}
   );
   gpc1_1 gpc2302 (
      {stage1_22[79]},
      {stage2_22[32]}
   );
   gpc1_1 gpc2303 (
      {stage1_22[80]},
      {stage2_22[33]}
   );
   gpc1_1 gpc2304 (
      {stage1_22[81]},
      {stage2_22[34]}
   );
   gpc1_1 gpc2305 (
      {stage1_22[82]},
      {stage2_22[35]}
   );
   gpc1_1 gpc2306 (
      {stage1_22[83]},
      {stage2_22[36]}
   );
   gpc1_1 gpc2307 (
      {stage1_22[84]},
      {stage2_22[37]}
   );
   gpc1_1 gpc2308 (
      {stage1_22[85]},
      {stage2_22[38]}
   );
   gpc1_1 gpc2309 (
      {stage1_22[86]},
      {stage2_22[39]}
   );
   gpc1_1 gpc2310 (
      {stage1_22[87]},
      {stage2_22[40]}
   );
   gpc1_1 gpc2311 (
      {stage1_22[88]},
      {stage2_22[41]}
   );
   gpc1_1 gpc2312 (
      {stage1_22[89]},
      {stage2_22[42]}
   );
   gpc1_1 gpc2313 (
      {stage1_22[90]},
      {stage2_22[43]}
   );
   gpc1_1 gpc2314 (
      {stage1_22[91]},
      {stage2_22[44]}
   );
   gpc1_1 gpc2315 (
      {stage1_22[92]},
      {stage2_22[45]}
   );
   gpc1_1 gpc2316 (
      {stage1_22[93]},
      {stage2_22[46]}
   );
   gpc1_1 gpc2317 (
      {stage1_23[73]},
      {stage2_23[36]}
   );
   gpc1_1 gpc2318 (
      {stage1_23[74]},
      {stage2_23[37]}
   );
   gpc1_1 gpc2319 (
      {stage1_23[75]},
      {stage2_23[38]}
   );
   gpc1_1 gpc2320 (
      {stage1_23[76]},
      {stage2_23[39]}
   );
   gpc1_1 gpc2321 (
      {stage1_23[77]},
      {stage2_23[40]}
   );
   gpc1_1 gpc2322 (
      {stage1_23[78]},
      {stage2_23[41]}
   );
   gpc1_1 gpc2323 (
      {stage1_23[79]},
      {stage2_23[42]}
   );
   gpc1_1 gpc2324 (
      {stage1_23[80]},
      {stage2_23[43]}
   );
   gpc1_1 gpc2325 (
      {stage1_23[81]},
      {stage2_23[44]}
   );
   gpc1_1 gpc2326 (
      {stage1_23[82]},
      {stage2_23[45]}
   );
   gpc1_1 gpc2327 (
      {stage1_23[83]},
      {stage2_23[46]}
   );
   gpc1_1 gpc2328 (
      {stage1_23[84]},
      {stage2_23[47]}
   );
   gpc1_1 gpc2329 (
      {stage1_23[85]},
      {stage2_23[48]}
   );
   gpc1_1 gpc2330 (
      {stage1_23[86]},
      {stage2_23[49]}
   );
   gpc1_1 gpc2331 (
      {stage1_23[87]},
      {stage2_23[50]}
   );
   gpc1_1 gpc2332 (
      {stage1_23[88]},
      {stage2_23[51]}
   );
   gpc1_1 gpc2333 (
      {stage1_23[89]},
      {stage2_23[52]}
   );
   gpc1_1 gpc2334 (
      {stage1_23[90]},
      {stage2_23[53]}
   );
   gpc1_1 gpc2335 (
      {stage1_23[91]},
      {stage2_23[54]}
   );
   gpc1_1 gpc2336 (
      {stage1_23[92]},
      {stage2_23[55]}
   );
   gpc1_1 gpc2337 (
      {stage1_23[93]},
      {stage2_23[56]}
   );
   gpc1_1 gpc2338 (
      {stage1_24[249]},
      {stage2_24[59]}
   );
   gpc1_1 gpc2339 (
      {stage1_24[250]},
      {stage2_24[60]}
   );
   gpc1_1 gpc2340 (
      {stage1_24[251]},
      {stage2_24[61]}
   );
   gpc1_1 gpc2341 (
      {stage1_24[252]},
      {stage2_24[62]}
   );
   gpc1_1 gpc2342 (
      {stage1_24[253]},
      {stage2_24[63]}
   );
   gpc1_1 gpc2343 (
      {stage1_25[117]},
      {stage2_25[65]}
   );
   gpc1_1 gpc2344 (
      {stage1_27[73]},
      {stage2_27[61]}
   );
   gpc1_1 gpc2345 (
      {stage1_27[74]},
      {stage2_27[62]}
   );
   gpc1_1 gpc2346 (
      {stage1_27[75]},
      {stage2_27[63]}
   );
   gpc1_1 gpc2347 (
      {stage1_27[76]},
      {stage2_27[64]}
   );
   gpc1_1 gpc2348 (
      {stage1_27[77]},
      {stage2_27[65]}
   );
   gpc1_1 gpc2349 (
      {stage1_27[78]},
      {stage2_27[66]}
   );
   gpc1_1 gpc2350 (
      {stage1_27[79]},
      {stage2_27[67]}
   );
   gpc1_1 gpc2351 (
      {stage1_27[80]},
      {stage2_27[68]}
   );
   gpc1_1 gpc2352 (
      {stage1_27[81]},
      {stage2_27[69]}
   );
   gpc1_1 gpc2353 (
      {stage1_27[82]},
      {stage2_27[70]}
   );
   gpc1_1 gpc2354 (
      {stage1_27[83]},
      {stage2_27[71]}
   );
   gpc1_1 gpc2355 (
      {stage1_27[84]},
      {stage2_27[72]}
   );
   gpc1_1 gpc2356 (
      {stage1_27[85]},
      {stage2_27[73]}
   );
   gpc1_1 gpc2357 (
      {stage1_27[86]},
      {stage2_27[74]}
   );
   gpc1_1 gpc2358 (
      {stage1_27[87]},
      {stage2_27[75]}
   );
   gpc1_1 gpc2359 (
      {stage1_27[88]},
      {stage2_27[76]}
   );
   gpc1_1 gpc2360 (
      {stage1_27[89]},
      {stage2_27[77]}
   );
   gpc1_1 gpc2361 (
      {stage1_27[90]},
      {stage2_27[78]}
   );
   gpc1_1 gpc2362 (
      {stage1_27[91]},
      {stage2_27[79]}
   );
   gpc1_1 gpc2363 (
      {stage1_27[92]},
      {stage2_27[80]}
   );
   gpc1_1 gpc2364 (
      {stage1_27[93]},
      {stage2_27[81]}
   );
   gpc1_1 gpc2365 (
      {stage1_27[94]},
      {stage2_27[82]}
   );
   gpc1_1 gpc2366 (
      {stage1_27[95]},
      {stage2_27[83]}
   );
   gpc1_1 gpc2367 (
      {stage1_27[96]},
      {stage2_27[84]}
   );
   gpc1_1 gpc2368 (
      {stage1_27[97]},
      {stage2_27[85]}
   );
   gpc1_1 gpc2369 (
      {stage1_27[98]},
      {stage2_27[86]}
   );
   gpc1_1 gpc2370 (
      {stage1_27[99]},
      {stage2_27[87]}
   );
   gpc1_1 gpc2371 (
      {stage1_27[100]},
      {stage2_27[88]}
   );
   gpc1_1 gpc2372 (
      {stage1_27[101]},
      {stage2_27[89]}
   );
   gpc1_1 gpc2373 (
      {stage1_27[102]},
      {stage2_27[90]}
   );
   gpc1_1 gpc2374 (
      {stage1_27[103]},
      {stage2_27[91]}
   );
   gpc1_1 gpc2375 (
      {stage1_27[104]},
      {stage2_27[92]}
   );
   gpc1_1 gpc2376 (
      {stage1_27[105]},
      {stage2_27[93]}
   );
   gpc1_1 gpc2377 (
      {stage1_27[106]},
      {stage2_27[94]}
   );
   gpc1_1 gpc2378 (
      {stage1_27[107]},
      {stage2_27[95]}
   );
   gpc1_1 gpc2379 (
      {stage1_28[90]},
      {stage2_28[60]}
   );
   gpc1_1 gpc2380 (
      {stage1_28[91]},
      {stage2_28[61]}
   );
   gpc1_1 gpc2381 (
      {stage1_28[92]},
      {stage2_28[62]}
   );
   gpc1_1 gpc2382 (
      {stage1_28[93]},
      {stage2_28[63]}
   );
   gpc1_1 gpc2383 (
      {stage1_28[94]},
      {stage2_28[64]}
   );
   gpc1_1 gpc2384 (
      {stage1_28[95]},
      {stage2_28[65]}
   );
   gpc1_1 gpc2385 (
      {stage1_28[96]},
      {stage2_28[66]}
   );
   gpc1_1 gpc2386 (
      {stage1_28[97]},
      {stage2_28[67]}
   );
   gpc1_1 gpc2387 (
      {stage1_28[98]},
      {stage2_28[68]}
   );
   gpc1_1 gpc2388 (
      {stage1_28[99]},
      {stage2_28[69]}
   );
   gpc1_1 gpc2389 (
      {stage1_28[100]},
      {stage2_28[70]}
   );
   gpc1_1 gpc2390 (
      {stage1_28[101]},
      {stage2_28[71]}
   );
   gpc1_1 gpc2391 (
      {stage1_31[129]},
      {stage2_31[44]}
   );
   gpc1_1 gpc2392 (
      {stage1_31[130]},
      {stage2_31[45]}
   );
   gpc1_1 gpc2393 (
      {stage1_31[131]},
      {stage2_31[46]}
   );
   gpc1_1 gpc2394 (
      {stage1_31[132]},
      {stage2_31[47]}
   );
   gpc1_1 gpc2395 (
      {stage1_32[68]},
      {stage2_32[38]}
   );
   gpc1_1 gpc2396 (
      {stage1_32[69]},
      {stage2_32[39]}
   );
   gpc1_1 gpc2397 (
      {stage1_32[70]},
      {stage2_32[40]}
   );
   gpc1_1 gpc2398 (
      {stage1_32[71]},
      {stage2_32[41]}
   );
   gpc1_1 gpc2399 (
      {stage1_32[72]},
      {stage2_32[42]}
   );
   gpc1_1 gpc2400 (
      {stage1_32[73]},
      {stage2_32[43]}
   );
   gpc117_4 gpc2401 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6]},
      {stage2_1[0]},
      {stage2_2[0]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc117_4 gpc2402 (
      {stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13]},
      {stage2_1[1]},
      {stage2_2[1]},
      {stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1163_5 gpc2403 (
      {stage2_0[14], stage2_0[15], stage2_0[16]},
      {stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7]},
      {stage2_2[2]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc2404 (
      {stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20], stage2_0[21]},
      {stage2_1[8]},
      {stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8]},
      {stage3_4[1],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc2405 (
      {stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc2406 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[6]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[1],stage3_4[3],stage3_3[5]}
   );
   gpc615_5 gpc2407 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[7]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[2],stage3_4[4],stage3_3[6]}
   );
   gpc615_5 gpc2408 (
      {stage2_3[11], stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15]},
      {stage2_4[8]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[3],stage3_4[5],stage3_3[7]}
   );
   gpc606_5 gpc2409 (
      {stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[4],stage3_5[4],stage3_4[6]}
   );
   gpc606_5 gpc2410 (
      {stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[5],stage3_5[5],stage3_4[7]}
   );
   gpc606_5 gpc2411 (
      {stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25], stage2_4[26]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[6],stage3_5[6],stage3_4[8]}
   );
   gpc615_5 gpc2412 (
      {stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31]},
      {stage2_5[18]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[6],stage3_6[7],stage3_5[7],stage3_4[9]}
   );
   gpc615_5 gpc2413 (
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36]},
      {stage2_5[19]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[7],stage3_6[8],stage3_5[8],stage3_4[10]}
   );
   gpc615_5 gpc2414 (
      {stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage2_5[20]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[8],stage3_6[9],stage3_5[9],stage3_4[11]}
   );
   gpc615_5 gpc2415 (
      {stage2_4[42], stage2_4[43], stage2_4[44], stage2_4[45], stage2_4[46]},
      {stage2_5[21]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[9],stage3_6[10],stage3_5[10],stage3_4[12]}
   );
   gpc615_5 gpc2416 (
      {stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51]},
      {stage2_5[22]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[10],stage3_6[11],stage3_5[11],stage3_4[13]}
   );
   gpc606_5 gpc2417 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[8],stage3_7[11],stage3_6[12],stage3_5[12]}
   );
   gpc606_5 gpc2418 (
      {stage2_5[29], stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[9],stage3_7[12],stage3_6[13],stage3_5[13]}
   );
   gpc606_5 gpc2419 (
      {stage2_5[35], stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[10],stage3_7[13],stage3_6[14],stage3_5[14]}
   );
   gpc615_5 gpc2420 (
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[3],stage3_8[11],stage3_7[14]}
   );
   gpc615_5 gpc2421 (
      {stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[4],stage3_8[12],stage3_7[15]}
   );
   gpc615_5 gpc2422 (
      {stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32]},
      {stage2_8[2]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[2],stage3_9[5],stage3_8[13],stage3_7[16]}
   );
   gpc615_5 gpc2423 (
      {stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37]},
      {stage2_8[3]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[3],stage3_9[6],stage3_8[14],stage3_7[17]}
   );
   gpc615_5 gpc2424 (
      {stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41], stage2_7[42]},
      {stage2_8[4]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[4],stage3_9[7],stage3_8[15],stage3_7[18]}
   );
   gpc615_5 gpc2425 (
      {stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46], stage2_7[47]},
      {stage2_8[5]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[5],stage3_9[8],stage3_8[16],stage3_7[19]}
   );
   gpc623_5 gpc2426 (
      {stage2_7[48], stage2_7[49], stage2_7[50]},
      {stage2_8[6], stage2_8[7]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[6],stage3_9[9],stage3_8[17],stage3_7[20]}
   );
   gpc606_5 gpc2427 (
      {stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[7],stage3_10[7],stage3_9[10],stage3_8[18]}
   );
   gpc606_5 gpc2428 (
      {stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[8],stage3_10[8],stage3_9[11],stage3_8[19]}
   );
   gpc606_5 gpc2429 (
      {stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[9],stage3_10[9],stage3_9[12],stage3_8[20]}
   );
   gpc606_5 gpc2430 (
      {stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30], stage2_8[31]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[10],stage3_10[10],stage3_9[13],stage3_8[21]}
   );
   gpc606_5 gpc2431 (
      {stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36], stage2_8[37]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[11],stage3_10[11],stage3_9[14],stage3_8[22]}
   );
   gpc606_5 gpc2432 (
      {stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42], stage2_8[43]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[12],stage3_10[12],stage3_9[15],stage3_8[23]}
   );
   gpc606_5 gpc2433 (
      {stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47], stage2_8[48], stage2_8[49]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[13],stage3_10[13],stage3_9[16],stage3_8[24]}
   );
   gpc615_5 gpc2434 (
      {stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54]},
      {stage2_9[42]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[7],stage3_11[14],stage3_10[14],stage3_9[17],stage3_8[25]}
   );
   gpc606_5 gpc2435 (
      {stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47], stage2_9[48]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[8],stage3_11[15],stage3_10[15],stage3_9[18]}
   );
   gpc606_5 gpc2436 (
      {stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53], stage2_9[54]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[9],stage3_11[16],stage3_10[16],stage3_9[19]}
   );
   gpc606_5 gpc2437 (
      {stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59], stage2_9[60]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[10],stage3_11[17],stage3_10[17],stage3_9[20]}
   );
   gpc615_5 gpc2438 (
      {stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage2_10[48]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[11],stage3_11[18],stage3_10[18],stage3_9[21]}
   );
   gpc615_5 gpc2439 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28]},
      {stage2_12[0]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[4],stage3_12[12],stage3_11[19]}
   );
   gpc615_5 gpc2440 (
      {stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33]},
      {stage2_12[1]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[5],stage3_12[13],stage3_11[20]}
   );
   gpc615_5 gpc2441 (
      {stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_12[2]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[6],stage3_12[14],stage3_11[21]}
   );
   gpc615_5 gpc2442 (
      {stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43]},
      {stage2_12[3]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[3],stage3_13[7],stage3_12[15],stage3_11[22]}
   );
   gpc615_5 gpc2443 (
      {stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48]},
      {stage2_12[4]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[4],stage3_13[8],stage3_12[16],stage3_11[23]}
   );
   gpc615_5 gpc2444 (
      {stage2_11[49], stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53]},
      {stage2_12[5]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[5],stage3_13[9],stage3_12[17],stage3_11[24]}
   );
   gpc615_5 gpc2445 (
      {stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57], 1'b0},
      {stage2_12[6]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[6],stage3_13[10],stage3_12[18],stage3_11[25]}
   );
   gpc606_5 gpc2446 (
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[7],stage3_14[7],stage3_13[11],stage3_12[19]}
   );
   gpc606_5 gpc2447 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[8],stage3_14[8],stage3_13[12],stage3_12[20]}
   );
   gpc606_5 gpc2448 (
      {stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[9],stage3_14[9],stage3_13[13],stage3_12[21]}
   );
   gpc606_5 gpc2449 (
      {stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[10],stage3_14[10],stage3_13[14],stage3_12[22]}
   );
   gpc606_5 gpc2450 (
      {stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[11],stage3_14[11],stage3_13[15],stage3_12[23]}
   );
   gpc606_5 gpc2451 (
      {stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[12],stage3_14[12],stage3_13[16],stage3_12[24]}
   );
   gpc606_5 gpc2452 (
      {stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47], stage2_12[48]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[13],stage3_14[13],stage3_13[17],stage3_12[25]}
   );
   gpc606_5 gpc2453 (
      {stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53], stage2_12[54]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[14],stage3_14[14],stage3_13[18],stage3_12[26]}
   );
   gpc606_5 gpc2454 (
      {stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59], stage2_12[60]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[15],stage3_14[15],stage3_13[19],stage3_12[27]}
   );
   gpc606_5 gpc2455 (
      {stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65], stage2_12[66]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[16],stage3_14[16],stage3_13[20],stage3_12[28]}
   );
   gpc606_5 gpc2456 (
      {stage2_12[67], stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[17],stage3_14[17],stage3_13[21],stage3_12[29]}
   );
   gpc615_5 gpc2457 (
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[11],stage3_15[18],stage3_14[18]}
   );
   gpc615_5 gpc2458 (
      {stage2_14[71], stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[12],stage3_15[19],stage3_14[19]}
   );
   gpc615_5 gpc2459 (
      {stage2_14[76], stage2_14[77], stage2_14[78], stage2_14[79], stage2_14[80]},
      {stage2_15[2]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[13],stage3_15[20],stage3_14[20]}
   );
   gpc615_5 gpc2460 (
      {stage2_14[81], stage2_14[82], stage2_14[83], stage2_14[84], stage2_14[85]},
      {stage2_15[3]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[3],stage3_16[14],stage3_15[21],stage3_14[21]}
   );
   gpc615_5 gpc2461 (
      {stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8]},
      {stage2_16[24]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[4],stage3_17[4],stage3_16[15],stage3_15[22]}
   );
   gpc615_5 gpc2462 (
      {stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13]},
      {stage2_16[25]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[5],stage3_17[5],stage3_16[16],stage3_15[23]}
   );
   gpc615_5 gpc2463 (
      {stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18]},
      {stage2_16[26]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[6],stage3_17[6],stage3_16[17],stage3_15[24]}
   );
   gpc615_5 gpc2464 (
      {stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage2_16[27]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[7],stage3_17[7],stage3_16[18],stage3_15[25]}
   );
   gpc615_5 gpc2465 (
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28]},
      {stage2_16[28]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[8],stage3_17[8],stage3_16[19],stage3_15[26]}
   );
   gpc615_5 gpc2466 (
      {stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33]},
      {stage2_16[29]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[9],stage3_17[9],stage3_16[20],stage3_15[27]}
   );
   gpc615_5 gpc2467 (
      {stage2_15[34], stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38]},
      {stage2_16[30]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[10],stage3_17[10],stage3_16[21],stage3_15[28]}
   );
   gpc615_5 gpc2468 (
      {stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43]},
      {stage2_16[31]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[11],stage3_17[11],stage3_16[22],stage3_15[29]}
   );
   gpc606_5 gpc2469 (
      {stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35], stage2_16[36], stage2_16[37]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[8],stage3_18[12],stage3_17[12],stage3_16[23]}
   );
   gpc615_5 gpc2470 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[0]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[9],stage3_18[13]}
   );
   gpc615_5 gpc2471 (
      {stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15]},
      {stage2_19[1]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[1],stage3_20[2],stage3_19[10],stage3_18[14]}
   );
   gpc615_5 gpc2472 (
      {stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19], stage2_18[20]},
      {stage2_19[2]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[2],stage3_20[3],stage3_19[11],stage3_18[15]}
   );
   gpc615_5 gpc2473 (
      {stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24], stage2_18[25]},
      {stage2_19[3]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[3],stage3_20[4],stage3_19[12],stage3_18[16]}
   );
   gpc615_5 gpc2474 (
      {stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_19[4]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[4],stage3_20[5],stage3_19[13],stage3_18[17]}
   );
   gpc615_5 gpc2475 (
      {stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35]},
      {stage2_19[5]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[5],stage3_20[6],stage3_19[14],stage3_18[18]}
   );
   gpc615_5 gpc2476 (
      {stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40]},
      {stage2_19[6]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[6],stage3_20[7],stage3_19[15],stage3_18[19]}
   );
   gpc615_5 gpc2477 (
      {stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44], stage2_18[45]},
      {stage2_19[7]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[7],stage3_20[8],stage3_19[16],stage3_18[20]}
   );
   gpc615_5 gpc2478 (
      {stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49], stage2_18[50]},
      {stage2_19[8]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[8],stage3_21[8],stage3_20[9],stage3_19[17],stage3_18[21]}
   );
   gpc615_5 gpc2479 (
      {stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54], stage2_18[55]},
      {stage2_19[9]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[9],stage3_21[9],stage3_20[10],stage3_19[18],stage3_18[22]}
   );
   gpc615_5 gpc2480 (
      {stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60]},
      {stage2_19[10]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[10],stage3_21[10],stage3_20[11],stage3_19[19],stage3_18[23]}
   );
   gpc615_5 gpc2481 (
      {stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65]},
      {stage2_19[11]},
      {stage2_20[66], stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage3_22[11],stage3_21[11],stage3_20[12],stage3_19[20],stage3_18[24]}
   );
   gpc615_5 gpc2482 (
      {stage2_18[66], stage2_18[67], stage2_18[68], stage2_18[69], stage2_18[70]},
      {stage2_19[12]},
      {stage2_20[72], stage2_20[73], stage2_20[74], stage2_20[75], stage2_20[76], stage2_20[77]},
      {stage3_22[12],stage3_21[12],stage3_20[13],stage3_19[21],stage3_18[25]}
   );
   gpc615_5 gpc2483 (
      {stage2_18[71], stage2_18[72], stage2_18[73], stage2_18[74], stage2_18[75]},
      {stage2_19[13]},
      {stage2_20[78], stage2_20[79], stage2_20[80], stage2_20[81], stage2_20[82], stage2_20[83]},
      {stage3_22[13],stage3_21[13],stage3_20[14],stage3_19[22],stage3_18[26]}
   );
   gpc615_5 gpc2484 (
      {stage2_18[76], stage2_18[77], stage2_18[78], stage2_18[79], stage2_18[80]},
      {stage2_19[14]},
      {stage2_20[84], stage2_20[85], stage2_20[86], stage2_20[87], stage2_20[88], stage2_20[89]},
      {stage3_22[14],stage3_21[14],stage3_20[15],stage3_19[23],stage3_18[27]}
   );
   gpc615_5 gpc2485 (
      {stage2_19[15], stage2_19[16], stage2_19[17], stage2_19[18], stage2_19[19]},
      {stage2_20[90]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[15],stage3_21[15],stage3_20[16],stage3_19[24]}
   );
   gpc615_5 gpc2486 (
      {stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23], stage2_19[24]},
      {stage2_20[91]},
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage3_23[1],stage3_22[16],stage3_21[16],stage3_20[17],stage3_19[25]}
   );
   gpc615_5 gpc2487 (
      {stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_20[92]},
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage3_23[2],stage3_22[17],stage3_21[17],stage3_20[18],stage3_19[26]}
   );
   gpc615_5 gpc2488 (
      {stage2_19[30], stage2_19[31], stage2_19[32], stage2_19[33], stage2_19[34]},
      {stage2_20[93]},
      {stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23]},
      {stage3_23[3],stage3_22[18],stage3_21[18],stage3_20[19],stage3_19[27]}
   );
   gpc615_5 gpc2489 (
      {stage2_19[35], stage2_19[36], stage2_19[37], stage2_19[38], stage2_19[39]},
      {stage2_20[94]},
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage3_23[4],stage3_22[19],stage3_21[19],stage3_20[20],stage3_19[28]}
   );
   gpc606_5 gpc2490 (
      {stage2_20[95], stage2_20[96], stage2_20[97], stage2_20[98], stage2_20[99], stage2_20[100]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[5],stage3_22[20],stage3_21[20],stage3_20[21]}
   );
   gpc606_5 gpc2491 (
      {stage2_20[101], stage2_20[102], stage2_20[103], stage2_20[104], stage2_20[105], stage2_20[106]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[6],stage3_22[21],stage3_21[21],stage3_20[22]}
   );
   gpc606_5 gpc2492 (
      {stage2_20[107], stage2_20[108], stage2_20[109], stage2_20[110], stage2_20[111], stage2_20[112]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[7],stage3_22[22],stage3_21[22],stage3_20[23]}
   );
   gpc1343_5 gpc2493 (
      {stage2_21[30], stage2_21[31], stage2_21[32]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21]},
      {stage2_23[0], stage2_23[1], stage2_23[2]},
      {stage2_24[0]},
      {stage3_25[0],stage3_24[3],stage3_23[8],stage3_22[23],stage3_21[23]}
   );
   gpc1343_5 gpc2494 (
      {stage2_21[33], stage2_21[34], stage2_21[35]},
      {stage2_22[22], stage2_22[23], stage2_22[24], stage2_22[25]},
      {stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage2_24[1]},
      {stage3_25[1],stage3_24[4],stage3_23[9],stage3_22[24],stage3_21[24]}
   );
   gpc1343_5 gpc2495 (
      {stage2_21[36], stage2_21[37], stage2_21[38]},
      {stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage2_23[6], stage2_23[7], stage2_23[8]},
      {stage2_24[2]},
      {stage3_25[2],stage3_24[5],stage3_23[10],stage3_22[25],stage3_21[25]}
   );
   gpc615_5 gpc2496 (
      {stage2_21[39], stage2_21[40], stage2_21[41], stage2_21[42], stage2_21[43]},
      {stage2_22[30]},
      {stage2_23[9], stage2_23[10], stage2_23[11], stage2_23[12], stage2_23[13], stage2_23[14]},
      {stage3_25[3],stage3_24[6],stage3_23[11],stage3_22[26],stage3_21[26]}
   );
   gpc615_5 gpc2497 (
      {stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47], stage2_21[48]},
      {stage2_22[31]},
      {stage2_23[15], stage2_23[16], stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20]},
      {stage3_25[4],stage3_24[7],stage3_23[12],stage3_22[27],stage3_21[27]}
   );
   gpc615_5 gpc2498 (
      {stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage2_22[32]},
      {stage2_23[21], stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26]},
      {stage3_25[5],stage3_24[8],stage3_23[13],stage3_22[28],stage3_21[28]}
   );
   gpc615_5 gpc2499 (
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58]},
      {stage2_22[33]},
      {stage2_23[27], stage2_23[28], stage2_23[29], stage2_23[30], stage2_23[31], stage2_23[32]},
      {stage3_25[6],stage3_24[9],stage3_23[14],stage3_22[29],stage3_21[29]}
   );
   gpc615_5 gpc2500 (
      {stage2_21[59], stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63]},
      {stage2_22[34]},
      {stage2_23[33], stage2_23[34], stage2_23[35], stage2_23[36], stage2_23[37], stage2_23[38]},
      {stage3_25[7],stage3_24[10],stage3_23[15],stage3_22[30],stage3_21[30]}
   );
   gpc615_5 gpc2501 (
      {stage2_21[64], stage2_21[65], stage2_21[66], stage2_21[67], stage2_21[68]},
      {stage2_22[35]},
      {stage2_23[39], stage2_23[40], stage2_23[41], stage2_23[42], stage2_23[43], stage2_23[44]},
      {stage3_25[8],stage3_24[11],stage3_23[16],stage3_22[31],stage3_21[31]}
   );
   gpc615_5 gpc2502 (
      {stage2_21[69], stage2_21[70], stage2_21[71], 1'b0, 1'b0},
      {stage2_22[36]},
      {stage2_23[45], stage2_23[46], stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50]},
      {stage3_25[9],stage3_24[12],stage3_23[17],stage3_22[32],stage3_21[32]}
   );
   gpc615_5 gpc2503 (
      {stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage2_23[51]},
      {stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6], stage2_24[7], stage2_24[8]},
      {stage3_26[0],stage3_25[10],stage3_24[13],stage3_23[18],stage3_22[33]}
   );
   gpc615_5 gpc2504 (
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46]},
      {stage2_23[52]},
      {stage2_24[9], stage2_24[10], stage2_24[11], stage2_24[12], stage2_24[13], stage2_24[14]},
      {stage3_26[1],stage3_25[11],stage3_24[14],stage3_23[19],stage3_22[34]}
   );
   gpc615_5 gpc2505 (
      {stage2_23[53], stage2_23[54], stage2_23[55], stage2_23[56], 1'b0},
      {stage2_24[15]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[2],stage3_25[12],stage3_24[15],stage3_23[20]}
   );
   gpc606_5 gpc2506 (
      {stage2_24[16], stage2_24[17], stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[1],stage3_26[3],stage3_25[13],stage3_24[16]}
   );
   gpc606_5 gpc2507 (
      {stage2_24[22], stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[2],stage3_26[4],stage3_25[14],stage3_24[17]}
   );
   gpc606_5 gpc2508 (
      {stage2_24[28], stage2_24[29], stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[3],stage3_26[5],stage3_25[15],stage3_24[18]}
   );
   gpc606_5 gpc2509 (
      {stage2_24[34], stage2_24[35], stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[4],stage3_26[6],stage3_25[16],stage3_24[19]}
   );
   gpc606_5 gpc2510 (
      {stage2_24[40], stage2_24[41], stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45]},
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage3_28[4],stage3_27[5],stage3_26[7],stage3_25[17],stage3_24[20]}
   );
   gpc606_5 gpc2511 (
      {stage2_24[46], stage2_24[47], stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51]},
      {stage2_26[30], stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35]},
      {stage3_28[5],stage3_27[6],stage3_26[8],stage3_25[18],stage3_24[21]}
   );
   gpc606_5 gpc2512 (
      {stage2_24[52], stage2_24[53], stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57]},
      {stage2_26[36], stage2_26[37], stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41]},
      {stage3_28[6],stage3_27[7],stage3_26[9],stage3_25[19],stage3_24[22]}
   );
   gpc606_5 gpc2513 (
      {stage2_24[58], stage2_24[59], stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63]},
      {stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47]},
      {stage3_28[7],stage3_27[8],stage3_26[10],stage3_25[20],stage3_24[23]}
   );
   gpc606_5 gpc2514 (
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[8],stage3_27[9],stage3_26[11],stage3_25[21]}
   );
   gpc606_5 gpc2515 (
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[9],stage3_27[10],stage3_26[12],stage3_25[22]}
   );
   gpc606_5 gpc2516 (
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[10],stage3_27[11],stage3_26[13],stage3_25[23]}
   );
   gpc606_5 gpc2517 (
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[11],stage3_27[12],stage3_26[14],stage3_25[24]}
   );
   gpc606_5 gpc2518 (
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[12],stage3_27[13],stage3_26[15],stage3_25[25]}
   );
   gpc606_5 gpc2519 (
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage2_27[30], stage2_27[31], stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35]},
      {stage3_29[5],stage3_28[13],stage3_27[14],stage3_26[16],stage3_25[26]}
   );
   gpc606_5 gpc2520 (
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage2_27[36], stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage3_29[6],stage3_28[14],stage3_27[15],stage3_26[17],stage3_25[27]}
   );
   gpc606_5 gpc2521 (
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46], stage2_27[47]},
      {stage3_29[7],stage3_28[15],stage3_27[16],stage3_26[18],stage3_25[28]}
   );
   gpc606_5 gpc2522 (
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage2_27[48], stage2_27[49], stage2_27[50], stage2_27[51], stage2_27[52], stage2_27[53]},
      {stage3_29[8],stage3_28[16],stage3_27[17],stage3_26[19],stage3_25[29]}
   );
   gpc615_5 gpc2523 (
      {stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52]},
      {stage2_27[54]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[9],stage3_28[17],stage3_27[18],stage3_26[20]}
   );
   gpc615_5 gpc2524 (
      {stage2_26[53], stage2_26[54], stage2_26[55], stage2_26[56], stage2_26[57]},
      {stage2_27[55]},
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage3_30[1],stage3_29[10],stage3_28[18],stage3_27[19],stage3_26[21]}
   );
   gpc615_5 gpc2525 (
      {stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_27[56]},
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage3_30[2],stage3_29[11],stage3_28[19],stage3_27[20],stage3_26[22]}
   );
   gpc615_5 gpc2526 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67]},
      {stage2_27[57]},
      {stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage3_30[3],stage3_29[12],stage3_28[20],stage3_27[21],stage3_26[23]}
   );
   gpc606_5 gpc2527 (
      {stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61], stage2_27[62], stage2_27[63]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[4],stage3_29[13],stage3_28[21],stage3_27[22]}
   );
   gpc615_5 gpc2528 (
      {stage2_27[64], stage2_27[65], stage2_27[66], stage2_27[67], stage2_27[68]},
      {stage2_28[24]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[5],stage3_29[14],stage3_28[22],stage3_27[23]}
   );
   gpc615_5 gpc2529 (
      {stage2_27[69], stage2_27[70], stage2_27[71], stage2_27[72], stage2_27[73]},
      {stage2_28[25]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[6],stage3_29[15],stage3_28[23],stage3_27[24]}
   );
   gpc615_5 gpc2530 (
      {stage2_27[74], stage2_27[75], stage2_27[76], stage2_27[77], stage2_27[78]},
      {stage2_28[26]},
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage3_31[3],stage3_30[7],stage3_29[16],stage3_28[24],stage3_27[25]}
   );
   gpc615_5 gpc2531 (
      {stage2_27[79], stage2_27[80], stage2_27[81], stage2_27[82], stage2_27[83]},
      {stage2_28[27]},
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage3_31[4],stage3_30[8],stage3_29[17],stage3_28[25],stage3_27[26]}
   );
   gpc606_5 gpc2532 (
      {stage2_28[28], stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[5],stage3_30[9],stage3_29[18],stage3_28[26]}
   );
   gpc606_5 gpc2533 (
      {stage2_28[34], stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38], stage2_28[39]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[6],stage3_30[10],stage3_29[19],stage3_28[27]}
   );
   gpc606_5 gpc2534 (
      {stage2_28[40], stage2_28[41], stage2_28[42], stage2_28[43], stage2_28[44], stage2_28[45]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[7],stage3_30[11],stage3_29[20],stage3_28[28]}
   );
   gpc606_5 gpc2535 (
      {stage2_28[46], stage2_28[47], stage2_28[48], stage2_28[49], stage2_28[50], stage2_28[51]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[8],stage3_30[12],stage3_29[21],stage3_28[29]}
   );
   gpc606_5 gpc2536 (
      {stage2_28[52], stage2_28[53], stage2_28[54], stage2_28[55], stage2_28[56], stage2_28[57]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[9],stage3_30[13],stage3_29[22],stage3_28[30]}
   );
   gpc606_5 gpc2537 (
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[5],stage3_31[10],stage3_30[14],stage3_29[23]}
   );
   gpc615_5 gpc2538 (
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34]},
      {stage2_31[6]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[1],stage3_32[6],stage3_31[11],stage3_30[15]}
   );
   gpc615_5 gpc2539 (
      {stage2_30[35], stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39]},
      {stage2_31[7]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[2],stage3_32[7],stage3_31[12],stage3_30[16]}
   );
   gpc615_5 gpc2540 (
      {stage2_30[40], stage2_30[41], stage2_30[42], stage2_30[43], stage2_30[44]},
      {stage2_31[8]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[3],stage3_32[8],stage3_31[13],stage3_30[17]}
   );
   gpc615_5 gpc2541 (
      {stage2_31[9], stage2_31[10], stage2_31[11], stage2_31[12], stage2_31[13]},
      {stage2_32[18]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[3],stage3_33[4],stage3_32[9],stage3_31[14]}
   );
   gpc615_5 gpc2542 (
      {stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17], stage2_31[18]},
      {stage2_32[19]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[4],stage3_33[5],stage3_32[10],stage3_31[15]}
   );
   gpc615_5 gpc2543 (
      {stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage2_32[20]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[5],stage3_33[6],stage3_32[11],stage3_31[16]}
   );
   gpc615_5 gpc2544 (
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28]},
      {stage2_32[21]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[6],stage3_33[7],stage3_32[12],stage3_31[17]}
   );
   gpc606_5 gpc2545 (
      {stage2_32[22], stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[4],stage3_34[7],stage3_33[8],stage3_32[13]}
   );
   gpc606_5 gpc2546 (
      {stage2_32[28], stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[5],stage3_34[8],stage3_33[9],stage3_32[14]}
   );
   gpc606_5 gpc2547 (
      {stage2_32[34], stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], 1'b0},
      {stage3_36[2],stage3_35[6],stage3_34[9],stage3_33[10],stage3_32[15]}
   );
   gpc1_1 gpc2548 (
      {stage2_0[22]},
      {stage3_0[4]}
   );
   gpc1_1 gpc2549 (
      {stage2_0[23]},
      {stage3_0[5]}
   );
   gpc1_1 gpc2550 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc2551 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc2552 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc2553 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc2554 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc2555 (
      {stage2_1[14]},
      {stage3_1[9]}
   );
   gpc1_1 gpc2556 (
      {stage2_1[15]},
      {stage3_1[10]}
   );
   gpc1_1 gpc2557 (
      {stage2_1[16]},
      {stage3_1[11]}
   );
   gpc1_1 gpc2558 (
      {stage2_1[17]},
      {stage3_1[12]}
   );
   gpc1_1 gpc2559 (
      {stage2_1[18]},
      {stage3_1[13]}
   );
   gpc1_1 gpc2560 (
      {stage2_1[19]},
      {stage3_1[14]}
   );
   gpc1_1 gpc2561 (
      {stage2_1[20]},
      {stage3_1[15]}
   );
   gpc1_1 gpc2562 (
      {stage2_1[21]},
      {stage3_1[16]}
   );
   gpc1_1 gpc2563 (
      {stage2_1[22]},
      {stage3_1[17]}
   );
   gpc1_1 gpc2564 (
      {stage2_1[23]},
      {stage3_1[18]}
   );
   gpc1_1 gpc2565 (
      {stage2_1[24]},
      {stage3_1[19]}
   );
   gpc1_1 gpc2566 (
      {stage2_1[25]},
      {stage3_1[20]}
   );
   gpc1_1 gpc2567 (
      {stage2_1[26]},
      {stage3_1[21]}
   );
   gpc1_1 gpc2568 (
      {stage2_1[27]},
      {stage3_1[22]}
   );
   gpc1_1 gpc2569 (
      {stage2_1[28]},
      {stage3_1[23]}
   );
   gpc1_1 gpc2570 (
      {stage2_1[29]},
      {stage3_1[24]}
   );
   gpc1_1 gpc2571 (
      {stage2_1[30]},
      {stage3_1[25]}
   );
   gpc1_1 gpc2572 (
      {stage2_1[31]},
      {stage3_1[26]}
   );
   gpc1_1 gpc2573 (
      {stage2_1[32]},
      {stage3_1[27]}
   );
   gpc1_1 gpc2574 (
      {stage2_2[15]},
      {stage3_2[5]}
   );
   gpc1_1 gpc2575 (
      {stage2_2[16]},
      {stage3_2[6]}
   );
   gpc1_1 gpc2576 (
      {stage2_2[17]},
      {stage3_2[7]}
   );
   gpc1_1 gpc2577 (
      {stage2_2[18]},
      {stage3_2[8]}
   );
   gpc1_1 gpc2578 (
      {stage2_2[19]},
      {stage3_2[9]}
   );
   gpc1_1 gpc2579 (
      {stage2_2[20]},
      {stage3_2[10]}
   );
   gpc1_1 gpc2580 (
      {stage2_2[21]},
      {stage3_2[11]}
   );
   gpc1_1 gpc2581 (
      {stage2_2[22]},
      {stage3_2[12]}
   );
   gpc1_1 gpc2582 (
      {stage2_2[23]},
      {stage3_2[13]}
   );
   gpc1_1 gpc2583 (
      {stage2_2[24]},
      {stage3_2[14]}
   );
   gpc1_1 gpc2584 (
      {stage2_2[25]},
      {stage3_2[15]}
   );
   gpc1_1 gpc2585 (
      {stage2_2[26]},
      {stage3_2[16]}
   );
   gpc1_1 gpc2586 (
      {stage2_2[27]},
      {stage3_2[17]}
   );
   gpc1_1 gpc2587 (
      {stage2_2[28]},
      {stage3_2[18]}
   );
   gpc1_1 gpc2588 (
      {stage2_2[29]},
      {stage3_2[19]}
   );
   gpc1_1 gpc2589 (
      {stage2_2[30]},
      {stage3_2[20]}
   );
   gpc1_1 gpc2590 (
      {stage2_2[31]},
      {stage3_2[21]}
   );
   gpc1_1 gpc2591 (
      {stage2_2[32]},
      {stage3_2[22]}
   );
   gpc1_1 gpc2592 (
      {stage2_2[33]},
      {stage3_2[23]}
   );
   gpc1_1 gpc2593 (
      {stage2_2[34]},
      {stage3_2[24]}
   );
   gpc1_1 gpc2594 (
      {stage2_3[16]},
      {stage3_3[8]}
   );
   gpc1_1 gpc2595 (
      {stage2_3[17]},
      {stage3_3[9]}
   );
   gpc1_1 gpc2596 (
      {stage2_3[18]},
      {stage3_3[10]}
   );
   gpc1_1 gpc2597 (
      {stage2_3[19]},
      {stage3_3[11]}
   );
   gpc1_1 gpc2598 (
      {stage2_3[20]},
      {stage3_3[12]}
   );
   gpc1_1 gpc2599 (
      {stage2_3[21]},
      {stage3_3[13]}
   );
   gpc1_1 gpc2600 (
      {stage2_3[22]},
      {stage3_3[14]}
   );
   gpc1_1 gpc2601 (
      {stage2_3[23]},
      {stage3_3[15]}
   );
   gpc1_1 gpc2602 (
      {stage2_3[24]},
      {stage3_3[16]}
   );
   gpc1_1 gpc2603 (
      {stage2_3[25]},
      {stage3_3[17]}
   );
   gpc1_1 gpc2604 (
      {stage2_3[26]},
      {stage3_3[18]}
   );
   gpc1_1 gpc2605 (
      {stage2_3[27]},
      {stage3_3[19]}
   );
   gpc1_1 gpc2606 (
      {stage2_3[28]},
      {stage3_3[20]}
   );
   gpc1_1 gpc2607 (
      {stage2_3[29]},
      {stage3_3[21]}
   );
   gpc1_1 gpc2608 (
      {stage2_3[30]},
      {stage3_3[22]}
   );
   gpc1_1 gpc2609 (
      {stage2_3[31]},
      {stage3_3[23]}
   );
   gpc1_1 gpc2610 (
      {stage2_3[32]},
      {stage3_3[24]}
   );
   gpc1_1 gpc2611 (
      {stage2_3[33]},
      {stage3_3[25]}
   );
   gpc1_1 gpc2612 (
      {stage2_3[34]},
      {stage3_3[26]}
   );
   gpc1_1 gpc2613 (
      {stage2_3[35]},
      {stage3_3[27]}
   );
   gpc1_1 gpc2614 (
      {stage2_3[36]},
      {stage3_3[28]}
   );
   gpc1_1 gpc2615 (
      {stage2_3[37]},
      {stage3_3[29]}
   );
   gpc1_1 gpc2616 (
      {stage2_3[38]},
      {stage3_3[30]}
   );
   gpc1_1 gpc2617 (
      {stage2_3[39]},
      {stage3_3[31]}
   );
   gpc1_1 gpc2618 (
      {stage2_3[40]},
      {stage3_3[32]}
   );
   gpc1_1 gpc2619 (
      {stage2_3[41]},
      {stage3_3[33]}
   );
   gpc1_1 gpc2620 (
      {stage2_3[42]},
      {stage3_3[34]}
   );
   gpc1_1 gpc2621 (
      {stage2_4[52]},
      {stage3_4[14]}
   );
   gpc1_1 gpc2622 (
      {stage2_4[53]},
      {stage3_4[15]}
   );
   gpc1_1 gpc2623 (
      {stage2_4[54]},
      {stage3_4[16]}
   );
   gpc1_1 gpc2624 (
      {stage2_4[55]},
      {stage3_4[17]}
   );
   gpc1_1 gpc2625 (
      {stage2_4[56]},
      {stage3_4[18]}
   );
   gpc1_1 gpc2626 (
      {stage2_4[57]},
      {stage3_4[19]}
   );
   gpc1_1 gpc2627 (
      {stage2_4[58]},
      {stage3_4[20]}
   );
   gpc1_1 gpc2628 (
      {stage2_4[59]},
      {stage3_4[21]}
   );
   gpc1_1 gpc2629 (
      {stage2_4[60]},
      {stage3_4[22]}
   );
   gpc1_1 gpc2630 (
      {stage2_4[61]},
      {stage3_4[23]}
   );
   gpc1_1 gpc2631 (
      {stage2_4[62]},
      {stage3_4[24]}
   );
   gpc1_1 gpc2632 (
      {stage2_4[63]},
      {stage3_4[25]}
   );
   gpc1_1 gpc2633 (
      {stage2_4[64]},
      {stage3_4[26]}
   );
   gpc1_1 gpc2634 (
      {stage2_4[65]},
      {stage3_4[27]}
   );
   gpc1_1 gpc2635 (
      {stage2_4[66]},
      {stage3_4[28]}
   );
   gpc1_1 gpc2636 (
      {stage2_4[67]},
      {stage3_4[29]}
   );
   gpc1_1 gpc2637 (
      {stage2_4[68]},
      {stage3_4[30]}
   );
   gpc1_1 gpc2638 (
      {stage2_4[69]},
      {stage3_4[31]}
   );
   gpc1_1 gpc2639 (
      {stage2_4[70]},
      {stage3_4[32]}
   );
   gpc1_1 gpc2640 (
      {stage2_4[71]},
      {stage3_4[33]}
   );
   gpc1_1 gpc2641 (
      {stage2_4[72]},
      {stage3_4[34]}
   );
   gpc1_1 gpc2642 (
      {stage2_4[73]},
      {stage3_4[35]}
   );
   gpc1_1 gpc2643 (
      {stage2_5[41]},
      {stage3_5[15]}
   );
   gpc1_1 gpc2644 (
      {stage2_6[48]},
      {stage3_6[15]}
   );
   gpc1_1 gpc2645 (
      {stage2_6[49]},
      {stage3_6[16]}
   );
   gpc1_1 gpc2646 (
      {stage2_6[50]},
      {stage3_6[17]}
   );
   gpc1_1 gpc2647 (
      {stage2_6[51]},
      {stage3_6[18]}
   );
   gpc1_1 gpc2648 (
      {stage2_6[52]},
      {stage3_6[19]}
   );
   gpc1_1 gpc2649 (
      {stage2_7[51]},
      {stage3_7[21]}
   );
   gpc1_1 gpc2650 (
      {stage2_7[52]},
      {stage3_7[22]}
   );
   gpc1_1 gpc2651 (
      {stage2_7[53]},
      {stage3_7[23]}
   );
   gpc1_1 gpc2652 (
      {stage2_8[55]},
      {stage3_8[26]}
   );
   gpc1_1 gpc2653 (
      {stage2_12[73]},
      {stage3_12[30]}
   );
   gpc1_1 gpc2654 (
      {stage2_12[74]},
      {stage3_12[31]}
   );
   gpc1_1 gpc2655 (
      {stage2_13[42]},
      {stage3_13[22]}
   );
   gpc1_1 gpc2656 (
      {stage2_13[43]},
      {stage3_13[23]}
   );
   gpc1_1 gpc2657 (
      {stage2_13[44]},
      {stage3_13[24]}
   );
   gpc1_1 gpc2658 (
      {stage2_13[45]},
      {stage3_13[25]}
   );
   gpc1_1 gpc2659 (
      {stage2_13[46]},
      {stage3_13[26]}
   );
   gpc1_1 gpc2660 (
      {stage2_13[47]},
      {stage3_13[27]}
   );
   gpc1_1 gpc2661 (
      {stage2_13[48]},
      {stage3_13[28]}
   );
   gpc1_1 gpc2662 (
      {stage2_13[49]},
      {stage3_13[29]}
   );
   gpc1_1 gpc2663 (
      {stage2_13[50]},
      {stage3_13[30]}
   );
   gpc1_1 gpc2664 (
      {stage2_13[51]},
      {stage3_13[31]}
   );
   gpc1_1 gpc2665 (
      {stage2_13[52]},
      {stage3_13[32]}
   );
   gpc1_1 gpc2666 (
      {stage2_13[53]},
      {stage3_13[33]}
   );
   gpc1_1 gpc2667 (
      {stage2_13[54]},
      {stage3_13[34]}
   );
   gpc1_1 gpc2668 (
      {stage2_13[55]},
      {stage3_13[35]}
   );
   gpc1_1 gpc2669 (
      {stage2_13[56]},
      {stage3_13[36]}
   );
   gpc1_1 gpc2670 (
      {stage2_14[86]},
      {stage3_14[22]}
   );
   gpc1_1 gpc2671 (
      {stage2_14[87]},
      {stage3_14[23]}
   );
   gpc1_1 gpc2672 (
      {stage2_14[88]},
      {stage3_14[24]}
   );
   gpc1_1 gpc2673 (
      {stage2_14[89]},
      {stage3_14[25]}
   );
   gpc1_1 gpc2674 (
      {stage2_15[44]},
      {stage3_15[30]}
   );
   gpc1_1 gpc2675 (
      {stage2_15[45]},
      {stage3_15[31]}
   );
   gpc1_1 gpc2676 (
      {stage2_15[46]},
      {stage3_15[32]}
   );
   gpc1_1 gpc2677 (
      {stage2_16[38]},
      {stage3_16[24]}
   );
   gpc1_1 gpc2678 (
      {stage2_16[39]},
      {stage3_16[25]}
   );
   gpc1_1 gpc2679 (
      {stage2_16[40]},
      {stage3_16[26]}
   );
   gpc1_1 gpc2680 (
      {stage2_17[48]},
      {stage3_17[13]}
   );
   gpc1_1 gpc2681 (
      {stage2_17[49]},
      {stage3_17[14]}
   );
   gpc1_1 gpc2682 (
      {stage2_17[50]},
      {stage3_17[15]}
   );
   gpc1_1 gpc2683 (
      {stage2_17[51]},
      {stage3_17[16]}
   );
   gpc1_1 gpc2684 (
      {stage2_17[52]},
      {stage3_17[17]}
   );
   gpc1_1 gpc2685 (
      {stage2_17[53]},
      {stage3_17[18]}
   );
   gpc1_1 gpc2686 (
      {stage2_17[54]},
      {stage3_17[19]}
   );
   gpc1_1 gpc2687 (
      {stage2_18[81]},
      {stage3_18[28]}
   );
   gpc1_1 gpc2688 (
      {stage2_18[82]},
      {stage3_18[29]}
   );
   gpc1_1 gpc2689 (
      {stage2_18[83]},
      {stage3_18[30]}
   );
   gpc1_1 gpc2690 (
      {stage2_18[84]},
      {stage3_18[31]}
   );
   gpc1_1 gpc2691 (
      {stage2_18[85]},
      {stage3_18[32]}
   );
   gpc1_1 gpc2692 (
      {stage2_18[86]},
      {stage3_18[33]}
   );
   gpc1_1 gpc2693 (
      {stage2_18[87]},
      {stage3_18[34]}
   );
   gpc1_1 gpc2694 (
      {stage2_18[88]},
      {stage3_18[35]}
   );
   gpc1_1 gpc2695 (
      {stage2_18[89]},
      {stage3_18[36]}
   );
   gpc1_1 gpc2696 (
      {stage2_18[90]},
      {stage3_18[37]}
   );
   gpc1_1 gpc2697 (
      {stage2_19[40]},
      {stage3_19[29]}
   );
   gpc1_1 gpc2698 (
      {stage2_19[41]},
      {stage3_19[30]}
   );
   gpc1_1 gpc2699 (
      {stage2_19[42]},
      {stage3_19[31]}
   );
   gpc1_1 gpc2700 (
      {stage2_19[43]},
      {stage3_19[32]}
   );
   gpc1_1 gpc2701 (
      {stage2_19[44]},
      {stage3_19[33]}
   );
   gpc1_1 gpc2702 (
      {stage2_19[45]},
      {stage3_19[34]}
   );
   gpc1_1 gpc2703 (
      {stage2_20[113]},
      {stage3_20[24]}
   );
   gpc1_1 gpc2704 (
      {stage2_20[114]},
      {stage3_20[25]}
   );
   gpc1_1 gpc2705 (
      {stage2_20[115]},
      {stage3_20[26]}
   );
   gpc1_1 gpc2706 (
      {stage2_20[116]},
      {stage3_20[27]}
   );
   gpc1_1 gpc2707 (
      {stage2_20[117]},
      {stage3_20[28]}
   );
   gpc1_1 gpc2708 (
      {stage2_20[118]},
      {stage3_20[29]}
   );
   gpc1_1 gpc2709 (
      {stage2_20[119]},
      {stage3_20[30]}
   );
   gpc1_1 gpc2710 (
      {stage2_20[120]},
      {stage3_20[31]}
   );
   gpc1_1 gpc2711 (
      {stage2_20[121]},
      {stage3_20[32]}
   );
   gpc1_1 gpc2712 (
      {stage2_20[122]},
      {stage3_20[33]}
   );
   gpc1_1 gpc2713 (
      {stage2_20[123]},
      {stage3_20[34]}
   );
   gpc1_1 gpc2714 (
      {stage2_20[124]},
      {stage3_20[35]}
   );
   gpc1_1 gpc2715 (
      {stage2_20[125]},
      {stage3_20[36]}
   );
   gpc1_1 gpc2716 (
      {stage2_25[60]},
      {stage3_25[30]}
   );
   gpc1_1 gpc2717 (
      {stage2_25[61]},
      {stage3_25[31]}
   );
   gpc1_1 gpc2718 (
      {stage2_25[62]},
      {stage3_25[32]}
   );
   gpc1_1 gpc2719 (
      {stage2_25[63]},
      {stage3_25[33]}
   );
   gpc1_1 gpc2720 (
      {stage2_25[64]},
      {stage3_25[34]}
   );
   gpc1_1 gpc2721 (
      {stage2_25[65]},
      {stage3_25[35]}
   );
   gpc1_1 gpc2722 (
      {stage2_27[84]},
      {stage3_27[27]}
   );
   gpc1_1 gpc2723 (
      {stage2_27[85]},
      {stage3_27[28]}
   );
   gpc1_1 gpc2724 (
      {stage2_27[86]},
      {stage3_27[29]}
   );
   gpc1_1 gpc2725 (
      {stage2_27[87]},
      {stage3_27[30]}
   );
   gpc1_1 gpc2726 (
      {stage2_27[88]},
      {stage3_27[31]}
   );
   gpc1_1 gpc2727 (
      {stage2_27[89]},
      {stage3_27[32]}
   );
   gpc1_1 gpc2728 (
      {stage2_27[90]},
      {stage3_27[33]}
   );
   gpc1_1 gpc2729 (
      {stage2_27[91]},
      {stage3_27[34]}
   );
   gpc1_1 gpc2730 (
      {stage2_27[92]},
      {stage3_27[35]}
   );
   gpc1_1 gpc2731 (
      {stage2_27[93]},
      {stage3_27[36]}
   );
   gpc1_1 gpc2732 (
      {stage2_27[94]},
      {stage3_27[37]}
   );
   gpc1_1 gpc2733 (
      {stage2_27[95]},
      {stage3_27[38]}
   );
   gpc1_1 gpc2734 (
      {stage2_28[58]},
      {stage3_28[31]}
   );
   gpc1_1 gpc2735 (
      {stage2_28[59]},
      {stage3_28[32]}
   );
   gpc1_1 gpc2736 (
      {stage2_28[60]},
      {stage3_28[33]}
   );
   gpc1_1 gpc2737 (
      {stage2_28[61]},
      {stage3_28[34]}
   );
   gpc1_1 gpc2738 (
      {stage2_28[62]},
      {stage3_28[35]}
   );
   gpc1_1 gpc2739 (
      {stage2_28[63]},
      {stage3_28[36]}
   );
   gpc1_1 gpc2740 (
      {stage2_28[64]},
      {stage3_28[37]}
   );
   gpc1_1 gpc2741 (
      {stage2_28[65]},
      {stage3_28[38]}
   );
   gpc1_1 gpc2742 (
      {stage2_28[66]},
      {stage3_28[39]}
   );
   gpc1_1 gpc2743 (
      {stage2_28[67]},
      {stage3_28[40]}
   );
   gpc1_1 gpc2744 (
      {stage2_28[68]},
      {stage3_28[41]}
   );
   gpc1_1 gpc2745 (
      {stage2_28[69]},
      {stage3_28[42]}
   );
   gpc1_1 gpc2746 (
      {stage2_28[70]},
      {stage3_28[43]}
   );
   gpc1_1 gpc2747 (
      {stage2_28[71]},
      {stage3_28[44]}
   );
   gpc1_1 gpc2748 (
      {stage2_29[36]},
      {stage3_29[24]}
   );
   gpc1_1 gpc2749 (
      {stage2_29[37]},
      {stage3_29[25]}
   );
   gpc1_1 gpc2750 (
      {stage2_29[38]},
      {stage3_29[26]}
   );
   gpc1_1 gpc2751 (
      {stage2_29[39]},
      {stage3_29[27]}
   );
   gpc1_1 gpc2752 (
      {stage2_31[29]},
      {stage3_31[18]}
   );
   gpc1_1 gpc2753 (
      {stage2_31[30]},
      {stage3_31[19]}
   );
   gpc1_1 gpc2754 (
      {stage2_31[31]},
      {stage3_31[20]}
   );
   gpc1_1 gpc2755 (
      {stage2_31[32]},
      {stage3_31[21]}
   );
   gpc1_1 gpc2756 (
      {stage2_31[33]},
      {stage3_31[22]}
   );
   gpc1_1 gpc2757 (
      {stage2_31[34]},
      {stage3_31[23]}
   );
   gpc1_1 gpc2758 (
      {stage2_31[35]},
      {stage3_31[24]}
   );
   gpc1_1 gpc2759 (
      {stage2_31[36]},
      {stage3_31[25]}
   );
   gpc1_1 gpc2760 (
      {stage2_31[37]},
      {stage3_31[26]}
   );
   gpc1_1 gpc2761 (
      {stage2_31[38]},
      {stage3_31[27]}
   );
   gpc1_1 gpc2762 (
      {stage2_31[39]},
      {stage3_31[28]}
   );
   gpc1_1 gpc2763 (
      {stage2_31[40]},
      {stage3_31[29]}
   );
   gpc1_1 gpc2764 (
      {stage2_31[41]},
      {stage3_31[30]}
   );
   gpc1_1 gpc2765 (
      {stage2_31[42]},
      {stage3_31[31]}
   );
   gpc1_1 gpc2766 (
      {stage2_31[43]},
      {stage3_31[32]}
   );
   gpc1_1 gpc2767 (
      {stage2_31[44]},
      {stage3_31[33]}
   );
   gpc1_1 gpc2768 (
      {stage2_31[45]},
      {stage3_31[34]}
   );
   gpc1_1 gpc2769 (
      {stage2_31[46]},
      {stage3_31[35]}
   );
   gpc1_1 gpc2770 (
      {stage2_31[47]},
      {stage3_31[36]}
   );
   gpc1_1 gpc2771 (
      {stage2_32[40]},
      {stage3_32[16]}
   );
   gpc1_1 gpc2772 (
      {stage2_32[41]},
      {stage3_32[17]}
   );
   gpc1_1 gpc2773 (
      {stage2_32[42]},
      {stage3_32[18]}
   );
   gpc1_1 gpc2774 (
      {stage2_32[43]},
      {stage3_32[19]}
   );
   gpc1_1 gpc2775 (
      {stage2_33[24]},
      {stage3_33[11]}
   );
   gpc1_1 gpc2776 (
      {stage2_33[25]},
      {stage3_33[12]}
   );
   gpc1_1 gpc2777 (
      {stage2_33[26]},
      {stage3_33[13]}
   );
   gpc1_1 gpc2778 (
      {stage2_33[27]},
      {stage3_33[14]}
   );
   gpc1_1 gpc2779 (
      {stage2_33[28]},
      {stage3_33[15]}
   );
   gpc1_1 gpc2780 (
      {stage2_33[29]},
      {stage3_33[16]}
   );
   gpc1_1 gpc2781 (
      {stage2_33[30]},
      {stage3_33[17]}
   );
   gpc1_1 gpc2782 (
      {stage2_35[0]},
      {stage3_35[7]}
   );
   gpc1_1 gpc2783 (
      {stage2_35[1]},
      {stage3_35[8]}
   );
   gpc1_1 gpc2784 (
      {stage2_35[2]},
      {stage3_35[9]}
   );
   gpc1_1 gpc2785 (
      {stage2_35[3]},
      {stage3_35[10]}
   );
   gpc1_1 gpc2786 (
      {stage2_35[4]},
      {stage3_35[11]}
   );
   gpc1_1 gpc2787 (
      {stage2_35[5]},
      {stage3_35[12]}
   );
   gpc606_5 gpc2788 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc2789 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc2790 (
      {stage3_1[12], stage3_1[13], stage3_1[14], stage3_1[15], stage3_1[16], stage3_1[17]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc2791 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc606_5 gpc2792 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[4],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc606_5 gpc2793 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[5],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc606_5 gpc2794 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[6],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc207_4 gpc2795 (
      {stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23], stage3_3[24]},
      {stage3_5[0], stage3_5[1]},
      {stage4_6[4],stage4_5[7],stage4_4[7],stage4_3[7]}
   );
   gpc207_4 gpc2796 (
      {stage3_3[25], stage3_3[26], stage3_3[27], stage3_3[28], stage3_3[29], stage3_3[30], stage3_3[31]},
      {stage3_5[2], stage3_5[3]},
      {stage4_6[5],stage4_5[8],stage4_4[8],stage4_3[8]}
   );
   gpc606_5 gpc2797 (
      {stage3_4[24], stage3_4[25], stage3_4[26], stage3_4[27], stage3_4[28], stage3_4[29]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[6],stage4_5[9],stage4_4[9]}
   );
   gpc606_5 gpc2798 (
      {stage3_5[4], stage3_5[5], stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[7],stage4_5[10]}
   );
   gpc606_5 gpc2799 (
      {stage3_5[10], stage3_5[11], stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[2],stage4_6[8],stage4_5[11]}
   );
   gpc615_5 gpc2800 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[12]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[2],stage4_8[3],stage4_7[3],stage4_6[9]}
   );
   gpc615_5 gpc2801 (
      {stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage3_7[13]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[3],stage4_8[4],stage4_7[4],stage4_6[10]}
   );
   gpc135_4 gpc2802 (
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[2],stage4_9[4],stage4_8[5]}
   );
   gpc135_4 gpc2803 (
      {stage3_8[17], stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21]},
      {stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_10[1]},
      {stage4_11[1],stage4_10[3],stage4_9[5],stage4_8[6]}
   );
   gpc135_4 gpc2804 (
      {stage3_8[22], stage3_8[23], stage3_8[24], stage3_8[25], stage3_8[26]},
      {stage3_9[6], stage3_9[7], stage3_9[8]},
      {stage3_10[2]},
      {stage4_11[2],stage4_10[4],stage4_9[6],stage4_8[7]}
   );
   gpc606_5 gpc2805 (
      {stage3_9[9], stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[3],stage4_10[5],stage4_9[7]}
   );
   gpc606_5 gpc2806 (
      {stage3_9[15], stage3_9[16], stage3_9[17], stage3_9[18], stage3_9[19], stage3_9[20]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[4],stage4_10[6],stage4_9[8]}
   );
   gpc615_5 gpc2807 (
      {stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage3_11[12]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[2],stage4_11[5],stage4_10[7]}
   );
   gpc615_5 gpc2808 (
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12]},
      {stage3_11[13]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[3],stage4_12[3],stage4_11[6],stage4_10[8]}
   );
   gpc615_5 gpc2809 (
      {stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17], stage3_11[18]},
      {stage3_12[12]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[2],stage4_13[4],stage4_12[4],stage4_11[7]}
   );
   gpc615_5 gpc2810 (
      {stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage3_12[13]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[3],stage4_13[5],stage4_12[5],stage4_11[8]}
   );
   gpc615_5 gpc2811 (
      {stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17], stage3_12[18]},
      {stage3_13[12]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[2],stage4_14[4],stage4_13[6],stage4_12[6]}
   );
   gpc615_5 gpc2812 (
      {stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage3_13[13]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[3],stage4_14[5],stage4_13[7],stage4_12[7]}
   );
   gpc615_5 gpc2813 (
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28]},
      {stage3_13[14]},
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage4_16[2],stage4_15[4],stage4_14[6],stage4_13[8],stage4_12[8]}
   );
   gpc606_5 gpc2814 (
      {stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[3],stage4_15[5],stage4_14[7],stage4_13[9]}
   );
   gpc606_5 gpc2815 (
      {stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25], stage3_13[26]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[4],stage4_15[6],stage4_14[8],stage4_13[10]}
   );
   gpc606_5 gpc2816 (
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[5],stage4_15[7],stage4_14[9]}
   );
   gpc615_5 gpc2817 (
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16]},
      {stage3_16[6]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[1],stage4_17[3],stage4_16[6],stage4_15[8]}
   );
   gpc615_5 gpc2818 (
      {stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20], stage3_15[21]},
      {stage3_16[7]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[2],stage4_17[4],stage4_16[7],stage4_15[9]}
   );
   gpc615_5 gpc2819 (
      {stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25], stage3_15[26]},
      {stage3_16[8]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[3],stage4_17[5],stage4_16[8],stage4_15[10]}
   );
   gpc615_5 gpc2820 (
      {stage3_16[9], stage3_16[10], stage3_16[11], stage3_16[12], stage3_16[13]},
      {stage3_17[18]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[3],stage4_18[4],stage4_17[6],stage4_16[9]}
   );
   gpc615_5 gpc2821 (
      {stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17], stage3_16[18]},
      {stage3_17[19]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[4],stage4_18[5],stage4_17[7],stage4_16[10]}
   );
   gpc1163_5 gpc2822 (
      {stage3_18[12], stage3_18[13], stage3_18[14]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage3_20[0]},
      {stage3_21[0]},
      {stage4_22[0],stage4_21[0],stage4_20[2],stage4_19[5],stage4_18[6]}
   );
   gpc1163_5 gpc2823 (
      {stage3_18[15], stage3_18[16], stage3_18[17]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage3_20[1]},
      {stage3_21[1]},
      {stage4_22[1],stage4_21[1],stage4_20[3],stage4_19[6],stage4_18[7]}
   );
   gpc1163_5 gpc2824 (
      {stage3_18[18], stage3_18[19], stage3_18[20]},
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage3_20[2]},
      {stage3_21[2]},
      {stage4_22[2],stage4_21[2],stage4_20[4],stage4_19[7],stage4_18[8]}
   );
   gpc615_5 gpc2825 (
      {stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25]},
      {stage3_19[18]},
      {stage3_20[3], stage3_20[4], stage3_20[5], stage3_20[6], stage3_20[7], stage3_20[8]},
      {stage4_22[3],stage4_21[3],stage4_20[5],stage4_19[8],stage4_18[9]}
   );
   gpc615_5 gpc2826 (
      {stage3_18[26], stage3_18[27], stage3_18[28], stage3_18[29], stage3_18[30]},
      {stage3_19[19]},
      {stage3_20[9], stage3_20[10], stage3_20[11], stage3_20[12], stage3_20[13], stage3_20[14]},
      {stage4_22[4],stage4_21[4],stage4_20[6],stage4_19[9],stage4_18[10]}
   );
   gpc615_5 gpc2827 (
      {stage3_18[31], stage3_18[32], stage3_18[33], stage3_18[34], stage3_18[35]},
      {stage3_19[20]},
      {stage3_20[15], stage3_20[16], stage3_20[17], stage3_20[18], stage3_20[19], stage3_20[20]},
      {stage4_22[5],stage4_21[5],stage4_20[7],stage4_19[10],stage4_18[11]}
   );
   gpc615_5 gpc2828 (
      {stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24], stage3_19[25]},
      {stage3_20[21]},
      {stage3_21[3], stage3_21[4], stage3_21[5], stage3_21[6], stage3_21[7], stage3_21[8]},
      {stage4_23[0],stage4_22[6],stage4_21[6],stage4_20[8],stage4_19[11]}
   );
   gpc615_5 gpc2829 (
      {stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29], stage3_19[30]},
      {stage3_20[22]},
      {stage3_21[9], stage3_21[10], stage3_21[11], stage3_21[12], stage3_21[13], stage3_21[14]},
      {stage4_23[1],stage4_22[7],stage4_21[7],stage4_20[9],stage4_19[12]}
   );
   gpc615_5 gpc2830 (
      {stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34], 1'b0},
      {stage3_20[23]},
      {stage3_21[15], stage3_21[16], stage3_21[17], stage3_21[18], stage3_21[19], stage3_21[20]},
      {stage4_23[2],stage4_22[8],stage4_21[8],stage4_20[10],stage4_19[13]}
   );
   gpc606_5 gpc2831 (
      {stage3_20[24], stage3_20[25], stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[3],stage4_22[9],stage4_21[9],stage4_20[11]}
   );
   gpc606_5 gpc2832 (
      {stage3_21[21], stage3_21[22], stage3_21[23], stage3_21[24], stage3_21[25], stage3_21[26]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[1],stage4_23[4],stage4_22[10],stage4_21[10]}
   );
   gpc606_5 gpc2833 (
      {stage3_21[27], stage3_21[28], stage3_21[29], stage3_21[30], stage3_21[31], stage3_21[32]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[2],stage4_23[5],stage4_22[11],stage4_21[11]}
   );
   gpc615_5 gpc2834 (
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage3_23[12]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[2],stage4_24[3],stage4_23[6],stage4_22[12]}
   );
   gpc615_5 gpc2835 (
      {stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15]},
      {stage3_23[13]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[3],stage4_24[4],stage4_23[7],stage4_22[13]}
   );
   gpc615_5 gpc2836 (
      {stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19], stage3_22[20]},
      {stage3_23[14]},
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17]},
      {stage4_26[2],stage4_25[4],stage4_24[5],stage4_23[8],stage4_22[14]}
   );
   gpc615_5 gpc2837 (
      {stage3_22[21], stage3_22[22], stage3_22[23], stage3_22[24], stage3_22[25]},
      {stage3_23[15]},
      {stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23]},
      {stage4_26[3],stage4_25[5],stage4_24[6],stage4_23[9],stage4_22[15]}
   );
   gpc615_5 gpc2838 (
      {stage3_23[16], stage3_23[17], stage3_23[18], stage3_23[19], stage3_23[20]},
      {1'b0},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[4],stage4_25[6],stage4_24[7],stage4_23[10]}
   );
   gpc606_5 gpc2839 (
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[1],stage4_26[5],stage4_25[7]}
   );
   gpc606_5 gpc2840 (
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[1],stage4_27[2],stage4_26[6],stage4_25[8]}
   );
   gpc606_5 gpc2841 (
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[2],stage4_27[3],stage4_26[7],stage4_25[9]}
   );
   gpc606_5 gpc2842 (
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28], stage3_25[29]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage4_29[3],stage4_28[3],stage4_27[4],stage4_26[8],stage4_25[10]}
   );
   gpc606_5 gpc2843 (
      {stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33], stage3_25[34], stage3_25[35]},
      {stage3_27[24], stage3_27[25], stage3_27[26], stage3_27[27], stage3_27[28], stage3_27[29]},
      {stage4_29[4],stage4_28[4],stage4_27[5],stage4_26[9],stage4_25[11]}
   );
   gpc606_5 gpc2844 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[5],stage4_28[5],stage4_27[6],stage4_26[10]}
   );
   gpc606_5 gpc2845 (
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage4_30[1],stage4_29[6],stage4_28[6],stage4_27[7],stage4_26[11]}
   );
   gpc615_5 gpc2846 (
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16]},
      {stage3_27[30]},
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17]},
      {stage4_30[2],stage4_29[7],stage4_28[7],stage4_27[8],stage4_26[12]}
   );
   gpc615_5 gpc2847 (
      {stage3_26[17], stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21]},
      {stage3_27[31]},
      {stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21], stage3_28[22], stage3_28[23]},
      {stage4_30[3],stage4_29[8],stage4_28[8],stage4_27[9],stage4_26[13]}
   );
   gpc606_5 gpc2848 (
      {stage3_28[24], stage3_28[25], stage3_28[26], stage3_28[27], stage3_28[28], stage3_28[29]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[0],stage4_30[4],stage4_29[9],stage4_28[9]}
   );
   gpc606_5 gpc2849 (
      {stage3_28[30], stage3_28[31], stage3_28[32], stage3_28[33], stage3_28[34], stage3_28[35]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[1],stage4_30[5],stage4_29[10],stage4_28[10]}
   );
   gpc606_5 gpc2850 (
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[2],stage4_31[2],stage4_30[6],stage4_29[11]}
   );
   gpc606_5 gpc2851 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[3],stage4_31[3],stage4_30[7],stage4_29[12]}
   );
   gpc606_5 gpc2852 (
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[4],stage4_31[4],stage4_30[8],stage4_29[13]}
   );
   gpc606_5 gpc2853 (
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[3],stage4_32[5],stage4_31[5],stage4_30[9]}
   );
   gpc615_5 gpc2854 (
      {stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22]},
      {stage3_32[6]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[1],stage4_33[4],stage4_32[6],stage4_31[6]}
   );
   gpc615_5 gpc2855 (
      {stage3_31[23], stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27]},
      {stage3_32[7]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[2],stage4_33[5],stage4_32[7],stage4_31[7]}
   );
   gpc606_5 gpc2856 (
      {stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11], stage3_32[12], stage3_32[13]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[2],stage4_34[3],stage4_33[6],stage4_32[8]}
   );
   gpc606_5 gpc2857 (
      {stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17], stage3_32[18], stage3_32[19]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], 1'b0, 1'b0},
      {stage4_36[1],stage4_35[3],stage4_34[4],stage4_33[7],stage4_32[9]}
   );
   gpc606_5 gpc2858 (
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[2],stage4_35[4],stage4_34[5],stage4_33[8]}
   );
   gpc1_1 gpc2859 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc2860 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc2861 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc2862 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc2863 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc2864 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc2865 (
      {stage3_1[18]},
      {stage4_1[3]}
   );
   gpc1_1 gpc2866 (
      {stage3_1[19]},
      {stage4_1[4]}
   );
   gpc1_1 gpc2867 (
      {stage3_1[20]},
      {stage4_1[5]}
   );
   gpc1_1 gpc2868 (
      {stage3_1[21]},
      {stage4_1[6]}
   );
   gpc1_1 gpc2869 (
      {stage3_1[22]},
      {stage4_1[7]}
   );
   gpc1_1 gpc2870 (
      {stage3_1[23]},
      {stage4_1[8]}
   );
   gpc1_1 gpc2871 (
      {stage3_1[24]},
      {stage4_1[9]}
   );
   gpc1_1 gpc2872 (
      {stage3_1[25]},
      {stage4_1[10]}
   );
   gpc1_1 gpc2873 (
      {stage3_1[26]},
      {stage4_1[11]}
   );
   gpc1_1 gpc2874 (
      {stage3_1[27]},
      {stage4_1[12]}
   );
   gpc1_1 gpc2875 (
      {stage3_2[24]},
      {stage4_2[7]}
   );
   gpc1_1 gpc2876 (
      {stage3_3[32]},
      {stage4_3[9]}
   );
   gpc1_1 gpc2877 (
      {stage3_3[33]},
      {stage4_3[10]}
   );
   gpc1_1 gpc2878 (
      {stage3_3[34]},
      {stage4_3[11]}
   );
   gpc1_1 gpc2879 (
      {stage3_4[30]},
      {stage4_4[10]}
   );
   gpc1_1 gpc2880 (
      {stage3_4[31]},
      {stage4_4[11]}
   );
   gpc1_1 gpc2881 (
      {stage3_4[32]},
      {stage4_4[12]}
   );
   gpc1_1 gpc2882 (
      {stage3_4[33]},
      {stage4_4[13]}
   );
   gpc1_1 gpc2883 (
      {stage3_4[34]},
      {stage4_4[14]}
   );
   gpc1_1 gpc2884 (
      {stage3_4[35]},
      {stage4_4[15]}
   );
   gpc1_1 gpc2885 (
      {stage3_6[16]},
      {stage4_6[11]}
   );
   gpc1_1 gpc2886 (
      {stage3_6[17]},
      {stage4_6[12]}
   );
   gpc1_1 gpc2887 (
      {stage3_6[18]},
      {stage4_6[13]}
   );
   gpc1_1 gpc2888 (
      {stage3_6[19]},
      {stage4_6[14]}
   );
   gpc1_1 gpc2889 (
      {stage3_7[14]},
      {stage4_7[5]}
   );
   gpc1_1 gpc2890 (
      {stage3_7[15]},
      {stage4_7[6]}
   );
   gpc1_1 gpc2891 (
      {stage3_7[16]},
      {stage4_7[7]}
   );
   gpc1_1 gpc2892 (
      {stage3_7[17]},
      {stage4_7[8]}
   );
   gpc1_1 gpc2893 (
      {stage3_7[18]},
      {stage4_7[9]}
   );
   gpc1_1 gpc2894 (
      {stage3_7[19]},
      {stage4_7[10]}
   );
   gpc1_1 gpc2895 (
      {stage3_7[20]},
      {stage4_7[11]}
   );
   gpc1_1 gpc2896 (
      {stage3_7[21]},
      {stage4_7[12]}
   );
   gpc1_1 gpc2897 (
      {stage3_7[22]},
      {stage4_7[13]}
   );
   gpc1_1 gpc2898 (
      {stage3_7[23]},
      {stage4_7[14]}
   );
   gpc1_1 gpc2899 (
      {stage3_9[21]},
      {stage4_9[9]}
   );
   gpc1_1 gpc2900 (
      {stage3_10[13]},
      {stage4_10[9]}
   );
   gpc1_1 gpc2901 (
      {stage3_10[14]},
      {stage4_10[10]}
   );
   gpc1_1 gpc2902 (
      {stage3_10[15]},
      {stage4_10[11]}
   );
   gpc1_1 gpc2903 (
      {stage3_10[16]},
      {stage4_10[12]}
   );
   gpc1_1 gpc2904 (
      {stage3_10[17]},
      {stage4_10[13]}
   );
   gpc1_1 gpc2905 (
      {stage3_10[18]},
      {stage4_10[14]}
   );
   gpc1_1 gpc2906 (
      {stage3_11[24]},
      {stage4_11[9]}
   );
   gpc1_1 gpc2907 (
      {stage3_11[25]},
      {stage4_11[10]}
   );
   gpc1_1 gpc2908 (
      {stage3_12[29]},
      {stage4_12[9]}
   );
   gpc1_1 gpc2909 (
      {stage3_12[30]},
      {stage4_12[10]}
   );
   gpc1_1 gpc2910 (
      {stage3_12[31]},
      {stage4_12[11]}
   );
   gpc1_1 gpc2911 (
      {stage3_13[27]},
      {stage4_13[11]}
   );
   gpc1_1 gpc2912 (
      {stage3_13[28]},
      {stage4_13[12]}
   );
   gpc1_1 gpc2913 (
      {stage3_13[29]},
      {stage4_13[13]}
   );
   gpc1_1 gpc2914 (
      {stage3_13[30]},
      {stage4_13[14]}
   );
   gpc1_1 gpc2915 (
      {stage3_13[31]},
      {stage4_13[15]}
   );
   gpc1_1 gpc2916 (
      {stage3_13[32]},
      {stage4_13[16]}
   );
   gpc1_1 gpc2917 (
      {stage3_13[33]},
      {stage4_13[17]}
   );
   gpc1_1 gpc2918 (
      {stage3_13[34]},
      {stage4_13[18]}
   );
   gpc1_1 gpc2919 (
      {stage3_13[35]},
      {stage4_13[19]}
   );
   gpc1_1 gpc2920 (
      {stage3_13[36]},
      {stage4_13[20]}
   );
   gpc1_1 gpc2921 (
      {stage3_14[24]},
      {stage4_14[10]}
   );
   gpc1_1 gpc2922 (
      {stage3_14[25]},
      {stage4_14[11]}
   );
   gpc1_1 gpc2923 (
      {stage3_15[27]},
      {stage4_15[11]}
   );
   gpc1_1 gpc2924 (
      {stage3_15[28]},
      {stage4_15[12]}
   );
   gpc1_1 gpc2925 (
      {stage3_15[29]},
      {stage4_15[13]}
   );
   gpc1_1 gpc2926 (
      {stage3_15[30]},
      {stage4_15[14]}
   );
   gpc1_1 gpc2927 (
      {stage3_15[31]},
      {stage4_15[15]}
   );
   gpc1_1 gpc2928 (
      {stage3_15[32]},
      {stage4_15[16]}
   );
   gpc1_1 gpc2929 (
      {stage3_16[19]},
      {stage4_16[11]}
   );
   gpc1_1 gpc2930 (
      {stage3_16[20]},
      {stage4_16[12]}
   );
   gpc1_1 gpc2931 (
      {stage3_16[21]},
      {stage4_16[13]}
   );
   gpc1_1 gpc2932 (
      {stage3_16[22]},
      {stage4_16[14]}
   );
   gpc1_1 gpc2933 (
      {stage3_16[23]},
      {stage4_16[15]}
   );
   gpc1_1 gpc2934 (
      {stage3_16[24]},
      {stage4_16[16]}
   );
   gpc1_1 gpc2935 (
      {stage3_16[25]},
      {stage4_16[17]}
   );
   gpc1_1 gpc2936 (
      {stage3_16[26]},
      {stage4_16[18]}
   );
   gpc1_1 gpc2937 (
      {stage3_18[36]},
      {stage4_18[12]}
   );
   gpc1_1 gpc2938 (
      {stage3_18[37]},
      {stage4_18[13]}
   );
   gpc1_1 gpc2939 (
      {stage3_20[30]},
      {stage4_20[12]}
   );
   gpc1_1 gpc2940 (
      {stage3_20[31]},
      {stage4_20[13]}
   );
   gpc1_1 gpc2941 (
      {stage3_20[32]},
      {stage4_20[14]}
   );
   gpc1_1 gpc2942 (
      {stage3_20[33]},
      {stage4_20[15]}
   );
   gpc1_1 gpc2943 (
      {stage3_20[34]},
      {stage4_20[16]}
   );
   gpc1_1 gpc2944 (
      {stage3_20[35]},
      {stage4_20[17]}
   );
   gpc1_1 gpc2945 (
      {stage3_20[36]},
      {stage4_20[18]}
   );
   gpc1_1 gpc2946 (
      {stage3_22[26]},
      {stage4_22[16]}
   );
   gpc1_1 gpc2947 (
      {stage3_22[27]},
      {stage4_22[17]}
   );
   gpc1_1 gpc2948 (
      {stage3_22[28]},
      {stage4_22[18]}
   );
   gpc1_1 gpc2949 (
      {stage3_22[29]},
      {stage4_22[19]}
   );
   gpc1_1 gpc2950 (
      {stage3_22[30]},
      {stage4_22[20]}
   );
   gpc1_1 gpc2951 (
      {stage3_22[31]},
      {stage4_22[21]}
   );
   gpc1_1 gpc2952 (
      {stage3_22[32]},
      {stage4_22[22]}
   );
   gpc1_1 gpc2953 (
      {stage3_22[33]},
      {stage4_22[23]}
   );
   gpc1_1 gpc2954 (
      {stage3_22[34]},
      {stage4_22[24]}
   );
   gpc1_1 gpc2955 (
      {stage3_26[22]},
      {stage4_26[14]}
   );
   gpc1_1 gpc2956 (
      {stage3_26[23]},
      {stage4_26[15]}
   );
   gpc1_1 gpc2957 (
      {stage3_27[32]},
      {stage4_27[10]}
   );
   gpc1_1 gpc2958 (
      {stage3_27[33]},
      {stage4_27[11]}
   );
   gpc1_1 gpc2959 (
      {stage3_27[34]},
      {stage4_27[12]}
   );
   gpc1_1 gpc2960 (
      {stage3_27[35]},
      {stage4_27[13]}
   );
   gpc1_1 gpc2961 (
      {stage3_27[36]},
      {stage4_27[14]}
   );
   gpc1_1 gpc2962 (
      {stage3_27[37]},
      {stage4_27[15]}
   );
   gpc1_1 gpc2963 (
      {stage3_27[38]},
      {stage4_27[16]}
   );
   gpc1_1 gpc2964 (
      {stage3_28[36]},
      {stage4_28[11]}
   );
   gpc1_1 gpc2965 (
      {stage3_28[37]},
      {stage4_28[12]}
   );
   gpc1_1 gpc2966 (
      {stage3_28[38]},
      {stage4_28[13]}
   );
   gpc1_1 gpc2967 (
      {stage3_28[39]},
      {stage4_28[14]}
   );
   gpc1_1 gpc2968 (
      {stage3_28[40]},
      {stage4_28[15]}
   );
   gpc1_1 gpc2969 (
      {stage3_28[41]},
      {stage4_28[16]}
   );
   gpc1_1 gpc2970 (
      {stage3_28[42]},
      {stage4_28[17]}
   );
   gpc1_1 gpc2971 (
      {stage3_28[43]},
      {stage4_28[18]}
   );
   gpc1_1 gpc2972 (
      {stage3_28[44]},
      {stage4_28[19]}
   );
   gpc1_1 gpc2973 (
      {stage3_29[18]},
      {stage4_29[14]}
   );
   gpc1_1 gpc2974 (
      {stage3_29[19]},
      {stage4_29[15]}
   );
   gpc1_1 gpc2975 (
      {stage3_29[20]},
      {stage4_29[16]}
   );
   gpc1_1 gpc2976 (
      {stage3_29[21]},
      {stage4_29[17]}
   );
   gpc1_1 gpc2977 (
      {stage3_29[22]},
      {stage4_29[18]}
   );
   gpc1_1 gpc2978 (
      {stage3_29[23]},
      {stage4_29[19]}
   );
   gpc1_1 gpc2979 (
      {stage3_29[24]},
      {stage4_29[20]}
   );
   gpc1_1 gpc2980 (
      {stage3_29[25]},
      {stage4_29[21]}
   );
   gpc1_1 gpc2981 (
      {stage3_29[26]},
      {stage4_29[22]}
   );
   gpc1_1 gpc2982 (
      {stage3_29[27]},
      {stage4_29[23]}
   );
   gpc1_1 gpc2983 (
      {stage3_31[28]},
      {stage4_31[8]}
   );
   gpc1_1 gpc2984 (
      {stage3_31[29]},
      {stage4_31[9]}
   );
   gpc1_1 gpc2985 (
      {stage3_31[30]},
      {stage4_31[10]}
   );
   gpc1_1 gpc2986 (
      {stage3_31[31]},
      {stage4_31[11]}
   );
   gpc1_1 gpc2987 (
      {stage3_31[32]},
      {stage4_31[12]}
   );
   gpc1_1 gpc2988 (
      {stage3_31[33]},
      {stage4_31[13]}
   );
   gpc1_1 gpc2989 (
      {stage3_31[34]},
      {stage4_31[14]}
   );
   gpc1_1 gpc2990 (
      {stage3_31[35]},
      {stage4_31[15]}
   );
   gpc1_1 gpc2991 (
      {stage3_31[36]},
      {stage4_31[16]}
   );
   gpc1_1 gpc2992 (
      {stage3_35[6]},
      {stage4_35[5]}
   );
   gpc1_1 gpc2993 (
      {stage3_35[7]},
      {stage4_35[6]}
   );
   gpc1_1 gpc2994 (
      {stage3_35[8]},
      {stage4_35[7]}
   );
   gpc1_1 gpc2995 (
      {stage3_35[9]},
      {stage4_35[8]}
   );
   gpc1_1 gpc2996 (
      {stage3_35[10]},
      {stage4_35[9]}
   );
   gpc1_1 gpc2997 (
      {stage3_35[11]},
      {stage4_35[10]}
   );
   gpc1_1 gpc2998 (
      {stage3_35[12]},
      {stage4_35[11]}
   );
   gpc1_1 gpc2999 (
      {stage3_36[0]},
      {stage4_36[3]}
   );
   gpc1_1 gpc3000 (
      {stage3_36[1]},
      {stage4_36[4]}
   );
   gpc1_1 gpc3001 (
      {stage3_36[2]},
      {stage4_36[5]}
   );
   gpc606_5 gpc3002 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc3003 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc606_5 gpc3004 (
      {stage4_1[6], stage4_1[7], stage4_1[8], stage4_1[9], stage4_1[10], stage4_1[11]},
      {stage4_3[6], stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage5_5[1],stage5_4[2],stage5_3[2],stage5_2[2],stage5_1[2]}
   );
   gpc606_5 gpc3005 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[2],stage5_4[3]}
   );
   gpc606_5 gpc3006 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11]},
      {stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[3],stage5_4[4]}
   );
   gpc606_5 gpc3007 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[2],stage5_7[2],stage5_6[2],stage5_5[4]}
   );
   gpc606_5 gpc3008 (
      {stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage5_9[1],stage5_8[3],stage5_7[3],stage5_6[3],stage5_5[5]}
   );
   gpc606_5 gpc3009 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[2],stage5_8[4]}
   );
   gpc615_5 gpc3010 (
      {stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], stage4_10[10]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[0],stage5_12[1],stage5_11[1],stage5_10[1]}
   );
   gpc606_5 gpc3011 (
      {stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[1],stage5_13[1],stage5_12[2],stage5_11[2]}
   );
   gpc606_5 gpc3012 (
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[1],stage5_14[2],stage5_13[2],stage5_12[3]}
   );
   gpc606_5 gpc3013 (
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[1],stage5_15[2],stage5_14[3],stage5_13[3]}
   );
   gpc606_5 gpc3014 (
      {stage4_13[12], stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17]},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[2],stage5_15[3],stage5_14[4],stage5_13[4]}
   );
   gpc615_5 gpc3015 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[12]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[2],stage5_16[3],stage5_15[4],stage5_14[5]}
   );
   gpc207_4 gpc3016 (
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12]},
      {stage4_18[0], stage4_18[1]},
      {stage5_19[0],stage5_18[1],stage5_17[3],stage5_16[4]}
   );
   gpc606_5 gpc3017 (
      {stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18]},
      {stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6], stage4_18[7]},
      {stage5_20[0],stage5_19[1],stage5_18[2],stage5_17[4],stage5_16[5]}
   );
   gpc606_5 gpc3018 (
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[2],stage5_18[3],stage5_17[5]}
   );
   gpc615_5 gpc3019 (
      {stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11], stage4_18[12]},
      {stage4_19[6]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[2],stage5_19[3],stage5_18[4]}
   );
   gpc615_5 gpc3020 (
      {stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage4_20[6]},
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5]},
      {stage5_23[0],stage5_22[1],stage5_21[2],stage5_20[3],stage5_19[4]}
   );
   gpc623_5 gpc3021 (
      {stage4_20[7], stage4_20[8], stage4_20[9]},
      {stage4_21[6], stage4_21[7]},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[1],stage5_22[2],stage5_21[3],stage5_20[4]}
   );
   gpc623_5 gpc3022 (
      {stage4_20[10], stage4_20[11], stage4_20[12]},
      {stage4_21[8], stage4_21[9]},
      {stage4_22[6], stage4_22[7], stage4_22[8], stage4_22[9], stage4_22[10], stage4_22[11]},
      {stage5_24[1],stage5_23[2],stage5_22[3],stage5_21[4],stage5_20[5]}
   );
   gpc623_5 gpc3023 (
      {stage4_20[13], stage4_20[14], stage4_20[15]},
      {stage4_21[10], stage4_21[11]},
      {stage4_22[12], stage4_22[13], stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17]},
      {stage5_24[2],stage5_23[3],stage5_22[4],stage5_21[5],stage5_20[6]}
   );
   gpc615_5 gpc3024 (
      {stage4_22[18], stage4_22[19], stage4_22[20], stage4_22[21], stage4_22[22]},
      {stage4_23[0]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage5_26[0],stage5_25[0],stage5_24[3],stage5_23[4],stage5_22[5]}
   );
   gpc615_5 gpc3025 (
      {stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[6]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[1],stage5_25[1],stage5_24[4],stage5_23[5]}
   );
   gpc615_5 gpc3026 (
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10]},
      {stage4_24[7]},
      {stage4_25[6], stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11]},
      {stage5_27[1],stage5_26[2],stage5_25[2],stage5_24[5],stage5_23[6]}
   );
   gpc606_5 gpc3027 (
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[0],stage5_27[2],stage5_26[3]}
   );
   gpc615_5 gpc3028 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10]},
      {stage4_27[0]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage5_30[1],stage5_29[1],stage5_28[1],stage5_27[3],stage5_26[4]}
   );
   gpc615_5 gpc3029 (
      {stage4_26[11], stage4_26[12], stage4_26[13], stage4_26[14], stage4_26[15]},
      {stage4_27[1]},
      {stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage5_30[2],stage5_29[2],stage5_28[2],stage5_27[4],stage5_26[5]}
   );
   gpc615_5 gpc3030 (
      {stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5], stage4_27[6]},
      {stage4_28[18]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[3],stage5_29[3],stage5_28[3],stage5_27[5]}
   );
   gpc615_5 gpc3031 (
      {stage4_27[7], stage4_27[8], stage4_27[9], stage4_27[10], stage4_27[11]},
      {stage4_28[19]},
      {stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11]},
      {stage5_31[1],stage5_30[4],stage5_29[4],stage5_28[4],stage5_27[6]}
   );
   gpc615_5 gpc3032 (
      {stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {1'b0},
      {stage4_29[12], stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17]},
      {stage5_31[2],stage5_30[5],stage5_29[5],stage5_28[5],stage5_27[7]}
   );
   gpc606_5 gpc3033 (
      {stage4_29[18], stage4_29[19], stage4_29[20], stage4_29[21], stage4_29[22], stage4_29[23]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[3],stage5_30[6],stage5_29[6]}
   );
   gpc1163_5 gpc3034 (
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9], stage4_31[10], stage4_31[11]},
      {stage4_32[0]},
      {stage4_33[0]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[4],stage5_30[7]}
   );
   gpc1163_5 gpc3035 (
      {stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage4_31[12], stage4_31[13], stage4_31[14], stage4_31[15], stage4_31[16], 1'b0},
      {stage4_32[1]},
      {stage4_33[1]},
      {stage5_34[1],stage5_33[2],stage5_32[2],stage5_31[5],stage5_30[8]}
   );
   gpc606_5 gpc3036 (
      {stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5], stage4_32[6], stage4_32[7]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[0],stage5_34[2],stage5_33[3],stage5_32[3]}
   );
   gpc606_5 gpc3037 (
      {stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5], stage4_33[6], stage4_33[7]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[1],stage5_35[1],stage5_34[3],stage5_33[4]}
   );
   gpc1_1 gpc3038 (
      {stage4_1[12]},
      {stage5_1[3]}
   );
   gpc1_1 gpc3039 (
      {stage4_2[6]},
      {stage5_2[3]}
   );
   gpc1_1 gpc3040 (
      {stage4_2[7]},
      {stage5_2[4]}
   );
   gpc1_1 gpc3041 (
      {stage4_4[12]},
      {stage5_4[5]}
   );
   gpc1_1 gpc3042 (
      {stage4_4[13]},
      {stage5_4[6]}
   );
   gpc1_1 gpc3043 (
      {stage4_4[14]},
      {stage5_4[7]}
   );
   gpc1_1 gpc3044 (
      {stage4_4[15]},
      {stage5_4[8]}
   );
   gpc1_1 gpc3045 (
      {stage4_6[12]},
      {stage5_6[4]}
   );
   gpc1_1 gpc3046 (
      {stage4_6[13]},
      {stage5_6[5]}
   );
   gpc1_1 gpc3047 (
      {stage4_6[14]},
      {stage5_6[6]}
   );
   gpc1_1 gpc3048 (
      {stage4_7[12]},
      {stage5_7[4]}
   );
   gpc1_1 gpc3049 (
      {stage4_7[13]},
      {stage5_7[5]}
   );
   gpc1_1 gpc3050 (
      {stage4_7[14]},
      {stage5_7[6]}
   );
   gpc1_1 gpc3051 (
      {stage4_8[6]},
      {stage5_8[5]}
   );
   gpc1_1 gpc3052 (
      {stage4_8[7]},
      {stage5_8[6]}
   );
   gpc1_1 gpc3053 (
      {stage4_9[0]},
      {stage5_9[3]}
   );
   gpc1_1 gpc3054 (
      {stage4_9[1]},
      {stage5_9[4]}
   );
   gpc1_1 gpc3055 (
      {stage4_9[2]},
      {stage5_9[5]}
   );
   gpc1_1 gpc3056 (
      {stage4_9[3]},
      {stage5_9[6]}
   );
   gpc1_1 gpc3057 (
      {stage4_9[4]},
      {stage5_9[7]}
   );
   gpc1_1 gpc3058 (
      {stage4_9[5]},
      {stage5_9[8]}
   );
   gpc1_1 gpc3059 (
      {stage4_9[6]},
      {stage5_9[9]}
   );
   gpc1_1 gpc3060 (
      {stage4_9[7]},
      {stage5_9[10]}
   );
   gpc1_1 gpc3061 (
      {stage4_9[8]},
      {stage5_9[11]}
   );
   gpc1_1 gpc3062 (
      {stage4_9[9]},
      {stage5_9[12]}
   );
   gpc1_1 gpc3063 (
      {stage4_10[11]},
      {stage5_10[2]}
   );
   gpc1_1 gpc3064 (
      {stage4_10[12]},
      {stage5_10[3]}
   );
   gpc1_1 gpc3065 (
      {stage4_10[13]},
      {stage5_10[4]}
   );
   gpc1_1 gpc3066 (
      {stage4_10[14]},
      {stage5_10[5]}
   );
   gpc1_1 gpc3067 (
      {stage4_11[7]},
      {stage5_11[3]}
   );
   gpc1_1 gpc3068 (
      {stage4_11[8]},
      {stage5_11[4]}
   );
   gpc1_1 gpc3069 (
      {stage4_11[9]},
      {stage5_11[5]}
   );
   gpc1_1 gpc3070 (
      {stage4_11[10]},
      {stage5_11[6]}
   );
   gpc1_1 gpc3071 (
      {stage4_13[18]},
      {stage5_13[5]}
   );
   gpc1_1 gpc3072 (
      {stage4_13[19]},
      {stage5_13[6]}
   );
   gpc1_1 gpc3073 (
      {stage4_13[20]},
      {stage5_13[7]}
   );
   gpc1_1 gpc3074 (
      {stage4_14[11]},
      {stage5_14[6]}
   );
   gpc1_1 gpc3075 (
      {stage4_15[13]},
      {stage5_15[5]}
   );
   gpc1_1 gpc3076 (
      {stage4_15[14]},
      {stage5_15[6]}
   );
   gpc1_1 gpc3077 (
      {stage4_15[15]},
      {stage5_15[7]}
   );
   gpc1_1 gpc3078 (
      {stage4_15[16]},
      {stage5_15[8]}
   );
   gpc1_1 gpc3079 (
      {stage4_17[6]},
      {stage5_17[6]}
   );
   gpc1_1 gpc3080 (
      {stage4_17[7]},
      {stage5_17[7]}
   );
   gpc1_1 gpc3081 (
      {stage4_18[13]},
      {stage5_18[5]}
   );
   gpc1_1 gpc3082 (
      {stage4_19[12]},
      {stage5_19[5]}
   );
   gpc1_1 gpc3083 (
      {stage4_19[13]},
      {stage5_19[6]}
   );
   gpc1_1 gpc3084 (
      {stage4_20[16]},
      {stage5_20[7]}
   );
   gpc1_1 gpc3085 (
      {stage4_20[17]},
      {stage5_20[8]}
   );
   gpc1_1 gpc3086 (
      {stage4_20[18]},
      {stage5_20[9]}
   );
   gpc1_1 gpc3087 (
      {stage4_22[23]},
      {stage5_22[6]}
   );
   gpc1_1 gpc3088 (
      {stage4_22[24]},
      {stage5_22[7]}
   );
   gpc1_1 gpc3089 (
      {stage4_30[6]},
      {stage5_30[9]}
   );
   gpc1_1 gpc3090 (
      {stage4_30[7]},
      {stage5_30[10]}
   );
   gpc1_1 gpc3091 (
      {stage4_30[8]},
      {stage5_30[11]}
   );
   gpc1_1 gpc3092 (
      {stage4_30[9]},
      {stage5_30[12]}
   );
   gpc1_1 gpc3093 (
      {stage4_32[8]},
      {stage5_32[4]}
   );
   gpc1_1 gpc3094 (
      {stage4_32[9]},
      {stage5_32[5]}
   );
   gpc1_1 gpc3095 (
      {stage4_33[8]},
      {stage5_33[5]}
   );
   gpc1_1 gpc3096 (
      {stage4_35[6]},
      {stage5_35[2]}
   );
   gpc1_1 gpc3097 (
      {stage4_35[7]},
      {stage5_35[3]}
   );
   gpc1_1 gpc3098 (
      {stage4_35[8]},
      {stage5_35[4]}
   );
   gpc1_1 gpc3099 (
      {stage4_35[9]},
      {stage5_35[5]}
   );
   gpc1_1 gpc3100 (
      {stage4_35[10]},
      {stage5_35[6]}
   );
   gpc1_1 gpc3101 (
      {stage4_35[11]},
      {stage5_35[7]}
   );
   gpc1_1 gpc3102 (
      {stage4_36[0]},
      {stage5_36[2]}
   );
   gpc1_1 gpc3103 (
      {stage4_36[1]},
      {stage5_36[3]}
   );
   gpc1_1 gpc3104 (
      {stage4_36[2]},
      {stage5_36[4]}
   );
   gpc1_1 gpc3105 (
      {stage4_36[3]},
      {stage5_36[5]}
   );
   gpc1_1 gpc3106 (
      {stage4_36[4]},
      {stage5_36[6]}
   );
   gpc1_1 gpc3107 (
      {stage4_36[5]},
      {stage5_36[7]}
   );
   gpc1_1 gpc3108 (
      {stage4_37[0]},
      {stage5_37[1]}
   );
   gpc1343_5 gpc3109 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3]},
      {stage5_3[0], stage5_3[1], stage5_3[2]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc606_5 gpc3110 (
      {stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1]}
   );
   gpc606_5 gpc3111 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[1],stage6_7[1],stage6_6[1],stage6_5[2]}
   );
   gpc1163_5 gpc3112 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage5_10[0]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[2]}
   );
   gpc1163_5 gpc3113 (
      {stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage5_9[6], stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], stage5_9[11]},
      {stage5_10[1]},
      {stage5_11[1]},
      {stage6_12[1],stage6_11[1],stage6_10[1],stage6_9[2],stage6_8[3]}
   );
   gpc615_5 gpc3114 (
      {stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6]},
      {stage5_12[0]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[2],stage6_11[2]}
   );
   gpc1343_5 gpc3115 (
      {stage5_14[0], stage5_14[1], stage5_14[2]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[1]}
   );
   gpc1343_5 gpc3116 (
      {stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_17[1]},
      {stage6_18[1],stage6_17[1],stage6_16[1],stage6_15[2],stage6_14[2]}
   );
   gpc606_5 gpc3117 (
      {stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6], stage5_17[7]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[2],stage6_17[2]}
   );
   gpc615_5 gpc3118 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4]},
      {stage5_19[6]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage6_22[0],stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[3]}
   );
   gpc606_5 gpc3119 (
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5]},
      {stage6_25[0],stage6_24[0],stage6_23[0],stage6_22[1],stage6_21[2]}
   );
   gpc615_5 gpc3120 (
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4]},
      {stage5_23[6]},
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage6_26[0],stage6_25[1],stage6_24[1],stage6_23[1],stage6_22[2]}
   );
   gpc1163_5 gpc3121 (
      {stage5_25[0], stage5_25[1], stage5_25[2]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5]},
      {stage5_27[0]},
      {stage5_28[0]},
      {stage6_29[0],stage6_28[0],stage6_27[0],stage6_26[1],stage6_25[2]}
   );
   gpc117_4 gpc3122 (
      {stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[1]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[1]}
   );
   gpc606_5 gpc3123 (
      {stage5_28[2], stage5_28[3], stage5_28[4], stage5_28[5], 1'b0, 1'b0},
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5]},
      {stage6_32[0],stage6_31[0],stage6_30[1],stage6_29[2],stage6_28[2]}
   );
   gpc606_5 gpc3124 (
      {stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5], stage5_29[6]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[1],stage6_31[1],stage6_30[2],stage6_29[3]}
   );
   gpc615_5 gpc3125 (
      {stage5_30[6], stage5_30[7], stage5_30[8], stage5_30[9], stage5_30[10]},
      {1'b0},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage6_34[0],stage6_33[1],stage6_32[2],stage6_31[2],stage6_30[3]}
   );
   gpc606_5 gpc3126 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[0],stage6_35[0],stage6_34[1],stage6_33[2]}
   );
   gpc615_5 gpc3127 (
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], 1'b0},
      {stage5_35[6]},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5]},
      {stage6_38[0],stage6_37[1],stage6_36[1],stage6_35[1],stage6_34[2]}
   );
   gpc1_1 gpc3128 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc3129 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc3130 (
      {stage5_2[4]},
      {stage6_2[1]}
   );
   gpc1_1 gpc3131 (
      {stage5_4[7]},
      {stage6_4[2]}
   );
   gpc1_1 gpc3132 (
      {stage5_4[8]},
      {stage6_4[3]}
   );
   gpc1_1 gpc3133 (
      {stage5_6[6]},
      {stage6_6[2]}
   );
   gpc1_1 gpc3134 (
      {stage5_7[6]},
      {stage6_7[2]}
   );
   gpc1_1 gpc3135 (
      {stage5_8[6]},
      {stage6_8[4]}
   );
   gpc1_1 gpc3136 (
      {stage5_9[12]},
      {stage6_9[3]}
   );
   gpc1_1 gpc3137 (
      {stage5_10[2]},
      {stage6_10[2]}
   );
   gpc1_1 gpc3138 (
      {stage5_10[3]},
      {stage6_10[3]}
   );
   gpc1_1 gpc3139 (
      {stage5_10[4]},
      {stage6_10[4]}
   );
   gpc1_1 gpc3140 (
      {stage5_10[5]},
      {stage6_10[5]}
   );
   gpc1_1 gpc3141 (
      {stage5_12[1]},
      {stage6_12[3]}
   );
   gpc1_1 gpc3142 (
      {stage5_12[2]},
      {stage6_12[4]}
   );
   gpc1_1 gpc3143 (
      {stage5_12[3]},
      {stage6_12[5]}
   );
   gpc1_1 gpc3144 (
      {stage5_13[6]},
      {stage6_13[1]}
   );
   gpc1_1 gpc3145 (
      {stage5_13[7]},
      {stage6_13[2]}
   );
   gpc1_1 gpc3146 (
      {stage5_14[6]},
      {stage6_14[3]}
   );
   gpc1_1 gpc3147 (
      {stage5_15[8]},
      {stage6_15[3]}
   );
   gpc1_1 gpc3148 (
      {stage5_18[5]},
      {stage6_18[4]}
   );
   gpc1_1 gpc3149 (
      {stage5_20[6]},
      {stage6_20[2]}
   );
   gpc1_1 gpc3150 (
      {stage5_20[7]},
      {stage6_20[3]}
   );
   gpc1_1 gpc3151 (
      {stage5_20[8]},
      {stage6_20[4]}
   );
   gpc1_1 gpc3152 (
      {stage5_20[9]},
      {stage6_20[5]}
   );
   gpc1_1 gpc3153 (
      {stage5_22[5]},
      {stage6_22[3]}
   );
   gpc1_1 gpc3154 (
      {stage5_22[6]},
      {stage6_22[4]}
   );
   gpc1_1 gpc3155 (
      {stage5_22[7]},
      {stage6_22[5]}
   );
   gpc1_1 gpc3156 (
      {stage5_30[11]},
      {stage6_30[4]}
   );
   gpc1_1 gpc3157 (
      {stage5_30[12]},
      {stage6_30[5]}
   );
   gpc1_1 gpc3158 (
      {stage5_35[7]},
      {stage6_35[2]}
   );
   gpc1_1 gpc3159 (
      {stage5_36[6]},
      {stage6_36[2]}
   );
   gpc1_1 gpc3160 (
      {stage5_36[7]},
      {stage6_36[3]}
   );
   gpc1_1 gpc3161 (
      {stage5_37[0]},
      {stage6_37[2]}
   );
   gpc1_1 gpc3162 (
      {stage5_37[1]},
      {stage6_37[3]}
   );
   gpc223_4 gpc3163 (
      {stage6_4[0], stage6_4[1], stage6_4[2]},
      {stage6_5[0], stage6_5[1]},
      {stage6_6[0], stage6_6[1]},
      {stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0]}
   );
   gpc23_3 gpc3164 (
      {stage6_7[0], stage6_7[1], stage6_7[2]},
      {stage6_8[0], stage6_8[1]},
      {stage7_9[0],stage7_8[0],stage7_7[1]}
   );
   gpc1343_5 gpc3165 (
      {stage6_8[2], stage6_8[3], stage6_8[4]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3]},
      {stage6_10[0], stage6_10[1], stage6_10[2]},
      {stage6_11[0]},
      {stage7_12[0],stage7_11[0],stage7_10[0],stage7_9[1],stage7_8[1]}
   );
   gpc623_5 gpc3166 (
      {stage6_10[3], stage6_10[4], stage6_10[5]},
      {stage6_11[1], stage6_11[2]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage7_14[0],stage7_13[0],stage7_12[1],stage7_11[1],stage7_10[1]}
   );
   gpc1343_5 gpc3167 (
      {stage6_13[0], stage6_13[1], stage6_13[2]},
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3]},
      {stage6_15[0], stage6_15[1], stage6_15[2]},
      {stage6_16[0]},
      {stage7_17[0],stage7_16[0],stage7_15[0],stage7_14[1],stage7_13[1]}
   );
   gpc3_2 gpc3168 (
      {stage6_17[0], stage6_17[1], stage6_17[2]},
      {stage7_18[0],stage7_17[1]}
   );
   gpc1415_5 gpc3169 (
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4]},
      {stage6_19[0]},
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3]},
      {stage6_21[0]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[1]}
   );
   gpc623_5 gpc3170 (
      {stage6_20[4], stage6_20[5], 1'b0},
      {stage6_21[1], stage6_21[2]},
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3], stage6_22[4], stage6_22[5]},
      {stage7_24[0],stage7_23[0],stage7_22[1],stage7_21[1],stage7_20[1]}
   );
   gpc1343_5 gpc3171 (
      {stage6_23[0], stage6_23[1], 1'b0},
      {stage6_24[0], stage6_24[1], 1'b0, 1'b0},
      {stage6_25[0], stage6_25[1], stage6_25[2]},
      {stage6_26[0]},
      {stage7_27[0],stage7_26[0],stage7_25[0],stage7_24[1],stage7_23[1]}
   );
   gpc223_4 gpc3172 (
      {stage6_27[0], stage6_27[1], 1'b0},
      {stage6_28[0], stage6_28[1]},
      {stage6_29[0], stage6_29[1]},
      {stage7_30[0],stage7_29[0],stage7_28[0],stage7_27[1]}
   );
   gpc623_5 gpc3173 (
      {stage6_28[2], 1'b0, 1'b0},
      {stage6_29[2], stage6_29[3]},
      {stage6_30[0], stage6_30[1], stage6_30[2], stage6_30[3], stage6_30[4], stage6_30[5]},
      {stage7_32[0],stage7_31[0],stage7_30[1],stage7_29[1],stage7_28[1]}
   );
   gpc1163_5 gpc3174 (
      {stage6_31[0], stage6_31[1], stage6_31[2]},
      {stage6_32[0], stage6_32[1], stage6_32[2], 1'b0, 1'b0, 1'b0},
      {stage6_33[0]},
      {stage6_34[0]},
      {stage7_35[0],stage7_34[0],stage7_33[0],stage7_32[1],stage7_31[1]}
   );
   gpc1343_5 gpc3175 (
      {stage6_33[1], stage6_33[2], 1'b0},
      {stage6_34[1], stage6_34[2], 1'b0, 1'b0},
      {stage6_35[0], stage6_35[1], stage6_35[2]},
      {stage6_36[0]},
      {stage7_37[0],stage7_36[0],stage7_35[1],stage7_34[1],stage7_33[1]}
   );
   gpc1163_5 gpc3176 (
      {stage6_36[1], stage6_36[2], stage6_36[3]},
      {stage6_37[0], stage6_37[1], stage6_37[2], stage6_37[3], 1'b0, 1'b0},
      {stage6_38[0]},
      {1'b0},
      {stage7_39[0],stage7_38[0],stage7_37[1],stage7_36[1]}
   );
   gpc1_1 gpc3177 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc3178 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc3179 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc3180 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc3181 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc3182 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc3183 (
      {stage6_4[3]},
      {stage7_4[1]}
   );
   gpc1_1 gpc3184 (
      {stage6_5[2]},
      {stage7_5[1]}
   );
   gpc1_1 gpc3185 (
      {stage6_6[2]},
      {stage7_6[1]}
   );
   gpc1_1 gpc3186 (
      {stage6_15[3]},
      {stage7_15[1]}
   );
   gpc1_1 gpc3187 (
      {stage6_16[1]},
      {stage7_16[1]}
   );
   gpc1_1 gpc3188 (
      {stage6_19[1]},
      {stage7_19[1]}
   );
   gpc1_1 gpc3189 (
      {stage6_26[1]},
      {stage7_26[1]}
   );
endmodule

module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor_CLA256_32 compressor_CLA256_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he781779bfdca1d88d016625303c36a38afe0549b7efc33a1f9702065414655142aa1ead2fbde99db26e30c6a864c9ecc63df902d3eb37d14910a2e6d96300077eecca6d91e524b770a72b1abb6556ee285e2f2949ee42d53efc86fa8c6be1ee92eb6fbeeedb211e83e7531d83a44a8dfc686e5e43c7e494c3798ec15fb29006bbc145896a8a168e2045422f191b3b1979f6375a3b5037e0dcca6716b22ce639d4400e198758c652d890def9869546c7a716dd01b6611d303c75a9cf5fbca4076e0b4791f55d3b231412b2fdf89c5cbf9beba20a49827d1ec8453a2457ce3d1a556715da98ade2957b32187874504f8f5a9156251464181b6616c38f2ba193e2dd36759929978491b602c637111ffde5a13ee3d98ee3ef489c6c616e8eaf6f9892ab9e8d64baa9f9543cb6cd995d134af95d5596782f9847593dcc19725585a54ed2222d203202aba4a91e5ef94bf23e3f94e74ff2a55c97ff0a12f2824fffa6ac1b619216aa166c11a210deecba628bafb15130dc9b48b66cecec877cbbb801548f60a23e5edd6be9d7e6cb1ae3c6952d9a38698e64a26b763ff83abf8af3d80009278b3a29b438cc0fd229a297c7999e58ca712fb864d6946d094bc2fc7b6d41b84b36980320c8945c1f72394e0969e6e91d6e6759d762d88477b9f0bad6938b0b41a5e4d9dc462761ad5deb7fe4e3d74dbf77495f81a41d98a19a31f3414def4bbf1153c363b854dacdffa1686d55e401743045706563e7347e4468279b2516c3bddcab3c6c40666f07fdd4eef78deda9168c6801831892ce1f0a3c249621958f6e5c60a469e777ac7c72a80f240a4ad9a790d2655e71ed71985ddd6326f12a89628c8b5e09e9d3dcd1f9c270bfea749cea1cc67de8398bdb54ec1e4f4e302704ce04b5f841eeae57e919f7305390ba8651344b7016276cc0364f525fc7780a57e9e9f62e4f6a79cb56a27bd944be35972eda5225d67811185692e2c9c2cc3580cd45c1f97ff2ffdbf6eea72a8bb3555e519e5eba32e81a596b52fc55db884b0014c86c2c14fc0e522c26dc87dd7f2cb98573939ee0b285dfd5dcca41e9d6fea16f35301763f86cce4c83653735934722e5978507854df0b808bc45698ac4de7e4b9a2d37573da47239d45f1527348d93f2f8f2834927ec6d0d2113b823460af4182a84cf239da3d8d6d243c1911797dd5427f07d037474e39d66401331ba6eace0276155adfd554f63f39a0ca279b631e7f284bbd963d90ccca1d4f03232472f9a41a4c24f602da3bf771c98703421edf98e0eda516690c2941fadbdea97f9cff7fed9fc5b96ac0a29bcd62b6e04fc1b93526ad7341edc5a39637d845285820eee3eea2ce379ee4060ca51472a3d88264691649c08d0a6abb171c647dac15dc6a3d63b63c8ae35aeb93c44d89a53198e8371c7c7b2999d815b8bd93c46bdb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'had75d701ea71942e2ce9bdf7b364450c324b1a61c4bd5d443f037495d75c5b440dc1bed508a282828fedaa2c8e9bd852adc1c528e74019f364239bdb0c0e3fa68cf21d66db6ac5a3b79788ebf995f7de86547f8324323641bcf7652dad103cd56b33269000e2ceb5f59f5f850d1789c9608133d808a3cd034d597f863bb630a23b847e6c171adb9f7673a57db9c87b68983b8238ed998631051e4f44de252ca887f9169768740b02f296e3fa7f3948dd9c8de42e8338300d28c63334ca7b8660af6c9f88ed16d49b1dd1769b9e1b3ef486937dec6308b8785b57bfa0df821cd54bbb2a882b436897d4f0f58118d1a64e5eb86f2bb4977776dd2114e86163b277372effa255dc1ba126f7a901d0963272ebd84c8f6965fae39d11daf91babd98a67f10053bd9cc12a06c2d1c411f91687408f53da50b272648cfafbbc7a6d0483af7361591dc139a143ee0609318c4b729f74db74e551e56a00b78177e32951a2dfe62ede4170335cd4d1d09872d6d5481ee8f473297a04bea42b31f5817409d6717005addff74e44ad9a73d7a5016eaaa1b5a9fae6bdadc6d8f8eb9bfa9da36c83121e844bf1a8413729ab9bb4a8bfce63aff6a480d9d72a60b636972353703e70497a682b873851a808fd9d77eef946e480d6377e736d08419711e2e4d186b8589dcc7ea0d4011d02a26909506fa6f5d168c0ef43cb723a5c4144b741065c217b79f0e15b54f52bc8e4300fff4822eb4e33bc27d70139dfd09e886aff55ee6617093ff11f756159b5ca624c27e97eaf0bc0c26ea51ded4521de46e294969f5eca4ba9cee72ae77dceaea7b809fe0f59042d43a1d279301bb65fa27cd0a95174d1f17ddce752e43b83795299749fec682b18c18136d102a9f2b97d13f81afcda95dfe90de1bd7b76718c048eda0d01a783be83b19a670a3e47e2de6e14bde438cd821d0873aa596a53914785829c4e5873d1d14ac472588f566dd4cb144d59847aa5b21e56aa86c13f7bb4edaed6fc16c9aed727420440d03c0565f802ac8c17197f46e5bab692b70d74089eb6e98da18031a627ab4e8710b91fda67fcdc8aeab6e4818128e4ff1fb28a58ec4680a077c80a171b79f1c01ab49f189b07efed723d88da91ddd189774e053e637099e4a89e225ef74fae5644d9389c3c016d36825e6458863fb0bbd8acc3566438af9c2c1f5ddfe86c79c96c858c036d1e403be59c69e3e37171557b59870e8f1c13d5d351b2e15f9d0d1abb7a2403fbbc0ad98dff466091029936c29b85cd227febd1727dd230b50602e5318bc8827cd9572cec563d97b2175ae0f13bda93ddce748846523a8721ebed186ab3d5f7d566c8e2f427071195a6d2b90a8abfed7e32db1fe3b3b28ddb2668a5e2f9da5fcf49eedac2f9542f2562839eff0a91aa80892dfe626b134cba4eafcdd0fbc8f0c345e59fcf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8ebf3de4f466e574b23a185a4a378507fd8a76b2729d5af6a55d16a879d5ec95c2c1a6f7807223e6cdc9bcf49554cac01374544f5ca2782b218c6c27c02577b71055852ba884883339117dbdd17cca0d6cbb5d569e627948d826f5cc41e96bdb983b9e978cab633f6612f3b46b7d57509609bc56c8ec8942a0dd98e442047313125ad81f1ebc9f3f815b0c596c104565cb99a9477e0617fd8aaaf43b2ef7383a8aa6f5180a4238490f7221acedc9a4d986bf5e420f0f06c2ca12f9151162cccbebf8b6208e899b5e91c0fa710053093906a59fd1eb0a8a40f1d18e6f4f8f29ed0a9a55d2978c3003dfc3212ff3cd384a01dac0bcd8b4129332ed803167271746909eab119a2174afadf9c3e172678959916d4c50648e00e197f7729fb0ea637b5317f7b2147a6d0994f5e30aa38d793595603ecae34fc44d9f0df9009355f52a8de390f16fd5c5da295429bfc15b2607d5c3335eec9b46effa6925441d969d5d692cf0cd57f54c8d13ae0080e64864de11c0cfca66e8d41497c5a89e7b7367394e25c2d02d7acabe97a97ff0a6b74bcb629f758af5f4a5a1042c8bfdad2db56a03765325bb29a543830c8bb9f69092e2198766860e5bbb1b4446ea17827e9e848596e58dc085c52190b276f3db134e1b0b8f24764d81893ada24e1d49cce0b0fd0a35f137095715449c41b15331aec49bf38689fbca06cda5f97c42015dda1d4451352279ea956fb8b9748bd87a06f7c7bfd482952b5d47df158071f7849acf05f5c86dad0e59b80b5c6c3a2c9dd668efd4952645de74e32df1884ab00fd4925e1be283d02e6ff4e607b3078f177c1f45c0ecbf45d1706d41b5ece597c2921d99581076fc84e3d91245a4a48a7a91b4991046abb80ba76298457bb46d1f9791280cdeb3be4d0c74c4dcb08545149b0a0409ef5c4a698998d8adc4d003bbbb1052799fe72412ef146837aa7615aef058ed9c69b10ca27dbb669da1da1feecb9c9f81eae3f2082cde08ef9d35d296e456312bbe566ba86a42cda9469e9a06ac3913c46f5edf4a835d3d480835c60fa992ceff4cfc9501bb2a36a18cef79b78c8080a3515ef2c3866c295d1c7e8cb8b341652a1fb76d52893e369109fcf2c26fdec3aeaaa3f20180064b7c190318611cbf68b749159284612fd09b7b413edd7bacb7cfcb9b9a1389ed7a643ed9d59eb875cf61b07e83238208bedb0888f58634999aac9706961bb825178a4fc73d8d31579db10fa6d2096fa5018fb85ac35f849292c468962f39647ee894f83e9b52065c7603373e0811f5229c491bdce58b5a2be84b152fd8ea6cb047fba0eecda547f39960fc0ef0828231d802950a4dc55d6619db3c88477b5dd40cc9ec1a01071611a4dee5fe93fb3ccdb4e2e554deecc83e402ad472602dfdc9a81e9350fe6721de46333ab013984e70cdb03f8f9b92cd3c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdbfd976d112cf7558ecff0debaa0131a90c266a3a454a85741a72dcbc7299a9e3759b50e375a93ee34d6475bfebbf76de71f667d97e864795e62fff5e774af93a7c93979070a0abe02547adf64e7d382f74b9125f97962d5b1d491c9b53f86c9461e1d8b85d2315ab1404dc7a2c75795ebf6405c9ee8370eb5b8f959a24c6e655aa88160567eef5f3f413895b2f4ebd2c229e6264e5579de167de69be0dc18ac9c1c18e7d32453f2adbecb4ddb891c1673c4145b6630e0086697f89bf878dcdbfe004e983c5f5fec8750af90a2d4c1a3b363f5bf252d1f95a2d8d3d9beb36f725c476d64d6b9d57a916ede6ce96a849918e25f2803557cb34ba0631a20f279dc05e8cc21d90c1154f4f9cb5851a1660950e29e0c8951f2bc61e5d13908e0bce2907f76338cee5f798de8a5cd079f2ef84dc67b784596ebac34321a232ddaf08c01e7c6eb34eded494ce8738b0ef2fa8e15423dda633d19af50ed13d139718b255613235a2c9691eb65c9749b45070cb695ce6b39d40ee82e5eec51946c49372b9e574362f3e6de024c2c092628103a7ad7edbe7c0e5f2414c73262f17ab391c33ceee404defb60fd54e88af4e0f80de250bffc5059925211cb596d9eb377f2416a37cbed2023c38b55b726735224c60514afcbe0a7b995b08acefdb1b3f8b5232b497f8d54f0ae903f57d5be71501bd5b3ded272faa912dd1c91defcaddae7c458b1d08a90cc5c08648a80d5dc5859fb806d20cfea6adaefeb1da92fcb635610f04521e57705f3d0674c7a3934f7825d9ae37614c57827b3c66f44e39b2c1c8eaad213f99068a3fa5ec3fb9a74527252657ea1ad1780ac5323b18073f704b07decd0a317241b232630dae2bb31d936c098f1d790416c3dddbb09747137f2684816d71cccfde44d70626990cb7f8e6d1a5dcd72aca02ae8b91912f6ca0aabac948089e45247008726f21cb0b53306a477db6f0ccd1ceb0d9e24cf3bd2237fab581609193fc91507ebd5d4c2b1a0174f31f6d6fa5eed0459fe51862eb19f77c390f93348253b18faaad79ba2e12f737a50aa54ce262a20e795ca0f0f00d99af154236625227780b1fffa0c37d0e8a23ad4d1f1a0da38e1cf08096f25462aa06c1c1641f50c4c39aa2e6d63ef81d26c797882687f51d97dd6ffa6c1cceb3910a921969b3ae3372ca4b22f0d4581009cf951f3f77e441b7319293e0839f8c334ba0c33499714441cb4cd04de69799118f56f615e8897867be9bede89151b145372bc780d49c8ac9d218c59db60b783ee8b23b59ccaaf0aa334f822646b6be5e9e8f9b97cf6b214e467dfaa8354098642ff8ae13769d97d28ffadeaf1c1cfd3cb38b4e6e500cc9f3ef2d93cd664e8422a1d5d35cfb2bbe747a7df4c968022cb1d1d7b66640d49745ccbbf9af03ef45c8cf572c22e134b3649e32e1c21ff3d44f30702;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb9c2239a21e368bf5957a4d47c8b6313e5a4b8d28bd8d495ff74235e5d6868d2a8dbb022e3af94eda8a6b535a5f62f884ded74ae34e6040739d36b4f0bd0b5733aeb307e23401ac5b7aa0dfa765f33a1d63272755507af546c4677e2c36d84041e6fc7a739c70dc667ee1c455fed5e3199bf53fd196882a0d9b8f48904df0932b161f619088aca2fb1ea8ee45f4f8a38360b121ba6d70f52727812d22f15330fabf9ac189a487edfb0fa2d64eae61eb4e62063ed26133eac2e7d8a8586e631386c5fbed740adf630f7ac6eaa9e25de86418acee2e0115791eceed9cec0450a0e93e3e0f31dde0248fe761740ddb66c5a111114fc7eab820ac6424280b6b82cd7e7bd97f5d06b70171cac5b77b2f602ead42311a58b6737baab357eb14766234f9be15795f347bdca992b1be5d10b58f1fc721357951581bec00e905b7e07ed2973d448a3756b777dd1077a84097fc7b0d6ef89326b5e8e479da8362c5da675d266f2b89f2ca2b7ee8f6018faea3ec0a2ec7183161818f9462901fbebf7af223e57f603a4d397803b06d426def87e9c34ee7dadd35a606b0470f41a4bcfbf1e535fefa60e450f3f6d52459318ca8471c50018f7f643f48eaa581f3073a5e87255f599cce4e65365ef07fb2e9fe8ea46a352ec4e1497021ce4366fcb8b7a2448b1339fc1b9fd15dc4720d898f5f66a0d1f2cbbe55e735478ed7ac9e2dac8507b595ef2ad9359fa629ea26ddbef260ca1f4bef195975525e2a5a218e5f35275945e0143c68c3691ffd2cf396713faf5984e770a5095cf961a83761d1792e63b7aabba56107daf0b32125ef4323ee5d5d9fe573c9b6a2a934e3378655fac0c870b5e27b4d61f3f84a1c130dbb4fb49a70720881a78b30d90178cb9a800779334731d7e97ac8bf8c8a6423e1d3d8373553254ddea28792715192856e1b73e08de1a73523c1adec0c990d667dd7c7b9ec7a9840f27924f962cbeb8b30547ff2561a8624a22edbc495398c1c00dede25fe9c8e19557ea27b56284e58b23c612ec00be583a0ae6ba0fac7dd9b3c3bc7cc719cb62ac8da6ec8f7b251c40e5357ff02cba13609938ab58050a60658c50f4d4e6352a265e17d0bd05c6fe8f27b1009dd156da1dd9360b78b31a986348b33f6926adcda71c329c07c6550737f905196da963f4d3ec36c1108b4ee6e1c2f2850c79c20f37e6b7b2b530ca7e2430df57719a1d2cf1a00d8c9b5f93913c71fa63333f39f014a742f107867ce304b4fa2470ef6be74814c10497f4d7064ecd17223664dd75693b468a7d0103458a5fd19b3ede348cce7cf953ac954b404102f9c278ea88cac80f55a23d468b533561d2f085a18c45ea0f6e0feb872e5dd6d70093b2409a64e31292738e9b0c6e5481372e91f57a25f9cdf003ecb1559561fe324b42a6d1b4cbee89e11d92e32b047a611258cbf83c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2b82a69bd4fb5ee55109c1fff2f85c62fa4cae5c87a85f34e23d7974d6df5312193c2232c6f184ea90b09f03510502b050aeea966a6329b92a1fa4cb573dfbd24260122fbe8e9e7c0be38be2b86c66e4bcb825331052830532ea943102c13faae781eb0ea23b120169ca909749ed055a659359080c407dfc17660fd33546061cfbe2735cb95fdc30ddda3800e7da3838f1e7b24d57808c8f35d84469b3f212880a14012905107bbcd44237f6b9388af8b139b364727a4d37ed8b2d9cf2d57d057c604816f065483a4b5c5212027a4c6118ff5017e217b351325464af125b849a5c12d4dfc8eef7ca08dd79e331eff37d6e647370f42e6a6f1e512a4b6a211447499d5248f771a78e134da35cc271fe5407293c9bda5cb953ba18a63aaba7a0b54678c4d5a99e6885e71ab7740a71d6f4f080ba4c4979976f774d95c7a029603c2ba4c834c984f8a08e1a983a950e5d810c7333f1e5b9ea48885fcc53513a3a65d00f66da0b95646f77afd73ed17d9f664ec01aee5567a575262947cccf83cc6ae4579191fcc97c68a7abb437d3e7080181ec7e881aec0d6815a308a4059cc80fd6a5efc47edaae73cdaefa0133db7c429e32cb8f19e972d74e574a233ff82d58354cdc69342221978b7a36bca8b9d563a98422edaa8ec73b9e0e9d9ca215b34b6866337f8732c0a9cdbcaeeda88059cd2dbf5b246e267259f3e508cf4d6079e5d975a8bd9496793b76cd8b7b1c10b608aef523cca2cc3c6408906ddd9ad1ba0e8a4864fc74624b6f23f790c96b1e6db216c31ba62c23d6bae95ce8e306793fc0d9c9c50c1388fe868d9ebe54a68e9278a6ffe6d8186062a37b0c226c4ede1e344038920a604d86a83325052cef2350f70c7d32b73dc28eada959055ee7c04a0e3ac13ca281d4c75f9ba6a4f527ffb591914e3fd778ecaab47d49b4d60c6270e2cbfe2791342af7795b9de112d6f7fdaa7f9973e7dc05fb2405893540254b58348e314aaca3a9c60cc4e8563d60c7a46833c35d516b117d1a022c499fac4f3803f83bae4241e5741b406590e700cc341de6a9ac860eedfdf59cba4b0b6c5597bd294fdfb7d6dccd2f7623e119e16659b8e371d4e01dc02c7c7ba2dde9e063a1384d33dc2224bfd99789f38c64574a95fc4df899fc00d1f4d4282cf17b7d45405366eb149b9b45c2d8f988bf31162c8213587e8e6bca00a0da18e96883f3adfb76056026163dcc5903afbdcee80ada5a230c16c36acb2b765e408db947cdfab4341c27c8e7bcf1e65482a61e43393dc070564f84eb799b5513e18e50658a0ac6547790da1a290cc74ad3f4450e8cbbdc56d2dac0c59e9c409dfe44cff7a20e1734d9c66db421d0ad34233c575963a98f50e8777f4abf6e89aba5dfbfdee9b4c0fd8410d5504b9631089fefc41aebfa57e4811a605f84d8c30c6d1da2135865ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6dd0ba63566dd870d9d80222cd9a47b56d7b48a23d127d5ce05a89b3308cc9f4d81dd631227ef3f29bf339da96b62e1ed32f41e8f028886591eb52ded0473449432c125f0f951b88679d628a9296059bf9b30d5948f4e38ec0b447d5316cdd28971036637985181d97dd05aa683e9c6808a738bdcd96cff059127131c421bff5d5b03b7e32aad7e80cc58b5ed24ea4bcda1704add1cb2874f8152b3557af0cfdced4794965881061e3489225d80f38b0f2d720d8b9fbc5a6cd8bc9651819f4b28b5b1ca1f27407aa7f2334b438dc1de4ac9e2f62228e335874ea74397388ecff984f1f1058ed4c77e2396d37565cff7ae55523812137831ce320f1d226f6bad83826bfb7c69dec054adc493a1e78c9b350b70adabcfef54f4922e64df132e041c09c7adc4708bf09de9606237782e123221dc5c6101eadfcbaa9b5572302b98e99da046f4d4eb4d57b2ba02820bd229a639e6977d7e18dc2b11438b936bf7ddab73bfb80e5bb8cab98fbb36743e9c06171f7f9c5617807966e1fd83d21ef1fd50098f429a33b8e0ae3a0ff328d83b76c388c7cfa2c072c0945fb851d07f93dfa22f46c6be7355ff7937b34e011858a9e5954b9bc404b0a5ed695d4f63074a8f64c8f7ccfaf858bbc74933f635a8d1c9eea57f52de2e54781200ae6ea4e3431b257990c4852d9ccb23628c4caeafc4be7c92103702ac384b508e28fda3edf173b76595bf8dda8fe77e5728236b3fc025f84abe18ec6edca6b7bd61bba852f20ef2660cfcb0737b9a1f2105068f97be55f05a1521c8e4d844937c3947bac37d1c2bc4ba698475d0b99923fa127d46e565f5c78a2e07e8e5d2ddc88e4b124df6511402cc8a2c6ab959d2569ede2935eea4db9f5977630d8ad715e15b09fb7782fe9b1e5163e00428158ab89686bd226147e8d7bc09bc92fe19e003bf7bfb9690c590c194f1d7a5e2f74528378e3572b0a74cb3de3a6ced175d3b891e8089da2ba0e29faee4e041aff21c88601efb9bd32febc2df6a47db9d4ad216ce678a0ff23c106375acacad43790d71e26d191950250fb7451d6b70cd8d5cf01499903952822e8ab9e0c9e50e8340c210f8d6a8c184df1fef0f507d7bcf2a5d2c0fb05413b3b10ec1f7b567f5ead3e35d23c7d94b03759dcbb70645548f8d28e6fbbe6335384875222ab1917d8578730776c567414612bf3f4d096ca9e5bf1c34f4bfe273d443b52552fd3178819fbbcd6bde8d62ccf7eca86480e782422b9b7f027c73122782bc1ea95b06cc3ae1264a5fe6f8ce49952bbd3b3f6c9fa7a394ba9f3670855333fd402c815641754f9a42ae15efcd575f857a9a376e788240315d19bdec69ea194124551a68c02336c673818eef57229efe07d0983ec003a88323cb5db5cac19128c0bc71c32284da79fcd1c4fb7a99a817b2bebce5b1be548487d160258877f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h133d96a1ae1f791e4c66f41694d7e74d021363b15668a83effa481cc9c206c64fe4994f9effca509d22ec7eae0651d896621ab9dcd1e2ea35e0d7883299137fb5c7a58c6b7a2b3ec0e25e5d01c1637976d8ba81b517c269bdb8d8b0b1a78bac97716afeaf4695bcc7b63959d103fb4ce8bcd7213232bc5de630fbb1d5ac3710515cd764ee5d67586be206ba9a766188137cd1b70d848ecad66393cf4227b037b51e2498d68df59a90eb293922a20159527deab68749ce09bbea7ae94b1f8087724febaba05c9204db744be8524f5bfeb4af161aec2b82dc04940d4d31cacb0a96d0b2a1167a1d666ddccbdd033db849d67fec5cc4b757a45dbf1c10c3921e698fde3282ed6d54aa0c4ed4b692b58482fcd76ff6270f373d6d1d01bb48c15756098b5299effdeebdf144552672b716ff0499c60f58fedac5dead86af8268e9f82fa3953a916edebb4c413fbbbc1ab2123ebcd3b56147a9cbdcd0dea5bf27341d5b7688935936c3741fd784ff87a7d14998f6909229d6ea93ce8055a596c38ebdab6b8a2d0021db5912aadbc869b43e22029f6f35aca4c89ff3f5a61e9b5613e500ca8469d8e59f227e1e181d4e51dbce791fb203fa222e597380c6c110096e67ddf9d05acf0e97b3ebf9cdb0bc88ed139c54bc57bf48001b11696c38b7a674708c8b89a3148894644c7ab63f4e124daa4bf2bee4cc2479da5d529f730329c850a09589b2c366b2aace000ea59f5c3d1c64ddc62beb6e9d3d25552016f7095c80ebe7b860d9121ad3d67d4d4bacac1a3e9b64e2ec5c970233d0b7c51444b9f6afa634c1623d5745da0e902a3aba0a9e7cb0175f329ce10a9dd590fe6f44ebb676de7e41b569e10c87aa3737429d7712dab2a76895bd7744fc874810867e6ee2983c9a5ae42c030505377f596fefa1463c840ef976a140d4913dfc95f4fb47def65c5dc4eb516e68ca203cef70af8dec6eb44206d037371383b68280868f37791b59d61021253074b6429073cc63930339fa334f91be56edc014b5853ee09dbb487cf7b411f530f2c393c9ffdda97861e685cb1e3e7c79805e893d311468cfc33696e822b5a49f72c4a03f841a89346139ac8e17481983823ad64ed8a1253d10896e811b0825ce4b49a370abf581df581e6d5849d572a4574604387362f4f517edd163018978dfc04bb375b3846e39abd418be4cd79df8d8c37a968d9cfd9d0076a5c93ffb9b125499fbe5547f7fac983f56ff7d8c13d4c951073394857292962e3fce8aaff58461c7dd8603cf891d94303d1dac56f58eafbc0dece87e54b5b79bbff5858786161ff3ececca7e1c420b6cbddc375b63bc9cb1e37be11974b8c3bc42c0b7f128e769034d15f5ba428587937e04a41332edefe4dbec33cc857ec092c1e8bef730725e5ed850b3ec799240e5fee10bd99ad092535bead4c141460bfa6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3f138c0acc5930157cfecff1c2e229da0b7537bfcb3c2703321aaad7ae8139719c806bb36b32d5ce95d7bc8ac92cc7f286566cc05799f343e3941ee87de7af5e4fcc0660fe11673fc8b87977843628942d8eacd3e866cfa19b1c6a727d68a50a02de397b326e2f3af7ae3649d7c06575b893be82d384b1e210873e41ab9f40c6ab2a51def3ed5bfa48485406b1a752a9fe8342cc5d10729ad49762c9688e1c7bc64e31eb910fa6b2a8f3f8101094f1d49ce8f6c6b4746c7bd53297755e3549d0a5f22fe8d99578ab2ef3b0e6444df2a7d019d4cad9877079c419191834d65cfa7b54f49bd8805fa9f2b44ab2eaa0ccf6aa847f678f23d370fd26dfddb5d319dd98b5780887ba5ff5ca891b2803720fe380550c88c8e05b91971dc86f40714e0473c5faaa5f861900059d058a7b66b5f2a295d7157540b8dc294c8f424b3af4b9c81fc98f6851845f6d3dd52bbd3734ae8a13eb26462b9bbf59a00e983256fb9747f4f2c1a420400a0b485b78933ae237e566f510abe4762946de986a20a8f1b5a32f8f006ca14c8f38e2cf31121f8925823398d9d2a227012ae7bb1192c947426f8cd979572fb60e536c7fce64b8be3221714962df5f0ccd00029a8dd72fc60f4d5fdccb73a23697bc0cf3305eee69175d281b7005e5e828d45b31c030bf46ffeb5700b2614bab1bfe43ecb757e64476fd85362795e5bce7c270dc0c3c8fcfc371ead6883b7faab897d873ecfb3f417325e96cda517c3bbbcfa9cc2764f5d37152052443cf93c724af4701dfbd87d16662fa06005be3c35502150a901aafe867081f3f2dbedb9e14926f8dc5cc6f71d63355f2318f132f68a16d49a7015485faaaba246b46c7367c8467e907f6de82b71bf8334ef828f7671ca7e4143d4f2d7bbf1d6a97a59760e3a51dbd1e6ef5dcfceb82bf577b81b443a624df651fa810045eb3c7922c7235de42d9178ad2a49afb59b5c3501cee097263b1f38aeb075e2f4b1ac4a2fb70e005b81f38f1c824e7f29b81cb1fbae37e77f5dbf318d7b1a1f5308cde2ef1256424a0adc5166d7e051f60b0416f671c3807d0479f395caaa01563c3149365b3a91f7c27c7a9d63f897d5c0c72fb5502e6f57f5a5a494b6e5b8418d5b932d1dfaa950b3726a6aaa5d50104cd14215753a9b125b0c663ffd8c1e7da0ec90a0a4c690f635eba6a5a90604f69235c9ad13cc56fe94d67cb1896104f658ed929a301de2d7455bf9e70b6f8ec29f1306fdb4f516cf4aa51a1c83b5ad9226efd59d29f19e4fc72a19417e3479641e40a970dd7efaf6ec0b5eb55c321c92a1d5f9939771424acccfdea2bc460ffe0f28ffa4648d86ae0d6ecadfc5b10a539b41f050eb9d492a8f06edddcc0f10fa49bcf59bfd89c49480d802685343a9b403b8de8106b5981160d38a10c337ba415d59607ab954ca700b4a2c3173061d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6cc57c892f1c5bfc85ca583eb2fe20f536ad4b9545f38498b8daabd1535139dd69b576010f61b6562e3f61d48929021eb7df6600f83674c4f215700f027fa3b0b74cb7251b8b4e72cf51619e11b2a567098b26fe77983790cdaa0f103c4f1fa247002909cab67c9dcaac87965e2f32695094141d7c0f3aa410987348a9c678a40c06d5aa57e423a992e3ff73f97ed886d1b704219c1165eb86a220fee72feb4bfbe60591a423ecac4d6c526800137584147729bb3d1acb26c9ad613b75bd57ff1fe55cd48d59cfb9447bb554a44fb759366326570f5b65ce98849eebbf0bc5f3b1b248efed3d3285a5ae6b65dee35cf3338dd6d502226df17e5d6dc188458c3ce98201fe3c02e2d916f09ab426dd9a17b0a6cb1ba51ec21fe794613381980a30d6e93cbafdfc5216ecd4ddc381c50f32d69f40f22e8dcc0fd2353d0db17d709b6abd3bb1c84da0a4847ce94d6c78c5642407cca2eda1a1427fcec93a292aeceab02c37c208456e6a445511894d5b281e5c8b30897442917528296e539e460dc141284a8cf0ebee25b76803e8c14acc8bcc5125e790e19935df849df95d90eaed87ffb70202f18807f99a55252d946abaa460fadb90ac6eb814ea24741209a95720c0c612feace1c3eb7ec5273c4a9a9d73805aeabd1e0939fab437fe38f2b64298a7c6e15eebd92088649d1b8e910da0bbd6d6986e055f71f3af84be650fb1ca6ba8a4d86f797b175978ec3ee3f4f5bf53e99eb5042c54fc442c71371a5c42ceffcdba4f5aedc5784473b2781e85055bacf7aa27137bcd97e796bdee1365cc772f782ed4d1fb5e8d5581235512dbe7cdcedea0ec71b6faa2d63543f89791744b4a6440bc2b3130c35f89b0b0a9172ff0bc6eca7995109721572a008767f77d7840753d510c7e927874e6c043aa6336a4721cf75037cc9da8c4de238d29448813140095175331c284bda8162ea30c5cb132d628fab7aa54f29df8c0ca36239b60dc2d9b4c2713880245f5a7949b7a217659b0fd3a91c65a1abf08e1c20fc78926159700751c2d766257a250441273a0452f7971d3ce997c85c09f6e6457f2792f330a04d41e9b3d5ff0f5dd29a854c0a80d7635dee98d047f0edc3453cb46aafc30de535a9df84ad7ce76effb37de40cf934f075098d50e985fa9c287a0537a844ae5d7df216fb584a7be7a89f0d6a7b86f60d3a9025ab68a127426d9967f9d6056cfed2eba57aa7928357e80fb19707fb0dd9c9c579c0082c5f6905c5abed79aec20a6c8e18a38172ed4a87f78a4a09cc701f8b4f54b19b59f497c1fcfab5d2b8f93f4d936914b5c011cf29af7fe0432a9b12809facec58096ce745d32caeea163f6d2679188d4a62a69a9dfe676df6ddb22f959a60976f14c1e3ebc05c5ce1e85bff1dd9d9ac9c2969befc7f512be36b3ee192471e55d625eca4ff84b420dc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd7dcdf94f600c7eb88f1d1f5e4b0259cfee4f6cee21ff66c6362275c38eca4d49750dab320561922b661f4677f8f95510932fe7ce98eeb93497fb5a68f7c721ea8675ac615467cce101c34ec5c71206d89c178de8c7fad8eb2e6315a39566dfdff05b5a6eb8a0d6e90d1e055570eef1eae2f89e2c70762a79b97610b0b8d578ff2b01d6e205a622fa67980c9667198751e436d64fb5cc9afa81eed49ceb5371f00a7e87cf93d408292f2831916f3e141156caf3aa3e4414a679217f4b1f665e3bb8924b1762b3a5b5cc0ddfebbad0f3f09af61cfe29f0aadd3dbdf3336762d2ef93bdc1e103b9d3f3e871ae0c5c45dff7c00d90b212fafa69bc7b4eedc86c7d1160a706c22ea73e2f6899ec115b6fbbd692663b236aea46d1bb1ae339e753fdfdad976c94bbff1925b2bcae0d225cc8f47be522364d3f838e980891d2ac6e752b5628449dd3c0985f7a4f4c6fa34af79b7c83e08d5a3bff11e128254f5810412014f0009745c3b86f3b0dae09ed34f3ba8f2cbfe8f4fe868f2e9e2e6d38d2336b9b3628140d1c66337555454c60921885ccf19691ae8638babd09900a7118fae40cd20f78744ea2ee27d1f2383acaefe7638a811540098a51835d1e74c1ff778a53d68e73e674dd8e36b483335403df8f35add4bd9f6ea04b1c7a663dfcdc1f93bc8490b26ec074e8de641bc4f5a71402b1914502708942d933ed49f91d693c3128d0acb8d6850e00f130bb7353e302295ec9e7ffa9e3c6eff14f262370c4c76e322331c3bf0b69ab1d38e0d27fbc3e1c97dc767bb2dbd80d9f48dcfb74f5e23e01a9d207fc12057cd0af54b26b6fb16a27b44e36886431ebe1996a942588a3d4209b8f8e9a1bac398f86c72e161e180c00e7f965ff34d3d0a8c2daea3fb7eab8a4b5e510421365814ad686b232eacefba31d5f01db536e0e397ecb551cf527597b76c185032002addd1483d3ee18fd9b9d512d1d96d722c6455514e12b59215e38e3a4ca0f63c4ebc80ec0278f365a382a0fb1ec56fb334d4ca94547540a83feac4af1c1e6d9008801bc2dba9d38f3dd016e83df0f48580eb2222dba3289f15c797f961e19f88216fa6582b81d12a41149231d40ced179e339715dfce1a7914e83a17659d5bf428220a680b2dafde1de129bb598cce1416c3ad572a8736cea4054139932df00dc192394fdb38103732e751718696d4b4afcaa9c3ff93dcea885ca7c18b4839ca434df5f7a46abffe80fb11a76a5804b0ab2de59859a245fa748bb95022ffe5e682acec3b70246aacb4c3599af6db8b8463e0ec4c2dc1165d94a8b57a1a977480bfa4a13ad39099e2c3eef90704358efebb03bc5495e36efa386630c9c703955449a180f1bf06c65bebb12b8d2b845e7bfbef16c39c478a3b5fac9bb6c1e3e037d58d3e2330acdcf3aac8eb039fc2a0713f17061d82bef33947;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf2d62c92831d1bba94534bb1b86596ddb5a83fd29c2545c227a03e25e1342097f67e4d95b567c2267d4c2517125cae430512d7839ebfb9cd379557ce3178a161fd77605c102883cae2d15be1f5eeb53940b41787d0c6d7c6a3e4375522e34810912389728dce494dcee606b3ba15573ed7d17bf56ed3606b5aa5ff5e58d2f6fc2b2c079f3e0cf3546da7c32e93c23fea4bfae2fa84ffdb58c2458556da58ae122a843f01e3230080d18b53d363a2b7e442d73945210abb447a2393feb6fa4d044a7044a2f09a455094867fbc5fa3bb61b57d53f7bdbfa414e20b81fbd39a4bfaf50c0d95701106679b92b79dddc28893d5c7526e95af65067123df5891c602fb230823107451275a046dc32d2e0c78ac62397df58bde056e4183abb458c2370c8992aaa5de41e92a2b0d00bad6e09f701af101b0a366e9a522c047a941c6b7d3daea9890e629d9ad0034c68fe8e93ae30eebc37fbf7c2c9cd65b1234bb3b632c5cb8ffbc033ca6353fd5816760ca2c8528749509c1787ea2c82d2d98141b83adf61e63964d8793692cee98c74a570605b0d9599ad275e1d500843799d00e57cf3d6540c787352197d7bb2659930d87a5674b81636523a9e6ccbe4e713eb83f36777f454179b3720b6b0caf91e7e4b2639a718c07748b03d22563658a02f3efca82f6f4e628ca7ce87036d41f1e52a0212acb3d92855a98f2464d2d2f0511dc9d32f4234d564b2ecf0eeb087dc07e13ccb9443f63c25a977d95b6336b51a0cf2e95e4058a01d3defd07b089bfa60d16c76332782e43bc3d2a7ac5aafb5cc7b5cc2f63e2b36a3a5f8d356cada37bf07ee65126eda0367f9b06ce3de0764c8effeb3c299852c88ccf0e8cab48ab0e33e51661c10f0d9db79dcdce18aeaf72a90472df891fbb474835be42e150ab4daf3ca84fd005d2016f298074335ef52e22bc1ed3dbe0342545dec6b8a214c2615392207d6ce53221d70a0552c060a20b77372219ef155199a9e6808a76757652f67cfde2aa58d24bcd5c6aa3dd61e1ad734d7f34380a2e5d36bdce14474c0240d76b8ec86eef0d3424b2313531613f6d0f30ec05f9105d945ee3d105cc0d3c2e3c22ff4eca3a72f0d51fd0ca7d2f977de46e1dd41e66d0026bf141a21309da18f8e9986200ab9b9b24b524fff04355050a817f91ed920d4f8b245c7fc3cf2092567bf44f1d48c6d30ebe1ecdc768fec444cec1b616769f998604a0c064fdf5059a75024a73fdbf4d8feecc5a4c99353540c31d71b26eed178b2ff470a415316f0a6c9e8c1c7791ba4d4d74582f294c78bc91052ed9f4893657096ddc28c1e112fcdd7e8502b8b23f2c083e34a9934cc18884f1b476b26a08f3c8480f5209d6ce95d8d05d0760e42da239c29e45255b3d6d00462697835ba0cfd74c6656ce5bfd8a645538c7e3986e4f7d86199b94ff5b202829;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he1f0fb6b1796ba22cdf8e57125f07dac6a6e8025018e9a09bf9d525f259c55e6f60f7e152ccecab8d56c4aa78f75392b0f1b7199151ad62630658af82505e1fc2d225302e79f93f13330f09fa76317d04ee227675395663cd5ed3b80b588cc8e036f478e98a2a951263460156d4131c7e1117a2d07aa4ed0fbd2f41559e95ae325f36609f4c0f770d1e2f8b6a994d256b7ddaf3fbf17101d6cb032430139561bf68bb79de7ea2d8637f33b7db6abb51bef97d4e8482a36fcc12a0bb98efc81ac343a468e2cbf451afa41bb986c79c13deb625998aef47b186909fdd705a4d2992b4569a9fb90f6420c420e7716734cd9271c911336b653431785291a0a2741a033b6da11380d478927bfd878a939b9a9c73ba990f7365cfdeaf744d0d18962ac152dc49b72696d80778db9ebe2ce00e7fca4914a1e770990fc1ed721a35e7da4cd680ce53823aeef0273fd714d900feb7589d69861dd0035b1502fae45217ebca5406ddf07e25619dad622623468507f42947570a680da8b0de6adb5b4004d6bec81130e9f003d6407fb3e1600c8499bea0bc4dc80428b27b8c03a4c197c29f35b4c86cc5e7412712a88cbcedffa1127a2d315288587feaa64f82e07f245682c90598a554f5521a9cef301a50f7b077ecb45b3e64e273d6ff89c3647d247079b902fd9269efe7360ce3ad84d1c92ea0279cd384657d3a2c88e4fe4f72841c30426bf5adfc313b6a86379d45b40ed412bdd3d2b421d771f1e17bbf5339739b348f0a07bc3155d2e121e7a49f55009a7f1337c1523fa8dac3f25cc8f6a483c7aa3500e609eee7472e26426d288bf36edc8a4fe46cc1f0b2ac5a3eea64944a6141a9569af290b931d2478cd533d309ab397776d295fb2ca0ab4885ae399182dfbb3ecd89ceb34bffce358beb60199b625afce8759f7da8bed0f83c210441280e718f18bee8d75253e6aa1acc573ad999c1a21103088575ea9804d179bb8d57d5f26a3d88cf1edb37304bfc6d7fa880888cccc3ff58d6db03a735ef8b05240c9800c91a2a9b796ebdadecae24d0116133d89f9872ae456237499cf97fceffe494ee6b26bf9dfd1c548c6e4dc54baf0a94f42e22998d2ec1f60b737ed0b42d3b27f69c00438a3b91c9cf08bab207f9bb47c6ace6d6f867b1451f3a369fdb92ccf9262cf338ac2c3cbffb16243079539cdc4ccf6e0072ec141752a1e20b68cc7ce17fd62150c6dde4d81c64ab7ce3b77fafb988b97105ae9c31785e720f0477ff56266d97d2bcfc307473856472803bbbb8fe4136c8b95974326eee158ff0e73c6ae4e41d282f26cb7c8b3cd7309a9c8f88326e14be87801dbcf3cf1373431167ee1c17d8aec7e12056881c1eeb843eb1e1edb18a3aa94324643ffaa1787060189f934b6300d98e1b211397c469f47875c2f1705400949491b33fd8eed2cc326c77a6f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9f6a8e71bfd86f417ea19ef98bf199914fea9dc1414f5bd30cef7d346bd54288c375c67678c88944045b3dadfd0ea706499f716b25244b7c0a557b72f5b854547403009e2a45acca7b1f97a8e5727c8042306f68d1201587e6111963a8977480925e382ff93363aa05ad9e04dfca378bd523957010a145cf3ddcc92875593d24a1626ac5ffd9302c918c424b7fa7742ab82bcd31712ba17d69b4ee5e39dd19a77079102e7bc4de44e22cc906301578206de8a0aa94a92d51128c4b3bfe99b1a511f04180aaab9bc948fa4475408d1d680d8d1aa5f71dd0772092c2c46e2db204b918ffb8aa6bf2cb7f1ed7225f3116ea255479725dec29927cc15083c9518be89171c1b0012b528879e6126d417e7e7048048d43fb0aee565eb4278d17619696eaceb2b01237aed697543c7baf8abc31fea8b003cafeb67204862e321b7e151db5cfc693f5ff87c062bd5291cb1a246f9d1821517230f17550e3755dd8182e452afd27d28c00d80521f9950a298e7838e950181b94c467b8909e5dbdc285832fb9c6cdd6b7b61f685e262b4cd66b8a6abd0db3ed0b8cd715eab871827bd5977bfb2c12f0ce6fc46743a8ef8c77c20af6528b8ab52a364a2719f74d06c3011fc441b6c06c5311e767e4621ce855859ca6f42e7b1b6b2bcf3f42b20da0ebe4ceded5ab360af2f552431d1d1cef94b7c982cc2b4e91768a8e22dbf68649aa9a51bc8cc6cd0dc678e66db2432d6e9a433a973ba9908c00b6f9375f6f36b0daad38541ab1ce9b2d2503c28f9585cd03dc0f42e3e48e348603803a75247e29c2db513bc7ad411238aab28bf23f491e267dfe9402f5dfc1da31eaf87f005f2302211fbf9bea0b5ee3c31c9a1e8481d66324a9f2c39c4ffea9abd04f7a402e3f406bcb028e86c46953ab3dc1934a3da0b2087adf2609a2a7fc128a62fbf179f2e5403a6604de579a32db35db68606346b486a085dc59e48c3ef49fcf4518a741c313aee3817f8fe8fe7949a5191306a15970502f2379b95b63b22e3abbbade95982aa951c78dabce7da5c0aa09e05e373a67bb086d06b04f5d36cb6f5a69967cb917bebb4357ce9e42bb3105d9842042f6a3d45a356c784fd2d63697ed4beb000f3a1577968c0a3bfaa00691f82252a6069fd913977178424d157a65ad1014125fef1e1d440477d20a77a0bac066127284b59a17fc25bda4a529b93210ba1fca5ff133e1dfa325744888fcbe79863c48b5a94904a50936f93c1c04f61ab8f6954c6396eb42786296f6f7b3a3812b89d7dd1054d5361c4faaa25bafec0387025e28935d8b6c2b5ebe2353313d94a349c6f06e153e66994adcf85ce696e54892a2599d4832c3ad28ba70ab83ef4c84352223ce68b72698c7c6e3618529e79eee8d2c5433a2bb2e68c3f7ff4e0cd15972e386dea3a5e3b09333fe3ed6268616bbc6313a34b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6c0b72ff51fc59729c58f9335a96e03f636bdfb0365d0fbdff3ed75ed93831ee6124004f2fd8a58d5c619e10bb638423f798cd9c1b6b6612fc52dc266ad345ad13f7e7ecc714b7411a80f4e5527e21d34dce696ed04a83235e7deb5e3917e73847e2ff64da369025152d4c870b025e3c2f7b72fef1664cc73b4cbe062dccb0b6a09c1934d8dfd299e8b2e7b8380de44b9bdd949ba5862996f6d4057e9f1813105cfaafc36266d28323fd499eed4b9c488f78142c08f978536bc62218d975e5753d4c990402d8d1c7e9155cab8039761c2a4658f36899e7ef5780b419534667b15f8ed9623ddfa8004e9f7094e1f5eb920bbefa8cf3645b46e104090d1b9f8085f24ac2453e65d21122a963eb986a35d1545f2f48b4e66441f645922984dd2484a13052ce1f1dd9fbd089dd12d3f035be539ba6d1a5f4156da08342b8ecded40a23b9a1e625ad3637880a2a5bf5de0f64eeb93b0363aeaa2308b9b11630c5b28ddf530a12d91ab605b4f55abc52f030e06cbd58b6c5aa27fc5d7a795121752bea333f388ea0e6bba1d110fc323309a561fe8e52d526ba7b62b8ebc3fe378c0649a32c792441b65202b38a85028f8007ce08efafae13396fdbbd5ccc8abfce3048138f28cf6e1e0bd7e92ab7fddfce34767c01e94f3d9e6beb702ff68254cefbf5098a0e69384179214d30f8dbefa967c890fb3abbd11d93e095e33f09eeaba9daf62aaa8c83cd50304aed38b919fa7effdd11a72dc1774963f77c487a2212782e30912c386191a3b6b3509eaa9fbe1ae111b8eb2cd95f60de9cb2c691dade0d7537ed50b700edf4e72f98b085014fbf9f3be431d716ff438f1af99b9b5c028cbcd54c27a79b9dbed7f71d07ae104e9ce602f5d403dbd2075c67f8386655a36e6d29911a073eeb8aa57abff6fd1cdb449a168576d41b75d8d77c975e305632010dadee02917c94b344f7bb9dc2d516cfee0d00da2f22f187580cf1718da8f494889abbd3d53ae840e680b6ed1827b4113729e6124bf34bb33addf07c0d0760ec706de045edc1b979fe28416323d365c353e4ace498ad88c0ce0f4e1115dcc522271ba9064cf20caff954cd35cfc9995c879703b27050d32e09980489c4cc08fd97470432338a6abcdd5edfd2b70894994301efb38dc46db2aab8b997a2147befd7819236bab1b8110999afb70a6a96ce978d9f60206673cc5e59ef031df1250f9525648c083bcd4e5613c07ad12077785e2cb2ec94fc7bc534ae98ed5d2f8329c22f77ab89b1e5da78b7a4b39f120f6f87b173235e9ed5287928d5e85692f4a76e6bc32c8dab73d9f3e267e1473f260eaae597beaa1b5adc3e6e3030227857d3ac7be7ed31ee07524063bcd9b8dc427c92473db1947e47ba369703cf65f733b6a3f90b92f917c630ba4609a179f87173f1f9d0099bdcdae5fe9369f5e806976e2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd48eee95f4a3f0fa3717c3b0b24e7c61e455ff513ee0c58f5c5ead398787661acfe7a53df5616b778b5439123d8b1527df08590c85aeb09ce1ca320b8e580773d8105839e443ca7ecebbfec51eb5deac78da7ac95af393430f1d30d902456d9980e8064af6adcd631900c0f5977c99e5a50453769f0c84bcfca10955898c444181ab137571c8aed0320e36d91b7827b42767b550f93facc5e7a94dd81953ca010d9ab4d4a9380ee15d71754c5b2fb3fe4ec85f5527be035328e0ea6d9dceb3f15f6236adca0c6bacf4de042c91653d95b7216484d74aa197b743b66e4092378cfcd790c2d3460ff1301e4b2db2fb10a6a2d9ae1f9a3ec824c4c0dd281bf498cd23368e8e8677fdbffa76b560ffe991380ac8f3dcd309ea8b80e8907e14cbe82b84694d25bed2055eb9b3e792c0c953845d943f7295113d23764d04fe32728f62debde4ca55486b4928756757c47e8744f3d6a23444394e8051947beb6eb200e8aab9d41a73bd3c19d8fd81c85143516124a0582e965a3ec318a33ef3b2dcd4584ae63b3513a98e72dc4191411906ab5688f4d48723630cb369b3370b3063aebcf390ec2a41e5cb7a3762da4a5076c56c8c00ae6a41a2a266c3419b279d0377c52bd90079b7995591ed34c69751d43c2202579bef648c7e9dfef7fb52882577ce0a305dd83de8834d90d97cdab8d26e62c71a1a7a9c78631cd0caf992af66c18bd2c8b3ddc2c6219cc4fc40fc972f8f8c3a296c72601e4a28fc58675f15fd441e13c131746b706b694a29926d8367e1c4dc8c0df7fc07b18fb9b820a931ee1f141307426d23f4aebb42afb394a0cb0817c580e6c217eafbd1652e17f8d5ce18974179e6b18334e7428caaeb10229ee2779569bba5004f6c8b9d9648264aea23da24c18fc876d1542abccc05dee79f43c8d8c8cafe6769f0b3883b8d1284e48ec11b3502b13206e77891cfa1d1ba2c819df487931d3140ed285ea75f8b24c6185c6edd164610483bf76724b5d5cbcfa2b22b29b7aaac3fcc89ea01e3af9146c9796992b56ddd2abc3a727108f7184a12faf0933b5054c27cdb2883089a667233e27cb61a6d1ba101e3f4736785797c9a53681d650acbfb88bbf25306648c0ad04c95cd275579a8849f19b381178631246556ebf43310c072b105e479f2e59548ed32aef768fba88ac43ed5a384cd68a7ad2f94c214e44f7f857924bb7c586917a8f6de5d8c5d589afce7ecd6a751887499b7af66bf8c2629ba1acf5d46f019c11d6464b77d8cfe4d007291104e42c092c04e825d39165737502c078b6df9dde92416b760199d3b1bcb7f35a8bf5fedba96613a229802e2e64e18558752b7acf84b5ee11b0b10396390e9182aec8c3c45a782a706639e726ebda37050326727da3617bf97e9094819ef80c4f299f3c6cecf00d237a3d3640d00148164ae3373aa2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc5da5991f1c04b9302cefc22742637cd19657055bbe2cf41ca25eb43f450cd3f38ad6dbe8ff863d6be8804ae1c59a939a751d1ceb3d5aeb0f1fcd831f353df06f49f73b60dbb7b01cd0832820c837af93a52a33b56788f155022865e7b1e2c4727b7fc712f64aabfa30b0d61100f4a2480b5d6039fc769cad516093c60ba7f464b057b70059aeef71f6f211573530ab201d332d0553cc49af55a2f5d275c66c3ec8725f337067961ba64b3c6148ee31b44425d1e6b2e14dae1816e228017c58801065bbc01e12b04adc0fa172e407943c840548ef642e9e2ce5f330b8edc009141d006bb9d25556d98858464124130ec95115a9655544cf73d5e1c69dc8ae3bf95cd7ed2d6355db5a1f2a7151953eef8b2b09b1c98b9fa897743c9247386d70ddba6a435b26cdd65638a5e82901364270be065221f32b075606ee63a36da2cd3d6ac6ec68b7183b5ab8a9bb86971d31d799e9dcf781e14a13d4b0ba34ab8cbd8a897fdf491e91f10f222eb4bec098e0a7a297903ef688232999cf6baaa370202584cbb05fb0699b777730c4234b98fb369c330a20917b02c63b7310825b10f9e1483912e0ee4b4335c081cb76c0e5c42151cae743fb8c0e28e922a1b0dfb13e6beec7887696cdb441792a0ca0697346eed3006b92eb9fc6cd9b5679a2a603acb510105f73a6d3863c07dacae278d8264ce8c072b0cb479f96727a3e82c17154ea372d065b1fadce1a93d9e6e49200f7e4ea104b65295a62e0fecad085685c71f0e784d084a061fc5d5a7b1df8b1fa22f4ad198f482b0d910834e669da65988a7dca8f90256908f81abe6c860cce4f3f7d142d7fd061768df0af574231980bf8bddff5b90012eaf5a7f211d97aa9beb13635c84a0469dd75e4f6dc7e94f699a3ca980b3638c3f57dbf94e2e652c4253c694b4c20afb86b94ca38dc95da782cfcea2c4f14b15940b8ee44cf7129c9c143ca40f9c92b33475a4fb587f683c8d0edd02d67f3ec38b02af9b87874c077c0c164e8bac1b4127b444c982fdacaaf38b1905eca77fd91c3c3ef70b2a063c1c53a88390720b593708293753a2f35cfb6d8e5953c03858aa792c3f6b7fd1b6bc24b81c46890409bbba6a65d4554d8063f704f1155b7915aa32eeafbb4ef4de030cb7df614634dbbf0a17b7d4e62d090f5d48d8dc17ee936232dd1ac71a3e6f8c73d3c35bf7c05552b61882bbe858e2855f5f769cafea6f69184527e4552d55f204f426fffedaa4fb943a2df590c3229b06e2c8fc69488effba100969da03c9c9e058ea9e7c54b70f80e1fcc3cb59dd4eaaafe704937340f58a513ad67c208bd42ccb013b2ff164dd5f609f1463e2fe52857d9de9f26d00837fbb15812ab7a5308e58dfe07d18c40c65bda8ae0e8f85dfda8d0aaa078b819b7e1d590fe7c03d808889f9dc392754e2a6d049845070df0ac5fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1fc39eaadae9919c4b303a229971590e3d43c6fb572994e1bd4688ba8a285a2db2212c8e854ae82c903d5227497179f3733a218ad54c2dcba84bef96c384f416fa468f953b5a50ab395d086a73022230da476d9f80282c479df3daddf3a6d3ffc61d75b094709c6caf41a41bd59e91dd7173fa019132cab5f60606ec0b188ed6f0a56dd113174fc747d9e8767666f0252b36cb6a128514ca8779072e58d204808ea9c35904116f9c21dd4b5570008fd81c90443aae4e901c90a25d7136130dd27437760183cfb6e42756f499b303ed05f49e3934398ce879a7b1c0304cf69c588068a023256f20fb8ed0d753d1b9d9a510abf408d2d0251fcdeb99dd34f4094217ccd53d11b6d3d44a08d9dd11dca72e4cb783c77f8463c2910306e8d7c632eea19032f9d8ad662bbcee6feea9517183f734741927b7d8fa1dec3fbf19e63c57bd5e561a5bb8d2088772057727ee1a451c8623a8581d1368ac1414281682958d48e8231291b022bca87da5363e2220d3116177dc81543bf97d9f85fc4cb4bad039397b23e11c044277729e00c36e94ae064240cb620a73a0cc234029d1ec0f3f664a9efd3b0a271f0a5397034f4de06c8cddf67b1fd5121f83258e465ccaff8f95d581a71975bbb369b90c32cc41eac2a2731b0284926b48d1107d6ecfb22b459021957825b4af7b77fcf58ead984cc43b86a0eea7bcac5cdac89f5930025f23e6db61909c4cb1825ca67635f1a055ccd3f1c3b73445e0a1ff6397e64b555c7a131381a08c9081c863a474fe7444fb3963570fc3ddef3c40da17224f3d289327218a77efadd1b934417ecd97edf07bdcca06c40b58967536bdc6a85a57ae9fbf30fa61ac4320e63aff61eda4d2fbeb565e82ded2ef47eb92cbc9feaadc65e3f56779399a4eff2e4256c2d536c353b4714f89cd7bc3f5181133d3afe0760b4f8f2d4a26f0e68336df2ea3a10a671b2da3f565e85d3bda8f0d49ccff361c0370ac357e5d090d38763f31d1e1c161347f1b19d64d22a6bcf0a924be67919fb5c6eeb6c075c4ef7fdf3fe38e0181ad69a1ddae159e04ecf9653d61fbd169b6b7cb4d4513590eb8dede76779225b18978c6746957c5ce7ed1c4ccd3def043c676bd68bf0345bb79bbc01c8c9e64b6a5cfb44374aeb39d8b5de23522f13d8c78c701b3187c477077405492b75a6ce0ffb167f48c0cf8e6cf388d1d6eba73eb2a24081b58b35767b7fef9cf4b12717a03631590789564607fd2fbf6cd684511f23c74a917ae27b4d021f6cbc2cb74429a61f7c4c498dcac91b84a25d4f49b1f8278bf103e435efe7224ec0d0ab8167b9c70caa1294ccd48b6ef6657e54786d8de6321c9adc934b4e8aac77985af9da5056caab94e4be753bff64c2617c54c7c55c591ad415936d9cf3f4cbb933ce6040d6095366d33f3a32bb365796227d78578e54e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbccaae44ac2037e7d4d60fdde01b8cb242c571b5c71933fdca9892bbadf043d22776e1b6c336bb18d495e7f89938787bd81579f1d0d45d63f9e59860b1aa67cb4568b224bb6f295ef91f0e66f7c4ed77c438cec9e133eb7373266c62f9e6dc285f97f2be96ac9d3a5303fc8547403ba1f0b624245697e86aa6743d3551e4732bafec08abd87ece040ec4bbf3f183322f35af0747595a199921197da105f378340349d2d4e980ae15b12e52e3165043aa96a58639e66a0c739c7cf99500fb176bdecf34ec7f6d27e4bddc32fdcfb0a36942fa694708cf8810493836af82e3e435c5be1305784d904e9b2f56394da8fcb1345fb05d8e220940f187d97a7cb2f11494edf25769a721ed4c1743291bb900edf2b4fbed56c7950c6076d0b6b115587990a8e617df4a3c09c0a658c30dac4798ee9a154feaca211cc4a1bd46508dd9f51cfa3b9141f5637b120db4d31c17fe1bb362b50f56bae59df707f489545d5c8e4f0438c4cae78a790e19d343cdb2ece8b025052879469c1be5aa0c3d8b82ba6df8c900fb8b6e184bd586bb2ac52dfb6c72300ce483fcef09b95efaaf22458ad35e590a74240ffd4514cb5699579bf1d80998f8ac84dcb0b6f29caff7d16d12e763a185207d44977cb1991945f72748ad6a7dfc7a316d087c0d8580af97a8123e877582771c23ff8908b9ffa127c901912a80033fba82bd7cd736a8047ef4df2b1c5cb1c12a6a3e47dfcf6ed29eb922579ee23ece1a26f65f8ad9a04a99fd78db6c59ccd9038d3dc3817b993eaeafe96ce439cc1ba49b27ac1c957adc0ee2c687b97292cda19dedfbd85f79b1a582ace2a80e08586dc5a1d872faba2e6a413bd14c079f913e2f1bb719e606699ffdd3f25193830413927294468a0590681253bfde851b1dd0f127e5de5cb9b502dff7334fc208aea49f5155710af6dae148e71440f098322c06ea58d2b04fb93fb13f27eb5bdb0bfe451da0dcd9f7e49afcfb03fda98d797f5d916371470a2a23419334cca7bb27636cfe33b824c3c47d52ffb2b072b097d57f45785f115c521e08809c8ec52052bd021db85228497354006a7ebf4d1f98aa98aa83d91b58b7c071da3c3296fdf0b13b8041134f13f8a3691cf090e5ec867608e3d74cab8780307cd61033c1df78f58902d05ce6aa9c66567399a61353c9cf239ce4a7882c2c2f353b05896125008aacb9df749be066273215c3902c4b2bc64a05c2b0194215800994fba9374bf448548f8bbe1d849fb54e84413406e5f921d78f7a35801bc7afb25955a119a8ff519f82c3a1e72f1a921e40cce73120e07f3375f456d8ebebaef59dfe00997ec815f1fb4843d58bdb811fc8cf34eca67522ffffec744bb9bec31d9bd3804ed2c6e4c6b6f5fceb9fa07d874860c00ac424ca6ed4623bfb22a0ac9517fbd31cc7efc49bc8f52f8cf61047a98b08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9663a8f89369ed8ca2724cdcc453a6c609b3ee5c57a1880ee24a99e0e273c5a2736e9ea7cbe2cfe7048fdb3556ceb90d0e5c20188b50c5174e64f2d324b633a25310c85f23042b3127f7a3ee44976b97556f3e1b82a11babd57cac342b7d2d6a14a72c1906a9745dd259f43e76b478fa9929dd7201d25422f9e8e00b349ada45156fb08c8f8852e39b28954f5fa292251a04381dc589435d687b5c4c69168b6c0f1040e54b6546b66b0f97b2bbc01f383e948a7388ac8c6c49cdde629d3a227a0dcd7a66a012c5fab224a83eae104c68c3884047d1131d6459c09b7829822d511d5a7e047b64a7151f3fb4dd64c650686a97bc8e32f64b291a57c6416b7d372afbcbc9cd7c23e826f28644f0e043f3d04ef54840c194aeb05f7b2de04a32ad874118a89dcfdca42b534f9d4ec57b4729f55ea4857586106d11829c85ee0ebc5ff93f8fd3da835521fc4640e304398cf7862ff86e237eda8baffda06d50b955a4e3df10e0674ba9ecebd1b9723044a9096f9ceefe9fc4419783a7eaeab322e32932b3bee49da0b4f7a535ccc7299b7ae5d9f7e6979bc468f96faa9ea7f9195661ce28fce18ed732b6abb63d07963b9249e39753c6f141740ae62b58ccf28945fa7e7e2cd7ea61553c6b8e848943f1408f1f9a8723ce0f80b8a14667edf5dcc05541c3eccfde0f31e075d3bef03cfe27a4379047bd4a9108fb03a39beb63caba26c4068deeb6ed1dd32bfc315aa95b7dcd7bf14c61804e068892ff4c690f6d16090d26d05ffebe8c8f2f2a114c927f3b0797cd2fca17b5e2df04cc9dac0169de623da0fe5717a948fb5514f3a36885edf8aa0ce28f0f71d080c5adbb1b179b9f2977a361b183aca323a5164d29947af4797d48637f91f2dc5692854604659e3561255cca27053fddc3826d77acf9b6b92e95e4d285c9cd5ba03184d42cdff08db901c3a904836c150ce0b42f624af92965baccf7e02190f285d827ab68265cbf6e2dbdc4711339d17feb4ec2f56c6a83df5fc68d1c8aa0bf5aeaaf0da7a4eb32686bc0e2ceda9a5de5d9026ebd5313cd5abd95a3f2713d57713a6b51af57fd83bac00221c0b035546ed8978c121e4a6783bce21b4fe5d93f4399139f90b2d17fb1eb41590e00d5b5c61ec6a8c17eb95a59d8e62478032bc50194d48d6a2abff89ebcebef5546da14a67b66fe4d93e3689b8d51fbec75939edfda7e108e6edf004a11c58e9ad022b8dace6a5c9d0914909ff5eefe3c767f49da1c7d3eb5812cfa502c540ae49821f07d715292b44f92434d450bc5bcc0f1ea228f910ad21abd52801fa2bd16ec4079d0bcc3ed753a81270fcbe6aac843f17149bb2c3b203540079619c08bfd3a4d8661f90e908a4d5b266a0d8aeb7f0fc0ec2849e40620bd60de7f355327cee10c7f949fc3517e66eea82908d88bbf36139e37c3563aec0872fafd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdff658673a45d823d8a06ce2ebb2414674aa290055f261f7559ae5632513c053b09224031bc0ff0162a1d7bd094ea075b42cd8906fe39ba6149b11909abeda821d7ddd3cfb1224869f7a4dd6b79a1c7d9b23cb8228fbf64caf89719fef16634880bd51a4347be1a754013d54f21a78c9dcf09ff845edcaef0ae1eb0ade8590318df5a753adb38d97cf85131cb4a97244b9fb1cd037b47dd87ac378e8a3080ecc10effb4783070f4edffa059f112eb85a62b56a2b7cf82c08fed7d21f6c12e303be3232a7ba6b086a242c3a90f642a3df64edacd9d76dcaa5f0268ceb2f8f016ebe99e84183a68371fa413441c87a0a650be4392077c8e79dadb3cdd0efc5e6645203e5034470ee99074c729c00244d858ca9702cf5764ca9b146a102b644ca9342bcea68fc72504b09c68c49a6cb21ee74332af3489e6d543c5e2ecd5fd2855542c3bb4541a4e5bd0975a3da9d51366be12303ed70e4b2d7b3c516cce2d8b9fb8f46bde4830073718f156abe2386ad780d3a0d5e6dd17d03105ab27df02e8d5cf81e47e1b8667749465bd376cb5a1eacb102417bb287e4cce3c08fa4341f7d9b484a20e2682e03f23be79dabe07a7b1646b1cc71131167f9f44af73c59bcbdf17b26ad306065975af980f35311630386583c07885de6bf2b9482fe4fb1de0d980329daf64c0c132ba5c0ca8538825d4bf2780378d87c9c6d8c6698a47c29d50c02b51a2096bea944c36e49d596225b262825aa87f59e73c5831fd5dcef13d3b0d64882d01f6fb64f9b93c6ece55d87d76a5b0fa0a37b3cc1adf713c737abe4c42387e39e807990f73d83018e2118c506232927c98c42bd63ce664ac8d110d7cf55a2092e2e77822498026313a44177dd137cf7b97389f6e0b6a19de59af83b885fd371507f11098d4e2b4efeef9913be7a1fa0102cb2a23f7dc6449a45c453c22224ba34b0b7097162f128b0953a1834970323a3462c06b0253ebe79732c51660dc54e91296218658f2511b848412648a03f078de5a5c94bc81c178ff6376f34d8b19ac217ecd32ba1dc3c5bfa958967e8becbf3c303d251cdd0593a3b18ca4f603253fd8b50a7e131002b1c42ef36ccf6b7f1c1a892621814f4881b2e299f2fcab1eaf3d02742f87e19e338079ede1b1bf577cd48e73cf01ba20de6e2afd7a5545cb34b686a6c6a3f4d9b0a30aa89e9af1d736d56bd37942f4b5a4e27386f4f002c79fded600f98cb370e11038b5e7efd0673eda0747e1ab47df0f7f97c061f98555ed5637bca22e6c32d786ec2ae26cf1d5238a343e8e4fd34d6930b9aed8e54e47506d27a649ff12ee7d785e674c84eac2663269800fb7c962393051e043deb904889ce7e8f53ab06e237d546e0d5ee3bde185530fd45fcacbbb66020867c85fd5b76c108e4e092f0274e0fe9bc92a008f4c4993a53441b4d2d80bc79ac42;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdc512b64b25089a975e56c64479309c3fedc49810bde8befe4c3ab3d37e3c4d867034e55e80c714eabb9693b951fa3d557b3a47cd4737a433ad0a6c83419051c4b36950e364198ea596d4e1216677cc61f12375ec7d1157d9107989e39d86d4b399ffd5fd94f7f10e503ad6eb16363c3c883e6ea41f7f8dce5839fb48e2cd1a1ce977a7bb1ff6bc53b18c2ecd63af37dc88c3968856344dcad29cac25343724897bbde82a207c857dda1b4e661f2936e0261d161b57b676af67a289717f9c093b2b40703314dfa2a709d451731c235d925c1e9325d129aa97342e930f14d7d84f2cdf95183b8485fbb9ed7426c2d2c8145ffec89f19b4b591f2da138b4287a6ccf2a50c18e7c143d1d711208fa29a47c415fcb9a5a3991a9715e02bfd99d20b870e5b524182c956942a97673951447891addf009780472a20af6dfcec8a027708db7a113bbc8dd504d0fdfdca71061097875282b30dd6103f41c2370d6e5d0b852229901e32b8d445e9f8ced9b034f91f3b10f5e41877c9629825fd2226345d353c01fe8d17d81f6d66ca29887fd567839546d9925b79fd2a4d36aa1e1b2bc606b2b234509cbe5bef81cfa7bde61382a777db23fbe3d0019be7e9439349baa552486b53b2da1e207399d8ba7f67cf94fdf44f493e103cb8c9f703929d365d88aba063745b638d2d066aab6c749705c064858366d45340d345b82b0aed83dc26938ea0892017d5044ec6b6711b6f4d82701297c55850eb8ac0dba5eec60bd76d7601e1c58075b06e43f460c97bb7e06bb5081bff1f78e92754a1839d14c68b94b66266a5bfc0e8d9339acc670a9dbdd030854c93e7b4b3a62dd8879beb57912353bd9f9dfe55630ad36ba0703a44b9afe02a5966814f58054a41bf8332622489e2f7332bdfdfd5f1fb4e53e7b01fe852928e9f9fe6d2f8aaa005d72f5e55e080c32238e964c9eb0d13e462db58fe5105d97f0ef0b71ad66f5cfb18c93f2318e15a9941df45c1a9fb0140d7574c3c0a3205f2de0b482ef42ea6f4928d253e02a839a5b60b2f8610e1100bad7a1dc0a7bb9c89f0427755e4dd6f7a666b6fe13b4b802430801bdac3dcaa6c3d9013a730ae3a853d4806cce1c5b0bd4b2187a1c205cce2cc6191b08972010f85e6eb78436a7ad59af6da9d57387949616e584eaa8bcd58277b959ec02d94db10b45e2388457971e8bf54464860bb66a27644c2333c655684db74d271e92c334e5428bff3ec46e64b562838f0a9e21bc354da5cbb3fd706a8b473fcc9cde9d4a6a2ee2f59c85ca40c6cc68e277cda72bd43b5e42981548b59c2464e948e5ccd4dad1043d0592bf197092c16065685191d9eadebcc58775872e753f4b5d02605ab3b4943b20a426a4d0d251645f121178af4fd6e9b4f0f88b46970490e5ab198935538692129e703c21255629b4bc6f90c6434fd0a342;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h35270246801cad03813c032dbd67128b83e08b226ef53e6120a9b22d2a5fed8acb181955305846cd140d476f6a19c5ab914f9894d122b878e1b11d683e95ba974e5d6241abb2491892cd8b46645bba515e5dd0a50b18000276d83169ff5ae96bd640322a4dfea1e6bcf1f4e2a88231c8cedc2e8bb5207d007988b6dc534bd5321458ed471628b5e0997e06f186723ef76f623e20df251315e943fe9364aa5b0c95b739033a971a45b731f84bbc519f09db76d3e36953c6e4f3a843ac8748b6d005d5fa011d2f3ef3ea5587d2f9c64ffaee4bc88879d915020d2a30f363063318273beb9cdfb00af658ea1739cbfebe65337fc394731266f05d46395176ae18a314dc83906a5db98fb97c74231e3f2fd04bf0cf5bb716c17bc50de9ce0d514b5112900159bacda7cfcd5ce5034768f59b640d98a203954ae2d320b39dd956e825f2a1b2603485eb957a3991abdb42f3167d34b800f77a5a0e18481d8a014335fdf5f29f9bf59415a58fa29c76ec0f4e6653102f56cd5b237c4ddbe422e89004117ea5ab0d8450f38075342891cc2f108e37868f39aa2899492b86e69b3aa5ace6520fba26e42d717e2ff735325f0e31c7a1d37a961ecb026b753ec6e3e50d6ff0bd0505793e29adce94f133810d483ac5a9b861a1fdfd060f96162b220eb68153412c4515c438e82f7a2819c3a2034b7dd6f46c2eb8f3e0f46a930fdaf3a018b3cd573807d22ea78c4a0e8f0e61e6d94957713388eba0c547dc4e0642dd208837b8166b971760cc81d4f5874237e1d79d81cc5bc498affa4e72f18ffdd578bd7211b8a363b84ee8547191a3b6176037e7271c3d01acb6b445132eba371bed3b90cdc4e8ab682e84ef8cccf2ca5c15d3cbc382a5fa86720b202f406ff78498e8a0a15d2babe962793e18c78d192a028021484a20e7245864308f8986ded41b21b7b52176b71ed58297a9e696399f3005893976cdf6344d41831f48ac7429483c0c973e1741f6107ba2828e77d96447307059dc8660fe9fd7fccb6625b33216e0bb488042a0d90bf25ef144d791843e359ad652bfcb9c6f3420c0f2b2627fc6c5353b817d38ec444e20eda3527a9567c78387532b2f57850d6eba3e79a1a0da6e6c3d0c6b3ea508b8c90c5955357262950cc6c1d48dcc4937c543f97c99d4436e5758654f91f5e9c3289407cfe6b58db78fbbe94180dec13fd2d17212b9092219e84748a9f3b4081e50491e5790114501c3d24b09013d4f3ae9ba42eb5dcf29611425dd4e2a57782f55e22354add246c9d58b674ec7431a4994185db40167533f7933b44e984293fccb561216f166876f9df4cf65d2c146659d8da981a586bb620fc2c492774f5f057ec9eda9b4e7d97a5cc39211b7eda2772e7d9e977458af5dd4c378699615ee37e9a18965101593c2a06ac1e6684b814242eecfc2fdc5223624;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h146bc4eb03680353499ed35f3b5fff0b4b606fcd269e84ddb3a761a9cda8a1e8250ec9a66d7d185d82ce35e22872fb7d615a1f7381e0aaa123e69c733ba620faaf321649ea05c48577d990c0ad085214943e5b7021231a88788f1ceeb6a5e4ed0e9b46214b29a266c4c11726261175fb9b1f2b02d010b21136e3a0f3c2d2f366c4962a8b8723bd043706dc5d7982151e223fa3b9732c668de38457e0651613625fec086739f78674c1e83387bcdeae6437dfca1adead123b2c2dd91a1f3db4e0b5efd04ed6a34f96a79f0ee6593a8c9d22b2d5355e159fd8bed56afe6c793900098d6271faa53a96d99b2d61d4c39de000cc2377d6eb965c0b891e69b3f2299b4bf31fb6b9c75f1ddddaf427deaa49588a09f8b1fcf3fc08827f274e53710cc442db514bc1ba42471833c0427a7755ec84e13c842221ea52c9610f312a17aacf1f426ab3201e87f0435b43c9084f0f06f5c393313b72bd342f3afcacc9ca1b4c273559009ea4a5285b491168e1bfac75874ac7e26d5403435e7a6e91a7aa740a96f128adfb40c8bf729b1962a851823ad7f2aea7761fbb48d38369b4933c08671714ee559ed02cac42e4e7a6a0db6709930106fdb3c3c303fba5bed305fbfd8b65b35421d7ff21a02411e46b692f39c53248069a67d175b24553c17e976ec119137eae62083f85bded577254667cdef5c9a99d7576ab7196230d4c66049ff09c9c3a48bfc834896d2ff2b733c4a16376caa8b54b5ec62e9d9a11e36519d94d5dc08b7301a6e3dbc70a2940f9e0d34e371ed6680a2bb6fc5e412d90bfa48d52b85316743910a28c3e4df34ca8de6523e867388551eeab868a97dbad66662a65783284e83ad24257e1f7248c1c84b0437479a7e59d3ca57f94f0bec3d737e2ac7fa7dcddfb1f8fc1f51e3668e70f7da9b40015227543fbecf5673d15700703d4bf781f45fce3b6a5c5e6175cd42f468b6a9282027da982a364a6d84d2c920901c8a087985fed09f56d39d7099035d8e38b9b8a497135f6ff4b7aad7eadc9efd326c7d09568e60d2e8f4481c1b7747fa0ef2cb11ef4ecc9e216c04b46e02a7d48f01c7cedc277283f7186ef798a8285d671e9a8e3014891c1e903e66ed7aa9efb1141e199d0f5a5d5d3b45fec4c0b096e305b6e270c593dcd40dafde4eac6e95990aa292bc21bd82c8141064fefded2addc29ac990d5e5888f9c4a26b4bfd400bb7e8786d78f3c4577e5fd87f94eeccb627b920c89158b8dddb5be9c20edc7897003888b1ef9d802e629259e95dded97195b408a693077e56d460c34a8b002471ed95b1309d401b6208f490eae2ca1ba49164fda69522983defe45728f18be61c43ad34e1baaf26cfd7775be1bcd9a53d270e9c64ce350b513f19069521f018201ea59d2c56955be65b48081e528c3755b1cda3feeb3c4ddf2b43ee2898a3a92c71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h834f0cae58fdcce8493980c10aec43c3a0c7395430c6352beb265a90c7c972323c383a0169df251685f16ceafbfa6b39ea66a662834a32b74c070b30a3b49127afde14dea52e2f07abfb03000e1daf6c3e33c5db065ecb8a83a3c16cd1d966383329b35e5d7b70ffee87f936f0db851b312d7c6ba8918dfbc2fefc1bff15c6e9b6a3090bc1f673bb5ff1d7cffe4550c606907b9443e28e435ebf9405515e8ed43a8c746347a9e01a1691c4320d34ec9c962d0a0fb4bf13473e627d26e28eb8306c8619334e16fbd713967729fb8c9d0dc7898a9496c568bb687f07fd5365492ffbe66ea8af0c15da5b6a2b09a6085fbf07ece0cc083bdd27188f2e793df446743919679e5eadb1e9b4156005edd807f0edd4625dc8d4a3965c23f55c264d55bab41e9c0db3a31e1cdbc5a544252e80d911d1158a90249c6205dfa2899eaf9e25d7cd5039c313c393d4d5be11c6e97e323f31b6f1be901a491f28183f5eaa0f85ba55520bb05e406e3eaf95a20f771ec284d1e9d739e9a516bcae33b378ae3500d0c82f0848a056a757cce46597ccce63ffde387a13e09ad8306954aba10b790ac1971f96af08eb675c2651c64205acbb5215d08a365ffb8b09ca70da2d57d4b7100b9029268cf6063adff0c419975608cecc9dce3588eba6cad6444d4c0043efb8d9439886bbfc245ddb818d71ce4e269d8ac8edaa9c2f9bf2794c61b9d44b8ac91750679c476f8f4174fce522cd2a78813290d5a81a62f959007a1675aa3ee137111291ee2284e2e3604c67e658cce3aaeb35854fec6ba396c04bd480e19793b26b63efbbbb047ff586f684ed408abb98318c5d0042f4a98ace51b25ae4699fc7c68d0621a39c0d81083a7fa7e11a2249b15962b4b3af4248c3a098277b93a1e9d513c73c38f0a60acbb4fcf3a51d5fb11f8fdf81d8ef4e5776ff7de2999a0af4941cecc21bcdbc6b921e0721279f060aa34f3fcc4f9f71dfbb33a751fd3e4ab774f77a7633ce33c99b4c59052ee0a865f72ee43cb4b507c306ca35b6e0cd9ff2b44ee95ba7c540117bc8f0b672d62b2ef58b103a2403694f7c172856a3d9f7b30d9d683b6038baf371946cce37f337bad2e54e15f1390e7bf9b94722f9f47b940cbb13fc95c2e5b5e56646bbab0ea1364def9fd50fb80101773bf423a8d3e68be24beb19571a39afe5bb00537f233d298e63fa24b99bb938d68fc3e9002f6045593a0dbe15d55d1128491f2c67ed7f81c41f3a437f8edeeb927088c4fd6c008ad476a73012f09d446f2701062f53af893df5f73610269f9bdb22d6339a5faf0c61cf7137917d0084c37416d3b50a6b1ea0056094ea73cf174ce2ecb987bf980a72fa2c07cb122953f06da8499dcf9b4d6226efaac6390d8843dc6b592dccb5a760cf3c3eadf33ca3fc4c8e42e61ac786cfc89f6075fd7ea7d0a0de81b04a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h44711cbf43c843a00ff5396f7a7fa8fbfe3b68f7ded8d6e966c299646dd2051b8a2ead0c6d6461e34c317cfdd61bc2f92ed485d0eafaaca89ec9e38401110343512b03dd581bd6da4ca7e8ad115acbfcf2b8a159fe8e3667ea7782f92ec87b64818e42cb9359594530477d877824b8ae054669bd0654ccfb2d3244e12c4d45e1e9ecac55816f55342add7993aac286290392d25b220e6efd0e592e314f1e5e49b3e5aaadeeea4ae27be974ee9a6e9c3a38d007c930bc050bba7e6c2c5c1d744973ddad285757c2039908c88776daed6cfaaa7c3f4e95c0a751ad6537908193789f2597c510f450161e7ae876263ba7a0555c3a31f90e38561708a4c9cfd60cb4de8834133476b8d08f51c7cbc2ee7171b780f6959a481fda40e13fb730f0619d84c57e1fa84b85ae00102dfe7e3d78622f2d6441e35f8eac428dd03f3208ba7cbee727f05fb7bae47916f1f485a7193c4d7bd828e9aaa0ad714c047a14d86ded63a565fe5a5b3c2babd05c4cd1c6abbb125b57e6623faf4d7ae37f3b386417316e88914e8ee8ddfa878f39d6c8ae0e397df27d8df4f5826c3a963f51ec84a153a7adfe298f3718aa2e707d51f7853130b535c64b5d1e134da84b1946f75816ebc00342f976629eb59d1b9c656d912803cfc7b97181cdcc1774b9cb0da772ed1c84fd802674d5eab224307987588ec33dc31921ecd8d2d7529c830643f8f06a8811add61b1947ee16946dbfc38c2a92d34e81a85a53bfd77938f8fa5d22eb43f65d53b6ec214e45d517d4b2da83a4c777a7f53a86cdd450c68eea6a218ced317086e31646737b7ca6519e630a1e8cb08c3eb7ae44769b976d92ee82c296d7a15e05c10fc6c55cae2d0dc861d511079951cf7df0dc1858540a4544030db27f07248b5342eacb9aefda1d4baf939442697805bad034f68f1c5f7b437ed9da47d8802e6ca6619896a6fcfb7ea51568bee85b66951cf3efe68754459a84164d64041845e77ff83dd4f11dc2f1dab853d7e25989e3a5c455bb48f05d759291a8c2918df1903b0d7479866990924cab2b9755c408d05ba7cd3dec1d0d3d37d066177491092bb53e865224833e7ef830f7c97b67b4d7f4e9152fef089a33751ed683cf3c8afd6326e064a9a54012a7da0b0cc03a7e145edd54d894fd6427e66a5c34011656e0cf294a8d396bc6083c5fcaf246882509b17fa58b9ee7885ceca013fd5a1c6217e204ed9c5a010f0770f401ad76f9871bf4a9f11c96ee4a95a930b9a057d357d95e325985687e6f9fde4a38e3906bc47bba10a0fac5d3e69f8de2bfd6a4b84e5f58fb7c576cc2fbf74c2196343d752871b6d1238feb5c7e8b0930fee0de7883f8ced678f90e93b0e14843d0843816ac735787a3b392ce6cd7a647d3689d29067da1fe5750c7a6ca53a786f78786ce4db06edd5f44375b212eac1fd557e28b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h26412c826f83e6ba2150885e264162308d73d0942d20cd755c33e1c238b6d7d152dae72f532c2f4999e2ca433743d6ead836c5e6db927da4648c2a4bf7a4d857b9a163b1d282d21f99b9cc832df5676a5c02a7560350f0e2eec1b212e7c643d088b5a3d799d7c4d7dd438cf5fb396135253f46c155f24e33d3677302d1331be86883b9743159a911f100dea90393732b2f9db9a5aea61b732dc00fcbd1b4ca43a00eb219727d979ca1039e10f75120ee8497bbff223f571cef0f985a1ef67c4f52a02a5557a4ac4975bd973ef211b3f453bafd74b47f314c31b30d4693e812771b7fa64c2e5b9356a64d96bc45e90259fc9703ffb52b7cdfffa42d2ed58b3e1094517a6f7c959d14b68a22ba749ebac96b28bf39a257cb6f803d2b46b4e506606844d32f227e547bab14eb4c2ed59afee70b117c90218eea119d34a283e0ef8d49c2267aa2ed17e4c6f5bc3bc7790ac583302b95054f7c62da78bd0f689d31042395f5f6c8b9199b97639e3100afbabbf534e668359cffc45973143cf082f85b80a3bd046d78d5e8f9b0eccfb0bab8414e880f82044f72ce3513c230bda8cbac6d9e8a3ee131ebe5d10b32e22a1870189885458f316ef88e180d136024e370c01fec837e66b32b8586b79bd8d5c856781fe49efde522fd1db8ff6297db60d32a69e4bd6ef924bd932476f7f2bebc53aaca31dcf93d36793e3b0b45eb8c116d2dcaefd72fc298ee1205b33b637fb8b31c16a4cf8c4f45019e3ac43143e588b607483e804ef1f5a025d776bfc540cf204138456926c5b77a50903bb5509f1af255d08eb114ef8894f6f6ac770eda4255bcb7f2937c392c711d9081c4e4d7f852fb79f6c0b4d2349c1b09cb171a30567f24b2cc9c78ec6c3c9d282c4a57d9a898ca0c5a3ba0ccc44ab2cd9bfe9db6052ed9cb5790869e7919e0835c86a945ea5552758e255e7619c741b464316e8673d9bd03629db6a3e0e10e7c97208f473e11b78d7abc7b7c4adb0a10ffa07a910f73c1f80c569621d8f0cac6e687ceee918ce49e9682133a6502f562ebf86d9bd0e23c7d06da82dbb7311944f3cf4ef8d1887fac76cea06ebb1cfcfb0c4f85a6248578b0275450e291b3fe14788d33b3aa03e5ba0daf52d124d05514119b3de780e062cac6ea03449bfa9e96248eefc294e7bc3122bb854e405f4540a334df05f8c8a8ebb0792e20190ec028148104770f3d50e290966200187063e0a05be9d94feb604036545394c4f73b54b3fa05bbed53e0e632e4257536ded26c9c162491c310b6c627c37c3f8c15a50537c60d66cffc73cf989c78012ac1d569bf8141f1684699e1c536b6b7721a2d579dc7a6aa48e9f2925f828d1a7fc939647e8d867180f03cbd96edcb1230584b7a8de9eed434357713cf9dfa1a5dcd3d3858c17c33a47a836e79c5fd2527ef3e29a3649a03e50fc7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf35e0cd1f1283e1a68417dab38b7e160f4f75e08d7bdce66dadff1e8ea91efc4dde42d39852079cbb4054ecb48c5a07029726a347ecd0cede9d1bb93904638f47ecd8cc5698c0298e7f3536412f717497dd0c4e42b3f6d205055d1003bcca9c2b4066087513d089cbcd9083fe3a0246614100bef81da85777349fac6c62539aec059184c55ca1edf93556ef809ac2229d88db9985867585a0d7217db7ef7ac8b46fafd69e8888e64e702c5d7269a3d74bb440e84d3ae3c8f2b1b18de165c6269ac1f38ad6dcdbe036edb72fd31bb948e45246e3c2ee1b5b98c069ccf20fed6b0aa26a99b8b18ed793c2546869b0d82b845a8029d7fc1d8784d69d434e9564839cb7887210dfa6609b23fe52dd4efb2e1b6104e0bfdff3553d1647c159319011b2d317653b5f283a0fa71b4d80b70f3f296d3e31fe4dba20ab3e9d5d762bac90713cae0c3eee22b47a4b9e67714479ff8404f76720c99d2f50a31d15cb320f8af7e306542928b2f811b51e240bef64fed2d8b3c7bbec0dfe41fc325b7f98bc8ff0d39c93a72673c067bf1418b1c398dfc5641fb3d955988e8fd371420f8cd938905505a5f7cace4fbf087a32e552797e2d20a6d74c579ffb83cef71b1601661645de612a260a36ef04f09bdcfab17565faff53aa37fcb9f47d885e592d86799ab378d99bcc8c6b68aa9f310f6ff2031dde832010e59dc5e621087a9717f431e4046aa7f16e39cd60881f03cbc0d810fa930d9971d6094721e0583bbe2eff652d977a71b916a9de20052777f0ae360247d074eb4400bb120548ddc13a551c28188616d92eb40fa341e8982250b941a1c969a04e24a1b849a1b530a8a2eea2eb732629698ab3762d528c349571f3c7655b7cd1122b904ba9080a8935e68417ad08a314657a8300efbd6684dc1d911b7a3b1b0d3ac54b1115363ca1f6e4d74828790e0fe27050ee7bce9b6151c0f235397787b122376befcddca6a93fdc02285e483afd0decbbd179e306c7885d48777fdd2054a5fc71801c95efbfb1c1e66350d48bd4a11d029582421e6345fd2c196cf7b053e73da9e25b50e3e27dd24ad18a099877140daa3060502d0c04e8c819517d4511affb8a69b98de0bf347767be04ac8453871b0195425d82ce726b51153c9cadd10647cda3899540aa10c1780214d542fc243fe9db7ec36f79e773db57f766a20f02b665b7993823dcf25863c81bd2fc0d1019cd5d8bc574beeb838dc015f9bb6583c88a1516d69b2b7bf1b1cf2743aecfa2ea7144047a024e01ea99b1914456d1f00f49365eef59b026cb1387745fe32c24268b2d1ded1777ff8b69939d33cd3837afb3b343f67768f1b2e92de2b9567ad3230336ba232168ad952caca5dbe7b8a3b2189a64fab431df60b8b07e9fb90806feae5ccf0caaeda2dfa86833d24cb296ce80337d3626095b87708c39ed1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb1cceca16d4a3243fa71b6f78ccbc7dc5b7e5653e7e86e4c1b4be657323a3b02b55426a0cc4a23c0c3e0e990368a7249c00b7d92f50cea849efe01930b79a997a95cbfcaff90d397b0b62965d7a138821b89a818e2a1a44ad317a25890360f58623373b3ccf82c21b0c137439dc16bacfa2fd6d201b60681157bbae1f8b8f6f1c5b2ae38d840029d9833fe0a687e53c3bf9b0087e06c398063326d503124f0056cc392f65997090ae04e26951ef24aa7b6da92d807d3fa73f4cffed7e23a766761debe1298a38a36ddad66bab02bb3c37fc24d9908b3a7ff1ac80c3f8f6b450dc5864eb52db1d356c7388f6b413a64844fbff9b1dfa2c6efb0b8f0d4d938367507f508bba56882730f042885d7ee0e9f666adeb6af2573ef9e9ce181af09a7a2246f5cd720e1cd3276a776a7bc7cde8f3006351d51f542ccd11fd3dad7d62f259445495241f0731718197a741836ea021afe0dfd6fb227c1984c543dc0bebf28bf0b5ac8429b46bc3af2321367b12fcf2a49a61e2dcf35664184c0785381a66be8d48adf385eec1940ec811e3203795324376abf900f65eb51d179e7cbbff0a2c42ad81803ef6ab782848001403bb7c61db6bf3a59abc49a1ec3208ccacac1addb916daa6ac93f76cda0f6c5c3671cb04da902514a4ecf818c78b774c36338ec382787af8bc468a99d0f6a125838411b42b369601bd77ce6861cd7c0b80ef36e02941cb33f018d4cd0de00405b8aa8e04ba591e914167d8901659b31b46dbbd4948931615dd0fd845599442452f0f1d0a0ecb386a657c9aa46c6cd66c8ed45de6922d33a12abe20d1f94260a3ce6f67d23d3da994fad83960d1cbbf59348ffbb58552a089c717e106dc4039727fcbfc288912d34db0afdbf86fb63ac2d172c839d09042314c90aa16a1a2b451be1fa119949ecdbbaa53678ba2b621080f5bbbb9ab82e4eb6f13a0550b94ba015be832292fd6be57549b0e331c22d5d115dd540ae34368b05c52a25300f33c53e6af69a1072786976122d27ea656b925311f7998368a713b0417e1fb0df89f927366f17566dd9123630c05de6134157d960634e9cc27f2477ac7c9ad4f0d439b7e3d0cb7a9753687ba508825e1b4b0bcc2d14bde7cd591ff4ce7dc0403d24d55952b6eaba4778aa8781767a74dfa17d28efedcdfb0ceb3a517b2b9eabb93b7f37c44f4ffc8f9cc2696ca8b6040994950fa588c2648ed9f4613943dabbd7ac3e7cff52ab94f8e7d282b840506990b894be67a8fba9f5eb12320c7e72f2c4b13f70a4d7419440468d7af8d22532436b1ad01c2eae0a57a365c72e4b83a312172ef6ab2e0c8354951e3992b91c1da652245a33c0c8d1908b2f66711dfa6e35388cfb227f562fe2b06aada3cae8fe5328a0518b016697fc5234f362e92844b74a644b3f602d15e3e7a629a16c896a96c9457fadd768;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3c8ec7043d7996753e6128f74e08ee6d87092ab9b0639a00140a6ae91401ef1a5084ea6a5128fef854902846d23aeacf8ceb1b7cae70cf9f159eca517e6480e446d8e154bfe395fd103462a4c8903dcf374375e5e0a465a6020e3e0e20efdc1248bfbe281fb36a8db92f76abc7770089eaf57e45598021b48afac420b9237692feff34d1cc8caba87477dad5c330415b7bcb4d4bd3b0b0242842d8a72d58aece62ba08a108b0626adfc5031f795e17810a2eb3a0fc19ffd39723484cbc7782e3a66712067cdc00a45dd271cd65de07158cb9b8d1e6a3c41e8c5bfb0ddc49486ad996aa0e753fe04566b909d16e032bd9c17ef3763fbb8f8e287c14525aa4ca420db12685b9890191316c93219c5f4fdc5a0a3e51c4cae128b1b6372fa46c7cc863be9534498eb3cd572022c8e5b586a85bf7506b4672d03742f5ac2e0d66efa38d773b8caad6ea2e15756d7b3204ed55560144280269925676877e3a36f89e2a1a13e3da94d1ea32b1f6a9e28f17a1e218300d099f07e76ba0727c2326a97e8ea27934088286036aad099dd09c4f574d10559af6d2f39d8e4e58b5d0b6633f3bfce94e1f7443ae4c1bd579c20d514d69135e6196d5aba73c1d747c156b65c8288c3ef9cd2f7b9befb10a630a84827b1cfdd840c210798c905ebd0268bdfa1d0c272dfba5f458206656514e33bcf4edafca20222b953be2f6e2cd1edf2090f9ef2380a04e8b5e4a7dde15925f68038c3d191e6ad74f0fc48ace5c0a00d162a5c610469c158499ab685b85364520f659b6b14c1fd107f7a9bfc24585195206206ee933b276a92dba278835f3d358bfe4779aece7eefbcaf95f6c655ba18e0520f4e41373ba7758cf0957a17f6d3469bc3125ad707d00d77adc7730bc7d379a9d2f166dadd11d61d2bb6a79fc853021a3d3629d81b45d0ec5cc93aab152fa8017e5db5e11213d987eab02b5b29a1e493a63898130d1bbef40608f15ec341c39664871a7338c55c1e30e41d512910170f8755c8576befc6bbc93259a8a6e26d90af083e3dc37b8413ed7f94d38a6cad1f752ecb22416aa93d7ac06f2b5dfa63114b241b7a4e80cfb51846a242e31badf3d6c58e31b091bb39c87593a3255eafe384846c6db8c79b1d9f3cbe8a801ed7bba60385ef7e07cf478d4b870d86a7bb3fdd4f2e61c846106d2db644b46ef438f5131f09fc658165e96dfce503ddbf82fdd8e1b48592c718311daa66e582f5283bf8001d67605acbe14f342f38f9e60ebf789e39a24ec58fb4556bff00cd04bd2c7321f136e86d4aa4ffa502be6074465191277e64290808f1f6d432125b2b46d08cdeb0c3e8e7809d0adeac446770b03abfc883509352dd3d94530dd16ff019fdb4d55673b1d232da635c27be3f7f67be4b29e65629f3b07b312e0d88e95299f2f66dc531b0e1e687b95e560099af54b2696;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hccb7766da624c4be91b890a3c5284f2b7b9cf60cdd492b21dc537345dc3b01bb55a3238b114330deab3d8b7cfce23c8fd4f6d2be5ac6eb16242b33ec4718e1584667cab7e01cfc29faa72d986c7909197aee6c6dc53e678344dc8c12950b29024dca4efbef0ac54651e55bd4fdeb8303d8e8122310bff66f7eefb429c2a2c7d3dde371ced73cf0d44aa6296a5b06f9d1b2282d38f872b364604932a1c3b39018c1921c391a7b0161ced3d57b04eb0388a6e23543e7421f6fcdacfd52ef6eb01d67dacb20c5a223ce85dba5df45d4a65887f1046d230c03588cd75287db034a8038c1819b27a0be23720db6f06b656e05157d2467cdeda0966978ad9c9c3ad8c08bb5cc18907ba511ea8d04d0789d6fca9ce96c787878f1de949585cc19e96a1a3ca51bfc1d5ae44fdba66ef4bb221a27d7fcc80d96663f7001bdd294d383dc7ffa8e87665b6e10d58070db62af2b13ccfd76e93310caa1da6481c6cee1ee4dca449a9174610d161365e9e2c945a6f812b95ca4ec00f79cca1518db1b068c2bbf6beb31638c989dde5166987417454e616b3103c32f9b036ded97d3d68d1ab3cdc42888763290c17ec4f341d60b4ac1bb03c3f172e24d131d901ef262791c3aae1109cbc4dfe97cf0d2116b4656ec4f3643e6129739e03c3a9153ab9d916cdff618530e5ddef8e6f5d55d90e15384d8e53d44f97daf89db0124b79f922402008089d4c71c200fca14d715ab8cef4107f878e79aaafeba7652e95c3eed72fffe9d23ca3684a6609426d2d2e07244bf08a2f0cb809974abbcb98f773fe5d487683419e550a3f593ace0122a1741d875483e58c52704be117e5eb34759e97ce1fc6da9f7be122ea68a9baeafc115ed5cabab7830795a643e6c2d24b7d0071e7245c3ef4a6c25bbeece27333abd4047997849c939c9bc5bc71fbc3fc20264d20df78416720f9282ee8dfa8868f91030db0784809d9cd0a8af68c410872675ff0ffb9b09e9b4360145c5c5988b5c0ff584cbbd69280983a05013540a589641c6fe734fbd4426e0bd9250f7a051b1ea9c531fd159ed3967e6cdadd2e3e10b42f5726972f3bb9b0b587208df5f0802b22ce190ab784cef56d05b6afbe77da8947ee7819d405e277a8b1d3c41ef05713bb206cfaa76e029e9ba53ec288c88998a28ccff267f6863e30e6561a9270165d2c90f75c3c62a2abc3bcf49976115c9a863a1a75cfbeb1b90c673bb18758a4f929c91ba5f892799a0f5f585c2fe258f5d4e496f9ec1307c68cd2a7846eb21291b3b639e21da916fc32fa33d5bce449a822bfbecdffd4f40d226ff3221904529c445bd9e498261e9f9f8e28a7b29e9c57f4d5ab8c670897e45a375661d59b9c880c63adb1f63f4152d839403dc90fa8a1d15eeb6017c51415d794f7d797440dfeddac7dc13f168d8ee932f24423c0d0f0cfc7d5a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfb97b90991a6c58b4424d30cc2b392db03718d708c2d13cffefe5c122715262f678815d4f2a8837bb9bc8406ef8a88b84f52207eef5eb6a39593e2bff52bd5fc4cb609192f1ef13c8617223c0df503a205e0ee15120aa8c158d94b24a064c8d45e6b1998bd0c20fb135e092e63cf42a3785e7e37939c912810d7cd2dabbc297dbe02586d77682cf88a53c3adc33c8cdc837ac1ad0f0bec8f4fb1e1aed14f3ef15c500ad0a9d0b6132dc770bad342ebd5b8242c411c05d943a12ac5ad281ff6070a7bf299055baceed1ebaf73000715c8383aaca455007a49741de6bb69c031d10f4027ad09005a1265ddf2d43f51928b0c13ac1b6c9a31c353dcee24fb9f4fae84abe11b30bb242ea36f4de3bb603df4d50e841eb7e8ab877a149d5d559874167bc7705041238de75dd413d02d5eca9b940c990ae3e293374d54110ba2529feab939c5c923dc1d748fb717e26d6a34e15f5cc511a809e2d38a90323a150a1daf760b3ed0dd60839151521bb5208550087d122a372071c65db37c2a66e5ff8054287d6305e7535d38ada32a4062698b385e0434424b0446b9557e6d32a87d74d174aa88464a5ec2776af179e1d632e7140c2c3479a3a253bb07d49eb0985e2c06b9ef5f22be69130bc07cd6603e9472379f3a36cd74704f98fb61a5be86d4d0389badbc385f795046e66288bfe8e9f148ba42901bb2bc0433cdf55aaf39c96fb267de72eb18ea982b45024807a17298010e948c76c71ae8e391e0ebb39d19b5b92a86ef502e292e4829babce07ed0f346ced3b5b2232a445c20d08b457919087b70c1c34255a6e020c9bf63e22c0b21ea40e4d93fff0320ed5aedacc3c4412b49e6d2bbc0ce03d628d9a2328975a3b7c6e314445efafea38aea63594e44c6964fd5b52f519e6c8a9414467b1f12c2dc29009677403cf64e7d2fedd7fefb5a2f0a7b1fd5889a96fbce8e322da0e988c853793e4ee79d3d45ed379ee991b469a8f2f2c97417c311ec1ad501423864338eb13119c507fe6782b55b46df02a63ac1a41c2fbb68fc2d31e88f40aea4185e572e906fb16e8d95b2aa778c5527501594fb80ccdbe03b5b500b12ff46cecf31ec3bc32c9930853d762815ac23938cc235ee6bfefdf0bd94de3e9e9a397d00ec0756c1dbb3f574ce8830e52b41d8200ef8638bb3aada413a01008a6cd874ffabf9007c543ce7891c6cba222d01220c64ef97499ba3a56e50fbc5f0c123c103f582a43b2affc105e454b13c95882dd1ad6186066e4d2b5d3738f89453f0fe9ba77daef80eb2451015e6710c6efc8d447078e850ad860214bf93d5da419ee95370286424976dd7cd1a49dfee6d68768878430cb50d4424dca5b53b045be931db30766d34e6a8bdb50706dd46666c91e73a1f3fb1cbf31555fa7b7ba445db947fdb5f59b04d7aa01a3a2638794f09010aee6375;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h43b81817e807898c2d1f183b9e0b2e90103229aef407b2ad5902e1d18634455cade627521dd4b99590129cdce335c9b60ffb856ee2c347d1d01ded6aa111118b6e98573ab75af2f39e76bb20cc4be375d6bd823051a7c9634ba7d2a61a9bcbe085e057a2ac63c4ed1e54bb3cdf9eefcfb07350d340476158a62935031012137a04169ce4e5703c1887600f734853f488efd4bf8bcc773c5e82f3f80fe58b0191edc2666da8dd4054e0f179e35b1ae1099e54b32bee461f9b6571555800fbf0efaad20b310af25579ee425c6872b87f2a0d763d4d5bbd56bb2fc81e2f7a2cf52757c654052d430bf713504315d0265b62fd12410a7bd87cb4f58bc615f143c96f26ecaee3f8925afa23996a8640916e293fb25be775c3fd31895ec7e5d7a65766c8a7b09e5d1cbcadf8e5ea22c3870a3a33eefb4768a05f89e12e5330d9c21353b6efe90105916049058d4161d6d1d70f8d0a02aa900a5acab4451899a36a3950199957d0a6c84334d117720baea3b8377fa3a4d9b7fae7492a78bcd867788628ddc081390d521c46a82223795a5eeaf34cac8f21359944b733bcfec62a89026ecd1ccd2cb92005f46367baa1336170c2e744ef53cdda48dbef05404c6558496da10f0e24ffbf7749de2890ca10b4fc9aaad0efe4e2cf4d42bd647e176d77ff9587c5d911a780e411a8f3a2298860b80a7d00104b3ea31017b51dde64170c3a8406b2f71d34a8ac6d12570a60d935e6dd93c23921e45a40d59fc8f3fda4f33c848752846083acb24d7edbb6599138dbeb92e01366127b520b0331de88cad79c51d3bd3c50767588c887017445416719de043cacea71931a3a603ec2e5a5d463eb87def88ff3e4beca70ccd8e5c371d171391f1d3a7358a17285248df05b6eb3dbd940cb49d24d718f8323ad55233684c6bd156527251465804ee520ae1d4d2a45a829418bab3dfe238bef374d190528eb89c93c1af4176605895a288fa929850191458eb59596579b84ae0b579daca50ba1538c0b0491c805ad8149443cd77420ce58fd610d64cc881c2c2fefa62a04a7e664344714a7e87ed3d250bd7f9be639ddecb102929211af3edca577aa2075349c834e475bc808dbbcc4d78712337d4df2af23e628420708dfcab480738afe64129b57d328102eefdc5da35eba855f19e194aa42752b89a036a58295d59bda4a47889ea5f4d1e9e73a74700fa256283ceb9d55e1ef8ccb6cb9f6e488a5114145278999ec7b292976b282c8c7870c71b8f2d371e60e4fd7f22af0e566d8957640b391afe7241b22b64b90bd0139eeee0900d45c2e9e8824b3119d814b11e1ab0cbc8e0511b95671b6c8cd8b0601000f7794d6db577cb9fe06711b8707b91a405c2c91fb7df6125179e16a63a177577cdb4566e01af38d09506680ef889b9e0be25042c6ab613c4f2693ee9c4af8d3fa0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h75d11ddeb1118e30cb06a8e8e01d3c725884e444435ac5a0639c5d06f04fa94194b65f1a251b6d1b47504dd8d1ecd67e5fc703f55e2fdc64452d731bc64ccf9b51155c35852e2a6f723968e8fe93dffee47152a214db5c122b1c4bc06b9ffe34fe788fa42495d99d44a288f04c7cb40771e1e1444363c1eb057fa9ce559785bf314731d492d8091788dc41bab041bda4af83e0fdc041f3f0b1307d1ebd13ff699a358ebbd2fc72861367fbb78da030ccb62bda7709f01a1214d6b49c41ddbbc7366a9657c98302213954808d204734b8e37b6c30e6a0a81f7fed0ad3f58371b2d4ce0520adb210137321144d8ed62d57f41054bd9eb34c61bbdaa1c610b5f04a9cce5fa97e7c4cce9a48c1190f92d9db91a32a40d5e562935c5418395904d3cdcc37cc1e4229b48d135f26cb72a36974d5821c66bc277f46cf09116efb399134ea49e759b1d8f558ac3cae102286e388bf4a43a8282db6ae4c9095a7d02e44a34c84bb326a8cdeb8bc0cf7b0774ce68c6355685b97e9d5b76d597662ab28730c532ebec374a6336cf7caa02f27770f0b62e5a983b4d337a33551943220d6abf83e2555b1d0fdbc7ed0b6012a2e1fb1ade32a07e1e8ffc3adfd82c1a5969f43ebfd1aab6b6f79c13fe7a682e51a067b8a45d054fae479af13c1d1294190eafc2886d17b38cd8eef690abeb8bf819f5e5e0b1e7cefb3bf8ee5f06059c087f36f4290afadde68f55cc849fa021505886d5a58986283d7c210a8daba873adbd8e6cf6d28c486b054f06896b6b6c4d9255dffa93d32a7b40e7155b0e1c1df7e28e393f32ff879d4fda2df4390fbefddbcb9ac785daea8ed4fcfc918b184d46cdd73fd0db40f0423f785d613e5ec47ce1e3542df7a7af88d853f5ef31b06bd8ca1822adc075d11f0d8ac3b20c397e26f7fc75099cfaf7e7565e77d2f321dddfd2366fe97db128d452f0ed1eb91825c5d1386b3107d80ad5fec82e1fff499d17f9468bb3454fd9cfe8ba29da1d8a34cc2c40a5fd68a155eda49f32d210942a130fe73685a70925e6da0e4e5ca046e862721f9688f11a78984e3c7f69335c9a94a0ea3e2409b8877cf19535bfc5187a0e42b44e6d556f41c05fc008ca517dd0569d76d4f64cd29d297687cb89238eb6f0d7f66d404a5fae4cc65591f642ca19f75904e76840fb538ce5203b54b8db9bdcf57833c453fde41723c7f7ad5ab37d340b8c9ccb3de60ea8a68976cccbf6264d9b020dbad1a53115470ce982d3d5498db2e5a4ddadcfcdf309a4e8e28985d2e44f3220e5a890435c8cc8cb9d9701029dcfd5c5a666fba10f8bcd2e258a3ed50f7eb5b38b8a0668410a5b78d4e1287c98369d8122c462c0716c38dc8bb6d14f969138c37202abf541d4c70e1068c6687c84027ab61a4a09f18c6c81747b6877587722064d150f247d5708a67eba47d3cb70fbcfc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1ccafa207fc5bb337dd85fe8f8c278f9c02e0d137afa6b09c0a311d489bdeb049b895b58db2f575e70f2e4d634876d2a94a10e53c94848ac3d8f5d8092e0783d06d98e1d6c49cc7fbdc691470ea267448934bbbeb6e166554a1248e832c2a511636a2133124675218611e25471593b38d8483366c8b0f24363af762e1aba18f8bf8cd3bc3ce4f7d85cbfc9be36068dd5a0fe66bb21a4e758e252ca509a33f3b5ea9749d320c9721596e38da98f02f077584963f689250c816142dbbbd3d259611ac9934063a069b4a9d13e0234cb652ec5b3f1125ecb154011f7677b6b588a9c53b1fef2ae1d6345fc0ebf632fc166c436d52fb4fd8aefd944ea864ec2ceee06ff90c401309d10f694ec97de687456624e7af4c7d5d9307b283d069ae5615406049a36d1f541fcb40b04035a261c77e9fb8ec1b308c13041304e9e053f625616cf4064bb7ed2a53ed0c6bfe533bb18f641752740d80321e21a848731cca9ae3ee0f38fe0e8b395675ffc25bee64b27166a1056bd13d84b58b3bf1011440859223299326019ff660f3e6c8b31c725a777b39b842e17aa0e98730b55a22a91cde4cfe48f9c07f333d4b6dafcbd4edc83249aba5b7ab48e8210a809642cea96b94ed30d8bb219e3ffcf81290215d6ca08fa43374e975d75de6062d7bbcc335804cafbe0354b278565a64db3c6574f8614f130a115c9c1ba7af368bade218780fef4edc3f21723643ab898e77ae386f1c29734435300dcb746baac5951ed19f0b1ccd5d9ea9b6387bdcd5788f91ffdfccab9064070f904790a0a2859da15d2b9d5215318fed895a988437d42ef13199b387161c3a0fcff82b454ac9d65ba495536b9b91a1f477f9af313cc00fca86d769ed391996c6c8a37eeab80bd35f01e17dd97774c773d2b6a44ab44a8136d016a9a4083ae6804d8cdaabf4c53dfdc096a785a5024a5fc7262130777cbfa1ab27e4ba4f2a886b061b2f8af2a70611514d0ef96134c41077c4ca9c0ffbae00b8e04ab8dd5c202cde192ee40a661d98bd2bb571e8252c89e48c9a1641079688057ff9c063c4d27a214a26b842d78e4e9708eb0641c73fc093407f9c18669fc3002b768c5b410fb8bae4090ed1619fe5d195cc3a743e03f43a210388b5095a91acb635db78c2efc6dfa88c8613fe6a259454182a48b77f016fa5bc427a142d72f6f0dfdf481184e04044641985649dd5d562091ad70c9970ee10c2edd4869f00235b4c1622def9073af389cd8e0cf4a366952ad8a8b7b39f11e585a19600fda063d839a5e956d4c0dfcb8f8eaa18776e98e34360110e92bf781fc10a4b862041b9ebea198990bdffa83ab92f48ecb8bd700e1d7e2d6f951ca2df7043a03688620d2a10dc8e9bf9ae46d3987f76121957eda1769d0fe1ba1f568c3a8904260234171e5ae634eddf3e805be318f5108f764641e5d78;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hea4352a42dc9d997bf8e4c2f57c9f63a55d38213620a32fedcd064857b1242965e55438d5434a57014173da0c64f4d47c65bf9c249b12d788acef14d7ed1a7cb0af0154dbea0bcae52df46f10170fa5301393e8fb13a31af642c2e172486e0bae50f5e2d8a0cc4785f8c5b2398d217d2ee17f49f296e84bff64202df45ff646888d1e680907c59b8dbd7ec62f653a7151c3520ab0e75bc2a6aad405de85b57cd861cac4d88c26dff5e6dd998a1776a74897315eb0b264022e6157d55bf9993c0dcacfe0864a0975438b73c900ab4d67236395611d6091ccf666f004adc521db32ba2776c5575be2b5851a97dd2cdbb619b0429906fdb98a98250db89e5315124edab50d51d1f7308b3d407c0badda3b2963709848f1aff15a3cc6214ac4cf1df886a37f87947fc96ee80182f68344c354f17d3a3ff7d3540b9964047013122b9ee9b1886dcb642f70aa4aed51cecf55dea46f82463f75909ec0adfab1dd0609b1b0b314dc467bc4a96695447bce96103f5833b40c7d79226fd0cf4153e9261c39b83465df1980787dfcbb9f12f08f5a9385579876c6ef3f42ac0134884fde262691e0479ae4ae7d2171ba958930f482fe52e04864fb8e4b468e1c3516af95ce2e1f94abee450b378443f7efc34fd061cf4aae540299ee7fcdc30a8e526757f1d251c91e5b856cc961d3c6a48d8fe989369b26933440a461b11531ca7abbbe7dbadd4f88c346736f6288ccd17cd1fce37e5351a6a34a063ee905369ce8e618a945714dd1994ec8cb0b97b1dd19ec49bba5457aea709e8d4b84af89ad7f59b4743972a159571f7f35afe7c954df06a681e4f8f84ede0b64e634d0ac2988d873503675101f33d2005f5d0c7029584db8ed4d6b2c476de4609f9375d045c7c713d8cdf97cd9e798ab43717167e020d6c218f6b8ecd97ec41079772a102564f980c2ce7ad86043625cd93080153ce70908c4649c159072fe8b0c4b6442292fd8ab67e10b82510bfd6b3314449ba5809f8baaec88d004c48cb8f596b4e0d187c0ed17cdd9118fd38238f2497ab4c2c41e78ad618234424e8ea80cb9f6d177240f68391f66163a9c14f13113e96289e69f0fc9a91fe49a1af0074cbda38b0a45028fd0bd60c220a0ebfa8b10fd44a39b49a85f632511ef015be6d88fba71f3cf8d6639bfbfa3d4c182d74adafe8922fe0758a531f492f05a1c2557f147dae077266d608b01ea325cdba2d8a2d288e7c9c763f9218f6416029cd27213cf1b4bcb961a2d0436472c3d0d9cfbfae951891119a06c2dc048adb29d0ad29200f8d8d2df9a34f14fdd5b820b3c8e37580a56441db8eaeaa0ef0091458bac63e55f2ea4345c71cc4420d1fdec360b15f1c92c823e7490b3c0a6239430c4427afcbda312e6b33e36d321936756c524516473d3890f7c3573863867f39bd9e155f728e822d66eff4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hac12768fefdd4ebc293093bc575bf36c592bc885e03de4e07bf803f65e759c8a295e9f9990d52bbf0e6bc083a8281be8740d8fb4e7631ccfb3a2e263aad129d4835e98b2341589c2b0995ee9b0b46ed6d277268f2f44fa04a37e25f2e14fc51664a04c487c0607c7ca331c00b38f9f55c26bfefc577edcb3e1fc5b28cfe9a1eb0cb5a06b43853be857d63395ed6eb4e13e36e2e8835334679d4fc98094d1bd469a4936ed2ba90179e4c85a104333825148037f8dbadb991ddc9a03901ea1e562bba846763b4b2bf2e0533a152160cc070480f80d361c01b673543236bcb72128c86644d65ce625f22338fad4f671b6c2e99c4727cf9acd053b2a9523ddd1c6172fdeb1c11b51e9d1f38893dcfafed6e26950da42028a8e823aa2132db319e0defe1d93967a2b806a3015332346fd27d1ca832f125555eff5d8d567aa74a80b4efc4d13f8275fe7138c851f5d4f08770cc17336a457b36c57c7fc35060c2cc2fa83d16a2a8100d3f62ca61a806245c0d36e9e1c34a204f3b6504664905b6c81ee8ec86326f5235bd41e8a9f512aeefa8487779a22e09d35ddda1e28f75406052e868cf7615d4bb4cd5ca1695535368f4c65f28cd892ae261be5225daf3be3f6a6f35d8ea0610a72667f32f3162a067a6b575d9e7980e152dce22f881b6a8676d93ca3b95eeb80fb9dfa378622a9804f15450103f241e69e966dbec0401193af5915f357f00341c6808569c9a53f989d7a3e77354f8a1d9e275bd31933405d0cd24f1ea80c786f2ca5b4aaca0df94b3af1d0181c3f5472cba57bf864fa83536f576bc7803ba4081a32e2ff2a635cfb8889ec34b9210a8aabe2bfe8171c1068bd9150ec07461bc9632fe81ac112a5e6630c29a4c6e833c3ce6ef489cd48def127d51beefcfe6fd8a1db25705fa7d4fbc89e0903471cd4ee987680b79eeaa080c3089d5718d489b0aeeeeeb02acbece2684b1278e7a0bdc8e01e11d5973a25071e315bbfb7fdf9b7fe042a1942ea24ccc81898f5713cf446f2695b8b4e3ded44bea0b243b3b83fd46a71bab6c118d3abab8ffaed2a8fa1327c69b45c7bda4cb68bbe1caae8086e83ad235a95b4400bee6b10b6fcd0fe2e9a3fad83326a1ddc0b2969aa7c3a9324d5cff40185e6a6e69ddb932c657860cfae05d4f68e6d7bd4ee52bb2cd9552c2f0231bde65243292dcfa1c1425e1261793bcf3decd0ec97055ac3fbd994c1531ccd639698e63dc68ba5c9b861c3b79a02752834eaae2e2298186b15ec4a9e3bb25696304d1005aa9ca341fa15150bd026b389691ae343fa6e0d7457db6b9b93e0176ba91ca7e2da5c54de4cd10a963443c8d2e570be64d4f78428b508c9743177e594fa71341ed459ab5b486d3e0906b8f1a33013290e0b12d537d7c4468f600f6e97a3bef079f1670eb1a83a5cb7ec2cdf1263e3783dde9d0172b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h65f78a756b1f42de11d9d1f636cb717d168f1158e75c1faed840ca04729c3fa3f7ccb24b4fef2f308c5778b092eb3711d867d3a7b7810a4271a486daf1f504525faca544e3a8d11316dc35b1549b68306c4d8817b4cafc33f98f2eb3f817950c743680e76fa0ba7e43ed8c33b242d09289d71515ec296b40069df7a0d1b72536b584ef7010824ba73c6d4586d2ea10f3577743cf5b8a29552f6d605ed3fbb173ace9c2849ff6df3b7f0e1ec53f0f5a4e8782323c4b03a3f21a7ec4c2841f7ce40e387675487894e0e27b9fc4536924f29e044ac6f2a07887e72348c2307c2263f7788cd150a0156199dd97742d74914f2c928cfede1fa9b8389dfdd030bd2a147845286e388933909acb1f10204a41be76a0595080973d726734b493372173e504c0012e60e304c9edeb0c08d4a28446e72a84eab69f0a0eda909aaf24c3840611a847535e699698406ac9e1f4bd670f5aa42c22b5bf897eeedf078b5f69b33702f2bde3de0df748faa25728d4bc80482b0dd46c1d8f76afe005e25fe0ef9245433b470a748030d71a4754995d8bf41b474a49cd83eae548a6d1984b30e8137174a8a80235edaa99a52e55f1d72f153365b37e810051196bb1950d0985a99940682de45e80f52c7ae74e0c2646c288cf93829d9d746b08712532be895e5cce4c4b73259b7a0cb0cfd9cb1cf0c3b4d7100dc6825714101a7a5e2c793aa1e603204d27751b2c3cad06e65bed86a2f8cfca17ffd04f6366fef8aa9b201d7988e7a00c91bb62ac9cd44e9cc6c7a069f30571facb385a7d6a73102741c5dbd857748b6b802287fd58569325e82c8b2d6e8925c3bcba76143c8b96d722867134ce2a230f3934a45697d282aa720099785a0c8c4c141a7795b97bd943dfd3c77b559d09ef6f3a5971c45b5bef40b0b3105e97b578f59eef59589865cb1adb968600cd0170e13e6fd800ce15d715fc836691db8d28ef348bf5dc262c7854c47e177a29900e499bbd5d5d045e21cff934b2874a0337497edb5e08ca39c6ba1c928b6f122c94510d0b091a53ebce0cb76077e98cf1761f09d6bf497e21f5b6e269ca84ac977f7d8ad6455b4b927cedb61b82b0fe6be58f31dda04dae956d65662a9b4a1b5ed19cd8bfcd73ddd6cdcdf507eb9b78669ce591b0f86bbd8bac10d22607403a23ac63d234dfdd9241fcbaabdcc1b69d0ffbc797d591bbeefe81ab2a39fc36943f3c27e7508a565e3640435267b5d59a7f06f4114bcc1f3266af4480fe1441406d2b7b56da1d9acbf503a96469355fb1728dda3ad2172fb32c1217f12afa84766c59220e4148fbd63228ac88d3344a65ee2362f6ee804de0f6d63742f7a70b68b4835450342ed73a190a76a394f4b2150664e7607934a6b6f586fabc5d139553d697b9da7511216369df4bb1c12b0591c8a3f88e4c38fe0771d6c798ddace3085d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h725d49657390edae189593688d024b5d9742b61bb4eee6ac4cafd5813e1560a7e14052e86dc4bee766d895a0f7c015a8c7758cde7ffa86f166bf938ca69618dca9e5e58cc7cd5f644e89c72695d6358bba06e3b894f8b6a24815cb577e16f259733f18dd78f9094c03243036c374fada7cb9f29be00158f5ac71e23e721d28a38a0b4b202af88f6613a4320d1e201fb101262f2d1d5d29255df12217422f8eeadad70356e2542a79d2368558fe68e393476929713bf7d320c9d0856df4300366dc05c3c69b3b0c886d0cb69a61a18ca8005addf0942204d3d2af7625d3bf6adca5963b8a7a5f9cd191f9700dc80ca79e1202911ae46b39353789a763a4720fc05df348a2e825b460bf3e81e46696b65122c8ecd5cedace08781bdad2865f1b4249d41c9ad4afe8a0092ffaed2a38bbe49c733916f7b13ded1274581173a3ea6ac36232d8bdf68cbc737d3ac2c4c2d2091ec790e9d6e0ff10502ad187fb7570ea4e452eefa24bb068489e286e9de9d077e9ddaf931f108a66c74011f21e9495c60856d37eca5c7871974f02521ef95fda1e545925a89aba90d435d4cfa5e28d816be8039f2f838cafd4d768fa86f153e09587d0f9367045ca86e11eb5a3eec247e306e5ffadde6c1e2d8f7e161a194fca72f176469ecf4fd2c7544d41420dde6b501be69a446de07cc79604149b2dce174d6def71fc626f63b9432853f170ce4e44df2a74cd6262bf1f7277c7b4ba9664ddb4ea35b7b23d229d0998dc3ceca4ad214520c04d9f14e4f349ec92dc4a845fae5be7de0d9c1f903cc2e71b0eea2c47c45a1cf3a6e238cb1f9f873ba86506c83ebc5b1c2b99570b1af48ee73beb4328a2fd1f14b9c50eee03ce81b668ba6b6b00d6a9334d6740195d57845ac24693247ec6dc9f02a2a990b05a5e2d4fa90554fabb00e5763e85e35040478beb2867e6a566020c167b52330eaa1b2c3f4bf735d010d414f2c2f820f6046798a16447fda57f6d201329a6134c3f59bb9dfe3697efb919256a38c0e2092f44c36157dccbc2bd0eaa7702be8ed5f4c320a2506343f169afacbd0ec329a862a37aa1a40cd09878c51ef8d4aafe777f77073436e860034bc430836a59e4135e1f6feb8ef1f81cbb4a9e2370ab8a9ad70f3845c59a104639c06783ccf4a995620b600a82bbca4e9299fa838ec3c91ec7bbaf4c03c3727905913b702055a448b2d8659760317e3d6f2610eb1a1c05ebe6556774e2df860b9ce3a501703952755d963c5495e8cc6cfb3a94fb57b225f3a6e1ae72b56d69c95b0aaaeabcae3eab3b88b935f4fc1c5c734e782fae2977916b6a86a4a5b1e4cdd49c41b6a89991a4a8eb11c3c71e9d627ae119a7708d416d0bf6613735454e1c7a87d8137364fda4919e7398b74d19dbf69e2041c332d1c06d5b1fc92c6d0981cd6bd51aa23a36f8c0ecdddddddd36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7a72b734c0b81362b85c005b4407c2f2410c37170ff63b1412342786b8b1d14c5fb2dde93440f7317bc429b3779562e30c91abba4288a00093f284189a7266e9ce51816435e26ca3b62213b380d7bbdb3793f994e9f447ffd0693e4def87222752a26e20580c018d4cfab181dc0fb4ea0cd4c2f8dcfc7c44659fcab28c37f2423fc70fd3223201c1abb1b95ee6deb1cf08bfbb17aad2a9f082adfc64e0fa5a4e7841c456b88aba4762a00f3657955cd2bf9d1801a275dcdfb1c8be4885a56d4daac1ea03d4ddc3c44df2ff99954bbd9a750968c2e9f6b3cfc2028d50bf336c1b01649806f3ba2076d83b2c4164f34dfc8758cec72a2a0b1da354447090f23ffa7674d5283bd6f546562ec67df02176e0f09b39e60cb59d1e852f9d88370db99e392ce21651e7aa8930281872517e7b8432c77ba8073f666824f1527f28c47ad402acde065bbbcb2b5c56304ccc51fa97974a9797e9528c17f224705293fb6131c2ec28b3c92499f9d4cedabddeb818c856abfd0c2ae68e20d3dfcd843fb68b10e2c3aca8b025077d9c3d91bcd6a1d5c82ec5374364f70866c21808c32a6c4fa58d7ed895a2a3ef4db4cdbe634e9e83353f1701b57b98c49584032f273d6bd22861414bea468604d6e2d0b049755b7b77a20052292388ae660c99c34feb5be89d90b76530ec3029df993e421302320e34ebc489eefd3bce23b08b7afe3b7b3cea10a7cc486f4026d8d70d8b2b1982b4eeafdf217de7faffed25831fbdd9d91bdf5596858f2baf54d64d837b9abd023140377d07855b938370ecf2384c23b238f019791fc50ad4199531971e2d4feac8e4bd900f3d200c4ea7ecff43630bfb5c3e543db643ba97e90568729d3caa2d2a721b24fe5f576d696c324fd3425d6052e3cf8cdca72f959eb70db74ae5e88c4a73a89ec52e11b9520d8df5c726229a2167ced1be3f668fa22eb7bf88869c258e3a3f03d19efdf0f08352291242703173fe9463b33d8329b4be1e045cb85109608bad85333a2ccef5ab69f48dd8032802311736fe488607d796295357d0b98c2bec4ff3cce5e5e90265e688bb8f399c4cd9b4b9f6b244c493963f2165ede05c83037220292ec04113c39b205ff91e501564b1e3739d6fcd3d8a98593e03b9fbe0d0f0c95f6c1abbcca7d4e1c90615f5ee2ddb3d9e5fb706def612a2825806a5b1512350e8a3c06d06dc5abd09b2ad1310951d173a2d4acca20f9f0b62523e9d759bc3d869529a7b901f64d6e845b76cb82711dfad7697d91b0f6679abb960e4ea1c9611a6a9884dbc40c0584d9bf1abef65d670d4dde831926c68d158c393eeeede5a73c682efd4723a5a69c804703e091f32858361dcfafbe32aefa82757b894fdbf19ea2426d883628843771688ec5c4df4138e1c83d3ec13c12e817f5bc985d0a429b0f5eb3b6c56778a2e953ce3fafd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3d7d7e3197a23fb608b3d6e1abdafac6e91d2d31448c9b4903990c008388bd15e26dab923ceb93802bc6e865bc513f54f91ef13bb530e24bcab4d03e9e246d1998ab3cfeb3dcf0312253db810c9514b0a8860443bd56add1a72800436efc4f706c98d18c6edbfb289c81b9c5ffd16e4b5e895b4a6475263221e68937192fd323186aeea46a1b40e920d665df8c7854453f915896917cfb1889ae6a466a62c6207aa40b14a58106cb5615ba3bc701873effe2dfda242c789c3412235f0d627780c19e22b5d885058801a23dcbcef1b3604301d7427e6e13805e941ebba58b910942d932767bcc255e31c47f63064fff4be784ddeb1a91fa28b3b1c97d140e78460054d5ef4cda92029cb9158d36a811115e3d0e6cc44adb38dc069db35c3e02cfb7189b27ef3524f75df3e7554b3058cc2ba098f5eb7a3894c09e80bf403c5287bc10781d3e988b5ff9f755e1756d70208eb711912bb51d1f174943322ad7ccdc31596706b275ccc88379ce8207d9cab97a1ea340303ac24e94338500f3d277f3a32b50d8a21679716fa7cf555b840d34fc18bad0658976b085d139903e94ff21aa13732aa98d10dcfd066b8b10cd52b8c79c6905984fd1f06d188934e905c7a5a2ad52f5351aacf9a285e91932d742a3fd8e5c8990cb7e9e22000c2317a1da6ff69c9c21b7473b052979e2086d446a7aa22230fc553bd694d10da834eee80a54708a09052d0673b558ada4efa819065ee43a830c650bc22da801a002e2478e97f7f436fd8634ca3db54c0ef0d5ecae2694dd6749b34e05234312e916489c1e4ab3769fef2eb5c8f330536694343526538cca934d9711e4279551f74344c7ddc8347f1896c591d1b904ff26c32876e171e685e13a8a481cb4675ee9e5d0ff03c6f0be0b040d48260b9ede87ecfc7307ad0590efd3f8db5bdb39a4ef00553632b2b305a56006d6f0fc99aaf16d54763cb8ffb48dfb67a8c81b65703e7126cf35c973c6eced7cbb010ba600dbb12f18194916d503a724d466d3d11f927680cdf5b9afde4c58d768221643f9a67922258e59c964ece789b9f21d614992420d6a3fefe5e931d8f1e95fdc5609f50c5f7715af8c027836f41c479e64cf59000dcec132fe82c6a782b8f02360dd40d907b2e90fb6b925950d17e743c2fa514c7963bd4972c96b2133b60f9d52319f63317760a40bfe52c64773d4b0855af286b38862aa8720365944e44b86ecc7995410ee67274e3f207f081b24cd154b1b98756a7867d732d2e6a64112d590a3104a291a4a83d45604c47c5446cf533932a8d372785e59518e8d8a110e8dd401f4431717cff57df14dc547c22c10214611167849501d255f80e8862d027677e8a1ff6d56157cbfad50ecac0050d524bf26924c51990cff2ba183e700c8250787bacb562f338f1e085d53d43f4ee8a55de8e04fae9c02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdf53c3c28c289ba8f8d10d4d3cf2000b9bb9f2783e50d9fbe354a397c3117c86125c4a764462716824205a3131f9224f2e6a95d21fd93dd5c6dabb2e2a0132d4017535b90718f102c633703e65a5859e6e5cb21b2f289dccac0bd8536bbf2be2f9ea57a249aa07ffa800fceb1edf65dd3f30d8ef0c4f40037266d4d6501f4758baef379b5caa95579221749dcc22b86d1f5d5856218483887cfd16c6e0fcf2300392e795d998b0dd01ea7e5955cc158d79df92ade5d47625bbf53720486da75d919af454cf8d5f1bbf6d8c279fd012e8f4de25db4aeb6003a37f42b0db5fb95a4640f3e8da4b569ec09dbe64ff439113fb229d0b17f95107ebe0c924ed0f3f09aa81146067f7214c3458c6dd1a02aa149ea13afce81bd788c29305ac6f08f06c01401e3fe4a35c987ac628feb3a317ffd11cc849e52bb38d210b4aed264e32382ff29f7af7be8d885694b11f0094e9b6cb570c049fe4d42d78628eb5b4060f014956231192f4114ed8faafdf987d91893e433671c66804add8edd816ddc18edb799d71ef5c656675c61a1b592fe9bcdea34fcaf217d1dbcca86ea19c2d1e6e3ed38da783c392b5502922cdfc674b38091a3c77c5849fa479e9e38b1aaa2727fb70d881877efdf1c69410ee1e35791272527c177e4cab0c2c9323769885c916939b4b7a841206840cd08fad465504cc2b7bef66db838bd59866e4d20f81f4bf0c4a3d197de52d8b03060f39ad060c376dedf27016e2a0c062199d53b962e466343fb03cf32d8b1502ddeb33b0a2a586c45347072d427644a3a24bdf45648869c9cf6f07637c1b112f7c491033577bee8e2136dad2a786f48de893fcfe921925768c36856ef97bf4ca424b0debb6a57da56a9abfed1dd8ee5dd1030bb3256626403f9c3576015a7dfcfc5b3dae66ca00027a105352334cc830cc25f13d9f8d2e1c0ac09ed17fe5fe9e7cd61756690f0f5ee4450a53c3366a0a7d0c0d2881df46e7af1dd22925384d277b1870b65f7cac53dccca5c212c376ccea946e8f2f2502d52d4c486e99a30a01718e66efbf29d11e61dab279a88bf4c18540439a860d3c8e85b74184029e559577fbbd92b7805336958d09b8c38fdc5cec8b7d6f00259eb75a0d36148170f7522fde5e44835fdae187d33bdf1a907e3cbb499666e8d126302d9dd188c4e626c3722f2ddfa5b27a533d2684e12fa2fa70203d753ac2accd0ac14f2d14e5c113fff988c2c08ec01e182591708b583b9e6ba2180a748556c1672da305df9678689c935226365a3b94e0b6c0c0aba8589e9dc46443c8baf1e7353581829ab8e817f3e3a1e896b605327f43027a21323424fecf79f9e538742e3f8a1af90e9c30fdc14e08efa53cbb7aee63e91bc5d63e154a41ae3a863e70a76a28f8a113c29694916edfa272f58cc0cca25f2dca7c5dc636912f03a1d42cfbf0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h18f4b6ef5f845cb27eb61fbc75e91eca23a9236c3228f1e15eb9841fb0f71e6ac752cecac06631a6b613b6319de4b41eca979ff63c6a22a7733c910eb4d225414b0efcd10a3ffa4ba52a5f9d909c9f06c46f6ecf2412929575e79835349ee702c68b9a77f29ed454032f7a51b48ce7300036681cbd738b048a9169edf23bc95614aff087366d610aed6f3d11766ecd42b88ade8dfea5c6cccbfeda2fc5e18ca3840d71be08c5b0632ba9eae23acabb10173caeca53ca48136a4a0a75df9fc0fa4cf45f2a432d1de6ce6d049b4d94a4c2faa4a3edd23f4562c5e8b260d750fccd5b00b296118adc9e63bbd63f6ee327feb8658ac290b6c6de6b272fc11084d4b470a6d6b8eb185dc2588c2cbb49ade0d7b1b77cdfdc8ef4cf8041dcbe0789753f2ed903c4cfc0b5db50a13faea490b3934a99483eeaaae699be39fb0de7de5391459547346101470c1ea364940fe765e994297e6f1727387f02720ad310b48eafb2418b827d2c2742822d9512aa336b1ecc97c5c4815f0f5e62f71a7d2acb2b4df863e5bf952ce91173bfc0260fea2af5902e813f0d858b9a9895115a65933cde1ac6a3ee661d2f8735d4d25b816b1bc1d598c0f8e9c9f637a6acbe842055c53ee43716b967626d7f60d6aa8cc4bcf50dc3065e39820c19d2bb13e67ab2d7ae19363c03f9019c4b217ae19f248a48df202a9fd9d7d7078782d3d47589323ba718e5d54ccd4c735e950c2af2766c0e1fcdcfc5157c6ef018943ab65afdb98abcdeb72456b7838550e3748d279427bc30d55d0e44b31be4ade6a005c41004da8db3e176a21c2e3c446ba57a8533b9451729d4b370d493d352ae9ee74b0455b6b515cf27d7b1bd08fb6ab1468e9d22a9a12618c05afd6290575f42238fe51733ee2293538061b619a9a93da191088e06e91fefa90f152d7d97f1b7aeeb7f2301db239d4e585bc9e4999d46fb179bcc50f2692260668dee2c93659e6f7382f5b9c8d537a68fee18a015591dc70845392fed75b350cd0383bdf85aefe2ed9a3e5946f3d37b0a365d0d67ab28b6f45c1cfc099c4b8b125d25bea63049f2f24fcf5d39a33cea6f5c2dae5dc4c434f284397c8cf7318f773884418aa4dee9bbda5a574c84cba646418bcba5ae0d6cea98fc43b51946517f39b4c9592d85eaeba6ccc07f6b01e827c29d4988a0d0004fff13093e0804b61791da34b3061fc5d63d0b9d37429b32249a556c7cd7b7659b71a53c96298a03ab1af623aa46110c4565b648454eb5cd50adb47bb131902cf335f25e1b6a2502176b7dfc101ee8833b08a56e1ce8f4c1341f760e48a4ce768d33ba5bcac2956b99cde840b75cdf9e1f2b5315f8903e9697eada5b5a2bc3b78c88bf3767e2b7950833e179a8384bf450a5f2d9aa461241dfdf1e0f7571e8bdad3f3591ea546eaaf97fed6e7fc778967d30a7e60391;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc9b87894e5d8356943cbe047687f73c49321d6e8a8060c4fa4f6e3322e04747f1ba6cb7c17b61fb87a52ae35e54795ee2198602f4db18303f9289bc6288bd6e860d11bddc47d439bee1cb2f80e1cb5113f116831f916e32dd0b589c1caa1e535d2608ba328c9116129ed4727253a42258a296cba47e4f3a9b0bf9b62cf6bd812bf482f4cc7c806517b4586de719217ef67220bcce42fc264fa5a851b9f8949839dcb354db309301d7346dc6c339f53758a1db74403b9eafba7411e46e38138d430c137d57e8cb2177200548430d2a809d122f55b5506f8d53b0fb95735b9ab0ec22d19c2fb062b31d50c0da747f7563c41b995f001b490ed815169d9402da11b005e1dcfb3d3370c7bd94ca68018b1c03f5ccfe904942bc608ff916e0521873cc4b77a663001d2cd66b92c17029fb9666cd68fc1a15c7b4d04df7fbf9187f973875df535d62973caf3ac56e8ddf7c920e7400457956aa2d7d97b768fe87d52a9b331e3a161d092a76a2e415d893c5749f418284bdad9a1e8ccd3ff75394050119bc804e9074d6771d1348d90d1e731e6142dae09e982b5886b9e3c93e970a89cd356f33d4d29c9abcf968caa2d20c2c82b7aefbdbd070c05f69483d1451322756f85dc784c8af5654f0f339237b5c42e2921519a710121ada328bf01adae4d06915b510e9ccfe56050f5df08f3423a4f8bb74daedc1ca2959d57540432ce2967e327d13757dce591a27493c3a2449875c2252addbf3f0ea24936f69278d36847b253dcfad0398974f1644371754b2b1e9d8fdf6c1e9fe62f5f12768eae91b0d8fdfba63595f765123a03881f4aaf043362d0fac8eb99cc9b3d48e4d850ade07f4bef89e55c09b847e157f604114ad5f986c85ffe2a0158677e56fab8710e3fdbc7b59fb5022f64dd16a1972080607f535b3da16d00900eb34e4e71fd51876291d62fefb3b4415ea947301a9d7c3d989f92c95d0696a2e6a73c2ee6ff9f1414dd341d7772a46920a39af4e3eb7b86619db5128569cac13bff6cada750f0a2d4f2cad27ff8b7f64c8c099886176f1ac5b349d157a8ecbb9f5d66f37f915682ac70f60f844712f2bd8a9b74cb8cc2bdf26b6b97b8e803e95965a4e5facfc1961146cdb0d5764e06b2a90883358be408176ac2ecdcd7a99abb929d9a5280e2c3ec60109e0a329170a417b7adc0d2bbf264ece9984364030cd9bef70d360e0f9b0044347efd8d8632b868c14aea697e71ac94eb9639682f370a2817584f5799a8888e0f5e6a90eab5b9ef60f3cbf0fc84c180cfc9d45118e6e8920227dfb51b4064ccec6159f3c2bcb64cc57ecbad67427ccf2c5f5d201849d9398217138dfa2a2f33aa8b95ed8c606e89df742a7ed89e27b9cc2935023f210e92d647e221062e2fdcab6a4522ecea6740bcf7a2a428b70656d7eae56c5d83852fbf46899c1cad8a60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf5965bd2f899ac1767c13d6c73020daa32e8a8838deae17037b6f8ecdd57c8794f18428a5dbf0312573e639df7675063e49e7d1c2b85949a0f06692f9d878478da0358e26756d6e732ef4f657bfae650f534daaade25aa17f20d7869d7ab1b10f26f171e37c300e548937f2ff0c91d64bd34e83963466c8dc9bffdc1d86cbab58fd93645a253930712cfb191fc98b1411fcb930f129dc166300a012beedc2a5748f8d87bb78b3a438fef078ebe9e51f43494cabd34b9b1824f96a5ca922e692909bd256407b6018d9243cf1202a5d792b05faf65e3cced1756a4ea5d8e78bf72c6974e6781fff81773f1e3fd60d985e2ccc17dc6b8876fbb34451071a360d8781d00f2b8fc21bacfb4aa8933c4927fc16689029e25edad80bfa181c86263f425c818c6e87609e4e842ad8dd316219da031786ef5a57c6a13bed51bc18cac0300c1205a23dccfcfd7ac837209b13d3d21ab29bfc937b38a08da8376bd100fd89ec4a4645e71a9859b9283fd3f52504309478e1b8970c98903545238c10ec0a65e6af0d72324fd1dde69e51de3ab5c7fe85b9afb8735c93e705d49f1fc1a782b443be33944377c2df8d63172ea22084f336bd5e4f2c62d1fcd093705d5e1fede7249f3175160208f4612dced1702749936af2a5985d0167aac162c5111738bb1e4525de5f81afdbb2d75d48b68ec75945d3e8255fbed37c6927cc70f49c23f8da6dd379936299b2a9feb8052887d3aed415c048a6bcc1046b61f064dfe5b09fe01dfdc8c42385127f11e02159b60d3725e02e8ee7ed2698823c9714a5dff4abdbfad150c5acaec7afb2d585db06100f6fad22d9c1f5675bae355e7ea5573a6898307a6912a3a5a6f423f5046e36f0447e4cc2a69ae67a48197e3254ddf56ee00264c7a5595dfce135331991df881db69b13527b86f7e8610c36a5148bf46d38169609d3bc4214e2f259dbbc44d5349420bf1ac46a4d877a991b5ab8d3fcd4f0586cd9c5d6bc14f14b4a182618166839ab8f2e9447efd0e30296e1b6de549b510f47bb5a71d261d66402946af530e705fbc36fb0a43c2394040176bf6401e971c2cbc6252702d425226ceddc76380d273d91d2ea758cb3d0c820a596abafb17ea6864b96882115f389c9e84c8e28bef7419d17d74f9a4b5784f517e8e81dd8dc8c9228a629e178e34d35d9d725d060127eaf109989dd8dd0e9cda00c2f95a583383c31918db1240c2ddc43a78ffa42f8ed95d53cf44c09b4108de6f8cb2e92b5058b30b976101558609fd099cca30ce68aff32959e52e1e7407fda6d4d9e73f7b2c8992603b8490beb43d72fb0cac0012a4c4f1ec9e8cccbd37d8a19460a49ccc7631e837cf89fb8f80b57c3bfe0cef51f1983641c89625d61cb33402bfa3bf298ced8d8343e4649b5d86f74808cc808478f30c0ffebb5cf2cb669b8d8627ae761e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1f36546c506ad944b19ff86480a1f7f7965d97f88b9b1ef71cb59efe281351354ce5c25d9b1e2bd872e2a41f11dc876e4b7ce87deaa75808dedf9911fc92e7c282cee4e7c605c585a03a6bdb0489c2aa41c91f9717a1b9be917049c6d0f49258265c83bb642e830b958af8576e6658fce8f8e2780375b8baf5b04285201a2e5318ab0be552867716cb8883b4355764c31cf8f7cfc7335b5ef6474010d57807af089d94c94b7e6b1c8c54c4f9109f871feaf0a877b8ab60e6148ed9ac5d738e8ccdd752989558505270b45453cc879ba9f758ccd20b7f9c9c4fb6804bf0cd54c9c69ecd345ab53e32cd9033269699f28dbdd88ddce71f3a29749e16536e619339c42fab4a518d8f666c192c9350d1ced819bd73dcd29130575da5f780bfdeda6a72273de4e2c7787d70cf553392d92176d4039d5477f53ba16dbcce12e037d082157a1e92303f1ab920b9f3a28fdf57b49bf4f66f6ff1bf9b226c17ad945c583fcc410833aa47d78e2b2e06a63708f41bb701c45757a7ad8888f7d1e07dd7113b97471c91056be947c19c6287c3012e159a780fb437239922280385ee2077531ced0f28a3fdf86741a0d8a52b8bda752be79e1ef06b4760aec1299258d14a9137f11c66cac242280bb3eea6d4c3ab3bffb24f551d791187ae84b0206cf3ac3b5a42e0ac9693760b124381aca53b52ecc7e6c73dfcb8fe7fafc95e032fbb8ca5249929ad1c84456684f7943081f7481b298ac28960a601affbe09b2d4501b9fb0bdeddd58e83c4e184c2c71c0f1003b1e6e62b8a47a2696962c3d5bfc286a7b4506c7f8b60d9ade3b5cb4e541c2b7a37e2e2d1d6670ca6020682c5a6e85baad68d2a0c10be7fd4f49f8543c6baf64b4eb3a34f44c03053a644f202ec5f7fb348c855e5b8e05549ac89115566fc092fb7653a118dc32d77303c3a9ca493d8635df3d3a806bc240f5a0d2ed599665c4edd1cf9a767ad48b5e488f49a0a86a3318e74a29392df1c9317e85d7b508249afbea98ed40614f12eea59cf3d691fb1bf151654cac2f3a565fc1aa2371e7c22b0a2a390167b72a76c77b77f946db372817e789d41e3f2698253abe33d2a7bef50936ff6f76c119b740132ee81d653fc17f6f05ec76e9a5481e60139a9480be4b0cd816168426cb86484210b706100f65ee6a180792f68db267f1bbb3d72fa7b94a50f404869986ca6f72d61ab48ab22b73d50e4884e714fadd940dadd5b57b3c2ffb7590f75a9c0f70da35e4ce453b8de08298d8225c61d16fbe451a1dacc00fc00749cdad8ed0fc185b553c928fb8d2c8b03c068c592fcc5a2f710d882a999c30d496cfbcda5de5bcd7b1a9304ca92cbb11080782cf11cc72e37bf1deeccaf1591f79c7d926e2e9ffea62fec238e86a0a2714aec57904893f230e90b5f5b54a71c15fe6aad4585c3cdad6d87489e13fb110a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6979cee2c81d7ea3220ffd381833e726513eb903d17198373e097ebe87d26b02a0c833b74e89584c710aa4e112159e9f6c3bda64a606ca2c92c0625f1e200403d1fe3f5be5f434c2228ec3a0b9fc5f8e283d7f91037c37c74df6487bb2617d5e43cffc6664eadeba6f912b53d47fa97c2263b9998ecd613b6bb19356d59c0e38dab00228340077fc8352e9f85c67f5af4cec8de20ae119899f4c02b7acabca7b7b4c637149b63c9bf010c99500d4f38298e84149b9f900feb3952d8900d27b6697c42740da17daf595e04d469fb349af984407c985c38ba821f067ee6824df55414d0b759a3eb3556263872c75748cbc6ba5615243586ce0d6fcfc59355a533fe858269238cb0bf6bb4c253761d2000bfca8c0c21c7e35f51523a8556e45d9d62a5c52ce2788dcb57ae73b610283351cbc45f4173984b093ca938b522bad57359e62d69ced8e7ddda553123f45c66fe5b1975faa7256efbfcc56c8174283625b069d3eb11010d9d62b3400c53781b22ad8b53e9e3ed675d62bdb2608fc071250665751a1135d6caee23d70b19729ed6438c0602cc50727b06ee005df4d4a2db5f4bd8a4999695fa58370691edc58897dc4aaeeb2b1e982ad71d5fbf7aead91bffdf76ccf154ee2b9d9f52c7e80de97cb1f88b0a79fea7f88739fce7cfcf9cd25c951909d7214c30fc02619851f01866ac6a301898b47110d2f2debd29abebdd8473e6390e540eeea6f17827ce1963b262c5e76b013ab0aa994317f59e7ed60ffa8476b04657bab285c17b9ad8e24857648a0d12b6c8b7be689131b7bcabd12bb7fb404984f5446f5acdda92a710e919e77138d4df6f6cb3b1e3333ffd0dd8cad4087bdd9318dfccd65b4d019f8ac7ec94d2bf9544bc2853d97477ae7d53a02f7170aab57b6fd7cd46ccb732d7123869f9513e7c250b1676d8fa8f337f6c157475a5a92406194782ef1f8ff497dba9ff95e7c4bdab13d5301b7887751a643d6ec81bdaf4917f94a55c816e6b21f1af258260863b813ebffed2bcd1ef850412c5e73c20345e9918cd23454cba603c97190c06cce4e7b5a5a82c5318cbfe2dd8787d1ef9401447ecfd7ed1d295e0dbe50fd6ac3347a3392a2e15fde10a6026bbfd84d5e58c1729cd9a1e92d167e8188898d48dd27912bbc663c286e7729a279a8a0b96c6bc7df6196945bc8a2c42b9f1fc945300200e9c02591ff6d27f01288ceb391563a50e38c69702519bd0b189dbfa1e868685caef334bdb6365f4530818d549406ea7da0635d126c2b547b6407c2a138f0d54d5706eeeaaefeada56d38ff4456570ef7beef470915379b2371c01f3dd52b2b31943fa7c8535f4e9900963c68b4c19e6327fb5b4c3cf485052d2fae3192c7290d1fa1a869cb4a20702b15b975f2fa32df600019ae1102344db5ff1166d965f3ba8983f92daf1f925a653516d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hccf3c6dfae78c83e11b8d65f27eb13cc99b05b7bf71305d45b5741a074713ca67626328daf5ffcbd8ea6017253e83cf147ec1345c8b0167b66b9cc578c7b81de7d7a555a1a03eddd1a4b35f8635f2eee5c9f829c61445d147a814334132b86896b5c1e17bd2da1d24aa74183fcd839a2e96d2856ecfd5a9ec6c530d533b26ed3ff6ce632e2e05f0c52d532f83c7b9d02f8e66b8e9ebcc4cbd76a06dc56010a7aed8fc9f37cb92aa4796fd4c1312087e93674920b9fbc862ecef7d762e6cecffbaac4c557f3e34053d0c9e46417d7efd842d78993c165f11964c653111137285fb2f79fb886bc5faec3f2412876c09ac75330c1bf71fb0e5cc7e01fd9946ce4165a9ab8bbe312320c3999e00c5223752e83b4dd98ac0804b9dd6c7252408cc6597d482508fa39ac69cacab5bc32c926779a70046d99f61c198559ef95ded1dae0ffc312c053106a333420e8af85fbbe56f1edb2cf7dbdf9e45c0581120d383b5618fedb1bc205fd43fa99e2468fb536abd9adaf1acbace862ed3e6eb3cde45f549a9cd05515648d48b743cd42e8296711843b7521597d5311445df548837af5e22f3009daa96c48b4f9ab3bd56c21ba4fd9fc2e2f32a26be33b48d6184c27f6191c40149faf9995861ac490bfd0376314e2ac5ca111bae6f3115783ab86e9e7e85517f18743c5aa50f9cca3cb8677240a63cc8bea081f6539d78d0f204b1a4ff13a15667761887b4b08717032e6ed334ec18fd566e60923021964dfe79a529964b27ea11936a44b39fdc4d361ee51c3d64883ae5fc5e5b211c6b95daadaadb21b4792cad2fe12084249bafee0cdee758cf675e4da2ff41325281f586ccfe06d62aee53dc59ddf0abb9882c477905c34bfab45da8d19f4928d9b5ed2f88897aa91c67a0d9f889f05a907f3503e0ec76116d06dc11b96fce700e1ad7da487ff581ad655a0e4064aea56d3a22ef4b41e95973712f87b9bca8e30a195f89711aad85cf2b3170a3c0fc45b24de8331a99246b6b1e4a2efc95e91fd344d8b6ce16e386f9d5ece48ef61e75a0c0f8093e69badee83b5863df59c603bd5f9abc34573711e71a0ac03b97d1e1f46d74abc89e2eb63b1743e9108e21dd2c7c13b1b2b9e11905d5e8aecd7a1bc22fdcce796dfbb0fb0fdf2c79d7711db6065e296cfd79f3cbc8afc790e5645ed94d1ba319b2a152edc68a2ea711b2cac6fda3eebc3b314461f1934c83d68ddd6d1ac728098f3064feebb7fb12273cd1a5db6ae4358e950298bdef6b1b3b2601660432a7e3fdfc1f226956d20ac1c57dfc9e1c21259d5fd330e07160e101d1a92b6f8d1bd470d28c447f344ab5298ec3169a286431725d375bf9eb64ee334f0e42d5194af876b2762f79319321977de0d73a11dcff50a429ff34a32a0b01b0370e2dacc1d68161cf37e8ecf5937eca66ce762e20249bb2b95f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2e79d1194acc91984ba734502cf9dfa3bedbf44c07eb60daf28fafe1d4f04c36642c9da0fcd2c7aacbc107273a8b9f44b25887bd7b5af5ece57e42bb66c79609549131171d1c42034f63438d91f75df3315697baa8b99b4d17c84c62d650a96ba0f4d095929c663ffd50484ad3af2046ea47e65168978594c7e2237830764a1193b550c9ee7b7e9a09b78adc4fd60b109c451ed478b873bdb2882736e140984eefe941cab366feb0c7f26c861b4aa0ab6a6c6eb9e7a2c0d38d97b365bbb248d1ce367d045dc39fedf7f874c9c6b25e54867f4d405c97e43430fd0b4d6c52a55bfb6c26db32662b4e94b985986c6fc66a11956e925716ff2a1f5af98479e9c20c054b58e747c758ab80c7764f708025871097892383d27b19bd3b55bf8088cc1b163413e2993e561b930c2df725d6834028be961bd7f28be6145923b7e672df9ff4e051f8a32228d09741ddd95029677303b454a6f78cbe7df6e0a73f669a5a7a51660cd3608f93dca5c08dc3a64245e902f628ba1bbfde42d6027445b3352e31ce66db8bd3a086cdaafd06c1049718dce8c60aac9d04a1a5886bd6a76ffca3be9d9249076fc912468419e7a6fd14ddac615dc873ea50389724b3be070cae2cc8b2008ce9a6df0ff3c2b679c61e3fc456c8c2ed005105e79f422d80767ff7e5100ad454c08dc04c4dbc3d9d556d56e6e19c0cb2d1ec117fe6198cc866cab7ff5a32df63747d372f637d71a01f4b8df625858f1daf2f30e4fc43dba49ef653f862fc4475eabc0ca47c55a7549bd947b1349e870443ddeae54a2546b14343841aef67ad85cb0a491ad6a9102242c488a77eafc6b45b2be98cdb512b6be201503fc301ea3961d81802023421e0fa94928745aa2ae01c7c08f899ff458e383aa6f3d1880ee17fcefbe30f6fca958a3656d0b0073fc1766cb20c4b564b57a5dc29066d0d197181edff3cc8428e1874d2f9e4c29ec6a831c219e25e090b9d310cf23b5ab246e61f5f9db04483385eac706f9ddbdd2f4f0712f2b4444275a086b39b0338a4e44fccc4e9fe6aa7d1d451611b3ab65b4d4cb85f75e82988fb2e5a80725962250cfadca26e3a4c8a9e502109c8ef39b1c2379787703ed5c49ffffc9117eca9c68ebde986c93350160dbaa0f4f012143520a941eb08a77a9570e9a5beef96a03ee0d667c8e9e2ac640db7adf3a966462eb070015f4e3d5ba45deed77ac18eee957550bbdc1c0efea083b1101df54d51f1b7f40f94ea0ab4179f92df0b4a89becf5066a7324f68f45a62c1273c7f43b435b507ea160895b37f2f561810aacda9667fe771108f8de4fbf675722164f8fc58ac50ca3e5618a2ef5fbd995bb868d51c3d1ba07b37776be5159b31ae43f1bc5c2f0aa71f2914c44c9be251860536f39b47f26c2e91da0eb3a9f69e46ca445a93f6b273e970bbf356d4f31208ae0cea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h19362f9378e37e82b8373ddd229e99e924745ca971f6d44aab2d7a91a01ccaa801470c155ebbb8f69480a76aabc90cc7b7e1504537514e31d871ea68f19105010944d4a650cc520070fadd97f4ddfd09e26d56f13624da8a0dc567a98b3b7c0090536a14438eb8cc2b801b076bdd2be95a5263127a5e7d2001fac0c0f0a96d22b3206b3ed6ccffebe7021bffce066fd5cfa0d8c522550c719b3bfd9f31f36774cae53a792c9e6022bc6f7df3ac664fa54a69f1bc29b81a33cb1cee1dd32240ea36dd900abc1e46f0c59b21cee2732989678a15640591fa689d1987489410fe046e14636349345ff2a1752de89fbe92fc756b491cab7531029bc0d07745ab203f4cb4e3160aff7b9e554232db367ee539d214eca950fb0a251cd2b88ba08bb94820e7480203145aa63ac89bec8f5884598b87b09523f3d348f4d8feb98ee603dbe77bf9075af0df6e1f9070edac9e95dc3bb854e83873c5a244f0ef7301392dfbf847a4452883b57703275364920c2b5bf552604641788245a45c82afec223ddc1ea86a11c874b2e209cb0912273659e159d351aa8f9147eb8bc478d852383a3bb44fdc0cd0519cb38cfbb4d75fde277d65235bfb0eb69a37a4449751a5dfc408a25058b90efb22907d520a1ed4b944b71afbaa0e8464f9f6f895986ae1ce8455acac249c09e91a88f3e4089d3a62f16a2dde3efaf61dd50d5f288277794262e9b9061353a31409296ace35fac2821b6978b9b31b5eb29c642d33e7f2e6c1ea6b0cc0341c1a81dc3fd2862e5466653a0844cc8da4bb52c28f0946e995830d8e3883a80fe29dd7f5f8a6293408c66b4823ea13dd01d4c3d60dacb3ed480bf2ed5a8da2ca79a5ce99869e2264a0fb55866ab48360ee8d7f88d4676073b6700ecda15cfa84a2d71723a1dfcfbd83eb9534b57ef58fd74df556657c36418a513f286c0f2cc424c0e4e4be42e0f8902410ff9c1fd08d86368b11e9762e60be7410230a49bfb22f3551b6d1093a911f516a5bed95876e7dcc0d524efc91a4592f1f268401305feceef5b16ec3c9772e6d760fbbbc9996ce071dd3b39be8f1021ffe0f972a307bf68a80ff25c806c05e61fab1740ffd9af27d2a98b8519f4e4297282b62d706b80561e4adec6e3fb91f3edb9aaeefc11c4117a622cf23128fa09c80bef86e5ba6c424cddc2b1b5a9483feed8e85638fdab6dea82d10d2c568b8bd86ec2b142cfb5437e6a15d93f33c53e74fb19aa4112ccde32f910689170694fc29a9ffb91584b215b0ec152c34e74b4f2faf6842f804fd81771f43b2c79be8b296b9d3d67bb5ae047eddb260c986bb1d0557bc3fbce484f7af12914cae1c84607a13ab64ed076dadf2c99d0e15fa9f8c28c39d16c050c098da0369d41894291a4ef527cfc0fc5ea185442393f42b700a7ddfc6064a9221311a7ad400689a761ab116e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h55ec228c668f11c0c4f68e032199904094f1d3d1a271973fd89bcc103db72acfcb9e96b85f2ff6936d609b39ff112d457f0b4edd510985ab61f03273ce58cc5b3f9037a2b4855b2f048a3d4c8443d7361272b0d5f6ee2e4fc3a97914097e705ff3e42e85779bbedc331e5ca5d2fcda69370845b379b51afeca24a1a5fecf6331ece198b9ecdbf2f1fe6abbe0fa95e5cbb302e1b88b4010b52c2e5961561548c1d14c5d49a9fedb9e9a2e013d73edf21ab87ce9694ecfa0af7f2a7504801626fda7a2df4c91e0b1bbb21fb518489ef99ac0bb65a726700c6e154499ca468555924b97a438c2358d4868805b9cbcabe43e2e77d071f396a90f69fe7dfec7aa093bf79517ffa775c6f0dc12d99a102a916089bd622fddaaae9a5d4aaf72ed05282bf28a0a3651288c3b6753189d9060cf3604566e673dd1ccc46a73ff10a4650052e2b97fb57f8591c6016c6de2b942e953f95c57bba2293e00760db6493c3616816a40a5a84eb88059366b84aab94fb66052dc53c120d78e318cce8c9c63c8c6de54d01063e4d8abac080ab72a37dc2ac3aae358cc8fd64c485b18d2ab82e8db06a0425d43627e2cf011159ed718281ecd516f4221839e55542e92676b424ef0b94189c46543f5299a82be661f759780a2581e63bbe142e6b3b38a18231cade9b63688ef1e7bfa3446a44a85489f13a661684ff1c164227bdb299cc3872912b18b253d6474b4ef7af968414e13287b3ccf1cbc8055e59fdbe827dd1cfe0dfd4c0ea6267667b3e94c42496587d3eb179108e8dbd16a5fabdfe67e953d7c45d15a9d1434cc199e1df9c4be91417dd0d75646986bd7055075734bd47e328424fe26e359cd13c7d6027169258a6658815215bd90df58395a25c66300fdc6ae9f0658078066b32f0b221a0682d32f874bd3fc796ede3a236ed1268b2b0e3dd7742eaff83db2a9a69fac5a421f55eaeab1885cc8668b3a7b3e2528316d99110517b701180f5d289ec665bda4787d247df8142eecec21efa838066c532763e4ce55d46c3c541a0f78165e779b4d9e27d1d313c97813eb83d1183263fa8f116b453ce7d6c83e65c1d360d79dbc600d26b7d55013c13fe4fb3580dafe8405855b14fee6def42326ab18000284bafb47adfb791bfe0d14601f2c6076f74e3f460a03fb971ec59e56eea04cf727f1015f1dfad967441bde884a8ef39913c38aac66cf79ce10768d42fb0c4f84563e72dd49dd4dd8f82d8e81d394023c4155373c0ca44f9dcb0f29556aeca9cb01345f56935eb49c3b11e3b156934cd43673013625562e88aa24f8e0ddeeff10705e3a6808a0fdc6c20866342deb83084495757e19a4ef7be5564d7b4f1a5743f94c819534887d6768a7ae681bd6f7996ffa6bde0bf024282cd485bb48b29bb179b8de0aeae463dde45a7b41aa9774f2d225b5a0fa03c6794190;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2a4dd95c29a052570f06a5e5d900dee9559b2c0e4eef8665dfc9f3e78664aa0f86b2a35a0efa0971c2123f5ff497121e457222d54c8fba745a0f4fdfc22ddff154a463e9faef8d700acd637afd5d54bf4ba27126319a693def719587afa8f109a915afa49a7f2b5e837041b3f2d99e261af9d68abda0f4db2a1259c788142d0556fb6408d5a5ceaf1a7a0120915c643dead75c2e119e5334b32c1eae98a20b58f9c53e7c20652591a9500905468aebb8521aaa0e3b3b4a07944c50161e16f15346458cf22a127130fa1a2807e688ed998de776daa637d2b2c2c731333c5a110870c7fd20196b2b3cfccb2a21bbfb1e29504f47b1eff9a24b5fb59dcccb582c92dd71664fc0eae7f39fb61b6e9f2e33b96162e97aed923434996843b14cd186c372a319444660956546a316d5ceab3fbacc1322739c29949ca4dfc1d639ef1b1d81c2295f0c636d8f0820e97249a9fc3ffa359bbd71622d1dd363edc5161561d5ea88b158f2cad6d137a237699a1ca831e4a035b237650825c244b9967f73f1fbb8a5ad285468ee30a3a213b3bc403eb37e8b772beb622fff28bf253726a8498faea995c9903bab6598cf9b4775e805b64fb7ad5daee12218f28c65dcf9a51f0cda7b660ef2e91862cfbb08f386d5789a0dc8591ab240aae06c0ac94bbeb490ddaa9384442914cf15291ca6d969d404dd880a219e3a79f5e2d0b36ec0c7c80b38c34ed0498b2826c70fb50236aff1ea56d902a8b6d0b5ef2a6ffe63b35b3c8f4e735991fcf713b084a96b65fe2d6a3ac7f2506a6c30b781cef84e16336f8874dc32cc706af62f4b523ec101bb772c23257c59217358e56f7101f970b35d6e068dbcea510da1f9a3d477000a802d751b6dc07fe1818272085bfc3ded713e0d5eae78f0dfd2c2b7703b968bb4e9c80916c0f233028df82ee8c0b4ad0d8cd4d1f2f2c2fba76bd9c72fb935d89ddc097c50ef4e7a18a9519523b03f525636cafa68585c83c0a0478d275413ddd9eec71b5f8570c02367a480b2fb1f2b9ba9dffc5546c908a9a35e405e5d848037de1086e7c0685c90e38cf6d4f490c346521105339ccf3553913c8535ec721dbb4ab09f5e557e1098bf3b690dbd81f6912ecf08aeb085be52a098a5601b135972f9be2ee0fb32af1f86333a9792d8f2ec7b6177ed6df6f2e99efb7bf6ae35455d0aecb8879c37ae48d7c9e43bf985d51d9f9dee90eaa63f83329203d6b5bcff6d5fdfea81f56a70dcf4d41455ef1fd48c8a4ee05b92336b4397a3cfab69ffc3ed2c21feed97cd60d5fc1bb1db0037382e4cc0e1c1057b8df41f0b721f75466bd35e37b183292fa167572d20c0d1d94a087f7c5362b2113fb47e4a4f246c1e0280e61bf730a920685ba5a2bc5f5115a7bb66d53f903477ca09170becc6e293ccc71a8b1785116e517770737806b7790fca24e7135295;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8b4cff4ccc16171b351dae245fa3e6ac62aec269095f079d2293a102e47872417d9a44c2693546e94e4ddff0e4c8404f7a93051a3700a027961cd5677d0082e358709c25832d93578bcb1eec654daf917f13a7a3434632bfc084b555562a4ba501725bdf112e9c4c85a2dcb7d6c87917712da3f144a5214cb0ece5c8d268adc3362e9c037a8452a465b4d9a462b443d9354d762426e00f1fd426839165e205ffc76fae3b363dbac66530161f1cb8e679cd4fb031568d52a4d279c96cc1463ab5da487ec1002db9da2a9467c7be896506b1e41aadeb36158b53e04e25cb556b044d08db8122dfb42d02276b2aa5762ec761b2a9eee5c5dbb4fce1be9278144f70022208f49550937a2dc63375aa581db53e57a25d55a42e16835dca611fc2377f595af54befbfc11b42a974dd035ee966f47004f82c95e6a256f31570871bbd943da796a7cd1257aba5f82b4d3b736df918467f4d11c2563c70b923bd99d2a45365916ae1d80e5e79489d796e16d1da896dccba88248627ec3236c402849264bf2494419f7bffecc5934603e41ec1c7816e21c81d7c25d66ca009fff900590046eeb2466d1b09f162383384e8575150fb55fafab64450e757ace9c560aecfa0eea99503d7cdee164cb81ee9f53e707a2c645a0d8a41aa5d4d7121d357fea604e2d7a35251a58cd6e339442d074859d6509742bda76b3b964286b94b98859688447ae16caaa0c7c6a2d2c927f87d09e539faeffe101e3141192144b4c1bea02b6aee8839e932c30a161b977d002d1f6ce2f3027217cb19c119b725ec17472abaf5aa8bf73e8b0c5c7accad3bd6948d6a4a620e4de613a0c4971cd47a1f5cbc567507dc0e98dd5f9e1b8238b343e81218f9eced5779bdc05c5ffb0061d2e9eacb146f1b24aac677f5491d9d9d6a07d0278445a60b83790f11c2d7bdf3ce80e849b5c1123aaf938ad5ad795081b96eb50c5ac7f00743995fab95615dfda2e547c3308190b9e17c6c90e6435243acd8dc6968c98632673d1bded1f1f29bcc2bd297ba2972019d9c39b71650d727c775e3d34a6932d0cbea3861cc1989dca43387888cd39b772ac5df0b9a797b7486316b3b3ef376256158c7ee4177103a8b519b2da2986062d645e0772bb337ffccbd4b28a9e835318473684a570b0c9b59d9cf2cbe3668ab3ee3f354ea351b7083b5895fbc2ba3442376d86385212a1bec56165be0348c95861567806925c1aea2a9516ff9e97ed42700f2111fb677e87fb32cf67b3e5af4743965a555c0d8753d6f896cb03041b494d06151a1d621d093ac629a4a78578e6ce4fd769dbe895f2226af4aae0dd03ff0cdf0024751a1f38479888924c77902e99dda2ad8c295e5010e9d70de4d05ed850fd9042d9f2dcde6b00e0107ca5e5fb0265945f14841de14990eaa7ffd901c37fc47243508114cf3de0bd8d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h42314e39da2931b92e16335b3027e4b75c920423b2a470bffc5fd571dad29e4a3e4b2336d1a0d5c42efbea0c161a4e9c138d63957fb8bef5e6a7ba08394040626ea85d2025fcb0b11dea356ff160b663df581df8d46467f32416a59b06dac212630632b9bd677c83ed630945f8428e8dd864a7dc45108afacf3376d2eacd7f8e2b5fb799a15f1b53b52e5fb19acdd8c32b82ab56dbeac8c3fb34b980f13312bd9b8c3281611ee3bff6e34d68ce5dd6dbf35897c4665057ee8aae77594ec051c6fc66957b243f16dcc4691a03b3055b90a4290ddfcd48ef9c58fc502f47997b26bc9d4b5fbe5b2ecf61334dd4a52d35aeb6c0f8829492ec6466f0f9fc5ddde2a51fbc95499af7f232935516d8f43073ef03e9c108c6094bcf0839401144cb5964f6cae92371ac588f93811083b0793c971a34fcf42bbeb9f7f27f85aa10a476876cd58b0e4bc6e6a313b1912fef3cc815c6c0417293bae7d5cd4b0a67f2ce396ef5cf87ba1f5863c6c666c1f18c7a2d1592c08333a56cf69b5b1cd8b148043cfcef71bdbbc7a02f30f67d30929444e57e1a3e381c0712ba211e97e74d97b199dd0a750953ed3a9269f0a3ed77f0ce4fbc085c3b086101cdfc35d61e2ef84eaa2028aa7bb51bb5e9e974ae722b1cbd15a4b2302a383ff9cfb2122e15476131a099715a7914fa16bf7e5d896ca3f881b4b262380292d1fdc8448a0d5963d68f9856d72db77d4d45fc4d6bb701cee87e73981155fadcf1e5924fc80256bfce6e29b72827a9914055da8043a3e920ef96eafa3f1ccb6e4d8d172b621801be624abcfa92b818ec0a1e1766c64261312a4e62b91f86c61e9c82d8fd208ec4056ff7ba8e9ff73ffab7e6b4043e4eee6817242f650e33a25c60d46e0f4c904a1ca74bcc73a8d5c4bfe125503141651f08469ca6db846490a7baf046e65dde1f3435b0988722da23f678db42b65e055b8e4d2b50f1eda91279cb0687320626b18c37ec422fb4872c67ba1519deb9bc0d11df08f165fc3a38097795066a20616215ee594f9ff9a60a45eb8c43ed65710c45d6cce55773696838b6b8a4c81e4841138645b61f9ecefc16e74b75b678bc70dddb366406d88a54d615f9215e8806a71dbb2576349c0636cae4367aafb29dab4d9701009ba759438469c8636e440324de6ded828a2c7a649c951f7e840e7a21d4cd17a945b1821714d62b69d18dd5372895cda45549e5f92c4cdfe021aca1fc4ca24543396d20d57b2264714a28b31ef1fb628561dcc88e544b2fc480d168fddb4ce47415de2861c64f4217b54bb6761b24dabc5d3beeaa2360e9e242d224a943c5d897a380924da5e9180d0590c1805ab83b7fd07269ce4ea9e85bc6b66fd22e57abf3de01062df900e3ca81880bfcf4a342f4f16dd29db384ae05e0b1849d3efd3799764b036c3c8a60c94cb58c13ebf4d8ef1a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf9ec1bda4ed2a3cd7b8a858e515a9d2d53db0b9e5d04ddcc8c0e92d709ca8c437a05b35c4fa1c23a573093162e625ae743fbed536799133bcdfb87a2b69db3da48b072c05dd7b0307e56ff26403a2caf973670b76bef78010d861d890ed4728fc2cf270fee3a7a4f7366de7a2e5f6c5900a92cfb769efd21fab252ede105e50d0fe442b04b86365896f0b46bd169bda9d6c22daad064e160eb3f98d9c358371820201730ea0d7db998584d634ecb6552cad5ac178cf4f291bbbbd6b3ff1ace6a55d7af30c3092f08a1fa145b9749db43bcac18d30ba382d559f445bfe4ab3ba7b0a55c481e9890c3f3f5d674c8f6cf1d518a5df63678abdc45e76b48f8253531577e7d02eea81535c5c9c297efd02501e908c6b0ad76f6f79c5f94cf714ac7aa3437c91142045e30ac3979f6a2accf8f21623e238309baeb78be69b51a59665862af8a68abda62716879ce21acf138ec470606cfff46464ed76e8cd152a928b73911f296c80f65959e5b586ab74526fe30d30f4f72d80dfc6623f6d1a085bfbb1c6e27a229746a32d1b923031dc5e9c05f1b17b003e3270963c23dfef3d7962e2475a04f32940a3120ed61b162c77aa50510bc98320289198e4efc4c70c1c198fbe7a47aa6cdba8f96816577ae1d44e3a8261a64d7ecec0eec86ad12e9e033ac54a607e5a5cacb58b036fd447f70dc16eaf73a36604ff22333faf88128632c6d05cee937a10cf493ae4ad1f294dd338bde25218cd964b50ca664a60cec73d8cd86e80f9bbd6ad44dbcd25f431f1d1b92ffb5d755ac36835eb1afe41c47d199e38dbdc37faf94a0d9945ab2d10566165a85c65dd3e3a681e37970210c621330222f5961eab12b19b7c9f1ef2a0a070bb8af1ef9951b11bf96b65d29455ed803f75c3180e2eec6d35d7952cc3a191ad6049be79c6f294e4c1325e69f0cf546ef79390c62a538004c3be045ca1c6b9cbe57c992b1ecc5d743bdf4494827ff66df7035946d97e957a62fced87e6182154d91b71e34bae76e14cbb1375a154d8f67626b4699eedeb09720ee2b6f61b79cc42ce46bc164e0d4fe198a69a9f82609cd3eb4fa5d2b94b92076e343d2ac0aa1f150bc19447dcf16f6f4cf77139da464e60d97995eb1e1dfeb93ed3af21c43e4af85d5e911b78a9aa241b836c102db92595d6273fab3c9fb754311daee218f3226612e9dade3492b88aed200cb646dd774c207aff1aa35145b403432c692440ada16e63f51b1d2ef29426a95eab7fb0725e4cef77d7d95e01eb11a7788590858204c40a32d2a22e3e2ce56f7f80291cda5bba6a330dadd297bf3d0d802e335d6d2418b192e65eff53ab49296836e4e462289ee5c3b103e986a581a4ccded18ee51fa4e20735c958b91513ce28d008c00454e27c9bfdbe72d3130ae66e36f9ba683217c95ec099f8d232f240033dc077f3fbb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf47d1107a10003ff1d979be7ec6d4736b3b62876cbc711d59265cd77b639c2132eaa3adf5798a4b62af9a15633cbb9b6a05f75ee157115931ef4ca6d25fc910831561346c1e9854991bbd6beae08e14968f9bf102f1dcc7f478ce406bc584dec75e96f63328eb163bf3b8bde07d40cf76f63347eccc770503ffb89b3f0dbbef48349c04f4e09ca5b00c06328033d21681ceb06ca991ce2813c1cf8209b742c649d5801e8711c5e0813907de6392972d0f006aee4670e0405feeab5b9ad33a967401ecaacf85e6b81c689cea47449cfda91b4eb892928c3238e99666a764e340a49e0e6590bcdb9d2020ebbcbee14e1b2350dc3638ba76bdbb4b4a43f194a7e186bf8dd8519350d8b06e01e4c9ef452482c0473744c06a297e99ecb9fda9f42512e1d8c8e19869013b0b1c77398fd22183530f8e729548d77b3d51c920689bdf7b487df1b7cec807c7d091b72b886676908f692e5e997e535c1a1bce0737fb2053c74f454dcc710da9bd6629c43bc0830be39eb9ff24624d9f1332f1e631ba02d61cc8a68a265cff2226ad208c6f4539613ca7fa07a7c743c77cc080bb2a1c3b7f1db9fcc340377446521b767562d813c07eb53fd6a41a36e13323900a3f4f4c3aa51a626d3ee4dd1916d4f7289f789e0423ea19a5b974ac9037e906a7c4dacff12a7293bf0c4c23f3397f774b91b6873b803a8eedb47b8f794beb233af6dff06e3ce1840b47402a5835584c6dd53306e54b823e78ece1737ac352870a48eb49b7968b10c2816d03d32b6ab179bf37104b2c9cf659d3912a08857886f6d9e69db3f76c55e95ba6e9c06c748ccee9ec3075b20ec25eb89af7800cf0494b8fb8672df1ab6bff0aaed111805da0e0548eb16d7f4cbeb19c93059f24902987b49172a3eebaa598084be98cd5f9a5a73fd0dfccb5c8814bca305a304bce14e0b29964c2da5412b1fffab2a3b26ee172ee62501cf3b9eabfadb727eaba5f68c81b0b6c9ae574d60fab9fedc7f8e3ddd7efb22f18e6d1e1e8557370b7eeb4bdc9fd33629131aee9d23f20b49d0633952098b7f3cdec29479fa4494853d5b748efd20a6a7556fde83fff20df250c45c9b2c084bfb66a59c5e64aaea34299ada2f1455ed9b43d80cf6bff63ab6ee1f0e8402404cb986c05db3fd38009232a8b077fa10cda5a47bfe0de120f1ca4b4ae8fa0a82a31e2b442dd477fb05e4ae741532d0e0813d0dbcee1b9f86529c8d55ece65245de4aba14a0d7663ba3639e161df25ce1eb2fba0e8f4ae6d8dd1db6d616c8715044726eecbde2b1c4e4dc1a03746fd86bc97ecf38626a81fd8b8edd303fcbe31555f7706b658cda52c7a457972366be278ab7dd80a3e111fc3bbc6f48e89e497784716826571e52693b50fedd05d71375a815ba2df91bab33e624456e2a8039d31544e61c7fe3726ec3e6f79b80664aa0fcb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h61cc37ebc54557d950a9b6e96b5fdf37ce4a13ffa449832a26b6de79d95c1fd12ec177b9ad64b1a310b7f8edf714d1bc30dc10e9ba0bdb24786eee7b051c1fb0be9dad8dc2a3c68e76580799cc08b367f495734b859214e0e6d93a5e53322cc93d3fa8fddb0422fd9475fdea17229141f554f5d2f847d466e9cba6285ef89915034e3305f6b82ea75831fcf51c95f019bbad5e136c24aae4145ea1150ecf78d1c3b6f3653826f544b968ef4b3fef3328df3535e2a748348ddb85299466ccd41fb157280463bd182da65043a3f8203ade29d45cd7a0650dbfa8a741e3e5f56fcb293530709e9b15f500cd411c8a129a97c7d7111d9d1bbe55a5be0ec7e0abda3a67d0550cc6a1fe93ef68ef70c06b76baff3a70a32f4d9287ef7ce36b7fe1cec816aff2d83d377bb443dcc4da30590e4da97d7b07e8f8b0e711ead9cae6c7ae2a8ba4b9f67147fea16ca10413f31be4d154f229d06c1337ac9254e1e17009a1d650dcbe2a714e5470613f0b3983dacecc985ce7c1d9d3a3cbdf6e9b03ff7aefa34edb1b8f2cc3870dffe635aa9cac67e0e94344d65a2a4604be4902e775d1bf570f889751d0451c744730fa0ade7a23dc3ae0a2d52eef0724bd32f82ac0b2fcfa96d4665348f160d94e16b164688b1b4dbab294bf379b6f609b8e416e56dafd8a9d02ab735b56a16129843edee341ad755f1a04e561645b30f61401bdc703a563a1d19dba48c44526ac21d08773274b3f8d10535f6d31eff8661d988e11d92a818bfba2ce89846f0452213780e97e947404621d092206f588053e1fb752adbc5a10650cf8596c51ff377dc08d0a72cb1fbfdf701fe450828a02d4fac8058edb10a3f8a45a3ca8d0f956560c2522d7e5552f8f943255e119451c014667a5d5b4c0766ccbb0555e0f34d410a5986a9cb042b5ec9c010a40bd06af0030d83918fadd6ac2c19d230fa59cc5960cb6ae9957f76816e6721f40a54c1c13fd9b9e85425787aeafbe3757f9b47555c2bb4973980f4636d1b7ef8c56c2dc76f4212e6f139716068e52230877c813f13b4529218f0236d32468a7e97f5e138c0470dc94469f4741e21ca0df044253a31506ac4e248c4126996e1f735412a1a801c6f114fe33c5d1b4775f20980c8a5d74d6790cae3aa6f5330723885d16cf8dbb916738bb4806c9cc8a6233942b19b0780dcc2a25f7cf62c65cc494c339f4d1b5d3656cdc474f650ee8ed0a7525ddf93e28f44289404a06f2d9761ab49056e7170b9f284e6dacb2798a44eeb13ef1aa66a3f298bc0fcdaa0905c1d1aac88f0bd2336871634f2ef968938114ede8d1bdfeed29cb9d0766452e52fe079479552693fd7823a915b38e2fba04dfa2fde73346c9e31358ded1b781c255d3afb161ace5760732a30ff1551ae20455509567740a5ebaf3d270fd7ad81ac126bb69f224e18b52c9bec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfcea37dc9b01fc423d7c37846057ef909efd2337f2bddb010a4072005fdb5343c16e18163f2305af4447f62856c6a14aab4db5ee4fc0364db2999e124eb3c4abc4fbfc876dc34af5186f152aac00adb0222fa2ebc770e37aabbbedb65f502763c4a2af5ddb88b2341a4d7cf1817b33126fd35cc557597570f04929172bfa01f412788c8c4770003ffc194017f125ff6b43580cd289eec8546f215c580dcadfa2c90c3a8be0681c07c9d3069f61066aae34a0233aab3808e68e7e9f9f3ba77f0074d91743f9a60dea524c71c0bd737f7c23b60e8642b86ba11f7531e77c5c27f5e16b11190c9b9f5774076b039b9b30a965e47b96e02e0047706605315d4d2d9168d35bb69838ba0fcb6b83c78ecb1fdfa26d2e62a5eed652ed0a6954b8978a132b67dd2e7ccda604d5284d8f371fc5ffd27bc8ba12970e5ab7905fc7f6452970f9605cf1691e0aaf9ad19ba013a80e15a425ae7bffc8bf05aba3697783f60ce35daceb76bb5bb87a15836be0a93fa9debf70a3c35a429bb91bc0f1223edfe8cc765df6337dc2357dd0447c7e422d4a572b2ddf0198e9623d836917bb6f683e576d064e8e3d5ca1e5c8dee8e0b0f94660b6c70edd5c90ed445ace86af8eefc3740dcb07feb6e5bcc38cc70a7d6d46293f1d8ed4e845633b329cfed00dc05e9bf98deabf5b14cd2f67420b4a2de6bf906f9f0e68b63e9b7e6bc7aea2384b891a2322fcbdcb59e961f77d6ab7add962c150a778e428df57cc187a7d9c8b9bd03339b5a201f8408b1c563191058fd6638bd0d4c0d632295a47b6060aac24da9017b87aee9722c0d72ee3a5d5659cbdcb6ddf07948da3c47ff76a280677afa7ad42fdd13d583c6a9890fbd78fb2c552e7aec4e1485e14837e6fb5021d55cdb0360438f39024d88be6b2852ead6fa1c59950d6ea3ef4f0177a01a51c8a37f905c83a9d482aa0701d964003df6d19f195fca604abf9d1f0219f05c1c8cc792a6f36b45521a21f7ccba130f9994fe69a4c14d9c7907e74f0e71522bff6742984a7c9c08a65e9a4bfbd841e72f71aba73a1312c1410b1c47035096f2e15e6ab4367f61201bbf2c32347f3902d5f70d5cf98014d2c194a5fb47824524cdb0e9449bd56d3fbf692eae5d80bac93985b387cebbdbe1262154c3b2f5ab2d0dc27c453688239b94bd5f41b95e49809ee405bb64f1e15c4b89832ed2a659186f6e4c25856da7f2a48d0dd75f3970ed2e46c04b09bbbbf2024c0f0ded1b3e10a952a1eca5a16f12053c2ddf4f5471689d60c7454150a7992e0238d6caff970ba8ab6eab89cd857ab6996f5566534f9532beea6cd03a95af8058e9b57987061d3e1637eea9c5cc6adc002797cc20ed92477fce546bfbb2cc4c5396e456f532282689455452fb40f18dda613064e41ce9ca424129ace7496aadf109aa5799446db88a8334d12f9f7da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h61299fb740267ea5ae4fd11d95f289b8f8ccecb69009a78bb28208b47849b755e5ba0550c1a35ad7b128eba75055d8ac80e2b10426597fb8ff9bc09c11861f4ee96ac58e90016cd9b64be6bc61ae1e70b4e89c224af37ac0a93b54292203390b27400bb1a86b4c7fa2e9ef7b39e99c802dd327a47f87b3327a88bb17c86d0313041adfd6b0fc3ac2aaa480becf200b8a08fe5fe3478052cf6f9f897086797b4a4e6a3f152e5b66173d121d66a35d6a355184f95b5b3758c9c8ceea0437248d4bd0356ed0f83bd2d48e5e7858b956563e8578555c0b1cca2056b9947a7963e2396d35321b9099cd88f72a10bfbcfec9365d1cdb4a3528a375d862b0c566b595d46045f31d989414cee797d4d4fbdbee5018f9617b5d4507dd1750318c25ef9109332a44be1b0ef484cf9e2c67f24d0f2fecf61e2735c49e5e5451201735a8fb139de87cc3f6e6e7cba2ece7385e11a48c5048a4373fdcd26857adf86ebf9e466bc0b29a039610e3934c64e8c0fbf97e82b71159656387c4cf4e11aa10103bdce0374d4c243fa19f4f75404569942878dd524f39b41110bf29266e27216245ee7354daf9adc8408136fa16dd586c0426af4af42c8f0cfc2d2381c7a7457ec01b899edbe97ca2a60247e2103d1d225038154e1ae19ec6df3d4c41a45111ceca48bcb3c2ea575119b142303a0ace4505083a763e616979a61b7c91ed38d2b573e9be3c9c97548e0ad2b3d918a8eb5268aa7ba42358f5e72cabb9cc795851a25dc399994d4987c823a61df487b529d51cd789223fe7898c86448322482e46af59bd2ebe4e5e192eb9a83f04145dcc4dd775693f618b3296a7d122396d46eded7e064b7845dcf23e1046eef9d0e7a1d53ecc26813910cda658068ea198058fb9f539e1be3f347d47ba336b6d672590fc6da5675e1da8ddeeafb006e79243592a0a59bbebf3b451f8e81a13d1c40b345f27dbf948a40554867e860d735a520162790c714dff6e3695e7143c6005e941aec8760f47c381b93c43985a5798a1dcd0ddaba2bb33a3ca6d761126865420f4d3632feeb5266b6a9ec07cbddf00ab2e40d48be81e4c80d09871378d6cf2a269b0dd6fa315f83ae65994459f709dfa6c0606acdcaae291d579f004fb82640652efba7721700fbae054f99bc96c2e0399c70d6a18a00bc8f9c84926bd176629b82b9cf396122a5406ec50122e8e2e54e059bf0ebfbc3da09ad7bb34c866be9c58d2fcefad57b48a402b506b0d386184ba07875480c5aa6c0b5cb144c9b980e7b4b5cd051c5875cfeac61875e4474448c74e8f95f371c5e202d9e29754e27fe116c4223ae6af9b4cc4f6ab301d1315a1a4be6558cf240ab7e23cfdf34ba0fdd2031877d465534a3b8699c58a7cc7e651df057e0439f82674e97411c43bdd68a68efc83ba7928eb27748ab530f1b287f3eedcbbc211;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h72b7702b0aa4dbf96edb8b7461f0e0a9b4881eeec9eee0fbb9532dd7a3e94f316d1688d476efbf616f0c83148ec9565d8cb5d5c8f7d58af6d8f21db21b29fa7747a0a6abd8f471e6c03d38603179bb1a18d0202f04ae2b00bd5f14d64360bb445898c59b5697b372df5b452f7471841660d7828f9088f2d1bf94d27057096c233cb46fddecc786860aba904871f46b5a3dfd73ba45dc1e6c641ef90ced2f9bb5f06c71c03a57a5b90966576d2a46de46f9d6dc5f0e794934b9736a4e7ec90fba11bdc1dafa3da7de2aa727d12885ea6e3f5aeb6423fe01a60970b4ecb89401ec5099647299e778b4566c0a92f55225c97960d7930c1cf2b628b4433a84fd97dc4d647399287a8f463958f4beeb98f85c08a01c95642567eac0f35fe34ac3db44dedf4bb6989b5ce5c9f1e8fef93d891ccb98f7aa78d2e8e4bd4c69af0c531a237db6978bbc6d0271dfcda4694b5df6d2c978915a70fe9faddd9041ccc7f0dbaa753e0f50bb1f52ea207b441b6124f14398d67fab241ebb340f40a67fbc2b45838fd3ad076705b262c11fa3b9dd6ce3a6130ef0318d7cef50819197faa508732b110977f43c28d869e849ff6e06e855906e8230bc448e1e3edfab13fee11d8dbe51c44d62a403fac1bdb45eb1fe70f3f6eab282fad54adab30534f72cc2c59842909bbf0a3b54164f2e50f76d1319880f437796c30b9568635c741033625d9efdfb0791d58801baf75ed3fdf30d4a4c925d25d4f085ac88e5f984312a36be20c9596488e4d9a647fb0881da853e71330fb994d32a278841bb32503eb7d3a620e0925807f3354e67a517e88e53032a8f46bd252343c0cdc241f1b2df9c4b2babba3e812884c7a168769156ff79e32dba0f86a9992b9d8abe59832fd50effbb77b7c934e9a41b8ac39170f0e73b1b34f91ba1acf3c33b2a0cbd3688a114129e1e67dae181d9ca47e70af4ecc973aa074cd88a26986dd5f69b912ba9449e14b861b0a2434f16a37b63715b4493bb26961246ca7fba1398f8e3fc5eb09fc5a6e131789b3e53076d0e5c1578a6c5d4ea7efde7b200a24bb2d77bd363134ae6fb6f41ebf43d30328bef561e34d0e245eb36468d5185469d4c7ff7d0a8bc5c259f50d20632b0b7be6df523c40d756995485f80ba7fdde3d7ea003b1ebc032ac6168ef772739da257f0ad258e3c92161c2ca239d308cc29e37f27e10c2348dd18a1be4ff63e1855875c68121bd5a5d66c84214f5f6b48b5423f2eea4bba7b4fa9be1277be4cc880c52cfb6d7c5e9f90526dc665f9017582de44afafb54ac8e8cb762802b1cfcaa7fedcc4f9fbdb502c13c19f394b6e21c5eea4bacdfe3f6ec5eeca1857e10bef53d19526feba62d5e3fb66711c5c1328c5058444f38f2341cf6dddeed0f184be985b9769596b72c45293e262be9c6c77ace4e106febff267b2303eecaf02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he783d262c3199d58f73d4fbda5732945002481235715a13aaa1e3864ce3b047ac6198f3fa46675a311d73614563944d151a9050730c8398ab7666dda86724409b67a01ed6881c780c81668c9cbf49102a758ab94cbbe5c27a9bfe88f26599e54d092a7e244022276a6535c2a4826219d20ac6b934a2321499823e82fc79dd50ef1988e9e0f47834db1ef3fab88e6bcfb4d57c17ecb866ae54918c6e9a9019a364a4dbd631e96eca29e771ac0f1254af11d5bc5aa1f80af6aaa466924eb6b4169f51ae602aaeb9872c4b9731a1120ea30d0a1c5a2322bba56cbd5f95f77e9e0e1ec9cd3ca3bebcc5c541238ab22a1083f4d71bb0fa644c5cb220e0631eea1b5591952320c3e060264c18c09eb0d2dc1ae156237e58d5dcc527a95a8ce96ffea2844d60a13644069e6b49c7ad9e542f2f61d1b00a176ddebd8a5edda3e86cfbac0273a50a1d15d37d1c346bbdca8e7fc3d5c51ab964a9b255d2c642c7f344fc7c01c23463353ee2706627dc8cdccf9a37728a3c618115a4484f8a06b57d50904dadfb530064a4b6b1fe6a41dc69752a1f813765dd46549876fbff93ea8968e599d5631a0a57d66ae25a778320871dfcf853f36c11050d4fe2db9b0f9cc68ce145dcbd1cefb3dab0b4a4ca54be3da77a31f839e0b6dc36f800f0d8c7d42e1c0e10a6de3a7411a15a3a1663558e9d48b2df05f2d639110c96998401d16316cf0c01288ab8f49624431d6f167650a4c37344186e7297cb7604ba42be85e90e1a4efe5f320e9c337ac3298ab03e171f29b89a466830aa7019cb28e17d63160966d7ef8e6ecd4728bd0594df84710ac696f8e060ead6b742d7dbdfaa4e8bb980aa9a81b3db04ede281d074a54b384383a5d143b1cf1c6c4f0e4d7858a8ab700353d7fa4d7900f746fa833f46c89aeefecb4f6f48421f1e0ce177b86e6b20b06573296da974e34b3db9fa34a7ac2650c4d618304fbe835a9431a8ebd47ab546624ee9630fc28c38250b08c403a641d096264e726bc319794e1e7427e25a45e869deca70d9411708f493b0d9466ab6da03b06dad9aef1c9fe5724ab105775cfa5934c78515bdb02a5d8abbab73fbb40d44b77a5226d3ada9f6a45c2bc2035c34ba9b92e49809f3ba75d4dd9f063f0c2bb127ab94b41eb4a6cf4b7c4e4fa4132ecb3a4340222e1ca9436756ca1d7543e3ea694161b83a11c07bec336c51053eb04c622b70d56d30cab46ed7f85163350223cc688ee1f8eb9b29996c4ff63407a2ddef4b78682f84c8b05a55d7e85fd89c2791868bcd27e2309aeddafdc11949876eddd9a4abf603442a0ee9199448f8fc85e6443c1d6a94cbb31746d0e60b98f3238db7fe46f2ab0e2b6052da412d396ae79f9354cf90cc3fbaa2f8c81f821b11cc7949a863ecec6ac2c9a4187091643411f4c21a2c8c82188dcc4aa519756928c678208f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h82114c9bbfb0e512e7b4818532880d0ebc8b549e18a898756c03d9ab12fbe69265edbd18dcdd11f5afd8f4b8b60ca438092f0630c2862243b5bb3df6a268cc6637042f33df8ed827896e9db22eb05ee5511b8b6a571be44bb9cb43d1c56d427dfa805692a5cb06da5cf1d77962ce4cb1354ca2f43456b05c9d73062dc4a0b3a06f12b7b124c25941c3f993605d4d716598a37d1969170e9429aafcb8528d7de6e1ca939fa5419bb5609374455f29f3ec77aba7a342615252200097287402b85e3068dec0b01a8ce103b0e9b293f30d2b88998e872200552383030d79f445a2e2da57eef399b89e00c0c5aac0d5d7c38cea9bc83b91e103167dfd75065a368365bc8322fad0cbfeb0c1db052b97d341d0abfb32fe7d2f7df5003f308136f57c1f6fa216febb2ab3d7dbd5374b0212ab827809ec37e2cd56dfeb1a2e5b826d1c2e04088d49d82d49024752c38cfce4df183f02802a244a01e43665c2e3563c6968bfc76136419de13c5d59dcaf33b9baaa727413d11ac36bf488aa816fdb986fdc97a74ca9436901a3d671ccd8ec82797556cb12ed866da7a6847e7c7c7b6346ea25ef861d2fb78f421684723d2311aa8638278527c159166c40adb603b9000ac17d109dd2b528893f980af70e42d4fd0ce79fa1a8aa6270171d1cceb2a46d7c42398b52ad605952c5930907b206f763658159e049c8c8cb3be0df5adc81181c412247136dfffcad2ca0fe42e671078ede63e77a791895dab630b9b9a25826d516be8f8c4d1973aab0fc7983eaefbc31115f05341c0262841d917447a11e0f69813d5150b2853af82beb95d3e899f5a122fa452264ab78e00aa040fa6c36cb60e4620b0a4028f69de0b7c1ee6b6fd900a1e3612a642514b6df9dbc1cc3fa5711d47bef3bfabc633f381f3e53e7bf8bd9acf60e8462373a2ff1d852dcfab9f7d9b3fc3dd55a033603f3193fbe77a2c6ecc9d98779bbef05abbfcefa90b72c9cddb4a559bf1dbb41e7e2c3f56d8b9432c81abdc0050cd7d11b65fe54584ff1786ca70f9d5d79beb1cef02d28cd1ff39b87f27b6a9af2921ad24191153053396c5622fa22bff384f2665ca6d017edcfd8a87aff8f7767509fbbeab83cf6102643386e97eeeb34a0a4c11b3523dc42a381c5b1e03a2ce80849fec042c173077121ea9ec81852f3d0849791c7abc8a046177266db5d9c810d47cac0ab37a526260757bb4b190a06cce7a4d540ca51dfa826bdd0f1a038cefdc939621174811cbb058ff4ebcc640855a05d138f6555bee1452542b9ff32184a18b459679412c7a6ded81b35980fdca6e041526cc68c5883cf69fa44112096f546d22224dca799eb0ca52aca85d9f14000b8719baa6cbb7d9d3689bccd4e6c5f6d8c250f1ff8ffaafd05b979f9e2d37f59b0d30ebde5abdeb2a4e945f0d928b0b533e796a9aea44eccdf6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hec21b31e6cced501c4dc5ed95b2c8270ba524fffc8ae1c2442ac0628a10e05fbe6165de761aef3e22ab4418ee1ce29c0e57477f2f8bb646061a49cb538883abbdcc60731c3d114b48052146888a1b325fd22a5181c12200c7f7e98a82ee9f6c3bbaf72d446b0062f73a6da8ff00d69c03d1f5ed76704650483d2cecb9166f2ed43515133c746a13dffbf2688b3c5d67d0102b2df99ccdad500b6fe42207bad94899ef9693aaf0fefd505023580e2898622ea1c63fcdfed1845b7c48c1897f433c1599bdf59fe7259cd4b971644caabc121994a81a4affee56a28f6498fbbe53d9f40518ba0a99c6e999a25a95a58355581f2497080a4d0101c08f8efce5a8e1fef21bb50e741d0423991ae45cdc23fbcfb74ed36e506cb958a5be503f20c16dfc1bd86311ad38d6078c2390751125e52ad60a0392a123fd0a5de7c73a648f1f49694e3155655299015cfac38226e38e318ffc59fcd6632855a12a474f5e6ebc39c1e041a68d0a9013d42fd418909ef4dcacf5a5f0c8636b36d0ee7f320a33ba8392bca1b686288fa74ef1c801c695ddf3bdba73c5eb2ef331321d6a89b9dcb48cee1bdd222f1237d442123f86c3035b5dd36c5818fce844a674ae9a60873460d1e75c30b34b2c99ac7061c65f4db399b09c3e5c58a128695b8f597b12cf94e53649aed524e1f065996970dc29db732153211981cfcb9fd7776de69d71342c79ef5fd154c04c2bf393d6807012ae18da9c4bed90b111eefc20dd072b14743a85609e7e6a0ec524edb2eea5d9a353b67d24e46bf69057f918624fd401c7d3ab94e25d1fb50d7e58901b7cbca4ff646572431f4c737dbef979d749cca4a174c6c2f1731739bb308babcbb6e34325ffc3c565427dee7a5af505ff348541153a9fbb9da4690f8057c45639946c24db8e48b306c54b8d8d6c669491279bc1a25b5d0c8f2a1bd60dc10eea7cc530d5791e21a33973808a1ecb2d8b159d8dde260379666b787b468e4c6d6c61b7ca4b8cae03cb770f7f8ab7f5a5e5d148db78dcc80a47558a172c261eea9bc0bc4104f7f947df641b5c1b49ff297dfbdc2551f0426e250e168bd32c19898dec073b333f71dcfa21f30b79ed1a25ec08744452610fa508a4b0dc1816d9fae9f5b82aa84008cf78c7302abae1a02628cf2c2fdef87472a40cac6bfd8066afa27e391e2b471831261de6bbc62e4fd191166127c27536042392ab23a86581e1ffb8c79ca5a9b27ea0c7bd61eadd216aca729e1eea3f0791bb14bce14572df45cc0858c2709591ee9955629830ad9cfadab969111ac9f1e4056ec6e133772837a67bde956bceb03ed747836b4346e47698c8cd7b26afc8702678dbd82dd65e429d62d730d5a660c98cbe857b7fff919c580085e65f2e78022d9464fd793022acc62e86076555c6f5b7e9c3d8ac498463a32d90f8bd908bf920;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha97f6f337715e3b947a54116967a64a1aa3bd4aa531bf567208741dbe9ab61706327af863f1ad789814cbe46732fc16e799161b2201477867c9fe0c5e443b1230ce0300dc99a9cce1b0a968121d0150270fdd72eb5a9418a8de6d3d2afb1612473977c0563e51278526163c5704d85b2ec731946eb92907a266b29e4bb633e95e36a6c6f6d2dbafe24e74de761d6c5af7914dadf82f977a388eede12811741c7948fecb2cf9e4b8b34edaafaf8e9ef36407b93b445abf6674be870d86eb0a9b6e3d130fe396f439d28fc053307aef15bf7d9b0d81be19b3b75860e05b771ed5d9ded9e8b3b757e3fede344069841bdb6a96b58a682b86490f37db7b47f59a9b5e21428acd7f97b92410260e0764815bdacd5f8caa9a26b0b03e01b0a1945da7b9d96db1a55486ca4b9317674bf6c5436a83ed2ff35a7c16b10e0df43a31d6dd89500d1a7698b2646f9366b56b0303c4480d41400651a7f0e6494d3cf436622dfcccaf8e15ed4f846ecc3ecdf582e2faf937b467055842abcdc1c91e61e0fffa04a641f3bfb5e234949fd74e3cc61690fb36c6c33d690826df8e8306e2c6cf70db3b9ae1521df7aaa149c73452a17b1b0c4b7668b9d2f0a3225fe4ab8815b990c5523bd9d37a4fc0efbafa64294464ab123372f1fcda5ccf147a2c0d99e3e6606a795446b37870d697542ce0847efb6364955282238d902fa5b689b12166d29b5479417cea46c172947ae558ae808516a140c7c5dd9e2d9ca075bd447d80ce9d068345814026546a7f6ee90947e1306e9d87cd293b8e8f079aa98af445e8c66c24b50a76b8ce5d63df422a9d5574e2f5e8f466df19dc6086670126cea1199e9eb572aae569bb80e3969b88b31a7d6863e228e9a3b4b5031b8796a5a4b815c4a64e4fe74ebde638dbbe170488091fa842f9d77729ae7a6a7696fc803593d385e2de6bf8c7823b01bcad26ddba787dc36b8de188b3a31723f92acf6fec561535162c7fa787801d0761615b5819c7ceeb4117f7c876fd852e5264857faea180fec22b66fba9403134f4e723e89ce8b1ac627442e7bc6b90fdc88b69431c4e476b7029bdbd1118cfb1d2f2b7a104eeacbd800b69cfe6e95aab4d78aee9a3052aaf36a73ffc3f3df49421b065b0ad6eadc235f2def198d9b5ac3d7356522e4f7459776acee5b6c41bca904d0523373cc5f70f80a9c757308010bed524c428253595660c3b2a4d23e8d0a877b87797165085a8d1172c5646d41284a7dcd42c6d8c313a11863ac2c6bd942bbd2506309a80825ba9b6b03b28705633e8430d1b1080546166aa7d28e78fb6d58179fa31ae4e5a2f161142cf9797e5ea6598ea12810cbca4d8b9490de294070de6182559cfa31c4349792f7b016d5aa3565db21b77ad05d45746850d6e1a8044e83e2fb7045144e65b83f4a01f2009adb614cfccc9cce3f56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha701a61e999d9d2b82029eb906c258932dcb4a821e1f2da94f268559227c432a9c4598cbf7ecc8597f05a2a508db3fa0758bcee9b3403b85451b331b258d258bd0fd127c93effd83364fc6334b97b02aaa34411d2f0ca509baa3581d9991fc5da43ee4f04fb4c34d472c6df54282cb6a78cb8be8b005cfa3548f1aa84e90e27eb31fbb52a4e3386f6208c7613cb41b048a27f6e640b47edcdc71534cbf36f40cbb122635d88053b8e920adfb4c271fedc6cafa66ffbc609b87426b8a80a79bdb40797368e98708778059151dcdd18ba38ec745ba29a649d21e1a46ccd3fedbecd5fc518bf8006447cc40adfe21ebdc04726dbdcbeefe0cda01080d42ded193186021957a160e906aabd2c7a626913e5b5f694e9ec608a12cab332aeb675bcc2ade685b01910cc1ef685f3658b006cc76046785e62a86a42a488c2b02f09b0ea9de0df0095d89dbeef26e1a7bfd6cc261ba8761ccdffbcad89ce90dee8049a138c7d9d3e420477950c12c6f2f5ce0380f39735cc9af64fa8588722cd4f3c9305b60118d6fc06d2e60fe8a89028b29065815a96a82e6571318cfef003c09c05177f6d2c1619ea2a0bb57e06cfd764f6ae4f67f88d7149d26992842cd53649b459d67474ffcedc826fc2b8cf10eb1803fffb46026b02c80be0b475660cfd70ea4611ee70e21125342109e6d2df45979a7fa18f02167180723192a52df4935a15d28682dec46f4f38df3937ffde684e05ae3f288403e954dac16353cb7fc7e7f7dc85794d17e95eeac2ce679f9dc42ded848b628c86126ae90d46055902459e26c80cf071462e90d7258f8c00f43747174136d1f06cfc4ba90e59a46f3088b28692ff9089bd661ce7479dd6f2c01046f387f0a45afdbc08facb6b14b83c738a8c25547afc4d927b61689bc6c60a2555a5951e197285a72ac34dc67f4ae5206d2d1ac89e429b4d395816f511b4909f7dd1031dc3f43b58e67e079e2f07637337426763fa370e902b17cc0ee26c95b5e46f84855ecc9a602306d773eaebb1d00c72f30c4e0ed9654cda3f4e64b79f3b410d55f8772e3883c3cb9a9bf1a2e91e095833c9de33b53d205ed85ffec961bb144d38530b8aa7477b7c78c11d20adf8990b24d0aad7e678fa939d8fbdb7e1a40d9110377a95c69d868000018f526542c19f1e2911eb03f0774ba0875fe1c3f0445f8b917157415c89f06e7622869a5317b097fa1a8ea56be52e04f215806b2640b73fbcf2ec0d3c20ee5a5034f583b795fbf750f5995a0f0381927e5018acc935cd7aad8cff5529f2e002501ce407d3112cec75aa435a717005d2749e24ba2bf8ce2471708aa72d98b02654960bfff757ab4d700586c63fe60e666426c663c13259811ba3c4c910461a59b1040bc3093dccd2d81fe98d0d736fa7ad675bba89ea15bc46282a01548521b9eda4abfe2dc243ddf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcb55b53c27959d6b2e22c40e0b4ad7033764f8900df8803bcb3343827e38a03a1795454817eae1c302822d377f03296bf439c2f13d4f54b4a0b95cb31a7ec3347a431cfbe9072a3020f3c414fea2445b0cfc296b482591fcedb36a4bfb81bb5995ed6195925f55bb21e9d9422211699d00b001756d3153c264c063ac5093cdd28f9b239efef0b90676726b34ae837774b1fadc6d0191da5f8d963fcd1036d3eacd95e66fb0cbe21d12360ca6d9f679e9e3cc5c3c1f9da729d6e02051d94f4e09d3fba1b2f921dac9f512989b55ffeb236fcf4cda245bbcd0fcb7bb27b38757b31776e75d5856275434407ea0c06f4404ba543aef785425ff45be4388e5d8cc1e2bd07a32e91b43b3a7d441da7406db5acaffc7625184e5082842e87bd7a7df7fc7e27b7d90a19250f2a4ccb419ef879b1f4a3d10a17c320592f947040c333daa582e1d19463d0dbe6ca2f0697420ee249136ef547c4a68271887cc54269b4b17456fbc65fedf114787e9d1d1aef07d0624248df0ecf355ed534ad2e05a976cca0bd84976b6bae2c80941e302be46e24b263277d4fdf285ce237e707f39178bc97eaf65730baefd737012ea184aed4c229162712b694a5b225f2f09f14b452d0245617de5cd30538145ce8b40285692d2ccc97c2258de13220bb1693e25461e6b1fb169436eb77efef8b0ee43da71b8254de27745c0caac828ae85b4232c98c89bfa695f8eeffaf7ff93b50b0a9362efa00e2bfde8c2afb183a0b7fd720bd00a6e1e80d393468c490b22f6d0d3744ea67a1c149b4c7604c89f4ccf1a6aa9637d001f8e5a172abf6a162206bf6973d87bd8f93597e774dc40f2c405cd652dbdb03838c5114db1ab95b1001278998e0c0e26701cbba41d838bf29d49f242177265556ccc25dead8e409d8872a16e0bf84df938471e2fc43bbfb8a80d48748382d97bdcc748427e9c35692a6fbbaeaa8838205d9619b898b5d8e203223843529c092044cfa58a7de0c42927984e3d0a6426dab425a7fb218aae4e3ff5dd87061a21d379d8efe42ce3b1cecfb1c2201a5d1bf8df121386ddc1e3c087f049f32da906b45212d4a23b5f907ef78ed8bb977363bd10e6f57d46998500579e060cc70467eb21b5de85748e960f7a4f3badf64069dc4a4e13f4f7470e88dfd6ff06e47b1f234e1dfbc0d4965a9e8336c78e39ed6d2de9286ff2d42aec45975b2360d17126cce3de72a035cb1fdf22b637689e486fd3e5cbf2fbd46fd6c6999d5a4efee75744eaac0103869c22cc7590e05653d05b5e601fd2c61008481c95302f07e65cf12a8d1e64b36ca23da8c3b68d74cf6c470395640b97f730a209362a336082dbe68f3969e354902b69fb359e20f172cdb6d45ea8c62dd4348eb93b7d5f14781b8ad617f8b50631f3f07a7e8ff43549b297b42a1432f7f5c2fbc709008e3120129f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9131949c10acd50eb435015bea0e8efed21ad66b82c450a95baf917129a2a479357e81715e95fa232f560f0180b32876f5b4b9b12584fbc234dc59c7e1d7bb0fd9681a950ca907cd074e57e9f98fab6f5deb76535b81582829949d291a1c2deefcf208dd581455e1d6cb4dd87ba346994c59bb3757f42c23006487931b4618f867e063ea9ca276a33c6af26231ef4d3a53036af6608b2c4951a4a656c39be9c9e971de3773655be10dd9846e8f3361e35202d437387c2dda343fec2aa6fc8d7b474aec8cff2949565b637b05289404b17098b9e68985288e4aa1cd831f1a1a123ca49588ef5d9b51b5c06816856c959951978685eda5fe6552ffcfd8850ad81a13433caeb57d7d3e88d24c29e0175d8b71502b6408143dd0b08205cdede287b99aeb8566d5557faf5a1e61705c6f9664abeb9c1f4edca1ed42557b880b3379bdab8b6dd6285e5e669f22fa4a21eb131138c459ff551d365a8cfa8dac78d1b267cf616f38900631f3432abfd4af57ba843cb4870d713e41f903d275189b1388487b9284b21b326ca007324ede6e734096ffe1b8efdb38dfc5740b1be6167cb9d8c5d586e87ff0d59e426720bf42b293745f73697b75fd8a53115e4ecd7eddaa03584ac785d9a4259845e0db888daf7d4a0f68d7442c30898435b80d00be366336140d6bd5390e453a0b1dde5dc2fd77aa561bd634a0cad15b11dad55d57a085063b9712e9b6ae7171a95b5f9d2ce51d9b2c86dbb56f32c44ee9854b2ba31df532e2c4095b526abad41cafc413aa15fef3a993e9303a351cb034660abc6903ae352e106fd8699ee5a28c9149e5982ee60e65e4b2627b1e4da393f5461b9a02cdb324a9b6c0cc4667a7a9398194a2270d6f10d78265c46eb4471f3e8dcfd72e462b8ee9827569a5add1a3673496306bae5777f5b35872d5dec441b30cc5e99ea10b077ffb752b5a0ddea9dcb96b5ea9b1c1f63181edad11f7444dd3df4b599d08610395012b1182fc76194c10fb333c6356554ed1877fd23a094672fe72f72ab67e7f6ebe8a651bbf09387e7d5cbf1b9473ee3c5f4ee314978f9e8418ca973b496b45c25862d06b806871a08a677c621ade14451e2154f0c5965d01f3319e8fb141109e4a49257f19b353553e606478b4415a2eb095c2c550de672f5f0c644935dd1b97267360256f553cd97480a9bd9d01d90b393b33cdcdc6abbbfd5cde93774beb0796ad162810abab2b5151b643f930f2217c86860523d388d7f2584ecf733f6819fd9fb5830eac65771beaafe733f180cb30a6ce1a05fb75eb5d2ebcc77bb34185059d494b0098370f9e1d27d1ab47a5f1ae9f3741efece9ad62d411ea3fc78932f12d8cd82a36913fd6b336530d47f16d174afbc6c1adc6177f6ac7bf152df16a1141ea21ea51d601073afcdbd82503ec6b3f37517993bab481ccc51f2016;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9b802908a55c64b23c0d2bd8405de561819de4f2251cca785e8d6df154c16736faa6307431d5cf29ccc3dae4552d4c289014953563dbc6e76cb61d287fd47f5f818ce64711592c025dccdacf3e30c9267b4a58fc93cc6aebfb0ce0143d899cebc0c7d7673b2337a781ae229b23c3a619bb41133c19275e0b1dedbefb400b63063a15b8afb81416156b6e9b662887677c6ff8b759b45e64e9c90d026c38685b2deb799d342c44324597702da8a6c384d0ddd4dbe763b4bf8a4d8a1bc1883c3dc2299d8fbfde3064aa6457fbb5508d8bfe2d36b9ff59dfe191eb9f25d745b510ee77370e61c815bbd0de029c47a0514c1d6f64239fa839e30edca7ba62be5d1e90d2eb9ee4156399b0ea0a3317e8c3d4305625f8dcdb2461d61f57e9635fd012a74b95a654ea5a76305b43bd3ddafc40a909b75ee11daabf513d151888247f80dbfea51be8e4be02e5301e938f71bff4d45e75d1f41937652f8f7d272a2039167d17cc63c2f15e6e8397049dec8df0dde21e070d38906591f762d0d51cfcb65d27c2b25581c5366fa9a7369686f53b699d52b4344a583eb0fb6e0a451c911646c5b15d4a3176971cf55c0313855f2caab787d123115ebb081d187cdbf743521c87af3c4088920ab4d3b86235493b9bfad4ed3b01f3821364136de7543e94ea54e4f56febf48f8667b9d701e3f640d698335c3a0a7e1d9753a9a35612c2f3bdb09e0614275a8f53a095fb973d6245c8df3080e59d3fd3fa96174d7012811892492fab3b831878b4249b09bcdb86e47537961a64cec3f1877cd8d5ad3bfe332f116ac521cbe2927bf867a43d45a7b5dc20c095b4858da59c1c0464e53b0d82e9eb5816dbbabe2f63683a5e758462092cbaf8bab3070ae2f4c7b2d70f0b6dea7ac876dd5921c66ba4b7f0dc2ec94e14b6b51a2af142072e2baa5540fb3d1111e48e5f8ef1f8d7a8ac89fa95794d778a66abe4a60fc88dc3a4efc463498302ff1d7bc0b2e5b3fb31b1bef64c010697c52fff1b7edf597e024287a1a0aee56dd50e010ed8b623d9f55fb3d3077cc27c231f655be33c58da9a3be421d7e53349bc4be31ca5965cd022fb63490edbe41c91289be0b1cb8afd77b02f1a4cfe49ae89c6afceaf9e427506a34ab24bdfe9b0dcc6be1e4fff05d2cee44348020028d54e9fef7a630b0e5b594facf1407c7f5eeb67844a2a03ca331e8abd544da481ac90111361b580a89fb8ffa56befdab4cf3a81cab1013759b2288c1769f5a5f6ed039212cc6fc0f778fd85ab9038b813736dc04347c68aa8c3ee7ea89ee43234389663b4b5a07567130ad0ffb684381cc70731bb1ca648f379ecb12d2c5f44cc59371de50b25131d98e8c5fafec8820a9ac9d425ecbe54079495da4c749eefbb5eebfb663d080e7377280e770590d02fbe149ced3079b1cf26c6a855a9f6d9f32ac09f4b6c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8c3b904e544073e9b1c68ee01948586f5843bbb304b8e8eaf778d9fb1880a100b6b085c0aa6293ba2a03dc9202bbabc32923bcc3342a58e46b508e9c1f7b0df727b1b828fea14cd7dd31887667584f1f62076667636b2d9228d5be745073f2bd17ec2827d6a89cce959b46410d427316b07a52e15d9ca149e587d1fc25f68308a7f05697c6b030af4e99564a6fb48c903231e1d6eb2e9b37aa9a4a95f02ce256f9d510f43a6ef28b233721c248adf2fa4ea2feb78b088bb624e5c9b85e0690eecfdd185cedda499df2f97a485f4975b8e9e85d6237a57e447023f5fbabfbc3332cd3e38725ee1eeb4e03a6debf1934db421ede8f4c18a4a1a49253725a4397a89ab98c744a6025330952d3f2b0f0cf0d2ef01bd37ab0586da44eae36df948881d6a695a3d5277dc827f0032c28b7b4a7f22d6bc14f7cb79e76fd7a1a932770c0c976bb599e085be111bdc6662512caeac3641bcc2839099dd52eb549797df78a8690c41190b6fbbd9b47727b2a75a7be855965497608ee2d44524fef1ec27008ee5249e507f9674df1c39c345044e6a97bf16382c078a83d0be9de78460bd1d805176fd638e0846a487d46e6087458ed64054fb67e46b59d2fbd26e543c94ab1430464059040e9383c7e2751f9d9a1dd39ffd3691dac810b908d943e4362d6316d2b206dcb0b023f3a2165659caa203ca5d2786b012e7fc7c2904dfe0b1725c5ea646654c3fb6018e0796df6104d6d72771ab37b560ffbe07d1b0cadc3f5d1e1cc911ad0403b8ce81fef7f6270172759367f52a9f6994f053d66e0d53ecce5b2c93af7da002ee144880bdd6ca21884d78bf4549b950a800713ad84a644a3e7473f9db1e733376d8e3ba6619d42f8373a28027f8070b4071f5a0a0737fb5bf87321c7a9d15a52a94743a7bb97a162c2c567a71f9306afd51392df7fb5e4d288048ac1238dc197a98a648fcbdf19932b2935e395140a9b92bce89e6438b02c608a25b44cdc05c6b0e075d69ed0c732f6b2de4b2c2f6b40b9376c5086a09c149407d2b4c080c42efe04a28ba09275da672e64dfed6c094bca6fd00e7056456be1dd71fa8fa0113e2193b7d829d6fa44fc2c01a106681fc2c6d1d1ff0cbaaed1aa2fa5b2b6ecab58ea55b3354a96b79e892093862f68c7e2843c7ccb2e0ab25ff4ec47cd205d83cc4d2503dc070448e668ed3bc8420b84b88513a8c7f8c2d32abc407f4f5ea1ada5d9167341e43aef40b75f3f05ad9f71189cfced6428d77631cb04e738c91f9abd01e10171a35405a7f2676ba6aee2d06dafdc07c5662216136ea26ddcba57a4ca819afecb8f1f9f656088820d4bef87ff7e1294e6f4e637500b9ee29bcebe371ff00f1a4b85d74b985e56071d1ee0b18ce279bb581d69ad144d14265720e7ad77fb095d1c21830d5ea4b745dd9134f710525d69a5b23b5dd76321;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb7c1d1d64ddb3478ea34707936a18092f1017a947484f5124d793a16b9be9a0a9553e3600af95a22a2fbd68af837a3eea05ce2285415327c2ceff313b6f05a9d2cbb19242bf80dc5674581862ffbe3b2086dac38660fe1fb167e92126daae9fa5908a9caffbf1a20f039541d332725414e069630e1a119e88e2cf86f37fb22085d13630446259a5b1288a45a302f74b990f1bb5aa56257f156c1cf3c71e41db9f5f6158811cc50e02b54f84c8f732e0fbcec89155abe60174a4c397fa3d2c5e657bf67409335414e82ef373dcdf27e89a660c02208b5ff45bfbeef49797eca9cafce7c6e974fd19decacc08285e7e932dcfc4384525103f7e5ebd0119b7cfa970b407027cdea05a40268e5ca305a5bfadbc91c44eec2e2707b6641ccd8d11494c6fc1276284536e86b635ee0ab77e79d100a3651b07fbf6201c45d6927af2718bc270c8c80e6781ab6ca87f5b9efbad7ea680573e2d5e615a4e37667ababf3b203a23a54204573218e6e9feafc9cd38f9c8001349a0fc42396662500896f494a65098970b148135afbdf73f4efdedbf67675835fb13b3c4358e1cdcc1f4c3f54add5925293510fe35909810df89b6c61c9d5dba62caba87e8dd6ca9328680387e07901151e106bf454260acca0de3687350a10838b5a7645e51bc5ad4a6c8f02234f51e7b938fbc025cf6e3bd08921e95dd6ecac75758cff633deff07865e5bd88fbfa8050a8358100d361654dcec1b2d1dec11073660823db88569130b90cd5578cc3d6a2a7128169343f638b0e40669d1495238ed3848a31196ed3825597186c0497c5316f992521012419720b7f97ba526047b6d4b96717aafe2dfcb07eae7e0a1d415915dafb69cf066908c583aee0bf6451c2cf4252aaea555d66a7e7ed0452ad94f90fd24614180a611d36ef1f6eb185e8dcecdd4a4e3cede0ab47398f0ae115704324fc7370b8348cfe885c69ec2c6d666aaa8ad09e0920753b4e494bef76191115d5e592b7fdffb61e08b3be5b3da5ea2d5c75ce2a3301f1b4e5f038846dd53139d4f18d8fe3612e6e2bcf88381493586fe346eefd0b470f5b64840bbb8e023a17dfc262cc6fb36da949f23e51c2c537cecd027853bb2a6b0293084f6af924cb499229590dd98549c54230d8baa7d9814f5dae767bb089f450d89d297e2c33cb4177883bc14702428b02bb97831573212e0cc00b7a4d2c82ad27175a48808141927a7b060894d1b23b12bb543c697e012c9f14ebd75cbe44e944aff109a3f6454c49ce1353edb9d01541ad708bd006b6f80d3c5f2e9558b45b1b7e867970f3c897d78ba847b60e8352ad89af76156d1ea24d78dae17951ee10744b1cd5a12bee827f9ebc85dc1b19c18f7cafc07188438b466906c5f2e616f379030eed1b11ca80cdae07f237414aa2ed58c23ed2fb4e0161088ca050e866f1c84e30;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb30490df9d6e93062344a947f0868480caacaf665678fa53bc5afbf526751e41808aa9da6f32524311b23216bd9d256542e838d32cdce82f9df75e37b8a72462ec081c79a27ed65cab2ac6c05829781ba69494d1fab6f4e1c082e4159d999d38761b33ac373676df7a0edc5bc23942c35502205c5f79e0f98ff050bb01fcde0bf6ef481ccf1980813f819ec07a6baf0a870ee0231538cc8af2d48b86fa06e9400def5dcc6b830158127479a8981d105258bb2b4e31f567a42841f85c1a9b47533d0a94f5c103915cc37ba70bc074f4b39f8da0b144e566fec1a1119162030594d2347139bab3bdad67f398b3eb00886a300c4ebb8fb02b3edbd97413564a23534775828d37720f485ec123c5957020c92f4521501f91cc6844e34f1d5c5eb104c6c81c1005b61e9223002f1ded226e5f8cbc1deff645a4e747cfd3699ba59e6ff2015f29bce0d0e2a610140d11fa3fd2610ee938246e46e50ffb5052cce50b2b7c7b2dda4bae559df2218af0c79ea1ed31bcf2e91f1db4447131985bc2d8352043c6e61dfd38739073770e3aaca11c80c8ee8fc0aec95b2e36a95f0120d94434de719a5324b3ffbb00a79c3d05d7aad73eba857bbf9a91b829a7860738f6a0d96d19c82ac0f6f66c19ba9f89b225099f50ee84fc3299e2927543ac9750ca0122b991bef927843a92a3b493b9a6c363ab123733071127315e85d5c52d1d860bf6189f0b9033fceb667105b0a51e594b4ffa89e1c4b8574f2e33fea28fce8b7c13d0c978fdd935bf8575b88923b3f7e88ee32547381f8d32d906b1e3bd23ff9735c0bd8611e3e9964ae85bbf1ac9150ca47a664a20fef64170abfdbda4b041058222cf1d231de1c5eaa438a1bd315bef780d94f7614b6ea9849062576b54ea00e4f8aa93642a5445605c97b7892d6485240d60ced8633304169ed8a1a76acc9ee58d4b5e8f5a440211a465e9702ed89dc6547cd6372bd73d9a09fa9f9cf885a76e9cb349412ac3529399164f0020739609e8f4e588527d5c30ef80fc27e6d3092f83655737558647e51a18186e5f611f21a22ee6ff526b905b81a77c1984d2e3e4dae0f43810a14e393448fdc27810caf84b80254f4c5da93a9f0a34f174f959517cf8f948963b1058b7c09c289c417ad11b6fb034a0d3ad3e99a97856c461338fbd75ef1064da7bca63c6748cf46149db731c75c022a5bd7b00dd97a4988f042c5ca42535f4bf0f09f82906f1a958848deb01f644fd2f06f99dfee8f185e3e47cd294819ddcf8d7f6d1ae5daeb49541403ab3bed5add18adca9818de824dc6b0e8e31984e532fdcd53d0a35d87f43df690ed8cb97c0d9dd4e367964cd0a8c75482ae95779f5f8e97bfca4fabdac9aae60be835934e30454f9e5fa09de45433d193331464f6c339b896484f01566efefa25b6e43eae52ef9d4f3e8497e8c22300;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbd422d2c3c63b16177f2b364af6ccd3f7856dde2cda0b633f189e2e36b47f8252537923b9878f63e738b220d950476dd874506ce305482ff4ffc861f81ad2e7c58cafa80144936d602bd76f982ad055110bbdbf6793473b4e5d2091f3da5d9d33fd359d79028fdde8fd0dc4d1bb04294df924d8a7e29f50f87065212363d9a79e22f21c4afb9e86e5d1691564f7ef2412100eb7880f9c72f631fb5db602c273a272d58457b482f18b0892fac5320c758d012b44f18a3e0013670d7ad89388f5442fafa07270cf911611e44fbaa8fe10efe2cc18a7e86ee77a19b0f64c5976dbf216f44470c56fec626a12f9fefbf6f79b02b55e39539f878675aa3a95a717a972f41427fb2cf49914573928ec651916e88017d89f876920586ff834a7a887a820cb75ff2700f1798234ce88cd1c67d1017f7dc6c1cbd17db903d6b356d250eb6de1955f0d601d8acd9169fd926b08db56cff42e39165197ad3bc95829da3233babee3b83b45961774634b45aa207733fe7ebe50a20f5498eb36e192a329cab1acc4896c501a31bbdf070beb2c272ff4dbc1eef5628b26984a41282b5d26750dd923c2b3638e8a223e28e7d864983934e357873f23ca55caae0aaf991eabecd1f8195d55b5eff810cb7a2e82fe1a1fa886d66e1ea86d51128e24d7baf4f8d087c2b21b18150a8e5ab57939f6568d1238fe1d007124ca23c0f77d6285028ad066b9a19cfcc5bcf20181a217fde7747241bc238bf3cc3a0a49fe683a41a7c9b10e90b56273f21c3a0b6d7febff3d7cf0650d4dba7ead6f8793a07a33ca264aa1bb2b48bd09f39e9d1db7325352d835576b9dab413392105dfef141aa2a7653e6f166cad01ef720275793beef16e02e7698af4246b7763d3eee99f5c35a323d7069b7ac0c72dab0e180a86d99843deca108deb7bd8678bf54ac2e6c7cfc2e85a378ffed2a3de66c92f6e94a1bf5e301aaada69288576bf5c1a146e7103f225033f859078b5720cf52f5980250b29abe0533ea2d7a28ff0cbb2dd90b61ec903e2ffd02aba05690c5b1dd74933243e8866be28a25367b6ef8d9f680f0a1fc6e82d934114cfbde5dc508b9c0537d7d6d40a3f90aea70cd24547b09b057fd9cbc1fb8036925fbe97374040160c46400465ca2ab88e118417b0a7fc91f7a06671aad4e4bee9431e5738c35b2c83e7f5ecf1b644ac5a0ba2aa3baea90c558f02bc7877b8522281e19c1204246c31be8db1ea06ceb389aa6d0644ea148a0033d9bcdb55d657baab9ce23ee60fe443f623bccbbab438b6dc4bf4c7e9deec199dc98fd8df0ab1e38736511fcf2f63f2ff55a248f1728a12b8e77275bb290d243cbb094007e910bebc97a8dad079711ad0210f07204d2b6325681b381b39cb2c803a4c058786acdfd99ee7a03ab40cb2a3f961889442fb913f242b88e8413e5fccc0987ddc2544;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'haac478da0da6b735529d6caff4cf467836e0d659de265c952a784c34afce62a0914df1098156c5766dd36d65755672608f105a6d11983a9130dd5b1772c4c99a82e958a927c694f207adc42d3e606461c1aea80613810749e27c3b9b5282278c82b4b6443c81a460dc04e23958124b2d199c117c55cbc6de198224bb33a3ecf38dd5ab60865de7053dbcc4676f0a6b4437efdbf08ee74d083e537f9af8767633ecd19f204bb5f19e34ce1ce78b12e82e7436b33f44aaf047d04ef065876c8fea33168617577f17ecb49d9177b45cf6d2c163431460d0a48b96387e396af8ecd18ebb8a9cbe0c9080ca923c0622fc2712429212d672336217b32aabad4aa1c6fb77de204668f83abd7335f914baf30ec3c41a916eac9faa97fdc32c5b01a7a68b346c78fc82456b87e4c091d4b17d5d572b8334e4fa76d7b70fd71523075e861aa0f60e0c02948b1fc77a7cd8514bd4d0aba13411b36aa195e803c3208d02decb9e4aa06be3e971d12551d396bcd98db31ebf95a9264665a1edb399d8b5e6bb707dcf30b0e9c634ca65f5fae38c203da70a4df37232387a3fb625ecc1340d8f7c39ff60354b80b88b8b8513315153927990ce9122efece75b8936139ae5143aa90556ca9f85c102a53a4051193d5cb8bf0e679730073474ca3207ebbc875f873d5359056da70af6ab55e8956dd0c85ff157e301d546bb8b4c112ad90ae4956d68022bc91b7663507259ae6c36819372161d57291b5161105df4529dd25d0fff59963ec5e8b377ae7d16c297e7878701d4bc22bf5579f9c6e9fa0a769d15971363c5c4566a1cffc47dec869f4636bf105c9da7f0da9a90baf61981676d9bc107fabf34aaa40a098372f119454f3b39506f2412071e5f940899840ca3d139dc072078f2289927b059597db7900f7a83ecece797e53c670fb25550acd0a7ae2c102d716634711253d118fe96ed91fda35e10d82d2ca4ad4322a4db52f17795f5fc7e395a6653579456fa83f4afef93c1ed02b9592d6e1ce25a761297a0ea1e6559c53fc731f2210521176a1484df4a402c102705adb93fe3635f35cc639948a69eff70ae831555066426b67ec0afbef9bbe14ece6b4b3ac7134393088b791a2ed498fab6937a151a95cf857a2e297c7d23f9606da8899742936e9c3240145e969f5bfd83b3e1d094f7957b90314cd5b340af84c04f8c6eb86c5894d1d959d013a4ab45bd3d6462317d793096f97a14ed06a525a364673ac64c312b249ceb0889236b33a52b85a8f1181b51f0e8341964afcec3d88527ee9ef70b02372b2ae6e0efcf1aa8384c18dfaa38e363e2b7f19e63734dfe36fc248b7aeb6c1c739fc7aa8e2ff9c53e1f0a7af248b350db0efc937ace05a4d2ceff32d264d9eb0288d2e3f6f8b1ebc4641feb7cf0309bccc2182ba8f7a3f9b87eec8e05e4dbd9a0d4089a7345;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4cfcf75ec650f46a7901446cd46bcee8a0d29998db0894dcb630bcf808c424dd7346b3d63abe05afcd21e2064fa9b3e776fe39bc1a77bcf0f02fc864f3ab0096c2f51181eb0289c9d03250f911c3aaee3d78c62a45d2184fa3961013156efb8540bf57cc5983dcf702003050a3304373e730c6b08c08bf994aed9ce586e57cc5207ee5a860b5a710fa163da2eb86d36b8d162ef95c67ce776adaebc694e4c88eba43bde152ffb165253c708c635969cfc69ca7ce0087c44c158752f4db9b97a2649fae4d5935bc0fb15ad3938382a2f2de747e3b128fdb0f7ed6ea6100ebaae3629155980326715b5b35577f4f475a064e3c40fb57bb897eef35ca04f119096f6b64a214f59da12f2d6cc392664951e629fb8e4e9c9739fc227d8efa6bfc3103613c237c2e5b486982198b63227859386faf75344b0a5359c3e4fd975cb9ea0b343a4c19e330babd3701b1a75ba5c7b9b60e4b05d9142b917b241bf1e6ae62a6aef5b24b0f692d0b9a649e5bb430e6e3a5f74023a9c25743b9f13186c8d66097ae80fd23b51f428375399d5e894c58fa60198529c0f1b5f897c1001d72ef4d78e237e0d37be2eb1bf602c361fcb4d1551dfd115df465b6c242e18882b1ca0c9244be15e2c0e8179b55c962a30b1b52dc82fa6ded0fd8886c621b8f1801fb5c22c20a1cacd457aafac285c934f9e29b1a70ebe6e9e1b61313ce34e65b69da869eb7d159b3be0fb6e66f5dd8edccf452757bb7de8739256e0d1665ef8fc5f0b9f2ea0d377f6222561e4f3b25cdbae1e472843d7b5e7f50bf0fba4406fd821cac49902eae2575515178a44871c7c0ca08e1dc42180d005ca40e40bdd66a802c2e7ad72b4d48ce25a27499fab32a59d774871c22c0daaf45dbd5df5b883a5231d7b20e1537919caef6925f40a91e109310a4930f808b4fa94f2b739d0b1afb66af91ef71a8237f3abc9788b060d89ed14a5c65f8a5b1bab32d2fab693b5e3a6e489016ce9781e4f0c763d38179b809532a08292fb3b7aa7980e37b4a42b614e4015c0ee83c843196f8aa39924fbea17151a66842468e3848aabffa5fbdfb0370c7a37970f3ad01882303723b20e62729516e9954ef5b9f866733b6af64fcab976c2970fd78e11ce9be1dab3d3de1b6cdf63639bbff026dfd4d313a4e2df4e3babec03daf69e6e58fc5a2e2192b0d967d41b001e980c5f74ccf536ceac0c062f37f7f3f4294805dc457c5b35ac01c363c9fbe42a0f8c303d394bced3c91dbd022c849c9968147e1c655f5dec47d56917595bbafe4e70f81bb47171690eefc9343709573694da4fa8aa9ae7d83166be73cee86308739437e1ea23abf3af90ebddb62c9098cff8a328829eef80ca696d7bac97f306442a46d0683e6af2c24c3609ead3b97832167178c35181a0b975cbb4740b1abc1ecca581c5a6d7aa0e9c4f81fb0fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf1f4abd05ea6ed06eb92ab74cde326613df74cdf32246017860c11ad5fe73416d48d75da8ced7283edeea8cad17340e9fb4b14379550dbb4900a53aa4b972fb5b38dd91238ba44566c92bae92e39b8def9bdbdd9ea181e059aef285711ccc965958d4ad7d1c3605e6d981def3cf669ba351b373920548d5914748728947ec14d6185460ac785ee5e707029073abe1a19bba65d9fb6322ee1c982a22bcdd937b900fb7979ef378c76d1dccf766a31592c8580cafd4a81be837337fef09cd6aefb037486ebf52e6a80cc12c6693b61044725c3dfa8bb6f3056043a53d796d2e699fa8cbc63021cb1c0315b67e010d2f6f93752edc622ca3b66433f4a4c6666d4065e6e7ca4aed06fb36d5b55ea73a03c943f898fc1d79ee3d110dff883ef4209574e3e80d427149331b8869a854ca5bd05618d1f8e5207ef186e294c07e1e80d16301083094c5fb114f0a1e22b12540c8bcbba920ff4d260e99969aecf264cb626cf14db54182f3385d75562293cd8e2a4671f39de6c8cace140e2bccc6d208013db728d3b6789d2fff2d25851dc7a91cdc8a98aa7251e9ae62b3d5c5e7ac4906f3225e62aaa4ab83e54f30e57a915308b2f0cc123c4ccd69623f24a3c3439be7cefb93f9a4b822395f09bcb60007b9efa7a043b0b6121db5e2ce2952fbb5a7fc03c5785de7d0ff33aa3e94178f15ce1eed900a228e69918cdaec03b2770a2cb529033728458bf861d6daa57dc6d315d3fe227763422363cdad2bcae2a2577e12e98ca2997d61bc670732dae53c4ad4b89d38f0ac8f2effa3578f895859ee72e4317f83d98d2b1ebfa6715a6448c4859d08bb7d1ba9c4158ab5bd9cec41aa9d2d968ebbea08b225a5385ff1ba8bab3ea8c620116a4a25ca9ef5e55b1e7bf79ec06852c5b21f00b38145f608a858b9a35f7f647dc1e4ff13d2b80caf1215f35991d115cdd5438496ace32a1e396761607326fbf348ff4e38b77c83a9149c604c0717dcf037ec7211d34e47b8d94d45c8d9ba7afb393febba199044ba1a4fff4c512a7d86e9b2465c686dca9cf05aee1f5d6042d82a3a70614f3500214004cc28fe83c42408d244607169c56c32b64dd6352ec7b065ef35b5a2b5e457d13a65004a7dea2626d3961d176c64b0b51f060bb40eed17b5fe431e66679a3e235726063624540edc38b5de989555775d5410ac13fb0836ad066f3733f98aaf68ae5323edf14edb0d961176abe736b97f2cffd6c7fc988c613c585f0927a4a5ba10d131c1e4eea25a11b778a45a6a22bd334dc54a8268a7fad166c32791701e268bfebb41048f7290751cb08126a12cd5b2163a3994e667662110182409884a7d117c5d666f61facc8330ea04f1db293eb1d10d05d23e91bf2414baee92db20d7b96b461a1f558ceef4bfe816ffefaf9e4c135cba2416f4150285f37c92dd97c2a6e3e5001;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h25958b784c01096d2bafd2acc264b6c3a709a96093147b1e3da20cc769f42909e14fae13f4cae1508a6c90f6ce24d00a8f7c9340bba1224a90737bcdb5caded27e746f9861b77a68cb49adcf60bfc8fdb5149578ba13a806dff783bcf2b84d1c02da411bb553c65e72910842ee59dde9b0643f36faea113d2aea0715851b84eb0f37b5d6c6e6e6698ebcc34b3715f65c07eea51a4d471522c72984fe9ffd75260d509cd05f443d548e56bd9bff800b74461583ff2d6a7751e7fa47671879e7c90bb4414365aedfd68b7beaccdec8f4bcf9cb8700168c69608ebd2bda86e184c02d009896916160d697004ca2168b857d8f1fed808b66b46ffce9e4d10aa9721c7534effb02de2b377f74d38017283d72b49c25d1a9d9d3c1661622330d1618f19ab62999532837993e1d0e7b1ef9cfbf87b049547d93e1eb49a80afaf0bec4d9164472ce3ae5d309349a3f7fa905123eb36e89a6a2f8c08a02edc2c90471722b3126f9de1b554274e059cdfbd99d5ca31890181c2bac44ff719442448ad6d762f676d868473b5945c327a83ed8744e5e1c007690d43dfe6f80dd0d17e3fb51a825bccad78563048b015fdf2bc0b0f2aff77bdd7b8fd11b4e698871ece811c56b6f2ff9aa294f4d8d037dc9214ce324e89a42fc24a0345ad52cd0b41030d5804576e543436b633aa3a171f0f6932aea25596a388c33236a765756899d6994924308d6f5a880a254751ddd2fd225b34821e55f84e659526f98223fa3a6d5b864ca7fdda0b8c4a6644f82bba19baa4ac128e9e5e717c2551e072f85e504fbebc74ccc008088fb6a5b77004a7b8f7b65788729804216886dc1f0daa639a78bc7516b6f8efdaa6dd63b679c2e0521fef0ac3476ea4da085feb05c4184bf1597027a7399f46d583fa280eedaebc1c973ebba053d5a7541453bb1402c7f36937773590637a7bea1fb378fbd26c30e692493248a812c6cc2a5db3b64e33b348338523bd10476dee7a32db7afbcfb8f9caf5ce32380b63aaf6e19bc8a59cea77554fc0c15241e15a309c702db2ebac69b89aa75384e6b06355301bca1dbc07c1c3d3a701a6017a1d691925b63accf486346bbdd8ecbf237c2c95a7525212dad65123f2f550d7dae4f122a213465dace41290058296d2c8723599f5b38cd40e262a1c11763bea673e347e5977887a08e56fb0ab28b40c32801711d1e7ab2dc2f841bfdb018805db2b6e6898392cc44423dfa002a8ddd772bceed6c43e51bb2126e3616de1668f38e85e630f790af70249574fc85e64f54e27a90781a3c46c2089f3da2b9e6c5faf0d0652ed1625378e9a5dc74bc8da725bc943060f3f87a799fc1c50e6780fe23dc1a6b1ca8e656ff71e7f8b7df76cc84d0927d205aa6fb08be1b7564911df480e1591a9245bfa725886ccf9c293bac21b5cc03263af95e23537cdbf8247b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5aa2de535eb91cf725ee432a42f888e62df1e90df982b55063ba50e9da2bb60fd8e8266e04ec79ab76cecb91ef347fb60c5b20703f73a5cc3b16221ac26d74ede8303c82683afc4a8aebfd493abf6be260ce6f3d97099445b5a99cc5f69e5242e9941a23fc260d1e1001161300e465b7518b5814e89bbeb09a915a6ea1c973f00191a86985ea9503f13a2528fa3798057127909daeb4f0708964ccdba63abd87e3a5efe62b61bb724d3ba1b8200daef6783abf5b1d2577ff59da772292333169edc715fe46ef33917a428385540632e27373a079ba8b9ff5b14ede9883ead4b9606b3cc08d0e80285e8c13d28b9fca123eb823bdea3fd53584475d8af2ce6e2633c12cc8b6e2c68797f6b0f5ca46b55748e0369e010901814fa32b5bfa20118b4fc51eab770e4936cb4ede0d78f131ec69fed31ec4e0f13d0b78134a937906d88a16d6a3649ce9c69ab0c3dfa1a30cbb2dad749baa0210667f2db11d2debe99078713f45b5cd6801ffe66a88a8ecfb7842a5cf66866e70e08b7327e5059526a4b81bcc1bf5edc0105559f97522797b74acf992abe15a4717d09d0c1bd5246365096a0586abb47b6c3c51f4094b579d3bfdf92dabda95a08bf0f4215309242a53b0c80a336ec7b9d23b6a3f45a59c16f7257e9e2a463b29bd83faa97af4ea0fc8c17b599038224b9d7204bccb019b30f46f3d9ad9202ef78434570846a63e9674b87491613bd951d98202edabd5c8819c2c16ad67beb3c2f208f111e9f081edc6d3417acaa2b1b8b2838c9ad36f6d5d22fe34dbee00f658814799601a938a5d50e32f454838d2cd40ab69c5e708921f07a0d9caf4bab4e1cc73d3ae13724b85a6de6674cb0c9c45ad21b60c27435d3a48716eb6e9baf04cea8334e8523128083a1ec32fe47090be83106a0225427b32f38dfd0ecfd6227b33ab6eb944b6545d1f74a4e18becdb1059a16157473bb0931ac1ebf30cc57b0cc6ac7ed520ce6d039d6ac9e2c23049d65747930cddab99aa8b10debccc58c4ef6af81e5ea0e30fd8ddb744724d2918ba769a564249a78190b51edef74de46d67ca69685dc094911cd1bbaed1695d809e04e63aadb3f6a3269ae10d41ba129bfe755ecd313b95b6e1250b763198ad0a5e4116f411a5c977867b88bd157adfb846b2f9925ecb425d06d91a7e12a7a001f06b706f124db553e2818c45120a093277f817f188d3e7cc74ddca5113b5a00e51460b28f2b254d1d2b0775f68865507155c89dfb1b8f63e4191b1f3e99ff2fb1d587cac4d6a442ea4438ba83fb0c2e7e9719fe38c05f14a1511324b25937028a7b664f22977b6307d69d57675eb28b5582891ab7a449ec723113f63f544e0963d30d86ad12f60034d4cf114d62af0b8900268585f88bbf09062842aed30f11c66ed152b9fd84c09196b808d868cdca07e3ddc033ba044ff8e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2b4a6e14b378983744ef26c92325ac057cff4f8fa05469529884dd251109af2efc735ab657d9882f3e1806d49eab72a347d07b8f88ef8e47590d4b6854680b9a549e6887bd0c4d8631a1dcae4f83204ee52d8218e4b73b77558d04244ffed93a8d677451dde76b492fbd38e307296286af546a1f0531c18bd4ded5ac2862219ae395a6c0cf69a924587a542b3c17ff3bbca82575a330cc4afcf6f1ded34627aa3d9db279a8fcf9365dca60095c07bb8dd409a60f2af1ef6e06e31c14a0b5778d5da1a2c66dd916d174ec441b8d1e15c49bff7aafd2f84139aa3e7b7dd43797aecc7ccbb9711d7c90914d1a7937f22c1117969691ac4e844ee8a3dfffa165545341ade53df0a5d1271705f7e75d89a8eb49b41f7e28c677a0c904ff02b01f02dcb8f60f946d912d417abfe8af7166400033863e2109d930f2e4d510f45e25cbf5f91effe69814994474a29101e1f2fa09ec1e9e6881529ff19e7e8a8be67b49fecb898ddc144668895f027c6c2033507f903bedd13924c53bd023fa36c845bfdfac778d22a2e7a59563a728a3de0e74738c9702e7442505a607c30b41b61881d86cb894f479b555c9b6b7e6c115f72524d4428458dd9b2999c82783441c1c4e8038eddcfa9ba4d72c8805f4f773c2000b784a6bb807eb297936ff4786be380b87888854e4e3ab65e0ffb5ed9f7f5aeb96eb8a46e5a714b88db93a74eefe66a6e852f058c7166e33ca61b8a856155fcea3392865d0ec2e210c64befc7661a578682ca3aaa7303504dfd946dc5e1dc7206f7f15e2175c09c01107f5b7f33fe787bd923c4bc7c372ad16a11d007b733c28f97e5b54d1b351062573d573e854e7dfac7a33a9d9266c855d0fb4da6ba187fee72737d5a41831312f626b93bc1f26f46824268de99c69126d5bfbca0500393d3a585da992e354edbe6af417fa1b13ba6d5d24adf85992dc8a95b808178c965da5309045e1be97d6e0efd6cf29ba98c55b14e43b35a21dd3bae502d736faf7d1ab6abd8674092ec08eec82395802fc1a457c1d2f787a227d9ed2b853a94cbd77e477126167aa4535cb5bb7c4e16aa61c1a234641757e1d4770637ecf13644de1d654f66bd61d0a2b6f9e7582e8e11a267fd173d8c12faf903225b7a076609f9328760e4e4992060bab0f79a54bc26b1851dfb3bbff6d69dbb62ef7b4fa81607cc2d5e67665dd11ca86c1e11e96ee4c89ae088e41f6e442601e3b9af3fa99910a4311e2402544d472d024f744de063e2646468c7256c160612e38351b145c4b164029dfead9048cb0a6fb858614d0bdb2f0603a157fda41227c7538233112d2b93b3892856ffe5cecfd402003b567bddf697282a140a6d4df6043bdf9cdfa7d08a90d053fa0399746794de2cb11ca6653ed227a97d6c04225f855d74d282df2c4dbe142d9b459dfb1e0732304aa34de3fce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc54aa44ae2c73c4e3f38f56aa7d5c37e22689a3621bbdb5c2e70d5c6aaaec87f13d2b4d8c8069063bec5b3c5ece6996d046e55596c8f848ad941c56cf0dcd9beb7bae44ec3da7caefaf0842cbf4f9433b45b5bb1c3f7e99533db863fdb47580bd24ec2f250ef14baa2c51b838edca6b82999fa7b6608ac3083afac4a55b6b775b56accbb7e028e8f15920dbab44b28d6e58f42af794bae443f5b6e3dafcf590be22b1f3e2662cff4c7a26649f701c43a61f2becbc2ff6cb15b2a171cdd46b0525710815bf838d0481cb3d72a0753ea99dd1b438d7496c1e604bdd4519b47ccfb1e62ad028a0d9a9b4de60d5a9bc9b2f02547b1deba05977ee76c2a25d1889c0acf5a38c09b38f2429ed98a9e21723bc65f6008c5331fe6fa05a629cbf2667f2a6e001fd031c97b2173c4495a6538cc5a90cd17c56a404783ab5e35af5ece75c1553b00d3cb08d49cae6b65980c183fa9a17bc137d36089a33fd3c56f63c0979cd077744cf1731a04c563c50de0e3a50c336b01355b218ee97df6b9eaaf4b21b8ffa243223d9c29e8852d9d96e0330b978a8044024d34196981ed274717db2a7141f15250d3f41b642bc2dc43ee969ec9af48a9f1cb3698a310521e189c976cb4ad65d3b4d522b702e285cc753e18b8b70a5d085a764ca987daa68b7527855fa60472ef81eed276005963e7c1ddd9e36401ba7426278c44e8617a92fc0a23caa8b2cbb726745f633074ea73f995438f00e49b3ad2e7cc29461ec4410e618f6ae3bfaaeccdf8031a30217650ec9f8d1b31c4bac10ea370555050bd771cce3c84df9215a4413f49ad697ecd75144f34c45c6f2b87d990794c7f550e50338cb5f843b88de62c5708a3611974e077f505f740b17178a625313b21b7b6d106dd7c0274fcab339f292dde6066b5f21b74d5957128e18335c2b627e8e1e7d0829aeb08a5810f7707e57ba3c58b33cf9028ce89df4c1cc15e1e241f6041497135ef5cf1ac19a24292e776a41c9be572685e3bbd2d148203452a29364ea6a8750b40ed2a62571fd3b84bbee3ca654352edd4ff9d16407640a8cfb371b1f944b6f80e9e22754944ab6004f782e6ec7c2f4e3ca9364654e9d84687f44d1ecf903f54f9ebdc1a58aa3db4d94d4a9ae398d3e89997d8cf76b7bb70ba240527c9eb3bf23caf979951b2c51c9145b9c2e0a8c95ee8ace182713712e2e93ed1d596e858a419229940259c887833d4d7f42445f7f0b6c8e16938afef66084f1d4982d643d59dbb5fe890966b67309a66664da0e8b4c9f7e0931ef27fec69da5098582cd0e908abb924946bf59add7ffbb8e9638ad91bcd225e2a68f4ed14567e6c1254796b3bfe61f18c21491898c36a65dcd2cd7e0e10d28058e55f3105e25e5964e66d6d68f843f1be07a2f5bd6ce821efbd0478a082f282a883f90471806a5ba1443c592bf54a09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb5c92add93ff494bfd7c393b5afe43f6ac36d5f30b9d4c152dbf858371e16475d453530fdb62684e73eef1a7f845473215456eac59de55aedaaa359743666768df44363077ee455465bc943ca98939e18f4aa3f53079f4c65c1cacc60099f56a134077fc5dbd0037db517a9f84b442b60e2faf7b166019b42f32a78a28fd7f2c22729f863d0279437d7f47954b73f6cd8df797b9ba20cea5c099d7ad3c5944660567ee2afa1ecd282512f92666fb184c055a7c2e17c49205e202589badf112950313ee98f29d9fa1307c4f9ea2aadea7c8a426a434f7b0fbb6bddb2295066c1f0eccde7e87e6b452ad3393f51968161aa227001e9ff7c3c4478ac1b07bf9bc10801cf3a7e9d0e32eb8cd6e52285a98371e4f09c4c358cca3abf69ee75c4c66ae372c35d5885094d82fa6f5abf4fccd08a492fdcb5f25892b7dcbde5673a1355431826c482ad16b7e7d04ff7a9cfb68ecafac4dc56ae5fe9d7ceabbbb656d1da72ccd09a635aafe215ed39f6ec34f85dd787a8f53abc89ed2905795fe60aaa3b9f6692b923475453a25114165dddb325799982aa8c52134124ccf76f8335862c5e6705ea77898d2d13c2e4826b54cf626c3ae02dea48544086e0a0238193530158557e940216c680bacefb4da3b4e0495ecd88648cc0eff99cab6cdab3c0b12349b68203b50a87084fb6a2f97141f45f9cd08babf3f27a5731a735d76aec31122ec660378015965572d56151ff445f794dcd7d4e4e16f1bd86dd406a5d3fbca4202b1d8e6c656049bc0c199ce9dabe4ded5e7c019c32faaf845c71062ba55e6e199f681b6181367fa85007fe46dc3f5da258ac12227ab36c736fdb08edbcc52bbfde0e0b3602669ce891028e93cd83a21687a155dcafc255fa3b32d3e5d68d882da4c40e3fd5c30164b6533070ce3467f0c85b0f34a4fa73fcfb1d52dd08f5f76715662ee7eb660be6e94e6d7904eb91be74a114e388f89063548ae250aa92c676be593f9ecef2aae26e78cf3cf217bb38540836b1a9279be03e7de0b0ed466fc6aa33a84d106d37b704ddbc59ad4da575d1a99ef76b53aa56e888f6c72de712e440b69ec4bf7c2109c94c9f461e0d6df1213c0a73cfaf30ce520d68123a9b2b9943b4840fb72e868d1923ede5d6cc1d45706c75643ee92cacbe703319c8ef8099e9f11b4971d5633a67d6ab8b15b0af1cda4c2541c06969e47c099feb934d469b023077f6b3061f5780906457de2da90255602c13d1da643e9a57b36945c28e9aa468c7c0c3dcaf9f400583ea92eb41a8d5d42e5ef1609609957962a4b4fbd8845454580a018447b7fecf3d0cacfdeebc3a6459101f2a28a20e30315a91cdf2932642685ccad0bd6162b581fbfc06854381eee308d80976aa9e444798539e2f35dfec806c5134badf2f6e042df1c94b8383de28198a1266a91179ac47aaa2c42;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha9ed19dacad98d32d9ff8932d596ed4b32b795349f21b3a04e7bb4f56413be713fac0d1bf72b803e3c50665525daf6eb0e5379e3e9f3a29b5986d15ff95b71ce7e8b891746f8bfa842bc1aa5975b0c0c784c9a91cb47b51875720f5db4cc5595d6d9cca1f92b7150e3e9c3236388199a5cb7da7bf1be639c778ac8fd0c6daa7ad2976e3e3ffd9e33f9582319c104f27e62240e2b1609bd5089b90fcbd7fbccfe04cdc0726e154a1dc250226420ba21575ad4fe39c18249d04030f3de2f42e6c41179014bee391a7767bf94d4326910b9ca886054303d869a8bf65cc6e36f4b3d3fba973df0e6ac6d843cc4e836bcc826d840b329ba41e04f780be44ff06d9967adcc7c54b640f520e8108a8e645554d9e3b895b5e5ae6c79d7db06f18f129c33676bf79d6e5b184776a7d906d1718cc35bd1d06a6ddc92b26737455071d0ef644e9582da91c9879b7f7436ef055b8e85f3c1b162918a54751ca162a68c9968bfdb236abe3168f0f07f4d3349efd07c3e36c877fad3c1c7ea27c4b3a469946e81573896478198a230addee83f73c2bd19a0e026e9fbae4e7133f4c583c78ecb236f5bb916d43be74f6a64becb16eaa7ebc14690656cd0f1ab75532e29185c3867f9c33826a4353ece89f20ae48c007a510e227b575a06e393e052ef8297694c81182fdd586a0b7de9769e107346a7b6580dac9fd57f53de65fc8ac6c8ce6e3c1afe9095de84cc0b41a480ae9235a853706f9764cb586f1cf43694960da903f717a62e43698ff110d4b37a5b338a23fa050a5338c1ddd1d50fa111498fe70750d7457814dc2f804af19d91740cec521d9f21282c89fb1269048ff7714e9a18b7aded4f4a48b43ec8e8d64ec7c311623fc130a4d39c4d286069292be1119e18d3e49826d7ab0b179a9da1ddaa71dd8ef32d138b15e27e88d3320c48775901fc45c8fe8af186d1e24378c28010e483f5ec6aef4079b3eb1da7fa8d4784cae90478f8b07e7abc9c0c2ab94a40c189c7dc5bd6624f585bfda3a72ee9d6d45190b2a609da7cf0d4e00f05d6bcb81d11c9b7a0f1528c3ae2bb774e7a192513a9249a861a09c6a87d2847e0d1637a0b2e551c83aa3174a513417fc8e06dfe8c47672b377645e946ad5a482072dd69a8f97ede6507ce30347f7e1e3c0fe753424c4bf41ca03b87562c5ff30bf19a83f0e48ce3c55fd58dab9a78d6e5735deda9c328439067517d6c0e58fc3283853b933680edbf6317848707c87690edb306e3734b5eedb0718f16c98b117363ba3ab911ead63e773c182f419750f92804d4cbfa198a1208db1265c3bc350eb65e3124968c2dbf8c6858bfb6492c9f04788be75b50cbe45cd32ba8da59f9d489c20d427c176109f2bafba855b99bc6c51f2d32dba2c58e85c9bee4b063ec0448ed322b0f59136943b4d31134d6886bd097e431c45ddfd537;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h21b424f51212e70d5996941ef7014ef61016a53bec9da5737a97090d44a88aa1cb9a2b401de391c1a59c30d5b1dd91323885a692adc19309809116fdf6ce0ee24d99574c6e1b871a2c4cfd891f554d32ba9103ddd1dc502b202a6834504d1aca88cd3c9e122772b789738fb06d5dac39ea1cd13412daf603454ece3baff7f1f0cd7da6c0b555cb38a2b778331e633112422eb28ee2648eaacf47be2b716b10d87ab7024df8109f46da75e199ab3c00a858dafa0b02e515389700f1eeb447a3dc9c3a1e38ae1695a30997d7ba84bf99c58f00e6d4d06028e51f2dfc479fadd4982fade5866486812bf940c51dd29bcf31c3d4f40e1e44cece6b3ba7d1f9491bc4f313ffb9db75369dadb6b92cd2e863455060762900c7116054654297978a2d8a509791d5d701ec10ba133d82f631f8ae2685febcde1eda2f86236175e9bd17f528b424d012df56b6012c6f34ea43f35f465f2bca69a358aa9cd83d0fe991dd1b751ff1646e2fa530993d124711d07107c406466eb386de3b6767bf1c36a1bcd5f0ecdd7b26493945668ecbe2ae10fd8778ee3d886231ceeb4dc065374c473aad672e9f802625cf3aa506d03cfe0e19ddd48d9cd0a99854fecbb5f7fe88ef3d0caff666ffed9e3f5c71d89508389166767de80829bb48af112f2cae543863cdd661d2f293632190de1032aaae6d8d0ac80bc23604da425fa67691dabcff22a0302f7763bd1741babed6e423f3edc95397058e890c69407da915934251ccd8c0d24e6f5d867080a3169a71208e6a8d2aff3a74878f1994fda7e60c8e3970b00dd9a482ec74e558f160ef30e3505b453de04018284685650f390c4ff0e03079f4cfc9da7ce5dd6834d8ee8374fdedfb8c09d60cc3eb901e1f6fb5baa1730140993e3d8aca3ad35ff4a64e45370f31236a9afc875acac54a4e163d64c3e7aea677f9b393499d25bb3861c96ca9b20f85e58894897f9d77ba0246169ffe320cb8253b0bd1646eb1084d5c241746ee5a9c16bd1d7d4dc2c65003be26396b8ec32e78a608bbfab3ea00f4f16473973260c9f297154e6ff584e39816b48ec7aefb6fd3e2fcdaf8d9dfc50a391bf0aff4bc73713c92fbcc4a73bcde70fe8c442477408bfd515ac0cd3b29145c4cda05a54e8396789614bf1248927f6299fd721d7c176c5f0f8e82a69fbbd29d0feca5fabf7153a57d2226e462b1b07b0d65cf1aaf38188d8f025b25219d63edbbaa2094b44e97654440baca9f473265f73afdd32090f178283028c8b244b1ce8cedf3f7c98b6e751f2600bec5beb02cabba1a3ab96c5444dc4d4c4241995f2679d9791b5b6d3174d907aeb3f0f130aa072c25e702d7b63aea31f11f5246adf0a14778dffc3b02f5b29cb44eadd19a6e5ae4c0aaaeb90f6e895fbc1b12379a77e0c215b7ad11a95efc7f6cf524153f827ea8a535aa73c5f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdc33087ea49e179cf91e468dc50454efe228ef05c3a9dc950be68bc1f08bde1eac5976ee807fec8600e71176f079e6bb5e0e56a50770033d37d5eb2d9d9d9933eb0d3d30b97c93e243baf558c3727eec6a2e6359e199d835ea722b20ceaea2f51996e16b6c26757b7690c39d44ab1e015659115064e12bab5a96df2524c0178de64938dfa8722c3623154e7ad7264e6be4b967125746a33c75c753a063f5a50b067772d27737e07173fcfbd2da9654768237f04541b1f658d22b9ae85591974caf2c162b289bee795c07b0b37079d897f716d24c422d1b65dc4e2aef1a98682e21d5aa0b84266410abfdd60890ac1c9d3ff5c4b71452c7e015ecee1aced347ad1e677538910e72c12a9a9381e4c19ecec2ceef1e41c9773e44ab57fc774fdcb408ff38814f183320cd2bfeb737891382d63512689e3b5699fc57d95312ae6d542aa71a1bf04f311edac094f2506a53d498469f412e877c5dc097d293e54fb9071a64d0a2a91a12d7f61791e32101164e6927ef0a12051e6f09244c2d77bd087f16cd9918cda227f844f002323536932e12abe264d625f79698e7cdcf40ecd450590ecf28b4f06885235a3850bf187a5a28d38192cec5b975ee98abd273c026b0415cacb9fe294603cd5436f49c1ca06f9aca3a2e0215322256ebb2d1aa3c4812f56a759a6ffca623eeb58da29cfe4f6bfeb00a7561f82bdaef87fed68d422cce5295c4cb2ff9b43489d6c35c673f74d4738a2efecebd48888434916266e742fdde8b1d3b0bea6833a5807dbcb50bc2eb4c737fb7e0d22883631eb4f8d6e573d196c774158d773ed9fd030b602d9f7851862f428b8c5b18c3824acf4550da1ecdfe2b1d5c68e84f389f2256d52ce2835300a2840779bb5ed523f7905c2d37063251f07500a044bb05980e0cd60981852e511b3ba389153ca17e28f0b79622c243b44c08c9c80b8a08e2dd0f2593f4ceb3b885a44ef035a7a6e77b56ebbf74aa79f731fc3885d0466514b948b84e2a62b1fee9a4b8c585ae5aff59f420b8ea4da7d3b08183575feb482cf8ec6857e6a2f5e6151f0ede85aa0ebd75bbe142070eb69b2e27bcc0354e9bb1cda42313d37b4d3aec055e96d5c313a972c65c0a6422f47ee14fbe7e9a6f13d7af4669f1f54cd1cc130f72a6130d6bfe14bfecde511562fcd8da9248009bd804b6549cf741c38b9618901887c55dc7513a0b640b0bd7f549cc78ba808161fe27d6d4d6f99dcca727b65fde2da53109e35104383f2c6012d3b47e81dc03bbb1e6bc858402d1248a4cb77e96b7296212322d0f2428ac2630012af50abe6fd343742b805fe52aa1da2fa4d07f6517986d934392c6d666607d10b3791c337b2a13dec1ae9e6ffb6516f100267186b5f7e7965bc79695e5da9c2e3c25304da5afe7c592ddcd2295555e2cfd7edee2fde674dc8c6f0ffbe9fd6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6f8e646f12f207c2ba8c0453d23f3872eb0ec4a1671ca56e211cc4d613d68662c9036c2a23fbcbceab640928fc244f88d53bd2b076874c33099075db7b58b626dec57998a2342225abd5a07b771b9a572acac9c6111fa9d2cc3cb0e92f643b4598bea13b952fd2d0671864653b4f0c7bf5906f94263aa40c7f378584c1c1b43b3069c3101b78b98fdd316000b6f197c25d8f643602397ae9cfc48fd6aa4ea4e80bb690414f8137df77f4ae5b99486a5ba7edaca32f7d416a090a4ca0cd05c3edc8acc1f26b7d69d7e28df43dd7359026ad647b93bf353700f6e728ce3d6ce158acae81f28d6082cf9acd9d3bf403740f1d0adeb1f495e64f0e07b5d896598d90ddce0b54abf2b9ad795a1e15a9db64f33219dbe2d20b5562e9b24061fae6d38e3fae1cf47986060e6467bccffa386303e10db3bba1b8b8b739690819c327dd4e9b3e9c98aa52687a314a8a30e488e68bbc60d7cb47a19fcedc5bf4979249a54871906b526f217df38460d9ce311ff731c16965226b7aa77007d68379c976677e0d352d423b70f697be3706ecb15f0dd8c11c57409db92f17a90f391b05dfbe75423d5bdf436607caf68741cdc02a1c6f87ee7a5ac71a8c3eb456f311540bf9343b4ff6fd6cb95da86a6c463f32d7fcc43b33c2bb08e4068c7bdd98905f4522febaf258b90dcfd44bc36706819cc26c394182ecbaece1475a29424ffaf6db77afd1ab3c8dc57a8e85bc7a2bccf3ad5c9a56ba90d30d583615333dc510edb7ff3cd3477541455cb048f06a45c6362e3b5436b452724997839d005684ab617a7edc81c7e1de22a562d225f5d089fb7866e57794ac6a234689d849e61e0a87401b61869b4267091c0c87210070d58427c6be2bdeaf38b0a34b98189e0851abf9b40a065b565f27beafebf1e67fba666c17045479ac2353d5a1e3abb920ae6b8401ac1e10dff6cf165ed3b69a50a6b2ae6a1eb78ad0c5a0b3327ec3a91f225ee8bc6c1881749a851546030c98576155c5de275ff04bac1254ad919578b6a3259a4327a8acf09a1a64a9a78ed8c9ca5cc8d92e9adea825b1377b492dfe280eee1f84f00baf19037b8dad17ab7b4357251bcbc8809cfffcd93e5c9b741d0c6aaa460c94aef2c56e5d3c8cb8180f62f12c1acc3006191dcf577b82be799c16a7db6129e7da497dffef960f4c974a466f901bc24b6fb92d61872857b42fc0dc6047579a3b2d98096014afb7761d25dd61fddde15f4b3864c1782a8983c54a4b7bb60f1dacd7edbb50a83ec49fa42b4ead2d7ff4c0341fe2b448d4432681cf52579f095356fbda4e540cb4e498d659479b26fdd1ba32a594acd29673bf847b8d62529b7d2c14d61730cc1d71fdc5e3dd4e61912ac845287949aee9a9615b63496920eba3fafbfe751feee2d59f2147935bd1900ef815b2f72293157d90fb2ae7277bb406a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb34200b0ed46bcde2bad1cb478105874a57d7d09ed544763464d6ab8d6e942c44f27c71559ca5469bfe860808c4a3790d1fed08b4bb9f6807961f6bf7627f68cbe3c507a06f5ba36f989c2e7e941e59666bfef6a830110d93b1b803ea0da659ebda3bc4568663ec320989b897cae454be61f582a5d8ce36979a4a3af157e4923de998e4faa2aac465fb8f1e2a09fa424ffa0290c9cf9b6d73560eaaea1dc477ddae2913705648c3eebf33fe3ff96b607d2afe8eac6afbdea96c92f04b3bf94cd3d45e221d6f5e139d7d0c92202d214e9590f61a3c2228fd2c8aeb438fca91654f0d90fb373cd4cac5f88ad882b8e03614d1903f204b934f91c2358458a33dba455f466d581430d1f5c084d79a2cf8c7504aaaa04fec05025433a8fd0218c63d9c8d657bc919b4a8d6f250f0e5ec4c9cb150b955241070877c935c434c2d8fdfafb28f6b0237492878a30c68c0248f84c097f9ff312a5ab5bbf55603091f483be783934d278f9a5ba16e6e26ad820e42a7792bd86a3877999858205b580f741b8dca586c3cb83eff52fc386f67ea8d37c5c60227bf973ab27c37553b7a93804d8a889971af8ea53e1b7d402478d5206d8ee896be50227390c9efff37f2e5c1cb6d0ecb4f4ab725dc558384821649298bb0f8303acc947203ca22b613281d93acec4d410e02b13b2cfaba4cc46bffbae2789e0f6ef9a7441c01d5ce2128d6c88e4d9b43b6c977a0e707975a8d6e3c0dc98983e6ba0049244c1c819f2a7a7811c11272490cc3ae40cbcde23fb028bf3421c122e9cda330608f46adae4a72ba18728dc1eed2d2e986c6c6aa36344b428be5ec1a8445f6830d755a9f8a3802f6d51c3407f20549e8c3e1f9bfeddb29a38c9a0608979876ba2a49d8ad9fcd47ca0a225383d5c682320e5b14c2886e056b456e641e37bd27879218cce6823fdb5e3cab0bbe7b21eded51f1ab4cebdfae49a0f4898364adc6c17a414c237d841749b50652c39b9905f9bd77498a61a15a57b8c24c5915adc12500666c353a643fc28b33ecbee7bbfc0939162b54486579187dff0819a61ca5d678745f8aa311ffac277e9db74435d8fdf7af19716a7e50127fc26422157e62964a2cf2609d3df1d8babed5d0675692b065823ca5119347790de6f1e98503de1770f90a0297624b93178948dd11db1141252ea9a9494accefe307ec478115ed0833c1ceac9619b15d91eb3bee79341176569089bb99f91da3ddc30d0ad26fe9927a7da6a10383dfdf7f1642d53871888dcfa1c08873d402059068a31d6e5f824c831bfee4488766fd71829b4de831a188ab971d29f9822b4ef23b4fd5d87bf681ba62b9bba282e0932946d0411bf0f2d1d732d5628b4624d16ca0125b4f8b338fda6bf66e88e8666cce45bd1c032802f5edc1e1eada0b44b57eb99e2307830b370bc5226a9970238c45ad3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7e4facb184ae9dc06c766a890aed6e55d85ad81014510971098ac838ae21ae850d7e02de048e72be96e80347dc77f835e56c3a3097e871a68ebd68f6af323145108bbd14113b84672f0baaa79bac38d082943bdb4b29410b4d5b49f978f1f41c2d109bae09e087dc63b7344d6dff4c9893e3c43e63d20926a7d8ab367b390d35ed4ffda0e86c5b6c78b356c9d2bbe3d29a291364501cf164f9fbbdcca575c7dfe2df6b2a160c427ff5eb1378f9e0ab549642e56a74d1e0c236a649caca508b73759959d0cf4648ab47ffbd2df403bbe14b0ba44d46a26139c8d14f6c6130ea00fa4bd0f3a36d7fcaf2c27a703b374aca83f2a068f272cecb3311d82032d1769a5f2e90d44ceb241821f020c64b107ed99feb42e976ed046fc187f87548313db454a2b5f4648a6c2a815b4ffb5fe1716ad8e39fa4fa8e9a75f17b1514cb61712b981651bfb1517a5da6febc5ac8a1de6944812ec9d9275962c030bcc7489a3db88ec3708e277f281684dcd4a09388ad99b831c1449d3f6a462d428e5f0023eeaa8af0b8b10fde15c978d3a4b08bd17c0615e1b7ffd706b9891af6d55679eeed5b1457c223b35e7decd44e7cd8d20fbf94442c19e57c58bcabbe9e5cc0842e14235fe8a2cf83b9305d433a5705629165a0f45c9eeb75630f25a7399ff50900d87ff4d728f1238010fb55567f7d9a024528f1d32d01a825a1786b54c0b3a909d3435f23e323e2df34380da6197b684080aac9ee662d12f8934f468f173f020cf9806d6ba88e2eb2ba469e5e10c37adc29c9dba77f55a3ef5fedc08f0ef0d19576aa881de71e39c07c442518f41b0e54800f8a4c686ee89b15c23b99ee1ff3fbf560045c735c35cd09df49112035b0e12b391797968ec3495417206848c29689f91292f43405509dff39dac1b06a08008893e39cfcad06b7f77d0b72abb1f574ec84c071e710fccecee38b464fa04a8c742c44958e232fe40a73f63f48c9c84453d3155e801cf3d27818aff75a78b5e9743b6a89df64a35c1556fa32257f3b733484128b449838904b5b1cb0901af06ed22a98f14916b50d72a4bc955a5dd6168f2a9ec4805b827c459e83250bfbb100d9a8c148ef22642e0529dc52ea58b7304df7925e4e014b4a30f5c2561bc1d47fa2a0adf647fa0045239c11af056db93efd4e552867da1a5feea3c9dfbf4d3024c89dd7271e8a89794ced26cba15c42e827d4d3ebfb8458d3c94864cf497c20f83dba1e306eda81743528e106e24dbbed052a5327379d9a57ee5fa64e78e83b60b5311251621f48400054564dfd93646fa8d12e0e01310806cd5460610c333144bda67735a68c2ca559c1e7af6620be17d02b0c632dd3425b1a2a0500a10bbbb4d1353cbc8ce486f298c6536c6c209b4594b147444cdcc11cd5952b825a9e81e8cb222df466c90253ea8c5c5e6d32db88f666;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1da1fc26ff033dd94cd271e3df134ee1d4b372c1ef53d4b9fa9010d2b2e9a0598bf826f0aef68a58880b97587325105bf5ed4258eadbd06f3cce719e6996f79213275b2799c2464fc7af72cee617902f691701b2435683963979e7b854320d238c49486cfeb1fcdb0b5f0434872eede8a474aa60c524aa2341ec79f943cfaf980aac1f90d3c4f43bca3ba13ac87c4b08ec6d772ddddf70bc8302d32b7afb6e551ccc19a91015137224c76c64c70e7a741e706c876d2cc5a9672b8b3a6bf7954870a78d7b73f16176b2c15799f870830a2a9d76bc7c8a04da2dc452f11d9337d73ad3724f0b2bd4e11787b3e81e7078b21e3ebe9ea006798f9b5d00599d31ebff02789514ed560c10c425c6288677cd504e3527f5f08f6249903c054c52a28da013c8a1a5ec8cd239ee697721b596cd2d012ea48632e1ec490bd08b2b68cf29b734768ec278dda4cc3f17ee396a71a0ca176df96b6fa53201235a3a316b05d6bcc297a7eedb5615462236a89dd1c05e780249cb3628cb55491322d95b6f6d9aed99257d7aeb04ca5c07fd660f1ae322ca700b225cf558ff60349eef4a6f77759349f4d03efa0478c8fe9791d268128a419c1df5597878ded140774920bba95a73416b4721c238ad7a7cbd542bc4db36f3f2bb50848e3622dd29198916fb9aebf48642c7726cff0565a0233a9ff3b3656807b6dc8abcb684a6a370ce48769732c1f2e1991aa1274b0138ae08e266ddf548aba05c2ceeb2e90f0a330c85e59567297ca7fadf6dbb6d34fc1ad32e4ca8c7a43682122f2cdb25e2ff8fa11f89f6a5e217da469580750ec0835d8cc7943006496912a24f65fd140e91cb5a10879406c6b6222d42a6ff798cc32821a3989b9e21beddfff64428edc66a899574e40a1f4cf6dc68dfd8e54734260db066954826610731b0a3ea3c5e89a22bb1159bcedc33a890f75248df4c4c18bcb4ef79b7f2e601704b10e3525cf62f10ceca67928ba9bea62b62bce2d627c0cd55ad69bb0eb41c48b61647e07f49f0b93c636378fab31467d0536b02583c796a834a7cf50cfdda47b10710d732bf94d8d2c11184d30e6b344277e5ed45885118ad9eaf15dccdb5e62eac4d0f09d8804969bce432f7b27af6657575e4a592dfa11a6e0d601ea49ce55fb4bfefd3d64267052e90ef0496a7d12862c5d8a71cda132da420605444a8e8601d759e151124c158f72e26ad158c997d4e703980b5651ca92b8aa524131ad9d40324b6c97e323730c4e2682e264f0cf4f929d3ab4ecd69fe1fef711058812750f17be4276fcf7e2b49a2be962edfed6e30ed7b07980c6f912e1760f03dbd8c8e0b96c69f3b13108434223f812af4fef8b45f7327f4474b3dbb0e2c49f3c65eec451286b805f1e17405eac8b625fea70d9763b59b1427455cfb8c97049be7fba427f36e75279e2caacf714fa75f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9a2fa733799cd14d2ebf06841e423255a538c12ae684649f9d70eb186ab0a719754cb580ea0794f03d368977a97bd2623edb9278593f5c8d136c35ed37d34466a2e0d2dbd087828168da2ccbaf46c9473c21fc504ce092bf591aa374039dcc78f45bd7e5666f7228649ffcde7f4b2bb2e4d63fa59f7dfb55a6bb812f678a0dae7628c04a894a379f54b3a74eb3fac875282c0aec9e3763343fe3f526515262f25ae50d7827241c2568222128f0a8a63755eef22e76c6cb634feb77b0a0dccf8ceec8b38860d98e41a3ce9f50c423c2a62a6a9fe0466b415950dd417ede4346ca6da33705647f2ea5d9ec40f21c1a2e4b239a0cf4afc2b940130572c5e8448a89367c188a6700e1915c7a3ee4b5d1c97e3bfb81229e3235fca330e041b9574d90999cebee9dc7e857c87aed31a546321464c2a80192972748185538731b44c8aead6146677e402d3d2080a06e6a6ee7e6f3d49cbd9f852b5b3c4c1d84480980f7ff080eecf34442781a2f394370de53e02a083bdecf056e139fb6d5a4885a0f311feb73383c4d395cb262f392a7fd8ed2a8cc130dcab2401a1d26f8a565f81deddc1916ff848508d6f582579b066da3747396057bb2d51f3d3b500a0364517bcb76af99b9b87bf26d1453a56e8214ba808bb2846f058a9f4f2f47e1f9d13b85673bdd01dde2df17228edac1ec1abf485c201dcb9ae944be190861a745f2bf2f07dceaa7697d914174832d4b2d6ad0ec58b0eaa7e29ba3b1e1de6fa1abc18b804c7750eef9deeba8927b94149940086df6a6edb1739e6e7bf6e3f09eaa28fb830e4a699e1e556d8e2fb90bcbe2a62db4027fed22cf6cc86aaa07642cbc4284adfdd4835b8237842662795c7dd364e22315bfa5fd329de2def9c052fe442a479702628c9a39d66830efbb326ad3c4e6b80d7344d1f1fee535b010955d5f7352b67889d65fedb9ac29f6968d183819aa1a78a0ea7d15d70fe544a4ead66d2d646a21622f8bb8b4492fc6217e5ff0b611891b091e50abeff4afae5c6773c8b678bd05ff43ffd62c3b780ea78c165e8e4c779ca2512eaaaa18a83ebdc339e6b21a3e20cc22f99ad56861043b83a32cb8d4cede171c4b1f615f807e256f4a97cab58a464574a51a800cedc90eb9494ce0b6940113dca2120193f75cc53d2680f8b66e01983245ac38ba364fa9bfa7831729964992b27f0ef6a963a266e340501c2654df6e0cddfe8f522b856405ecb4b6b539fab9d7cf18ed82ffe984b3381a997331ccd9a65b697881341d927028b1dcfe8e3f472a07aeb800756e3e7f70d98c43aeb864434beb66c8a69ef2e93d23c995d6b6cfdc49398624a595c879805ff793ef2e90d40f57d382c34e78be4c41128a37f01808d00bca8357a3e9ef984bd5464486c9a892e0a22b7bb1a521a3a37215e307243b9ae3300f9b4c803a86820f2b6126;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he3456c23fb636985a46b7675d31cb2386416d8af20a4c6044fdfead064ea82ae74564804309890c80c21d4c39365cb4b061e6bb671af3fbdafece53e8f059ce94ec232d5640a039e81e5317e275b430ef04d58631c31bd4101e89038279b375f7b4df3794767b1ed22abe616ceb4421314b3dab3c637d42a32156b14712b0b61a1bb4ad455c71ae99e9f32458c45a82a67ea41a52772f9816e5e5cd7094dcb64f3069d9366e661c77fec1f14b08fd5b3a3805045e1b39f39d257c9a0d15ec108650aab256477b7151f1a9777faf364181d92af7fb582be5c1a4541fd54cc97cbb7cea01a9158d8c91addb63c30a388413b479c8f74960ff0cacd35bd171c16af3ae69177ec7af2c4bb502f01cfc416653fc6776e09fbc07c0ba8250655d3c33f4021271e20bbcd80d0ef34c6fd3a9c78f36eec2f88e12e2159c4ff40419ea7af27ee0747e66428cffe92f8db8833bb4c26b03bc7eb736a39cba4b473de7544a4b281c5df79e678497f8e772367d41e982dc9bce50b6078fd400fd2701e88b6397a0a2fb4eed2bea5df45abacf20a770ab90d1300d3572cf96605ec0a322d3be752700fe4495290c6a5a55cce10a8de8edbc4c470770fbd6c49e7fa9d1884c8e6e8ae2f28cfdc28fc39a02105f3361f0ed7bfb194aafd40354fd1f574cff4e69fb2b685103c35c289101e7188746e7b99865df30d54bed2470b62b15e7ad5083c3a73181b3947c5bf8a3f0f9432ab6c4fb650736a9adb916341008955745d7a4115f16f2306c1938ba8cb19840f84338df780b7816e481a526e187be35ff7161e4fddbd8818301656321741dc7edd3f17c4e89a7daef89d00c9ac4ff27f17175cfc811185952221bfc13c3003ce1a7c7132408ecb97eca729f5762fd79fb57141c7a2b7664935244d1e377b96701ec46318f7b5ddd481ee252165c8da685b0324d42d162a530304374629b1ed0964658c291fe89dfda4322c27f2174ca20d5bf2476c217388870ccc06c6b8b2770e3d8bb6251f62ed85c70e5dbf9af55a5721b3e9bea20285ec9c2a4361774dfdee4f618b4b3c3a30bd0e89580cd58f5e16105de140dab2a00f3caf2951b968baa5aec6ec5e8eae6d204c8d539a6134bf771b00dc6a9846cc5c61a2739a3b0a87d4daa90eab208219e11ef33f70fecc537ea68605c9a713e24929650ac7252322feea496dc10041785d38251a6a257dfbbfd6ed113e4abbba88758e463c29c520fe0e00ed99dd8267e4ab63e7e8175cc88921eec24628973f00054dc7a69fab9d30a56f8e0e788c0f8d362ac3c6b035454ab72d644910f0e3ac2b5abe173f6e99dca8a701e19ad1e19c2a251ed1db85f15376b1e80d2c4494b33fd9a8902881dc876a8425293efd9e926a2e98ef5773956022c2d0fc8deab60d535cd79eebe3143c132da9cd2f62065f3e9a55291db5036a6be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h374a64e6d8160bbacf00bd55ed73def69d28ec028add849219a6eed0b7624e2e9b318f50eac5c40837710ca37d64cbf3cbb77afd4061e8e85e5e29dddb8f9201cb2a42379be72a2d2106e3f3195a60d9dde4a3ab971ced3947194c59da1eea0103db3e9d0048259b2a9bb7415cd2e94d4b6520d5a11237db12a8ee98f4475107225615ad22f70180de29cf87cb852281b3cabb21b716043bdd3652c63b8210a294ef89bbae11463818edadb80a8ae0e91057c0a70ca3b21befe328cf2778eba64b6f865a52f9198bbd208336a824f0ef6f598d9409bd1ee7cd8e2bdbdba680c864e7fbd2fd2dd4028608854be5361bc82c9b24cc8a9eb49eae2375d4b752492734180c998e677c6c283b6729f6b682f90954668bc531d866a9a75306e8875fa81df0c621d05e72b28fa12cab2aada940620b19d33deb5d8004cda0c34e404ca49bd3962cbe4d6c1bcdf01bdf0a24aa9791cee4540011c9b8f2dc833fa04a834e8617f7c1e50f3c35c5c47d4e7f175744f48314b6e177d99fb25bbc7af70a7b4a8cba20454feb3bd059d0683aab30695b5b015f30885a415926ed2fda1df72f81ac62c9efbb1e1328e588551e2f0dcbcc06924c1edf23e5866c5b6428dc0c63467aa767e1b89a42534fa23ec2311e5e04cbd962badbfe8be635c00d6a90792ed3138dbbe060d5e1a63e7e397422e64e797760dd432ff4724880c1d6b0d7dfbee54bbd3fec9ac22c62012976a8ba3ac4bde449965ed8590053d0d815b442c8aaf84cc2128c42631fd21c33703d5957e52fc0b4bdc66f04ad66caf56e63f41863cc7563e98e3be8648e76a6d7f6aab234f87b91c8d83ff70c6f28fc89c0aeb884dcf24ae833b5339a5d7855a5da6d5079cde8d14ec5a3417e42ce9c09eeeb51aca6f0388e1fba38eb37aa595ab6fa6de3634883602831d54b628354a5c8a5ebefadfe8d12a2057bf4e4826007e4f73ceb78bd4ee8055d701ecdf759222bf295223b4609770f98fa2ea403170299be8e5a6aaf4c64de6b0da2235ae5e0e47ad93452dee6ff04cc275dbacedf2d603511e96167bfd2a81556d13fdc018f62b0e6c4d63b56e71e7b11c011f04faccd8f8e03499cc75e9d5b3ff2784bd7bdc3ceb84ca3778ee2385a4c5a4c506a2f1845015e16c60f4a2223cfe64ccc88eeb8c38bd46affde2b8409a4bee9ba56f6acd9f9cfd5863537669635639ab19784925a5c57293b4cc0433ce4b07277bf2789ce5d20eb3618d3934d84ccb894900e4e01125f27a8cbc1cca62dc359fd4ea378be883b133db2341421ef839813171c8ea0527f84817a77c929a254cf8b3e90da8079979fd9b155e1bbd9d4a2c3054be6e86f3d2e33d541a92dda9b410008e57da870ab5ac93869061d55d51a1201babb38d44a711e4ce90c6d651441c6cf280201a75fb5a864491808146398e9439172e403695d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbe96921eb7071a8176f60033f3551955fb3ca500066a4982a61ab69723f09da444dea75ea2b465e3a32d8c3f966843bb4e03c414e2dd1783f1b80637c424759aa66580bac8a12d7e5f102e2783ffca8e6e4444ed61442fb27eed0a13637e637df230f3aec63493be43889c78e9919f6bd0f5e89b6f70d69f383eae203d487136797ccc13d71532d4845b1bf5b867894ac7d9fdfdf7cf58045512fa9b7f3ddf303685664b0ae1a339477f7cf1cb746f063060fc7841305fe8bc3c423b6e7f02ee90c4b453a65890db179d8ff5a405044fcd88b995f57b1e1285a872f53871c846962ac33aeeaf847a82c70d7d138bff3d91702e0f1bcf863b4c8f27d5852337c49e2577ed64bce2b385a1f202f5ce7636f752fba4192afbb1ef5df192f403cc7088decee56973010f84b449a6b329f1758dc8d6ecbecab9f5c6a9821f3a9607826fa5280e0b2fe2a5b60e5b44efbccd42afc1e8e2649e3c9bdee50690935db9fc0e7b6f925fc17fb524971331d327289438e65ca09e2e39a33a54b75d54a11ccd11585af6478f0431358416fd2b617394a7b569d796ad921daefd82b07631a46a9675bdd7dc5701ce35e41e0895fecf9a7a9bbd13f39713e71532714b44c0aec0512d7db835035ac65d723907f09079ab0b66ff0557da9f65a7593af371f0b40b44f27715455ace9faebe7a4781304ba384571c473190e08d403a988674d87f25408967734b052854c9629d01bdb7462c28a4528e3d7e5bc54a765b4d9aceeca95ad80dd55e5dc5df355b4c483faa8cf4bd7d97d0a42ecc4e3e302764c14fbb6ea5a5d3203153c60dbacf7005f20b1f22cabb7781b4d2198891bb77d675bd48ac9966a3f05d5a545a28339c8a602ddcfa1f3cedabd052feab863a5591fa8faabb2f16a08343d4a542e6c28aded2629c33880d8bd6f812b1463d9429c9934f10262e8b7742f0bd1abcbecc6c81cf882ba0b997f653bce9fa405947c19f0ec0c7226b63571f7e653ee0bddf7a6ddf36ac3cc79d0e2094548551ab2910a4f1a6c1df4655d922af404efdea8b9e6c093854c945bb9f444f9555869ca198a5cfcda09473e842ad0c34a7858e436553eb4bf78faa6d57f67201f875cf7c99c748e35ff019e4802fb9c4b3fd65b2b7f4e3e284d816db1907794863a78da3c1560393fab5573d89d12dc2db221d3e106c6464c5d6bbe6e5aa5aaa0f2501c0a7e2a0a0bac373087b58705231284acac68eda911781c78f3f614872c983504330bf281cd2bed9b26c1d54bca4068dc2a6a44d61a59b061b55ba5a9371af31f65d866b45fd65663d704322abc8a9092dba84f7fc767967268e3ce63bf76400730caf9ef6008bf2c4775c65e7e94ccd6b19fd9b231361f1e3d21e87d8e800d1dedb550176dd7244fd0212504fe371ad6cc0cb2a53bc403b8a6192a31171c953f82d7f711a39e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hedacaa6e5a378a19cd9a17b81c83d73085569d4f5b39572d8876b357893338ebd83ee3d2a32dbed32081fc261bf103183e6218b60927bd6d5aca140102b36e93fdd67d92470e10f6d7f6717f5ba4ca406eb38754e7516e7bafef53fb0866e74db63d61f611e296cfa2125f78391bee9b967afaa747617dac1c87e6eff53217e8779ae6693ffc4befacb5cf413263b89c2ba484beabe78c27641674a7eb8b148781b96f12b8f3006f7c43f25152fe0ba5014ee4728eb48f50d5886694f98642e500ef238c94dc74be4f392e17802266b3cd964045fbe8832b4b8df57221d9d7c61cfc05911a604645e99020d92cb7437c248d45a71cf23edf9e6e4d34d63fd1184a741bf41732f8695b07ef8a7821dc37f2c114fa42f8bf986d8873da5f8420c72cd947297f265a97e9e6917186d2cd5e4a8327b565119e50045865818352bb61ba14e996c9f5fa1727feaa4850179c8bc5b98ac4ce550202d03859ee8ed7f95e2ae1cd978a8c485270fddfe083cc34aa61a58c07273b5eb8d31d7968244a8d3f028522114ad85f53624bffcc5ec15db5720e0b2305226eba128fbd3c1d8199fcdc7947eae7a6b86df757e7d091663256c6e9407676266ef6616d4a0b9c92f91d9a6a27008805d7f4d7984fa310529ade68a36b26241f09e3b6a740e1528e004a70e1d2c0843b7e87fa27799cd7c1861c91fdc5748f5e2c4d5e86385598fecda2658a0906d474822da5997e8e9aa30af476d70917335832be2adffd33cd94608d3c47e4cc08ebdfa7971704b595437c0b731636d15abeff79ddbf073a8ac8a12f44ced3d75340a6de642403e759091b07a91033dbbf5d1b5dd63d604ec8af6bc045cd1ad7125cdf58af29091fc7cce2a8fda857486c0c427a736ec4d49b85704dcc990f583e00ee48cc8f9ed5bb9d3ee3daff72b87851156f05c3678c3b8f7a2f5604392d9e0e8fdd6cf997954f81938af7ce4cf8799694ca1fd593759c86f488a73656c3027b8f05a5b7ca3be41ffc8799fc389645f0c066992a2110a9587e8cf7ec9834e9b7e733e6e3fb08774c5c06b6b90d5269b3cc8b0e918a8c2a0999667dd8a7987f2671c90dc95e89762b1268d3383809bf74b227b142d036f5474a0f7c4a95d37be4e81960dade44878c375c9c01dbe5e0fec548adf349f269a972aa483ea94ed6dbc478cdb90212ecb81295c39e60434dc941e811f58315d9562a2755a03187f330b5e4fff102f8685f860829e0cf06dc807c2091731226a043f1b449056db5420b0f1c875124b5823ab3c374f04f22b27bfef1e8f4d75dc3a193f89dc19037d547c71c0398c4e6b215b8d1c298466c73915450720802322055209fce4f090a46b6aa603056a803dd93cefeb5814811e1de693c777bdbd6ed89ead90fc9a2f805b6bd8d62d80d38fe6e7d2fb0e83b2cee832dd151ba548b8ff3d0a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h726ada41910e4f97ce3bffdbe93579887dbf7e3bd704c8ba5e3091eb338a2f42213dfa47e7651ad44340c330030401ab09eb2e43d112f6825da92c72e45af32d8042f603069a8a1d38061f79ebd4ad268037b5b96b859f489b7c520cb6573375ccf76165df645f55bd5146209ca7f4aceb34fef60c4c4e303dd605119aa1844b5a4e69f49f6c194f5102bab7e08788fb924a54f27efcf134fd46356f6f1084b48a75edd7c63788fe051da5de968f4b795754d2a55290cfc1ccfb386a4403a1c723820f9c0b41aa6105268194e5144abab55a5e832dc17e388b9060a513f1aba74a2900ae5328c7e36d4a473012090bf8dc5feaaf96a2745cb692da7660ead72c1b133bbe224ad0a9cec1f1fe3983344c0476066c7d1b927025f9952495d148754d9890a433e7580cd4e98ce5b9d35d38ab23c788c6ffcb24a6d238296d5f6b1e88358557b87cffb5921795605b3bd5f2a3528401dcdf366288717459ca308489a827d0f35e9d4f927084c9aa0f5e09069b270aeb257e4e2c6e72c500a7e617100741d6e44d5cd0a591c1dad5f913e7f1e9e5f4ec58b59dc72b7a1b388d22abe0dc93745839bdd05f9b4de5db6440e0ee258c6883144c9d2703b16381acfe7d793a0de91654e3f31143f55fa1b8f5c976048d8b9f5e254fe5a5fda6c065403172585d1e7a1e1b0741e4412009447b8d6365a6979ea111d0091ad6fb7e69787e5bbefd69b6d3251c1fcfca40868991c49eeb3f32ab524e38b048416427ed36f2eb3e5736d64bae0fb47df3420b5fbf7d079a3737791c0c194d171c4e88353093efdfa83948d6b9f22300fdc5ecd863e42d62fabd22f1a9c15d343bc5b8a1995bd3fefb268b825f799f246a92774aeec0163ffbca52f15ec3d6fe72ba00ab9127014c36d3c55cec01f5b82baf7641427685860f5a9df0abb998e572947918013c851400986d6696cfe91bc5f677031fe2862517c28164c1fd11a74b491a8d9bdecd0aebec878a0df2af03abe7bd728a3c2a9761e8326fcd273befd39f328f98d8133c3535dd068d2ea0754245945f9b4d90f0e462b8de63437d0a0389e8f96696e9988fe8cdcc3ba831d099d8af0e37ebf2046fb13d29bd58a78ccce987856b30105866af33d87d24ee71c6c258e4b253fc823df6e1fdd5d2d83b7dc7bd0d313d7ac7ca6e7e30eb76b297e35e4b4528a398d3bdaf5e1a3e335f3d417df9db717834fddf6151b9aaaa62790c9a81a7488d8028887f78a86365e5e24dd960218abd6a7481e3e645e7422c38d94d8413fc27498e0aee57e48e097adc190335e380c34525fded35cdf22cf3de5a25d3bf009d40054248ee3abc194063e1db278b91bb32a20dc90ab7b85710b5c7a5437e691324c28ca65663cc624debe9d56d3f4ce860be9c6444d63fdf5a52e0c354610a93ba8de6af6fd03015652976c45702deafd3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h764cafffd9e96718a70cf4d69314c410adea9ac148e43ee6f7c2edacb550b594b05113e503b887f492f5a8b69c6b11b72012fa59f9f2ab5202481d2ce706e323c272838b17de335015736a555fbd6914c379c8bedf32c08ee59440afc448d409b16d43e924fb8fa3b0766906467711210bd0cbf4e223365d492d12eb3241b68d3d62535e6c6d8343966073f96a77af703e22803a9a42d41acc5e2533a3dc71b5346562ec74dae256ed22480b35522ee4ef3505ba6ae9dbf7791dc5002321064415ce0079a8b41cdf780e339428b2d6c667d46cca1c36045978391cbb3dacd566d583ec0458f8821a0c02d0d2aa05094b6db6ea164cf2e32db7f0ed7d8a2fa102d7dff771d52724fe977fcfc6970cb033326ca0b74007741811f106f27f0992bb0196149a8fa08d84fdbb3572b6f633519ae3012a60a330a18cb4cfae537cbc00a06eede327e94182fb228c2175614c2b8a7f84defda71a4f7d57fa03e99a61963f2d406c45a317bd54537a7f19f68e202d9a0cbc6cbe79112c0747d148b0432ddbff51837488d1dca528d3730bd0e23609d2f4265079789a8e8442ebf4ba77adebe0484598ec5a0f3f8bbc8b112514bafad91c712f077c07bca01825ced40caa70ed167539fea0307d796c44cd9156dcca2a2b3682b81b0718a27cb8123eadf0f518bd81e176d824dd67070eff6f925a1c02729dfe1a0758568c2b154006e65284b61beabb762308dcfaae521fc9aef68afe52b6b7c510bd3ce845de0039004b1933d9c46003aeefc3dea736ef547013c27a64e0fb0ca8fd3f8b1a67899390a694a88c7d837cf8b45f87979c0752d05bfd82cd0b7f91be3c5ba9886ec7b8a164d98b1a836153b3f016955bfb34b4d172b58ba2c66e553b9a2548d4945a7291b67890723d2b195d55f763f049a2a5b38cdf3e1e7a9a2a0c75e2c9c8b030b06040d685f3c4fb3e6b6dd0c1111fb4916039936c5dabc108b0738084d37be00154a4d99509e6357e3aec574953d67232ab07e9cc4f17c7fb59cf58a13acdc16bbcd2af55ef76da53c32cd729e5d9e4562e73fb4b9b60708e6bc82b6e13dd9e5cae7ed0c40de420d103ced79fbe42cae7e792c269cccc4bcc0719abb189caf6c8002964c4e03dfb407ba447b493179c33c841bfb1376ca5dcbfde3e1f3492a2ff759db483ae1da254a83fb26a70f28d3d2cf4512013d7ba128befd4dc81be8931ff51298de790fd86ad80488a8559cbf1557b080956bdcded04106c74854831972a6b29af45b28b3440ae8339a4daec45c86751af58b6823d1270270f5f9ccc3b59e1c601eff14bd041cd6409699c78cf41bd36010085bb17be5fd7c96b60f1f65f83015ba8fd065d3a1eb78578f144d96f47ad6733db6fce67b806cbfc0dfc9c66aca6d56f049e8f44dd83c38d90ba07aaab4a9e02e1a02e604391191dd201d8b219;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h36550c444e78e25b8514eeef069053664798a5a1e3629eb41588b9b2e8626e5ddf8fd52e2b5b15571d61ee5e07f3a3adf53e54f03ae21d1ef93a4fdcad013d05fff281dd7a5247fea41da23fa8c33a509fbe73947810b6dfac12f9e085992058ecb6261a0aa312acd2c7888547eadbb12fa0f63e291a866d2dffb76b0bc6b2805e14ab246c72f31e7ce671ee6b88eae477943946d1af8a35e6b41735b518ac28d420f5ee46568cce0f10808b8f81bfe35045365189d591a7a9c286b9508a340f02e5aef1335fdf1d9ef07d4b470195cba223ec1bb66923350adf1e206e94bb2d1cb1519fe0c4bf5493e57661e099a3a70b144eb8176b9ccabd285190f50897eafd35abdcfb8a139b617c459f8f098a5ef8ed5de7b50e1bd607a80ecc46df23f2c29b27915fa3703860b400aa353c2eb1c6d8766fdf99913fcca6561b03d9cb0cd076dac08e7a7a21dda8c12f1772a4448fea0c5d673164625dea7654d0b31e70f0d4098ee456331859957288491b941a850590c3c2d8d098bab3a03154d4e12761a95dcedaaf831a39a64a468c7aa341a2c860772ff72f429ed1b3d82cd90f641303e5f297d84cc0e8f4a5f5fefa1dcdf27baf9324ede52a41c93bdd1982bac818c0de502b64991cc985a1b47d8595ddaddefbaa89f7dd3a9593bef20b31793976845ab7e6e315005d715d8168f5d5e2e93330987c62af24953c9b0348d674ef1fcf0b3759290925dd186549368d0df1d88317ecb89d56ab60f464ffdfe1ea056c68be6290fadcdf2f5ad09f30c6e151ce5692c75498e60c4fd239f07fccbe353f8952f1dda81ef1ba146f2b57cbf17802dcd8c33e1ee612cfaa604738d51eee9225f174e383971c07f4dbda65f08d3b5e2ad0380fa5057c5d1e3c7054b440cd3806f87881160ceb70b360e0bd998ebe38250b248f2dffdaebb4b1d986325d03cac7d7e3ac96ea77222fa715d202c0876bfb671e459563a82b174a28eab64a4480ee3bd25ba15c7fb9e2c021e489514baada2708bca650a0de5a84857b538cd4a3b783ca5090bffe9ae7a182cc64d5e7090068a31b9f21b4a2129291e1b0ec120f6a24baf2c6b366c0c4c92eeeead8e6de8d991fbc169b71ca9ba1ed2bc13b6d024e9c5ffbf64c0db03391550419f713e7994aae80229831e0e2310ae8a303efb2773d0c69512d6cecde947316794fa40d7138cd2e3712917bdbffbb7086a8c6e88695cac3ab79de77d962e969f36e1ec965cf776285f33b1cf7b7c7a1361e58cd23cb04f64e1135ce32571dfdeba2f40dc7277ad8be0be1dc4e4fad2560e0b25592d4b4cbc92855b580af82f06205baedc2c198d9b6ea156a99b39ea955bbd7cbac255bf0466cd38c01bb982c4ba94dcfdef4add4d3f5503c7614fc180fe0312a677fe8dcf1edcef345191d1dee5c447fa87d0103e010a77ca6243db1cc9a26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3faa004a1fac255084420edb7dced3608796b3adb225e8dbabd9f61ba173d8a8ad0481944765920647fdc38905edd071dc9ed5d7d3336aec2ed376319cbb1a7c2938c2aaede62c7001857f0d9643dbe9eb631adfae6cf0f13372d4b51b5966473c0ed1dc5de96802625c5c561f762d93a37828f4613a9df78303a03b980f35303cf786082dfc923f6b16922a4849951565c3241cb18b501095683bd97ee594842f22936bfb3472deb925fa7af912769b189f1e2ec18b49c1f8c7dbff9504d2f9cb6e08247db3c526fbf0b4db9a5e9c00dfe20a154dbeb0d999d79f9065048596b7aa4c280469e699db7c317667e69ae9091729491cff4c19325373fbc1dab8cca4c1fef61fbedac40cb7b8dcbd909b722b78a616a23adeab12f9df5daf36006d9df4e9230a6dc4e388fd337277b891e43b6734cc53e52d54739835d4e026559ac44708d3a275e1950407d9263e24488c885612b60b47fb829d22f3ae428f7c6dd87316f1db2835585a1e00f7ce32971ad602e1a9f0193e1a4387029677609ce10f0dc85e3e915ef24f40961d746d521994da42c5d178302f89fc2b1c405e31c860daff8d6dc5b7c2b267e08ed396ed4c6fe52ffbb0f705f3f768f44dcf0bcde20d06167183e02e435be0abd8a0cf737835a7b0ff110ae914df1c730efba1528248eef269becee2495974de21baf61deb385fc556532aa85e52ba4a0420bc5a5c8a6e5f304e67cd46eede3f0de798c1cc30dd45df4207fa5b0af6b5bebd0e3ffde4467d75c140a13c53d03eb5dc24a149bc5be886abc118e8c72b233f87eaab9cbc975d9dca3e41f93e43bfba4c4624acd3bf49daecc9f1597357bd7e9cd0405348f7b6fc92b62b6c8c8ff26dbc4d2f5af53f22f59a6b5606627096c6f2c5344340e600d3cb51049e331358b1c29d64d2f7d0723afdbca1f670fcd1cb6bffa780747159aadaf973b42e86ac56fa81ba7fabd5d8d3a1d502d6c86aa333716d875fa5daf49df35ddf4303523d076cdfc782f3062d38b2811a471b156ad357daa623c7278b4559975691685137bb9bba826f710b847461af1fe91215e4dc27b6970d939ffe1c2b6991c0c0951ce845e140f1849a12eac6e15b182ca4a233684e8f0aa0ddf45576f49a310df0f8134bf25bc478f3158c4b0d853f8a345821dacb150fd3e89f2973a37fec7521fbe3057a2e069a170a039f610983e57ac68c3ad45981959da469ad6f014330320c00a82706d4822adba3f600725759b710838236ce6793a721153c4a2f7ecf23bdd5f5572ddf9472a828a4e0a9f59af37e08b20d0d655952fa42deaae0d234d99c1cece51131c29aaa31ad15d04ce520b9e12889a4aea855d9defbeed5fe7f0f5d1f80c2c13b5adf3365cefdd6737864398a987755b0feb2f17043b55d0616ae7d7ed4e724402029be4956c6355b716db9d146b0d331;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hced71fbbce985857a5f7720ccd9eda01a224b69746b0950975356738a9dffbc2cae1af96b050c5a9fe8fbfc7ed83ec84df289ffc5408e1a362d5b95da99c24e3a8a519ace1a567237850153260e4aa403a08920ccbea5598b7a5d79692578b36645d3b4ed16a084b53b87aa06ac2b004b053fcf18b213192057b204eb1f4dfa6957e3b81c3ace8fa9b2995e1dea739b243f44954208764cb1d297f5a4e34e1684af22409c58980fe3607a695303ce5912f85dc9a61bdb4a701b1b36b9aa0ebb1d572cc3a9613a3a6928e831d5a545fcae80addbca1abc79da941852a9d7566ba33e48270b414da98140defe75d3ae1972ebcbf7db4cf8c4fb1882bdd15348fb48be5023093731aed102819521a562f5305586a179e2d3a930d64178e7639ef8b325b7268e8cb4fa4890126007aa3db58e6d9fd15288b52c7fd194b4680de0285e974825a46e0d365b04f6641041c3c488a738952129e5476dff5a7d8b03831d346d2512791c4cb4d8f45001aeadcdbbe5c0c6d14f97d1c09067fdd5add6a03d58218eb2b3827f206d65d81356432f6e823c2d1c62bf227fe149662e625fb168e84fe2cb5a9fc2793d2e54d1feefbd86f5f4502308b1a40534ef95d84ebbc44f0de0b7ee8b28b8f5aafc7f051c1faf14250612a64ab22700eb8c274d3c513801387ba58f9436d70db08670f0ccacbf10f61008ea4896f0fda645173912665c8f2c2ba1216119806b1a320e77a3b05b8212a3f1b0d1648cc0127020a941c4949c52828ea66250785583816c59e0640eea67cc9d21516901862d8a1b60e394c295d074d811c4c8cc5ab7a74cd613401a5c0488cc395079248f6a94fc1cbf45995c65cda1e1e99e31681749c7e01f80f2bbea9b4b77f0004557f68f95419316c95db15e598e4d41f1b736f11e43a7d46a07a9332af84479fc6833cea49d31577e2c5b15ee2264145ad30e9f3b18924812d75df642b3caa85b380c260046d6db0c544da99a20cdc6f47c51886060d1341e3bcae35a5a5f5c882390bcfb542399b57586240e287aeac7227ba06e66067df154a087566fdef1214867e20934a3d4444c3c6dec7399cc8e2a1333ddf623c1f37d8b64c772b164e4a5c4a06d075c66a2265f729cd629f1ff7b201ec7e476e207d6d218ff9b1b1af2134b18039abecb8ec9639fae299c602b17d8679852ec5168626a73385194aac64657fa9a163d59a9623e84448a81fa2e06cb88216d17415a07b8833d5ea58da13a913528b68c33648e82718d24217851525f005ac05ee10108b0217b763b5ac004e88c4bf6722005b759f7f3fd09ee0b5935b326f1ed266f29dcb4e732562bfad38219cb988da78f1bde48f7dac29f019bbc6b28f4277aeae391487c1044ed71f7edb27e69b78cf74caceb8894261af76bd75308640b53092538dedc4c2825ffd67154d74126bbcae3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd06407ccff49be0373084c7b524c3d88bea4c08d7f202977f6e184263a30e84b260ba7d8bcaf8b90a082756b4c1de536351c94a0a4b199aa45b593b25a68eda16527bf0d7e7cb858b2c4d9dc660cc3b17a867665034e23dd82b576d93f36f7e94ea0943a98ac2ecf5360e57001cadf20193aff8c3eecc7506be56dd7a031c435978c36d776a660f5383acca368c0de80e5f727335189c00bfcf821c7a50013273a1e865f04779ba5f301de858b64c11129b3296dd72a8269a89ba9c7aac496a6eac0acd84fb2f2387583ec5e63614f4f3fd2ab676fc4f661628978c8e87e852040f7e0369624418e0ec4a562e57ca5def1c82a2ed37ac93e337bc5af61a0e5a3c5a91fd04d223d87cf69e6f14cb849f15982fabaaa7b9252e80aefadc6a6d489bf26066e1d7688015872188499b576e39e48dca684eb3334462fbaed15e697896b368b7b3fe557832743991e5b25ddca0e9325d3168b162a9cb394683d7f456d12c8a64fda99053b2c2791176ad34d796eeb3ec34d384889ce827bf5b0232ea8732462265267290979077cd7569709948c2cc75ec3f1396c04603c4abd3bed1b2a78787a85473a81a2315ffc842cf8e93628e886994605e59457cb75395fd95e9eafca9b48a140d94ca2f7139d675d3f2ace46e9d51ecad4fa81d6f62a52ee32eaa39d0c8a9d97bd8ee465941e2b5657d49ede5e0ef1626fe96864f3743a7cc3bbfd079905aaa69a2d9d2417f3176dab3d5da91f284654c62d7716922167e3dc4792eba4c732505dd5580568bec41f4afec65af7d8cbb44e0ee4be2fd878ab4e8654d2c0131477bc3424577bcb5519bbf65b66946ca1569462726ede30daa09e114db7ec52444853b8dad2ba33d73a16890fa8e096622b7321799fe540ddf7880cdf60d3c285e61202d99834b0468aa93fdeaeba4db2298ee397845c5371ddbc51921c4bd6914f7698d66e29b711fd1d082de176fa9490a934895ef79f0471e5ccebebad247ecf0a84dc2b8b15cd281920d060f50b9adeb7f45e1694f056756f54366cbaeda03133c5d89f28b3e160b17637df10152673ed858b59d194a5e59ce8ac91bc5cf8057c8351edb89cd41c4e6cb29ae1301072f9a559d79c992aaca73e3e62f3bfde85359ce4b057fb4002fc4e4480fd66ebfd604747083767be31f8c4032a522b52653072cf99769356e6caa45150ade2c00b72104375aed137dc0f3255009aa6f53b0a547deaa559ec915bc1278f994aa64b9ada7018d8cab44e08d7f244b442dfef44e9cb1ed3137b0725b5aa8db071a86e8a37436253fb32da756bf23ad3f1d38dc69c347a8165ee4143dd19a1d9759f3bd0130943136b2a4c19053cc8f7539c0f5a1272bf0e5325c9c795cb85604541248ddcc19b1704629373b2d52166959cd2cfe4edc8a228654c66262f3a2ee38d39dd02ef31927e2422b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha348885d9d41d15faf84231b0c03d2d259b5f5f9fe12a3f1625da0e215591054ff9d6f2c24408a78f08b4bbbff414f54cf057c71d69f5cc5a0fae5b71e3a40b05a33a60d2772fa516151f3e525222bd91d8e38727c505752156ea919d9a449396c38edd4768123fa74a3829bd9882e7e685ef093f1c4f7c33ec333f35e18cd930ae43f68d4245ad8ec06645510490ad7dc5c3e79f2674f8188d491dc0d249e60ea5d117c91ec8fb2525017a660b67d20cbefc6955ca7221624c596574d84bbc2ceaba103897a52ff4e9c99ecd16bb23b7b57762de3cd2a9b5a3e808f3b0cbf9f9060157ee746307863a6483b54b6a7d7d41db520512dee8e11afd79db4d1940b2c2ae02f7c29d1f130ab09ab4cad0899fe8b33d2b8f5a783d5ae13555af9802a2ed2fd1aae9b82b5e58292f763043fbb950b757506d43b9d67fed880502a71ac851877105d1fda171bede2e6987799047bc5b797ec934c9bccb5c403f3401c5989adbb12ae0b77f4ab63a7302f58c1a2dae4e7065dbbba7e6ce96a51d4dee60b5b337c32a0cdebfc3f2aad179a9219b5f685513d06a9c7a40c465fb7f18e6de6682e643d6236f7f39818d9c9712c7bab700850a6b14f01e33e1eb208552e9fd5be145f4fa8519b6135d87c07650fbb07263106582461f653a2d6f035c6f395aa05ec42683f220034afc39caec669c798e6bd897e2d873348c908341ad2d1fac1d567958d42ed306cade79c41ee1e2823e4bc73673d877a5e67acb293286a511991b93016dbe6ee3800211d10579a804ed29535f8d75f535208239e7f6432fd0aa008d6385fe3f866a2da8407ef6a140b77335cf12e39f3d81800e77dfe7d8b033b34c0c8d89a5e7dfc1f96fd63b922f4702a52b9281a5373c57b15f190cf7e8e5f147413975bfdd1931c3c0bc84cb0f3739f4ea1972d0a6c83db8d30d20d74b414ae26dcd3b3cd566cdab742bc9abef18a72508f8768f6ff4e8443c5b4a832bf723a3b85ab5e6d1b1048825569d11b2bb7b722caf9fb54ac9bf45de8f4c03989cba94a311b642c85386fa890a55169cdfaaaf56dfafd8c8471faeefc40da224e82b63b535c8eb0f0e4d614821e7a8513c39edc6b7dcba347b13d46a4fa72bf7470153368be59b3d9c56da81619c654e70e2550b1ff73768cc0427bcce545738f508b283dadb00e37998862acf30500bc7edf719b2ca193b82235bc529714d4fc9de832f1b43f41b668f5d6bcb2a3c4d58ee3047a80eccd25078ca705aeace7fa6adf0745b2cab4bee1533e52865efdc2d1d02d4b9783a6de0775bfde77d94b5a3f30182d6c3d07c98de004d74553afdfb0e09bb2bf6303924e160c9ae42fe8b617ec66cf045a3131c3db7e3411a0858981fcf4e678f5942a089fed859750e07432075a3690347978abb543d0e4e4f548cfd1d2895c8b3c13576cb5ae217b9652;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hab53801930828539ad1698f9c07bc7d0864dd29e53a5d38dbe7bcbe9ccc2ab946d872379c92ef27454a07da2c71013fbd6e0f5b652e513e3410864b151e21ffe5f87c64c91d8ee85ea604c951a573c5bbc3e7ba4aada4296d73dcdb1799df2d9fbdcfd523c6f08a414dbb7e38b9afd06f56753418a90bd3c85b787ca908464ab775d76877742da7d44dce7b19d175f3c556855ec1c57cfaf5d49c7e0a9ee8b50db8a846f7ffeca320d6b2c6e74ca9b94476687a3554a38c24ac2ad6cac961884f3831a8d897a74cc75d0e23b110ce7e5d9e9b32a3c89ac173bff4077415fd65a958e1ff948b1232f6679748110ddd23b7e6d85f65351803c3d2b2e454c79e9f7e5e8605813b5587fea837da1f599e4290d86def16ae6898fb4170471ed49d4fa37fb56c8c5ed3996b866f03e7326ada2a4287225e217cf7ee8eacc2dd06b2a03ed651e29dc25945229744ecfada9c7a83351a12446656c196e5aeb0bda46e0bbb941ef442ff4ac9defb91ea569918ff4901c6e9d2c15c5d49db4e5bf4c2123cdf44e6ced0213fdda16f6e2ee3215a90b4332aa0eb2c78f53e6f4aeb14334192ebfef9f729e7547c45f3a4c58176d18c36d69eb0cc198525f090b59e7a00c30146e73bae1789a3447737414fcc1172e0d3f37c39c9c2751c7f70b8525f2d32efabd648dc552f0835fa74c43c1b09550a7233108216ff1e2e27191aa446042681a10aa9a75be0fdb6e476d173d90e95f5898e9fdd4232ba0c36f4f2feaba007f8296027df2f50052993b960053459eeeb2b8929b07b6074122315d383ec0d9320222f927d1e3ac8c83c2e164b2808f47d5955e6434afc4ce06bd54485a15c5af89b03d708a2694e9384f0dcf14f4ce67b9a47439a196423578ffe4c14847583310b3b55bafdc80080e582b88ed024ab1b9909e4d7d4a8a9ecb68fa0db086094d93bdc937081263147e48d2a553eae8fc64e7b85799b05ff56374b0f3c270f8c8890f8da3336d4e4837500f7260e20f1a8936c3a8574e2e19f026b0afbf78fe383c152732146aca2795c2706d13fbc9437481e274bbebf55455882a54f726e9d05991ca18375d1186b59b52ed22e4a7b80c11042ffaadc6bbe55192828cece1f9c043603f6c0fe155ae6a66c03ff03f0c3ca417a1a49c6cfe048c8b96c919e20fb489366f6d4971c0ba7f3b5d5891eeb5c5675ed91ff825e95e8f75d95349d8d5cc1660e1feca684a2c6d76f38d6616912e2e15715df5c61da752aef95028aaf17786cd3c9eb751f297befd9a49b8ace766c9eca8822ad63be0ec6ded9167a100e63c66ede6dda4597266ddc22d271ae90f30bcde84b324ba99f9e81fa31dff0dcb1d69ad68c27da588c6114ec2589ff2ae64435e31ec06e5b91019500f59e2d899c5516ff68af2ff403d9d628c3843e22d4091b6b0fa2ede7b4ddbe93cde9ebbda;
        #1
        $finish();
    end
endmodule
