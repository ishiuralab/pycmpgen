module testbench();
    reg [25:0] src0;
    reg [25:0] src1;
    reg [25:0] src2;
    reg [25:0] src3;
    reg [25:0] src4;
    reg [25:0] src5;
    reg [25:0] src6;
    reg [25:0] src7;
    reg [25:0] src8;
    reg [25:0] src9;
    reg [25:0] src10;
    reg [25:0] src11;
    reg [25:0] src12;
    reg [25:0] src13;
    reg [25:0] src14;
    reg [25:0] src15;
    reg [25:0] src16;
    reg [25:0] src17;
    reg [25:0] src18;
    reg [25:0] src19;
    reg [25:0] src20;
    reg [25:0] src21;
    reg [25:0] src22;
    reg [25:0] src23;
    reg [25:0] src24;
    reg [25:0] src25;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [30:0] srcsum;
    wire [30:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd34a5eed79da82e92f7b79d1a791a4b50b08ae1e461b3c1d47425c24bee63d788a70dd0ba6061eedcc27b4ea5273b7ba80c5fa84b2c84337110d1c82ad8b26a98e234e5253db0b7f762b7312d886132beb679f536;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7a41b32b57b5b8315c47b68ab3009b2d80d5a05acaaa55ee51e42858e3b9c3ca8a3f333352e88986ddbf8207b2c3e0226f10d37f7798d3eb62eba91c1a722891e47b3b7fb46986cd80bc7a4922815752f1236c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb023f5cc67daa6576cdd515a1e42b945671d5eb1f1b96b7a25b108c5de523dd3830057480d1eec0ea0d587ec410a7763f313862d60e5b3c4e6b85256c2d6e3a30c7d03e72a12c10f5a96a8cc3d65068ac713fbe70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26ac9c52d83fae9bda919eb375f146d7cb5e5df375f531af10ff2ebf89f65945fe65c59bff1bd13bb1e6a6e6282805e98f134320ecfb1e891253bf3875bf7b537c18022ad0fffc63f6b0a60dfe42dbaeae602b783;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h667dff3991eda17f8b0ef6a2ba28bbddf8e0a04622479eae8893c15c46adf0ff3193b734fd9de897e4966b28a02604e7c1749f0be27655dba1f4e054f73a08604fe654591dca82ba0b70eb5ef2db0b8170b35c229;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h667d5630c30c8e6422b3d6af1f03735bcc4374010d837c194f32d512b9bfb83e2720258bb02fe739e505a6de51bfced7c0a65934e4fe2767911a63b179ece85bc3bfbefd3747a7fdcacaf81a098287e19ec9f3c4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd26bba19b584dafd8e22a2758ffeb9fbb92b7e54628f3a8ad86df1b5d96e9b7052f2cf5f1809207e2ac50bec6e63ec15d37236fcaff7b8c0a85ac8a504e2dbf47d835a571c55e3f1db30396cf19eac0f602514da0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94cf0582bdebc2b2778632d9fd231389149c9e51ede5d0ec74548ec4cb60ff9b30570fb628c620239f0e48e50621ea3c5e732d19432321f27e5217d6a57aa659d9d0b78c1432dcda82375babf08ff712cab55a25a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45f4216a385f8cac28073dde2be354b24bf0591d0f39cd69e8394f513e7b432174c0b9fb6794d8dedf75af33e6f32c1d6a54ea65c2b1d17e84ac4807b8ffe2b799eb2a34279fd3a11f33b97091cc6d5d61f76909e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e2b5f48edf66ec713ae183d39abe8c78002e670b0270a9d05108432bb17428631ffc98e504dfc724a876978a1c50846e96feda0d62638b2a34f188613a64b675869022c3f9d2ef7c7ebea9d5c72c1adde7ccc629;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b95fe9ac2a383eefafdf9a72566ede9dd2ce066a8062b9226d8d0505384096fe2ba4c7fa37cc369328301f029d2bd3859ff2895e19ed3ecb5fb6d1b752c691e3b16d0246989a9d660474a02800deb5d4d8560c38;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2b67178598c6b70d35cc7d6aba284e681fea4114da9bfd6ffefdd9b7900b8340102aab3e5f83a17292d2bc826f20a8f17657202df44ba0e9149274683a3043c8792b19df50809d8f41e4796b17aa18db9932f536;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h808d45d4daa72e2cfddbaddc152cfb4b1f14d3a9422c0b265b6c729bb94072d72180ab4746bd3d2b9fc7e511158b2a1b6e649a13be81bc4cc21101b62d84062bf5090bae4821d2aab96e47412d8203b60086c4d0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63905cdf112de0bca106f9a6526cbe80a615897b54b3820fe09ed153a2cee49d4b0244ae1abc36ae3801487945b59faad4425699a04d7402687a76aab1ff001b310774aa7d0b74a9dc2d9ae489fbb28d8def066ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13ead8bebf06bc6b4e89d57397c72f24f084dd2a4f86b303fb396fe7cd90c2042a406418afa64afec1acb2239dec3757c0204523408b3f36f79fe4a0f12dfac0622712fd5c0e80906250352fb2fe0f88cf2930ee2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35dec8e925fe2572bb45eb56a0cbb4b97c9544b777bb25326a42d979b378526909a768ddf2b05be2713d7065f1e53015f3040747dfdbf5b0f26eeeb9006ee1a21a7f264abf1c37e64b194647b3681b31be21d7289;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f23b4a360eae06a8542b62a4fdf477cf5c41f5120725da6ad0334a4d204bf685c46b5c3d0a0865559ac4c29358be49ff530c243317be4c9eeac6ba492fe74f93ec2cd2cb9bda9b54747012f5ec6c6a9608cc4926;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd59bb5eb76393775c94429374d99fa9f0d262ab38c4ef65cf65fba293f4be7f2d31a63176454c43cea2f2b4d0eeba10dabdc7f78c67a8594d32c9b7aecb770127378c8697b4a6ae0e519846825cae2fa6ee55fd79;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3fce28b8ce131e36e6d1c991e41eb3293b133b8b94732aee8f33a078bd61736b10078878964505f7ff35d30373f573183b4f487e31acfb4eceb071bb2b616ba230f9d6119a6a2313df8beec58d27b010c0d139e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h387231b6f6e091614212a0b86a9a316ab2f8245c27309d52e6497d1af0f4ed8a5f2e3c04465cdc09ac8ae679a62eeac62a9f5d680422ab11e0d70e73cae5bfafb4fc95618450e2930e0cb8c38e22622b30eb36539;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha943651d6590128c1959a5cf780c3452fe7777c67085b0b918662a2eab3e23a424a0ad8a1da5afa200986d49ca2a082f364849f246c0cb77582559fc6c10e50f0528ed8553ab5edb925fea1a6eedffaa05fd85a7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd408fa747a816ef13dc60d9048c406000537291065ca0a20f5eb972301a609e0e78dd8d6291f42bbdebdbb519224a82d91d4585c7d1d2925171e75e147dc52789383ea0b846ffffad64f1a5bbf69dad8e47ea6148;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9dad2fdf28e83527454695e0c972d3402737d6721698da954f3d9b4abbb0631fa1774ed48d883be5b4c693f07718882412bb9ddca49f88d1b36cb318e67243df2da31c54d37484864a8a124542bdcca489c3228a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11ca17c8a112bdaa5ef9e97b381ad5130e4ff4d1c565d45290b54d18def90c6cf44bb44f6b28b7c496473accd358950c3eb669d1b0adabb7760ba4b0fc15f12faca08aa03d4b3cf83105bbf820336470872384867;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9384fbf34d2250e2dbc73c1765b3b43915ce8a035545746963477dc9b368076b31fdcfeebcc93397bafef368d12f9d652364f95837b43105f26a68a24fa3de3eec9ddfafc433cbc9510619d7a17253ff19e1be29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae1922f9a02e22a1e83744e0d1ae8fb82d6a432ed485cf869e558c938b1c6dcdf3a54d48f6531732c85069a61ffdfe933f89bde7aad6d3751422d7ca6c46a64029c106c4feb7aef537e9c1553b670068c6cdf5de4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ecb988d4c419b6438f8f0e9ec8d4cb3885d024f0148cb84bacb9d7f07c906396a1938a3f4d83e7b84f0ff206046235abcde71e81764b95cb65a5fe9242bdce3a5ad2ef450e5619009d1aa34d7963a79bbd01848b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb91f9f55730689630bbe2e8ac3bd61b76364d8cfe8f43d32df35dd4680f15b6d8088db18c6bf80808e302ec3f83de6371501153aaafdf667484427f1f89dbf8e2f08102a3b6c08f472e3a3db24cdbfc5b05a1a540;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97b85c90ec3adffdaf193ce634ba19af045add6a5df57e2b0f6ff4e8e1bbddb1070468f081e5efe12aa9b25d717ef0dd95197871233c5f66df3de12777b9ebbd0e2d11cfac0b038b241aefaefa288ce97ad41d163;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b581c614d2bcd96660eccdc865b7e21f45031cb27a721e8c2f4a625b4e4f3c1909c4a209c109f9a726ab196d6e1579d0f80b71c5c6529648fd30fc7f63976e7f890f2bd9c5f84bc30d3db6cf94b898e58d8cd031;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8bf6b347ad9b9795e451bd0b245e89dd6b6cafd9223b4c23cba571be9cd9ebaf4cc464914c9f7f8c4b0275adb9a0f9c44068f39e43e03aa36ad566a5455129bbcfd73d325009281d5c02467d6d3a3ad92350d677;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb1cff82576f30ce756d45720872ac2213c5e57bf959ea16a7ba5b444faef5f9113cb9731ad9e77b236e3b8b3bdbb2c3cb38885ea64ed1481ee376003edc8d6229002aec68b90f3831680135da47cb13206f99629;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e8a07fbf0ab896f8885f5c3089e60259577abd48cc2883dfdaf612138f913281105f7ba4a92597c3f54648429060e8e96a8ecfb3a57c22be9a69187c5865eb651ae8486cdf2fe4e328ba199da81f0fc5db6788fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86a3cd52fd5d2fb4db6557cea0553943c393f540801e81b23dabe24123e6357ddb298a2114651dd4814c12637cda9f59ca8e56311b03c2dcc7cced889b04e44775da5eb6a8b4827ce289593ed10fe430e553ff062;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41c657746b14eb3bd5376b0ee190e80d50dfce8f88d3d91a9b4294e541386144eaa3cff9c8413648c902ef8c8f6d110c644092d047dd73219c1627c4e6f8dc75e91f08f2be3b3ac2130d969128a20ff92521e13bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7ba396e70ec3031158c7b0ba292eee565c3f03133e2fcac997a706064c3ee4e2c10010aee84d05741bd20e3216df6954c7573b5921800bc98ab5ae970810110c4a658961c456c704fefd0fb4ad09a82dda8d9414;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3cfc74427b20bdb6dc9ac055e3d9c4cb4667f23e704d36f04bb2837d005859456187a9fe502053a0ce32708b2c2491097c5814db1cbfd34b64502764692e6747a60f975f8f64fa1d32b10f80f685125febb4bdb9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'habd5af94314d59614cd469b5ec5623f494df7e84c08566814840672f70873ede270c6631ea6b62c3faf15b26deaee56e2aafe586df402b29e22b54b4b4d0e09b2e90bd7853baac9f6c95ebe1b4080d8b67ea3812e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a9b59ea6946126a3f2ed358c1acbf90fa226d6300009ad182224b53c664d4efe66acccd5108ab6ea4f1ccab5063e43999bbf6270984d2a9123a04231ab5f361a72dec978d08b139488bd92dd385eb89b5bb107c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d17c7439c3fc03ddad5f5ac9269d7f6a334a568a4712b6343925337774128d0b1dc7689e3cc410b5514ed34f60065c6fff33928513e0de0d876c9c211f82d4cdfb821c30ffc327d3776ed61dcabb170c2ece6443;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5178278adb88176a6da1683bb46e19a3de2aedc9c9ae26b8f9a20c0d1a25e37784db4139fbb2caf82ede4b812c291e38cad446f4624445d1f89d630cc9418c3e17fd97dae0fe57de5bd4245164299ea23e573010;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he81d647bd4c78b473c3644354760bec62a296083fa98035dd82e01f12d32e976229ffe28548000180fbbc450242fd1b74b54b695d0b675ebb1017ee5568149ff53e686bfd5107ef40585861f22d27d7c97745c46f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67c5b2e0dee3bc33ca73ea685f1cf1ef9190bc8c5261e2c2a263708082a6aa24a07faf7216860993962a41ed0e6e9dd0a4da82ef5fce82a8e1574d3ce9bc058a42a51f9f3a8e25fb178a8f1ce36950ef7379a2abb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h895ce176bb611cb95444e9b84a7138b012b19dcee24ddf66e62ba55cd2cbb2de97f1592f31731ebb22705888be40138b07636f874d0fcf90d0976684401ddd6961c59f798bf6548ae20b89773d4cf9d93dff2366e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a5549de1291696b3930c8502022199ddb520131e39c08db129748d18b3b4e2ad548f65b0d50ed031a2ec910c93dfaa2857d3077ea111642efd5c068d7100831318e3de02aa4522be8d7b0524304d899231c24bdb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dfc6d489fb988250bbad283138e8cd58afc9cbfeab79ed7b98d32135d8dded899612fcc89db0e48fc8b61d6df8c49ad55c9743ac22a836f9ba9cbc747ff946589adebdfecde3b17a73de47225d3a4733a9e7ef81;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3e5b30a9618ce198ad88702c4916828877720d269a6e70874b11acaf1856690a817d4699c9628d03b1d5b266132494d2dbcf43c3a3ef19003812b2d567c08f6b0ef98756a6a3a9b4f19c101acc11a794f7d7fc57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1e72d200296c147ba72510702668d215e699e6c5557fb4b60f9b85eb5a02ceed6a0cad6e6e352b43ac8632c5903e3c703b4582fd577d2d1f3b47177bf62c817fa3d033781379f54dd602a488e5aec3ef0d461346;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2e75e4dbfa410b9be72935a9bd75483054775b1c1d7a83dc6c63b072064ba0df418ab1c3a6e2f26dbcc45a195f5c069fa080f63ef88e2f2cd04a13ada5a602152e833ef12aa97574351160ab1a79b97edc30724d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53ebf5a0b4bfa61b4fd7fe9a2c2714ad2cb62dbdbbdf0ac9baee7c1170aa85e3257b25e81cb8c6422149a46eccaa0baf3fab1dd4c7fb4803556d42c28bd0beff8331599b7b5c1eae3c824c8b1496b7eca1c0378de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca3c6a9680601e9b6800c6526f6b719c8443a3ce853ad7c3664c9994c45d983f41ad937db7da68eea281abe13cbe9001cc869beea55398fcbc6df2db2219d7d4928e2a60d88075bd02742c8d562526b7f4e7c416;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h766495af25889fbbea0a153c78fab0f577d7009ca87d467d930ffb367187a3cfc429b253a187b344a2963cadcf72ad326fe705062eb356bcc297ba30de05f79a23c77724b3c73370d8efcd4afb58244b45fae57c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h992b4a025f925641b878051032e26801df6a24e695e0c4ee3ee7627817a3081657b4f8304b71fc4e4e1839cec88da2ec5fa352f3b816d0b60c4e8070eda652677ff47f77cef6a54475647478fdc90083977d693fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb85719cb50a56536cea2039fe94ba5e4dc1ee84eb92edf604932c66b8196b5eee3fc4064cb5d847f08a8489af1a011b4d18a7e8ffba062eb17d576d9247c6bcc384c23c567a62b8ccf75808b5990b82dfd94f31ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha36c4ced16089d31835560ac71deeeb37a8e9cc9a1825474ab32754f44dc46e56e17b8fea2c191ca04dbdbf6cc59bd0d938702700a9f6cf853f638da3b920ec1c3e6404cd66c654b2890a132e547cab94c35e86e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h489cfc265aaa28ff2094aef18621fa88a6472aaf0619a5d626d5bf4b48eabed03f9fc2b5ae2ff5dec2165be52f3cf07616a51591c0755e0baf378c129fb374713c6bb234e9ccb5baea5313846277dc8902ef1cba5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h569864aa6e57755947d9e53b5a57e9fe414dca0ac945bb6af875e443ac00f423dd2fc8d4a2db4c8c418d2f295baefeaeaf3f22ca6284e4ae1fcdc660625c7b02f6bdbede4d13d3ffd5106c4299851f63b94725c4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf4c8c006b344eeba1b40a2da1ef2b4075d3941630ee683e1f3c6a81b79a9843bbbafef3587170ff011190cf671d24fcc14789a3310d3f747065f3fdde8c015ba74ea552b1ca264e7dd282dab0b874996f8e766bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72b278cb406e981d95bb0434605f1140f06ced86563518aa5080c9f89e4c23b65e9e4c1266032db523d43fd0d084a12fec881c37d85a4fb70078c3e1553dcc8b104b2e45b030905e1e23b1067387dd1be9928d293;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f75fd042957b9705f7d87ea04d5d526c7779de4bfa8b5e32a0474ffb182ece0c8f31a4d4f18ba177ab3c2356ee07001069056bf51d88b369f4b7f478a2f7efd1ea204a2c629cc58b8d3cfd62038292a5827cee28;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4da8120e9cc8b509ec5af73ed02e05a6e5e2586cad34240dfbd8f0d725824591ea6f837135afd0be1922199837fb774c2ff2f4526792ca867fde01fff04884086748d9c03e8c2fb2a26a5c30ff427ba53f943b779;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9288d7ce95c6b641857cbdbe429abbd5f9d3490a827b446479226cfdf235f3b12110c928c617aed5c06c8e5b96d8c00828beac6dc7408ff1114c312b6a74afeaaad53d59a0042f9938afb1498cc8c8b29cdef9344;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0fc6a6e4a3f33ad4a809e8ab9bce37b0d3f90ac732da1bd055a6f840420f5bdfecc96ad15f646780ddf378147f886cfa829022b8ff1d79f784d25ec03c61813b65059f36b793a9d7e26af3548383c1111ae9f6b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75dc71b75c4fbebffb8c75891c5ca007b3e7c5c44640fbdd33108657103f44dc6ac158074834e070602d1c094ad7594b62cc8e35bf775198c5003e0c0f4b34786e565149a9e0eb156dbf8225a9eb6cafe3be821e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haef2f9d456321c6a0f0e395d4e557307e289a1d8a62bd87139f8608a8e4a549bfc585a3589ca22ee6967b78fcf6fff8581089783220f1c3c743b7297e2da5d14b5c43200f0f480eb624f0e3a16974788dbbdb55e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hade97c12e903ca7d63e3e20f82c31894b10c332fe5bc41cce60be080411422962ec5fbcd31d7325b200f8041ba759d7441598195dda3399300ea935f4da89f724d5e8682786c6c94b01f5dfa2361a889995f4cc51;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he986200025f71566850140b0f8d1f6cd3a7f544f31a6b9922837c5087f2e0e50ab81083eb9c116dfe5b591376a0cd8a18e7bf886ae358f6f4be58b5d41170dfa1380a0dd4be232f869a849d96cbc4fbef2b612d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d7cba7d18d41ad0f8f94ee4d0a25415f44b58721354a56b292017a9d299496b56a89502de011fd6bb7791e320c970f7d1c35cdbea1680fcc3bff2af1e43d20880a376621d38c73b0658f6fb2520b12b0a3e2010a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67f8d6772cd8bb4f4cc8c876d76047a6fb28985a5fe1efa138212a97f0189cbffafdb6235966da649555421bed4b99d8bd82f4b737973458d5af9ba27dbc4e6185e1b9ec1690d6aa4111879850d12e6a86fd1369f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1d0bd08a6972cfb45b8ad57e9a140d4478a3be6e4f878113002cf6ef9c711341ec84db62483756923ceeef86bd56f693c2d4055bf7ee8de8ba591f70cae5a60ce6900886113393be4628b0150cc0ecdeb461080a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2167b832caae5a9be813911a6015dd4535c908fa570c1c73c77a5212dadc4cdbf24e33ea94ba84d990d08858bf6a5c51d48d321c18f895d947169853bdd6822c28a90783bfe042b12fa0be08da0dfc55f9de5317;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99ea80cc20583f0c1fbb2dc7ad3d59b602a260fcbb9c5be03bff54febae2373add66207dc6b14c109ece1b36ab0e0bafe101a55c7f9ba71f21e589b79547f552618043c63b538575afbb1d7ab8922e5be79240b5b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe174831469e8aaa042cd0d62c99d5f45aa9a24e7dcd3d34928740f96f101add2474e85d92b815f89e1cef07f8003c72f05188dff6425844b3251e5ac20edb409848c52b8aed8f04d81ac48b3b4ef4fbc818f70d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h166876f40e6fd83066e30f5475de1fe85be8b522f7483700a46aa4d82f8f1705aca8d76cc82227bc9f1ce57b949dedd03731ef9c9701ebbb4f7dfdeb4c668aa796978f896349a810c9e8d54e22dc89f06cd28be60;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h778d1eff4e434131c06de440cdf9ef8c97d3f9bea582faab75cb0c58a961aaa2403b81968dd61da2607583f3620c0bdf634cd79b8fb8dd7c411afa86bd850d7491a8c39d20ad62327b8734c372a0dcb6699d84ff5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h999c1873dd9ef441924006896f7531dde3ba5ddf3968a87fc573fdf2ac8b5216772fafe8b1d60e83bda902c977490341a742e028617e4bde9bc9733eb1a8466e9f55266c0b5d4a00db179e0b550db18846e7b9028;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda2ac24865bda548f541b9568d6ace0248dc6305231ad981a02a1f50dffd1187dde9a30de321666dd19907b0acf948c777d3f1c16bda4dbde5655229a55f253ce877730e0ecb8e9a31e02ac521e734d2f42e6e325;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6d631ae1f541d5364f0df81b3ecdb045b048acdb6792c1ad6c839a805fa593ae50bad7c1a6cf3a98c47e8036f5ec7f023375598643972c9a3cd3bc08be40375c558aa64cf1918725ff691b85807630b812e37255;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90d18b1432799bf1d7bd2c77bdf867e0624da0e593c3facb889ff5ca0a46dcc23909ee827583a5df3ddf40a5440fc7eced75e18efbe3e461a436d76f80937d95b2fc05d9afc6d6bac493e86488c6572d770d57a97;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h513f93ff598324658d5c9493bf006806006dbb94684fa3f76582aa406e5bb168174050f090897f873f10704259dd10c3318daa4b0421eed75c8ccff567882cb6133e67ddf2d49790f5a31443233f30d656e496b7f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12bbd7f4d94f27972af86958879a1d0529ed52562074a87c33ac0475dcce2c2d9218a9fde824a17703aec47ecf3c5ff6a81f84b41df2edd22d8b0cb6f6e823949191f44c938dde3f0d60b386d73fcd4cd85b30cff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe6dd84b53ef75fbd8b044d20eb0f67ca80bc8d7b73c856940d8ecf92ddded891f757f9a10c80c5ac58d0014d4c9c325329c23a15968e09302e99596e0e2481ffff71548dc01029fdc52c0c35d2f4557baea35d68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c576d6b7bc95ccc0753815b9500a4920905aecfd7e56f7fc92a8964881ef1f3aaa9fee58ad620026801713cde2bb9107eec3ba0f939007ff6f7ee9075076f4755309db022bcdefffee2d855f90336ec3380a56f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bb48648409235be0badcc2c523899d9c9a03805b16454bdede3522d17838995e55d7dc30b4c82b4930bf3aa8576f94d342d99a466e3e7e6d64a65278929a54d98e6b8cbd9c4086172cecf325f98e0d50ce919aac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56ae4821c32546a013b260532dad89c724bc03785c9cc564114f30634fd0125c42492137a696e6583317b3a5c4a8b3919aa86569f28be10538988f59670ac54e1a660dfab1d3b3d21093a295a15b6e5addf3051f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd5b2a6a61eeb0e3def56219c030ad64a857a5ad163914d0dad0f8cf4d9eca99192d4c2a4cd0c0f590a3c410523c47224e7c6137a98d0ad984fc6fb7b4122724cfb4d830f7c34ff118cde3579e163bc8552520bc3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e80d07e159cae0335506b3428da0a27a2dbe2a728e03122cb47fc2a1f7779f86a9d042e2873482f790d574c7e4dbe9d10a8b7c60d4ce1ff9aa942fd78f1e4ccdc099e28b7e34ac2eb0a98a563f4c0c2a8bd639c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fbc82cf943f910816459a9bf5a89f3260117dea60b1f054805381c5b87d1f400d1f80723d8305ae5fbee764024e134b5b3b19b217f15815821eb6153ef5e5429f3521c89f37bd3a07c7305d9bdba67e271802caa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb53cd672275e9ef95bc85676fa9df0b2af6203952501c8cc88bb9197c706808c40ae8f960e8f52abbd67c162cfdd2cf002a0b2f267737164f474ce7ba522560a75999b0e7b23fab7c055eecfb331496529629cc53;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4fb304c56bfaf4b25de34d379ee8554a22ce37e9a4b2fd0caae6a21f0262f47cdd3fbf91e4450b9e682ad9c8e57225df94d9847d2b5dfca279cb8990baa99959503d6fe758c2c47c51df95b4f8f37a18e2b97fad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdb71c2e332b659f535399ca32343e8c7d584648c33e77cee91e70b1663386b95cfd12cb25b624df8a9e0b8b697278d0d19385bf4f158b8d01c81c8d2fbd5695b613a7e72f43c71b7451bb1dfdb86da199d55ab28;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b33eca9450d862c1ada622597642e1dc9cb318b89e0a4bba549649d8878932319c1168343ad4165462fd1ce7ccb3a39d367c570a2c5844b2cc42519f282430f3dd68febc8377e1aa9f999820d32e54345d1241a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h232990a3c5d1b253d4b5c70d6e25b1c2edad2c3d3385d540d125821febe76a1e267951eb881f6dcff73aa9a4e4b2b1a6744c66a7fba2b438db43e621203073f2fec38cbd2522f11bd7f64a26f6aebb62ebcfc5092;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60d40b6b20e4097ea6ea96cda5db0ebde4a3922f09b452c93445984bdd67719b1221776eec254e9adcad8ef96a87a7c6c1b9e89bdfaa11441d43230c337de9b201bf4cbb64480350b68f6bc843fa9478cfe2937de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5613e719d00c4857c8bc9278c7fe96cd2b802e185a32e0103ff3492795a80d361a5b8dc2e522011e3806102b8354fb0f47c93ad766c106954268b53aa1a060e3ecf5a579d7e2c52b90c43488e00a6331a6d0e04c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a96bb8224a34d666323e12949bf10435dc5f03835f2d9a590898baaeb26bda7f6c7f4af8ed4dcc549e1ba06130eec90a7acb575d377ece2fbed09f1072fb080953505e818374b15807f35b6a67186112760068ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f3085831730e432ede5253492c5e035a34aff0224ddd62fc99303df2d05caa0dd9c2b168e16b357c066d7c60dc1aee10b40a61eaaca0e698fdba0caea2d8a08656bd231364dbd4cf9aa60bd435064ff1400ac1b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8968df3dfa3f83b7c306e17ad29654c24a2cf467d9a4910634dec1ef51a8f64ea55741c07cdd77839b7b40dd5a5d102bdb7a6540427aac66ee246e2a8b8ae6769285b52d6e29e0dedbea41d24f4185904f11207d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h422ff18d8ca4230625fc4686ab5ec62927b15c87f3bc551514c9df5e1e847b6122ae2e664c0f23a355b88c5e94e027b57935f849a522c0c96db900cf238d2ba4651a9ea895707010802ca3054f6269d9674fff7ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf39bd6837c6d370b4b54c8a313a6ef2ad5fb9c322f0559a4bcbf411a47ab87e0c524726c50281faa04f64336df199cd070763c9c2d782085046ec4341b76e04af6394c0174d216476d186da90a589f6e00c880e05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bc49e9f860e920e3fd2486930329fe44d464977af95426919e6e9e70264c6e504ea830842a08a3a08ce82efbb730da60e65ded6c8a5056140f8877b17a5780aa9b7e8dde1ac8ae1ebebefabb74b7cbc036544d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ac455ecf7abe1ad4686889d3b57263c2660ec0b935a3d4501668a625accc770d715547f738b1bace316b5d31ae70c096173796cbda3ef89a66525cc1757c9fdd1f43135d07b6c3b84ce21f7cf07261920dfa566a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57b94b4bf575da4bcd09355d7ea6a3b5f9eb903b88d4d4eff618f874f4eb50a9025b0f7bda77861eaefe76e7acdadb45d4e9684c0be86f7e28a47585b81002e81bc4d73809ef0418351ae4447fc6815fa1e01258e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7c8965b7ebf1ede02d02602dfee4ebf2c8a2612e3f5276457605eec58c45e7e8d9bd025cf0361ba4f817cf520def6e3a9dd19239e51fe70f9e577cd60c503fcc337c60fe23faf02d7af69d93bd2183f0f9c7aa1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ba9992ae0503a7ea84f8a44dac64d6232ffd31ca4d53085d724419885bb01cbcc7785ee8641677e0a7365a30a68058e3b135a7408ceec4903cdf3cc340b362b715b8fc4230b6853542a3fecb97fb4b6a954b8671;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f16be56319523d77326e80637f5884ad5f630005f34fc8ec9617825fc095562f62f0dc6476594f5ca0f6ff296758a31028152e0684ba6836b0a7e32c4a4e0f2cf9d29cc413e062dcbeab7047047a8358e9f69916;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91164854e70d47946edf19baee6862baf5aa539bb1e3ebc8307a65467e315985e3610aefb3223d03fabe875d4b67d8fb85f1867f7154d977c4ded0ed76c6876f5d767db837181dcbee45a0e7c5493651000e89a90;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he161c9bb757773eaef31a0e9bf14bda1565b6f0f335f89cbc14fdd9a6bff9a9bd15ac37becb18aa260e671864c03ef0f17e97fdb2cb87211f6df048bcdba1d192fc30c88520a20630c8e0138095e006885aaf20c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7e0d99a8a1715178616470f1adb9587d6bd37f325428440beb6bbae41db72e802bb58fce624a872dcd7fbafcd3c6ee8800784204928d42ce7f462cb53933e730e970beaf1f0fc15d810fb064f5cbeb9ad13e71f1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he688d12c621ab838346a04b4a6378f05a8a5f4f94eddfe9cd002edf3189c2b6478734db9e2ca2ba9629b5c3c5d6ad3cf6f3147105b6e8c06bf9ee63b1dd64bf72b18e1efcd7d3b3bf4ff440e1fee89e131ca5ff24;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a9ff554b7ac2c989d0ccfc0a7c4dea355f0de7cf284bc471be62eb84ae9c1341a3ca61ed5f0f24227e1354c2ff2e3e7b4f790c7fc1852a91cc019c229ce69e8e2f8678ef977189b3c02d23adcea8e65a533ded0f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5347813062eec7e692c8715f827834d35cc432788f64d55df9f8ed9cea6cd84a7f591b2d83c16d13aad5430928659d8a6c76dbdf4355a7ba1526974778561b3e9a9a82f3f42f367a85f4f0ac64c00b7f1ed520d11;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7fbc22dc487385f0810e080885bcfe2a2b54a3f1e43cf9beba6ec3074870ee47870bc17942ec9aab4e126f34d83115bf17bef4745b0f15fadf43c2eac6c23100b7774612b7539b5ab3b45491000eb88d8437b1bdf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haae2dc90de1fe8ee7b7471383cfafff8e5f386c399bd6a5917f4891e5b6605f1c273123d0272ba527833d94a5e6dad2cd8bc68a0e6789e8981237475a9d913860f38e46786d0b0671ead92e17839e4fde312606d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f1f4b2f607ce9e574a81fb275e29dc387d13d3712b1f0eeb08e236854bc525f6bc8fdc531b3f5dd5241aff31a4b5231a784d20ecf7adb16d3928e9580315746aa52fd1f5bce9ff58543d30cea2f2224b757fdcab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81ddc3b8f3418b7d7ad83568530e26bdba19edbf214d07b38f71ebf3b3586288d898d6bb148d67f60e6b197f3ced25e0364b4238c4b1da63b64387bb11237d5fa23f0969a8f24f1fd114a97017425fcc5e0b525b4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h293b8155ef1237c3696ddd00ffa365b3f267d911dab8f1dea596fd4907212dcb069bd92ef8354d349fb191f8367deb161c7a51cf949c21d3b2621877f011a228e941dc56bfde2f0ee83deff5b02206980729d182f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5964a5b0dfda8641c7f2ed22cbb2e08aae68a39b3154e9e2c8f8dfb395883e2f8cb93736a7f6750db785e55e607f98d49bc7cd5acc74d4a5a0cd0c6d73d6808ad12af9186f4e2fdbbe8d83dff6b05db8f051c9a8f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59f3b6af162e6413d6f27c0c4247a10eca090bdae48ab9cdc92a17ce60d5e8f548b3f51ad428ec8ab538140301b12eed80231d758b82018458619a81e077fedba60b4cd35525adc36fefdcca7a5567ad667c3a80e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6add6995f6f836dd45b760f8d1bfa605edaad42f3d2b285b0ef3d8a0e607d475b06d0c216af4a4fe1289d9d92af4748a0ef089a17bc2c9df0eb671d2e9d4ece5d315202792a38391ec4bf47da8da6ad34b630dc77;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha153de108a4e190b2b474ee9d136cbe83733312d6be75ac5a37139e9cb1f41815ba6d3214b078886237b2e6d801376b960f0b124cd491f60c9880e7771f09d0e267e444a754b0a173c3e9b6e34296725eb89d4086;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53402db0d147e40e7f24825b74a2d6c6a1a97e3a47e8524826ebc8e6568e021674a9b6cecb6f0885e276c0daa5806f98e5ee19b8c31e466dff0de0ce14a33b94cdee0e6653a2d03e5efabf8df8090ea51333cc12c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f5f5e5b6a188dffa92bed52c3964a30dfb0412623c52d2c06a1a4af2529c0fab97ab7bd5967e4e030c37df1d7a3ff5b9634da2af02709e0247a54fd1e86b90b3d1e2b299ed0cbf818ea686a9f88adcf8667c5ff2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88e9fb0a45c6f1f7ca87c850b4f8ed4c641b06d35e9dc9624ad277268f35a7219be3791e650859d8346fb22d851a0aa6603e60c6ad0657297b7b7bd6b16590aba4888a7ce43da2c53683177be637d433e0b04a841;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd61a660420c95555f8fada5d846e8ee2502e20afcc4cea48a712e331635ea04586d33d45a757c81669cca12c15b1f34414dbc6c2fd7665af8a96ddfcbee0f38affc6e2af8fd48a592ae5e4964249d7be93d7effba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1614862e5496545fdf765985a54d8a3e919f3dc9cab9e4ca286d022379c9a4a89b9fad66b9c485138096c0b75a94769be7c6952f67fa462f2a38be822b01c378168e136bebfa3069e496f74fcdde4e9fb83e84ad5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd87519b892326b532eeb307bd49c8733d3d8c976a927f255042001543fe2deea9c2e03a0d69e49cfb9c00ddf49e057892b18c8df8250eeb4397f484e855b655ddb14e5dbb8ea9a7eff03a3cf4ed12b61a35e2b6dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1abda14db4b29b7d3d9ce9c48b7b95c9ef25e08a07592ac6a45619cf1a1abbaee122ff39a1bad793e3c3a76c604ea089b49201e718a542ea251d85f19463e7d31f6cde74bd51944f8938253c71cf01d172a8d964;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75d66e62a191f92592200800b3f48ceeb849348dcaf17d0f1b0431aed28b56632ae5b591b75c1ae52d40760d66e46d3311ebf7eaf5a9e915503b2966c810775729fb48531e7e7cd40514560998ce36abe527e7353;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d6e2cbf78d0dc4378e783ef308f93aee7affe32eec0f08fda1183263ffa2d4c41e8bf485949000184d159d9c99e1e9df87fb29f596c52bce8e48ea98b0d18b1435d390d7f32520b18aa393937bc04092c2192e68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha01e10284f72c0bad383fa34ac4f38f7e43a3d22edc60fb5302b6a101ae6b3634a46d6354381f63bae1e690abdd2c2de7c3be6bad2ab6a6c7cf4b531a2ea5e3e66024e8e1c47e736ec222a7b3b32c95676d191ac1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha44df961954d55ea5539a5f17e4913f9b06d55875316609561bef630d0c89430517ec28d423c6f7be824f1adca6ddd8844db14ba9c7cfbb109176299378de65d0b2ee3db8da08b704d60035ab7a428f7fb8c3bacf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h639766dda5aff60d9ec5f594f2506e4623872fa2bdd4bec10d0350a5129ca6e2ecb64e297044f5d4e64940ba4a8df61824bf64a041e022dc168a01c22cf66c9cd10fbce6ce40d26eaf49f19ba122a753a5ccf209c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85f7bbc7726818e6799fc5172be0ea3c6ac2e00dde061e49d99af25e6dfc76c8c36944c34e49ca55ea2d6b62ef948e21af1ff27bb8055a156ece2571d3cea0428a5362d03e3c0db92338d809b063bdabfebbf0c92;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40aa27c15dcfcf6db4a75bfc18c9f9ac589c6cdf94ea3c01f09172cc643a611ddd1669b204c60b24855a1fc97b8491e09702ae8f3b9a3174cb69b8fd5a70dc9a46f515e1e8f10a52d43292e84040b111b5657b593;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h151604cfc2ccc19255efa8bcf966ee063b04047f0d07177b47353ed847d5276920952bf4ff1b58f42711d9926a57ef0a1240ceb291625be187861d42155ca1afc3bd532ad59dd5657cb3fc00d9a48f2f1489f213d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3214cb33e1b4d4f305498b023bdf35b57c00e3c01f7b38c634ef59ef94b15e07f4490089c02ac3e94cad4d04fd35cd7544c0a689c461aa3c768692ddd74431ee23981f3ea02af13f271cc019c3d97f889f19224e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha85a821d7f3b71f2c4d84dd0c7c7c03e5a0c1e235ebff128af86f915c605736d62a98c1798d6a661488f8e5dafceed80e28c87f02537d901f9f36592b3d95eed7ec6fa403bad533721124cfd283b288ed9dbb0188;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a61e56f7fed71005f9ce91527ec9ad1fbb8748e5d190095f3ec9d14f8f60e7aefd38c7fb3392acf05db7eb8f1854bf6234a8bc85d9dc57f5dd6d52c837ddd10231abfa6c0376a84e36a81ec83d16c21385ed873d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac77b637564cf0891f306613f03dba276a81002ce288865b18f25e0885ca6152461a3c28bd78e889d3555382728b2fe775f6e2651386ff70112845cfdbd77a143f75fdb7b52cab26c74b23a1fff160337b2e9a6fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59a0df27837069bff24f36e581bf7637d5f0d074db5c624888602ee0f266b50f477ddff3ee91822303cd45b1421917b156818aea72950771750e2d0e68d6e1f217a77516f1685ab7ddb5d00693454d8f9cb7da690;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h460c03e446a78638970a50ec15b82b097b366101d5af386697fcdc2f9ba8119ed8a2c164d4cf8700cc7f175c6c0f8c355a8817ab97c1f4dead63b6292e099792feb76388b76113838cb3e79929354682c3afdbd8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51ba2c1f425a387adee272159cbe3f379834569f7877025603fd7e4837a60447b6542b63bd3442dd872d6460781168acab300b37026cc99a2dfff8e984f99007d2d605ad850320bc9aca1b35b49418b34177b8d62;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a3f2b010b5027febbb0555fb77d498b9a25e05b967d4c031b2f1908fc6baf6133941b696190c9804a6bc75366067f6e753611df0a8de8e87b40d5df946f9f6bec42211ff83834c6f7aaa73e55357d0246de6e3bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6121651f02e10c459eff9f4cb5eef86e68378dbf698d9b0727f94974aee7c6b76546c8f2f98309ed7adff8385c6d0dec47db8a43b5e29ccd313a5b701aad0d622cb3ec743eb6b1f2ea543a93a084fe1476e75862;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d80263e1fc36255361fe85d3d3f69b4478bdcd4e2dbbea0e10d71e85cf0cab84fd6a3beb38f5d0fb3be0c4e6d7ac73e2116ba9d2a29de8470e33c533c007d07189cc6e6b1bcc9a28f164b46761afb67453063218;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf922b4bdc57fb9ffb799cdbe3e7f0bb783ea1ec11a0994102581b0aab1aa1cd7a2b79cf452adae5f212c7bd3f7d69c8718d2682834a7b8e1f29caa8c258a6012e1a1f5180a673947d7e50c0e916d0d42b9868eb72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3347b87b5822b1be92964aec29b8a3b44622883e616a20f2e3daa1ee0348efd98f4d2a372fcea351942e0b891cf158ef9169ee6b5378841c5b38368a01c144a16adbe15d230bdff00ca277b9a7624a52d2cc06d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2787550df3b7cbc7f90e1ac63bdf98a7a082cab1b9bbc74e29eac3b68050106f4e785ca5b78979ac8ba45688d87064a4870089ba73331f27f38ed37f5e60311c7444a6ce79a28de0f85806411c158652185b9d712;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4114a4ee6f9197cfff525dc8e54350005e89ca5d978d17fc382bef112a2bf2f1417bd8345214913de1b4b19c8e0d0bb9ee736884c42a268e47eaf5a0deddbc9e1c4d8c7080bf242961bbe79f94e824db12ed54de0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83eb7ae49d161821de9c4dab05e19a6dbe3b70166795f78a83263b43d6aa25c260126294f9e64cec3ada81a43bc1a35c875007f09425a545063fae78cb7aae25ba69593c9e90fa753441dbc5f89b91402ecc67dae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h742fd22b5e97946c8456eb35a8e59e81c470713a5cda8a13386f835ba193c33d3797321c6a04896ec62d7d33406908e4b9309ef6159606c1a65f4b6afe687ac10df9009460a14eee36a520422a9bb795584df7b59;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b8f873210b31f75f2ec541d165b1884da2cb3a7ec187090e6b0492d57aaf9134a98fbc3dfb2e7c459767464d1636d0ed1b19eabba7cc60452b22e3f72f7eda5e397e43b9721e95a3d9be1be8cc3bf2acb89f1ad2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1376750c6e0776a007023591cbc9c07ef6939f30d4f9260639250d518926bb32b5f71f273aed43493430c26ec21b52aa056b4b7808d8a8524eca4fc840fd1ac4bab7d0f8caeab8158901646875a4f396d5c6e0532;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h347cadee9ac9ba8c36a21c0f0808d048e16f4d96e77defa4de3442c272c03e13c487002bb7c6171bd69609d9df4e602107bf304809d9ba5f11a9102dbc1792a367a49d1816ab04eaf81803ada322e84d5c702d5c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd83335dcda71b03e6565c926d0586047a9c291575bbe837a13a4407690e39d4d48311082343956830aac0ef48c83516de64f7254c0afe778dcf8e5e9e3a97031ae1e547346ccee64178d1f518f0f3e9091868662b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0b98a8459956c0cee8058dbcb9059cdc9ad1e526097c0e9987236e5737f299c63c6179acb2fbff92d028ffdc74a65e30c604fe39bfb077104fb4badad4d0cd5c3d2312d5a9f9cfa4b4791db631e5f1405acca551;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2986c7d6fc292aee0db339c754389e170972379710d855e132d81e03f254917c01e3bd4be0e855d79683bc411d45392624fcf99581a5276892a526ad070a60e4effe28fd0ce0a5f01de760652d5498c2a1ebacfa5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdaff6666e3c8db1c65a8cfdb5838274b5e1381607ee14cbe9022831dd04b7e9304f35a12d7ec1f763d3671ae4d35b2759e662a97f42a905ae15ae35553f49273d4993782c737cf4dbc8e1c954a93bb6af0cc3bfd6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3df0d79a66064339498323690c737ba51b5110e02ba23c16582af7d7ea425beb2de2ed8275497411814b22b0b1d31d4d07fda3444ae702765cb325d0f2d83a4aa256a17dbf6047085453ba002360d3e14c517e937;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dd2e7ea3c59325b00cb64eb94dad85ed508c793605ef1b6f53bbfc7eaa55b712bda9d601cf32de1b05214f5dea95f94798910f366b69a872473c50759ade11a982e638b55cfb644c4591eb72347e250d79d6eba8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6662e98b82578c43cc485d01e2fa03bc0fb5318b3fc4b0094327ae712f415b01082e410b366198234f9f2811c1645f54888f6ba9c065cb8ee5e76607c99fc19d635bd561ffacd9ced9fc464214e86e41f1ca8c37e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba3db9f58d54324b696f26e6f1f072307c79def60472a8f463378d9401512e8e139f67b4fb47642830291d3a9b4fd91da03558e7980fd6b41f223095a38dc871b061a8dbc553d14fd7fc32b49f092101b9c41d4b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he26b554ba45b90b1fde8abf13fb82bea5f52adb89f44a4a99022a257bf32d908aab44d8f6e92230eeb227b090891567cd019fa4191cb408a085d74806670150c44f810a18d87cc6bd4b5e2efddd2ddc77b3528522;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ad8d10d95b4805a2f5d5da49b1eb14ca072f2e59a9213a2a0d9d8dbb26e13f5d06696dd68a4252b3acf8327b042cfcc6d6b023f181c093ddf50454d9d915cb22f6d98e674487217de6ca7e16c4f05f449be9118e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3c21289a6c3c0501ccf51f39bc0335e055d92ed19ab7c65429b69eb5744d9cd21d3bbe7f470f7d62d72b2d6e138db0a11108e3e8111474a6d93d49f5e1b5b92036b4a7d6a4f74489c17e3d4d183d8a6f57667eae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h423caffb57800e8c575f3c5a57d12167740e21c09ca9049944d118e9e66826de977336ef66f073ef51befc2404bff11e44dd023e60eecace67d8f2e4186123259b546d39d03f1f55ef7adf6c459726249fb1af58;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81923144eb3a4dead869a9141f7d7351cae4fd12658238a568755bac9c8c4917ef08bcb9337709909c6303b1f251f55a54f7d7541ba5b5bd3736820313b6eae422e97e08fe051bd1a96ad1e59f7eea6ca369a7776;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fc73b8d43b658872c68ccc8df772eb5c1df3f0c090408316336078f40afc3391ee92a266d6c57f2b96f913ab389d1924c3dcb20eeaf84632cef3ea5ee2a09eeb8617e528ffb88d55f4448a32236f515629d0d568;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h520a55a678a238bc5c30816ccd24f7567db3213164ea2e0ada84f859e677b792beeb03a78b4dbb9fdec7e9a97e36d0c719ea3a2fc31596352e8f4838f87f75370dbf83470475a658ba25351afc26ee2adfe7c7240;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha75759a9a4133011f711db6a860ee366abce88ec85c86966b7dac20ae27d5320f44f746264cc0b98c40d5758731c89bf3a099a4fa0b6e838d0a24538bda167877b347b4b62266fbb43acf39d0fe0696fe48530640;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha063b75d3c91b87eeb93199cfa4697a12db6874cfe840575c85bb08d20a043f4c0ef1201b33afe5d106fcf65bd52ee229b1a9b403cd11d225bcb548c64b6a2356f13790aad5b589fe79b0f1de9c98952c5eba986e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h705f5e0f1d9497edd8a2f5aa23e0e53c5a8d11f2fc4b4f17ab6f905228a44240c8fac4fb4492ca449793eda9d48f1f374ae3a4db9c9a3466bf459bace21c126b9ac7bc90d1fdf856a21fd0e601d97c9c3fc9a6a95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7178fd8038e95a58662d88f07ac84f1e5523b3cb7d65c569fd19086ce3cf1e5e4154328adf46389c80df55f24f1b9b6bbcf5ea25e3dd48599dbf74faf7d293e8c3a92fecf448949cdeb032254b8cf9ca44798323;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd879890ec35be187757b240ceca17d93d0524c08260fd6d2da7cf38a876a84c3c7e5870ccdbfb482fefd01762383c383481da096bb8375dacf3ad5b3260c4d2577368e1e57614209aeacde4502e8c3deac60b1e2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hece5becbceb431c4c667c283cd92568073e2fde78f62d3a981d97bceceac8fe996e9cfe1dbbb779664465e1911c8946c089f405ec23cc3328f262a3eb28d03dad2852b0bd7ea536250d5decbe7dcb95f1bdb7057e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35823780de4aeff06c8603e821e77b65ececbd017148a5cce7d9482d5e5d6e92ced2ac866b27b4f36c118e54696c6b5ea62885d236ec232b5a0a6e2ebb69d6bc7239ce68cac831eb435f95f37d021bc65f6aee1cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd51aab03c88967e3075e8d25d6bd0b89f0dbf8177d22fee929a8a26e2a781c74fc51c4eca2f652263d8d7ee2082fb42d673b3591a0b5bf6640b39e3c05b372f9213ea0ab6dcd10aa57944113780edd07dd997dd6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1e2da549c45886843715b6c493606df29785672e7ebda986915a4ef7f78507be10e6e93266ae8f00c243886a96bc258b279ea036e6168bfceef569066728ee91c7e4668aaa70b425b168d00f6ab77b85aa9e76f1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0fc223375d80f72aa33b885c5988799e8c56a542920d13bd868d4a8e04f0f3335dd2215dd3d3baac1ba28614f889cec98fdb56ff7c70eb24573d30976e8ebd82232c1faa9aa0ad6036c144edb09e578957683aa8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32a90897db95e8ced40ca84095f923fe0d5afce4cc97dd2625edbe0ba3210ac7f4297475cbdb56af55d21141bef5f5749697d63ba77d89c4e74b4158c453a9d211f343cd055b48bb09deb7a6d15ec94f74a57646d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddc1f6861c5257109acc593668ef6d760be928f0a1351d530da60a9a0fbddfb4bfa26f253f15ce9c8dfc36b8883d8ba609069d7b328973aa5b5f789953bd59747fab1b57c4be5dbe96849d1bbc3a22f308ce0978d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68ac953244036b5b59cf83610a8e6f1154a3fffb61ee7ab1336a9d4e6a3ed14df72b4ef17dd72dc4f9c94cab924e458768c061a98f0186e380994306a876d43810e85f2c973c33b6ac2c95e6d44cea5b10b89bfe5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h128f07a8d8bf3f5c12bedf28e834c5acbe9767dfff2787824757e960b48aad5a06d0fe6eb60dc70af4958610eb3dac6d8a487365e54720b94afa6965d934427a0bff5995d1956f16dc0c117d0e2164368b6107875;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha81147753a0f2a90ee63944fa8df34cac788347d44761b77b417351973b0c24de9951a363a106ad3f6c01858efb4f2d77a729acc9282c3bc20699a1a41aa71eb2efa2fb6809ab2ee5d99b97cf3de84891c38af8a7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha28f3ce78ffb49954d9db6c0e0ad4425a983c78c5c27f6dd46a777a3971c357809a3c2d66a76c4d899a15b134c515577308e19c720d0f589f1ed52fb8ac5c4b0b8dc9b75a2831e19f3225a5e9b1fd6286270521d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3eeb7da647ef2211ba16e3b3ad62a2d93c478c93e5173c1035fd85bd68b15dbc784c0e0ed60a848ee8d676b1edb683629fd80d9e643ea515b62375000cccc815723d6f68d0256caca0a77491701187346f8f04abb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36d73cd70e341906eb32a7e56c34886cf1acdd5bee1e649e8dbb968970eef15cab6bf99e22d7856e471cd0a645644e9d57107e4112c1e74577d5fe769421e7cee75081322631cef281c27d8218b56357fe9e425ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ae41c9427f3813a94c7d94aeb8500d5f050b5759d35c80827d6030202463c1c7b141061c221307877bab4c38d902013b637fe0fab9da8c84e7504dffb93604a017b8cfe72e2829cedce3e4118c9c0b252b9ead68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5277ce174272bde518156961683a1563de93df29ac1c520aa0a6fe978093b84aafdc1288e37f425c11ae77821dea78db5c276767718333bfef46fd761e5094c9ce74089154a188bc78d01188edf27a3ea8ef4861f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d665e66bc54e5997192fc93198155736afc8af50ce04094cfcac9567473fde6e124d183ca28d7a9dfa64ae45191158951834b6d9c67c12d5128b38bdd563fcdbafa20c3f6d8d6b8968b017915a991dae6f1110e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h985bfb06f8cde457c1d0de1da33983d2ed4ddc3fc80a1a87429f3ad645fbc3c881b492c0f2033276b0865dee13febdbceea75e4dc205d3f9f610114ded664a78adffd5d554a2f991f61118b995485c5fad873e986;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65685b5e303718298a787b05682488cdaf233690ecff997fcf481ff440fa12964a692d96150b0c0e101c7a7277ce023948cb579dd67c26b0a711d58741b2d7140629bb91efdb7db8800464560e51bacbd319d8cce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13472b3826db96c2fcce72d16ecad1888581be350e8d91787a73ee6aa66ce9159f87988537db64674342ab9f9fd237e43849dce191ce3f649456fee6bb37803f347520ee2ab86ed3db6f36bf84eeb50ba2ad40e75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he97aaa46c2302994915cf8781170feb9a21eff498d1a01a7f6493c35acc299b7fd5ebba3d7a9595a9b6a317a5313c34abb38529b736cf06d11b28b984faaf16e2f399c394692fef828a2d0205d7674f76e174c09;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c2d0398e0f1c46d4c790e39efb90f24066831e3e4fc531c629575aaea80c2a0da42a29c42506086c8ddc1abecd37a5174640fe5f781e39f6728f71ac253f9436a724785af9e293921ac48b49ea7f5cbd4ccda2d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12a4e5f476ae3b6cfa2d82e09a944d76eb5858d570ec7505d3711aa668e2ca1733ce9789c702b1b4752fb7b168d4b156d844788f25f190fd26aef55d8a7937258560c30549ab71ffb08f0995586c424677ede2df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc3aa9e28ee77491b6b27c8984363aa82d34ff1a2e653104b4a92880f7f1c04bc7e4484d23e05abdd16230256395cbf184f7f2c5a1e401dc2023427d7782d49db94e254bda70f1b8ad5700e6b6d478181920d5abc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd84549c8bcb1b02172b701a11608aacbac0db55fd8987f5548a9b74c30511a8f962581ff995e924762faa1842b555ca8b8ea4cc939d2218a298635bfd34642c0d4de08227410d90dc97ddb853aa862ceb1f76bff7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3bffe98c4a9cfb0165ae04dfa9af476f0729f2b8f20fd2c89ac58c1d69b23153d5ed810236a1e070714c37e4ee0229dd004dec57397e07fda2be15c4698c676ae569508be02d35e2b388a43c2882c57ef1c7b3ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d9801c93d6ce47052be4eab6718c86ad3a2d5033de5f0fd63e2589024e9555079f53b9218946db9a9f0ac33d67f6e8dcc5c6bffd8c7114348fecc5751da97623e464a6df7e12d7989fc0e419e54da5cca74a05ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63b010841e033a196899a98891878ef3a3be16edfd7a41276e9b429ce1f16ccf92769fb6f7802dca42f206b0808f41b9dec5922bfe2c40f526c67668c3102194c1e8c025845bc1e8a9055bb7d9b152772c5df304c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2165140ea69e1ff4d5deb35169e9285e87fbcb11e46252339740c9aaa51187f01d0dacfd1cd7cbb0f25d6e8f96aff7cfdeb48d1373c774fbb78536d82cd730dd1e2bfe5567ef16a82861d1f0cb120ec3ca1dba20;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bdef1ddefda6f11afc3d3cb19fe1a1690f9f3e54f6b314a542291e1e1d7bac7b8608e702b3aa8bd1af2e70d46455b68854c03628f62e303069ec5f51a1c4fa48f8707934c6c700e4bfcee6c7824c2dfc5e5427ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haed1a65ffe5f90d2a9f7fde11b9b73b7b2f61f935e976fecfd2789ab231802ae66e5aba0b1263259a35620ec3b2bfcae007d1cc8736e0dcd6ba8a2c6f65619360ac762445bbcb45305a62031aeb4dceac18df2232;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h634548c6829ad33609d6bfbb3fbc35b27c5063dea5bbc82c700520af88fe15028ab46ddc48ee205b35adf27964d904c5db0a00c85fbbfd49a0e83bcf45b18cb1de467b3ab9366a2cbda3dfb8552437c9b93c24582;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa1f7847e9f3d82a366402ad83998a773d045ea7c5ddd1593c44695a2356cdb9ec8a06b8c99fb9d8270d80c48544e5cf98814db80029135926593fd083042b42aa667cd5c520285dd8b55ae492276af7f3f8cecf5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80df75b6feaf3b9f5613afe03a60c728b409f45cd8f27cce8071353d7e28b5792c5cbc919d41ee11c541095b918041a715c1dd0857478b73323d9af4dca3dab12291754550b8809b4bdf2eb68fe0872359583a57e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3057d09d0d12fc4bd89b152b74e252d36656b9db91d2ae2aac41b77c3eaa6e3df2ae96850ee49d9b761703febf2aa27976b6635426ef4da5eec81188f4530693b79d4115714dd4f2b4dfac6832b05358e371cb598;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1280e639acace5a39cbbbd23bf54097aa3f9df3817e158afcf796e8b4722513baf6df56d82f520879b624d9756f333442b5b1866b8b6034b53b86038cdbfa835f0f37964add37c3ea98a0b63ddf88598330f24d82;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65c0cd05dc9597b0d5be0a8e10a9b242f9f0590e39578e1fc50cb2d728f9df43259c926b34de4e6b5ee8bc5cc34b483d5e7962b55343c9e6d59df4c72eb7fa9272ea8421b046cd58095a9cd5e6c5d11e15d1ae9b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbaf7e0063a1411e6c08781359291a6f0b840550294c05cc5250ed9a336317364263f62a7a83af024d485bc4880ed8a8c27af9b3c9664c40e27f8c28effd201ecc4293eb2e370798a94b83f74881beef0f40a2398a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e21cfda3a81cfc5f36033bfe990a9ff2a030de3a28a1a85d3448cacaeab8db8fb5d8483418666337bd52c0d84bbd313aca242b8ffc05626a106ab327175980353de873a12a9df59473a5269b48567d6f5e6a6241;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67a8bb9903b8ba02f5b57445bba0656e38ecc8e1121882e26c9ced08d869b07801e6df1a2fad90fd5895843336fc8a0421b44903009b65f59627153cc6431c86448826862b188110a20b90d844b6ada7cc79caf0b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9d56c233f5411c38b71003ea7734acaffe137fb1bb72c87a1113c50b7fe156717735ad49375e6c8ad327bc56e2f2a6924b9c3d991212bb3572fe3330971e3236e7357dc07a0cb13e9b2ece817a6e9294426640b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75fcebfe0b68371095343e338b4d6f4889f7d3242d9b1260ea16fe648a4a34c49c161305c5ce61667b71b4446485e0070594a4c95a3ab2e2782bf86d749c0d1e896dd980ac26cd57797b5fffccd274e4010f60793;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7794324ed5b8c0b7cf5f17e541121aa526290b5adf1143cd2104602f2e34336717ba1af68d29ff82b153af12e95e684bf441c9d5bd1ccba19cd9006d41e039e80db7117249ad83298208e9c46846905bf125de0f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83507c797f7cce692ba41886183dd4f8b934b3c7719dacefedda67562d0baf8850ad2c986bca5fa1d96f98ab513f8f03712c5d310e1f88433ab0cb9914f5de3d7eca095b994ceb5d92ad27eb89668dc45e15f6961;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcb07796e28e262202f832e06357702ef1fd0ee0a3bbc2ed77968017d0cd20934d13ae8b43784f847c741f14475c8ceb5f6276cc21028f9052bf0ad7369b71f5b08c3d178de54604ce693a96244e7e38b4e2145bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78427ec680550d03ea068b88ec1907394c322881e5125732364b565bb6a0e64bfecc77132590f0b5462976fc7957acdb81654950b43bc932a39e2d64221a758b8196e1295993e737c8286e1b546f69b207ddc1e21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7354fe69d6263f06b60781ab8dbafa75eff06c7ad9c3da8f8e2c6adffbe003b339974185140f056eed5489afa804256f6901ead2d54363291b93204042eb038dd727290a776e073e8601c6ebc5806d5484fdef74b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h194ef6e8bdbf92746de92ad7e0c1e279934cdd8256a93166bbf33801e4288fc8ee546a60e685fd9eb14706592f56e5509efcbf8a95ddad1574dacc0c42bc0cc1e5afebc61cda781aac2c7b01965855a6b58ad48ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9483df54ef077b041da67f516b0761416d14c28a1f2d14bb17afd9f2c50965c36801b8e0efd6bed9e804e1ae095b8542f5b48248210fc96a03a2ce23f64997be0675e4f6cafbba2107f84cc9a2c325984f93b854;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h159ee43ef501f884791b763fe0c16a937aaa3b2a018ce56bcc81fc5959a0ce11105dc6f83891566f391eaa0dd0691cdf7a21e34a63bd0384ddc269dcdb2ee6216fad1faf0e5bee6ab1b9025baff31bb5ba2ae0c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1dada88190fadeda87c85fd02cce678112c57fa0e3ca441b5b648677f02518413d92e5acea6e8cc0ee4730ae52f00b6f4cb69e0dc2a03b3be4a38c90a460e5cbca9691dedd3bed4ed96492fe35638b67fd9de848;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb50ad764915b1424c023d7a4bf2081c461812047b07b56cd2f4893a82aaa162071b7fb8769c0f09a4fb930d3b3bac53b9ad1eb2d4e9c77657a76b532820ee1e64a37f92f9e8708a95a2c3cc6ab04f309037013777;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c2626749c4f629de4e12184c00d7044479c888a4b9fb0086c148cfb4afe6d418910e13d852ceff9931e4c0a797388b4217343ab5462c1d52b96010ca9fc9cf25ce215932cc7574dd2c5010021e121e473ab5399b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea7797b1297dd442a92497ef2bf16bd53e22f5ab51612742e4a9c0a471acec7295ca29144cdc2950c03f927d6400da9a91182ae4958c66c927ef3ed0a6763698f695b9328b5400c2239e4fcb3f6073d60820fb89f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb656f5405fa374377648c100c785d6b5441565bba7947de2780de8eaa898338953bba9b1feed32df64c33882ba2d74f915caaaca0ae3e263ce944eeef6a66c99d33b1ba9cf439657cdb2e4fea97ead99a8a5a702d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha86a595ba9a96d0191a0244abe2d33c374261b7a23c6bc90942549d4b7fa92b33c2988e41663715f3b09b5eb55213329a4aba254dcffa4b822c6db525acfe99f79341977773d8724f0fcd5c9777517bb6af3f58b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h531a0ec309f28441ab8ef457705cb196ca8ceb44c22620b430c589de97e93ee0acc25de122c48f236594a5a64f7acefb50703c6c7543f4a6ef79f2cd59aebc45f479aa10dce3bb6eef96adc1b464f799af85dd953;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h732f8bb1518ce57d4d0d1eba17095b5684ab5b99a1b57da988672bfcf0bb8f7e4924db9dea54edafdad987637552465770c0ab9d87422aabff7af67f84fe4e1a8e19a53d8d633bdb029232fa72ecc87a299639811;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c8d648733835a178e4a538cfcc68763ea2762e5ad76fe92bc696f129c419de99776240c63a92019b31f75dfad9832ae58b640b1769e2b2362020c4a4ee4ef6c5f396c0fe4b3618dd7796077bf8e67d2790fb3851;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5a60096d1be9c1f6a6cff9eb799e400a9ef5adf3a3ee9e5dde412564af6a382aff7023c326ffd3221db0f5fb882977812a55232c7f57eb74541f66bfb73dafe8bc8e8e4775f25d6d19e77e512821ed2476eafd1d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfadaef8e5caaedcc4ec6fdc2e70008da2f7fa835a01c55a5dd12d5c95f262e23b3599038657079d81f414c0acfd3b45a0d3a51285d603c69ce606c5d41d80736060d055c2fb2309ddf8877572c06ea7c2aa95f6cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35a956284db703d0e05c9be05b08e02efad6bd9e7f3c60a76dae3883bd0c09f8b273d7680644717b0e241b87237a8917411d84e819a04a961d6d4ac3ba1404664fd10034cc2b1c6b14a0891ab627e358e6a9148c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2c036a62fa0b0696a0f69ed9f67fe78be11dccc92cc0e6791b1d0d803face637f1bfb6dac271e7ac7151d8e99d7270329d1a55173e85d529fd2646d5d6cd7b103f3186eaf713fb1dd2460d5bfad7615d0365f2cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2342180cb3877b6f0106f513c9000ede96db0c259edd46630a5edc63dea1e4e08964111590d98393ae762e26d65af729c729cd580f45227900ba7ed85db69d49e04581a7dc9ca03c4c990b5308382082d2d3fb8be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb22a54d36ebed5bdc8147f1b11e31a755d7147a83d98d297f3352f90753bc7aafcd49221292cc52ddae8ce03c69b29ee01b0d8b49caac971c1f66d21f9ef95a596f9c1836672435d8a489d42cff10685be6da1356;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8dd9c74eb9598148764fd5f4747dfa1c52336d864340faadbe1db39a250cab4952afd0d2400593250bac730174a2cd0f96c4054588fdb603e63eaac322bbf45dac20f2ed48b7fc66c9341bc348530cfe575fd1437;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8011ea4d86c30a59ce18f2764724739896364c239bb7b61a83109d4fcee37158073724496f0f1d7c88d93344c89cc209b39632e5654996f1ed8c2522d61835182c1c923f67d9f0e4022d86f93e7679c885d43bd09;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb161ad43cb3f0a65374e31ccf44ae457f1f763d1e504f8d240e02561186ff15528d67a245d2ee841511f6cc66ed231544d310386b66721616b9c22a177fe7890aab848dfcf20206117943f18b861cde332bf9523a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h949774162a42a42ce090505081a405b83f42820bba09f77f574fdc0de64f618d1c1da3399af26a97f12d8e6e02af7c5e209fea3dadb2053228e7fe30b03e8bf5e50ad6a7dbb35c7bf1783b2cc8a601fd2158aa669;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87b4cfebfc5d9b3cc168f3d3b7c3d69190b7610de88b8ec952dc68ff8143f0256481e0684f0ea7ab140f60730097409e1787f37784190debbcbe8e2c9dc131f87b579de9bda9c9210dd0a3c9d1125d1d86a92c693;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5919a675486fe4bf99d059ea9a039220d2e4c2e2266529156771a81f43eac74237b8d9e052c2c4302fe46acf271579758d8e0f46bb33977870483e1bf961c4b9816bce79f2119053a1527f25831d70967c75ce902;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74ce956c858ae87895639a2aabda2e6a54f5ca027c409c7ad8bb590f7947c2192209b8af920a036cb74806ee2a99edc2b1c5a7b51f002e8e0a2ac5d3264c8a3acd3e788896a9e43a9bdcd502d6b466b34b36599fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc25c248303cedcbe0cda16f67051783105cf35577b72c12aceb5f47978413a8dab5ed47318cc4d7321efd3b2b6a8fa605a6ce396cad943238513ed049029b37b5b505d62472e1ff574a62c604832f9acc64ddc681;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h682bbb1b1d41d8dc84b492d6e97c94c14414ea08eb45ffe4cb945110396d070a929c65c6ee9920d4241cc197e969ae916351f42d9291bf6ac6c45e0080acc4437b1b4f352ba3f85b6ecb3988ef8381218b27cc4b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e57e2d970a8bfd26c8fc9a05d4203ed297df61ba1f095d5303b5965570b8c84bd396cae843442bb958a9c2883bbb5e89cd2ec7b5d84f4dbfa2a6a297280313cb899f6ab96fcaa9f245f1edbb278870488b00d1a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9fe465b846fa4cebcff6e772700884b8ff1f5729daa272b4db38e6c550584f67ba7e39f1fdf6c2c0b6296fa29648671e05acd35c0a7d4fb7a6f91a65bb7c51093b16de016cb1d9485caf2b1b2c58f807b4d4979ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b9de869af6cbfcaed34de7a11f9f03b003169510c2e3c2be960936a68ff2726792112d14b55a69930f5c5645a5821d41141721015f6463b50f29160c0883697ab288c3fab4f14da6b423b03421df0493d4490f2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4579cc2dbe7aa701c9f22fe0dda6fb33d4f3c177de7bd918b1125b918419e7ddfe699fcd78f5dee2de289aaba1fd1a5de1253d8e9f7fcfa31d1619dbf7a75717c3c2317380f115912d6129efe6af4ebe03ec2e5a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f8585b7d3ddffa11b0f24239d2ca2c09a4119bbf3622e9340c052072976fda73e5758801f22be4f61109c35cc8ce9c907536863e01074df3b0b50dbf4e964daaf42ea0177a46a67cb694026b244ac89f8994328e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68cd91f77471a20861315ac9e9245342eba6649269a4a12f0c952be29b22046b6c4d298a9640e1dca7c3644ea205831608e12b89c1416282e28c72a5af41c4c9549a493d1e8274367283d1c06f3f91bcb14b23b16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b76a6cbd350ee82def02ff0babdbe04c7c567f7cd17ca84dad0400aa3b5ecb50b013f8b86aa4eb42a0a80e2c42a3664bdb852695dbdbd955fb199571fc781120331cbefdefbcec0413a4a93cbb77f1b24f0ef4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54d09772dc5bed56b01334c87834097aff79a5f861e92eb5f7d195dda7e17d134ecfe6208b14300fa4fea244cb33ba11efb23db913fff1d93d06e400ecbea86b010ccb9cfb6a0dce1af86c5dd247c8b1d1558c24c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbaa83721f1c13eb4d2db66defbfae88d3c1d91da8131c879da00a824a56c3f5ea0b5bd1c7e647cba44b3e8b1fbbddf20b5195c7928ef40470aabe9636719c6a778ca242b4f26293d44fd5be3f680809b50101ccdc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h838a3dcf630c151847646499c860e614e08fcf0686fa92df33fd9d74b25f98e961a7b3e4751437fe13084f7af6f3f986f8b4dd7db4094cd6a7d28f0bd9706a486366fb2af8e09e1cd50bc1e25c6dc15eecb051af5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57f0c5e9f9488af60a8846c4241df316f68584ba3e1225ff56b19ac1c887d88ee28e6eb2a75b039e36c94897d7797c439058016900bc95c7a9bf2d5bfd176a9ddf73f50efa50b342f6c0d3dfa006f8677a8716721;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h279b3cbdcdf269aa934ace803784b83a733aa1e69606b8f9df5920e175ec827de4e6f7a53e536f756c4fed75f7bb41726c61f9236d4e3f6a9ef8197b026043a1bc4aa9f372f7aad613db04704a2d2e66d9c45dcee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27b508e7034e8fdaadb5387dcaba2124de5784833a451f60df22366f89f2602a4f907564fc6a2d3ac5ac1ef5c2716885f09ae67a4f1a45ae3021dcd89bea6196562a7329f3883e1754a15f58f95d20cf6fce662b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9428fe336ab4a49755973a0b9fd4f85aacdf491a86d0d0b9e7119f000e200e8697741b753137cc649d032988aafe51731f3b368ff143a768ceca9e8e1be2e8ebf4869a39ea6ff6117443396b7d1bc110508833df5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21a220dbc7034b8a6f8aa764cbb0de775c9b0e5c9242a6dbe27ad032b5b95f0f25d59ee2fde87c7fe7d67d9813513cd2fe2ae3e3117596cc58b512955a57ee1728f43de7278462f1aceb6e47950425d800d5813fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a027cf690f544faa045000a4ad2f065cd65faa2a500bc454e47fabc3a7bbdeca9d5f625f05fe4427be868e1d3603ad45167eede0a00c0c6b5d94760e9dab45c8d33c968be52d629a1b1ee72b350d94657cfc88d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc42bf3d5832c8bfdee4447ca1159f7e163096cb9d4be4f0cea3c8d7da348bc6d051f50507db207c914649a7d5b951c89648f9dfa8f2d611cd661b5167ea7480e247dc4090cf1e84bcbf868838ddf5cfc891add7b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5dac67d21fb38522581321043f3fb56f2dc9cdaf2082f0368699957a2c5c751400e61bb15abeeba60746627735ddfe67a12ea591142b8e7a4587228e149a3080d9bffe85162ec7fde8e838c3434cb6dcd378162c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47c11f114e2c46e31921ff13724c0803d5572da40578ed88f28b7268fb1e4a83e50764b7f95877c20122173060ed0184820f1f3b9dbf742015e6ff78f6c2b6b470dd2789af3e4fcc6251c96087c4407258a9e3e61;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d48f07b4536e7de00b1d32c18b8a7b571082d35e22415d925c2864d44dac6092d78394011a9400955bfabb5e1dd51e2aa72f64da5cfe3ffab2f78b30fa6af8b57a4e4d9881c3122c2b426e681ebba294dca4872e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13f517ecbab373183d55e35bbae0d9da70b88e69d0ebb7967091f27b037b7f150c9d759bbde14042e74f7caa52abd04e0c8a3ff5b72c35fe0e40ba47b421563b771eea03ecfa65c187f1dce4b11054b83d4e1cce1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9199c707c4e7a60bb63d7a8d0712338fcce1325a6678af46cc39c389f8242f64ebb23f3f2014fb457aa2d91be8606b60f1345cb23cdc9d86bf0269386aa6de820059aa369458a364891e119a7137e47c1e2c7b233;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1990b88664e6d48da5b574358a73086372981390f07765ee6eef007a8876ca8ae251cd44975c692c63e642141e659320a17b33d967431077e4ce07c3844c82cbd3bf4fcf462564fe5c3bae8ec55c7cc063195d9b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfc01736f97c6a1574068b65066ad243038bee592df4528ffa6cfa9d9eadf369cbad162f94ecc0f10f83a809dddfab7aa5594b75ec9c220121f9f73ccbe687c1cc4c4ff02cbc1bb5786de9b04111686ef24615ab8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50a3c6b1e189048c8fd20742dbe5ef963ebb3602bb9c90932fa2e3422d8dc7ed6c3dec9bae78bbb994cbbe36f4b8df3a1bfadc905709ec635de3b2a652ed467da4aa7ad97aee02799c68e364750ba0a956cd34aec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca1bde536ead6dcb32692ee556bfef58f14c30d484b346b852f0fdf7c944d372fa5cf6549a68d1561c63c58d8c73a936ed56c3e82d6660f0e69e63509dc901047ad75d9d95d89340b8addcf4c44092bae4cfd77c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h380723ffa00b4c95e66f6be3e904bc20b544a1b72152e68086290a9b09b3f80215adb2f84780097d6bd94ffb971cbae917577513c68678e0c25211e439fc0564caad531f9901bd4defb69cf4b318a8a3e45c4f85e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c607f83bb2903ccb6b27670bce6adb5894eef0793d045eedfde608dc7c08f135c1f832ae4bd955b05b33a75ced50c3579fe2b39e9cc925b8a041b25f1e0f0436b1cbdfbf524a6a0f17d72084f09d9ad6baa6bdb9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he14f932f4badb9376ce2ecc3e999858017d99e5fef19d673a3e14d37b400a0d4cb7b5ef4d38ffb1e48db8f6f4dac05db748436a6ffc1585de55522ee0040495d7897e02e6825b0160ea2e94fe982e3b8348c753a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c7c72eff41aeb2a569469f44ccb52a3062a292d00e168e6ae1084993a2f0f2243a2ce2fe8b87db9fd64c4f430d434912bd05a99eec6000f2ea12aa40a0b2e75a4e15148cf3c124b095d54ad5fc344d940fe70247;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h524cc31e671343081bf70e96cbd79a8dce5daa319a827976768f44c27c13f94819a66576cc282365c56aa4096955badafdc2c638567aa57d118e4168553b28e2c627b8aa9b2f8c383ebd8545ac4c36f0f3a8ad258;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8530b048a1efb0126438fe3dc0a8405c7bb66fb79031c44b3c96731da98b88aaa492ecf60a1caf75d3102aac98a550358d03129225d8c26bc7ab8d9ff356628f07775cc4d2c183934a70999049e24df0a1a8a7105;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40c50b2cfdb9bb745d0f76ade25f00daca38fcc94890a3a98aa18863369354ad35853b5c7148904fda01892d99eb946634e53b30a40915239a67933810e35759bdea566baf59b1def670a2aa2dd8fc02bf7998221;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe0a47243931f6a20df3b7c6db778081e13e6c001cb8869c6e4f45a74eeeac4a5f868391e85922a97cb1df7dc27bd48d97b4a087b7ae5f8eeafe35c27befd75639775bca4776b64a82c1d1660b8c205435aeb5446;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h645817fcdb35c99468cb64016955effc34900dcf0e320fc35c7430c750d4f18a49907eeb801e3b1ffffcc53da91d3b466700b0090157b7b2fe2b0d4809697fb92562fe50f4200171e4b6bd0adfaeec7eac73b5c45;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf45e86c27f984efb040dd6fb111a498daaf1a1558f6890a09a14e530805d75d13905492790968710da4312103934ddf3fa66ae2ef6063b0a11ebed256d24a5d04f205de5ed2275e9b030132093917c02ee66c0286;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cc332ad747fbac8c46ba1eb4e3f5e74dc32366145e38172dc5ca5b48141e5349a4184ec43ccfe5d2d8640dde62798acc2588cdaa755f3210c9e96395c5bc99aa4689115cdd185c361ea5381d7de6f70b6139d52f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha45649e65507912e5b7ecc7aa4e718ede9613329754b08be1b646153ed8368539d726a3b585b4aafa1d362b6726c1efef61f54c105c46f4cc5b1b0ab0e48155da537f7ad1db1b015d75e7d76943a9b2be0ad70390;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h129f419d12502f40a5fbe16072d8e385dce39473fccc2706db5248fee6089187db0fa29e500a7c014534bcf51e6ad9d0446597ed794b32d77a609e63797d6864d47cdbdf0703c429457ca8b5c50098f78a7660a6f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe29d726885b7e1323210d4a3584f07956e1d614c98dd6b618252b69e4b8b002aa55b0c6106237cb5f2d545b559940fc7350e2a58d566b95fd1e09ab9df1d76f6a2bc6ee13abe7bc36a31e13858e0e7fe956ae86a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha391b2981a3dc38a1874db8e0f7ae4ceb036530ea510b176e055dc3e68dd8cc26fc293b83a60c9e51b8fdd2b8ab0a470e38c221b508f6b35ace08943fb8ece402ec1cd92d798123941eb644fac5a7f7abc1c840e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9388ee7a935b7ec4a43fc3cbdd90fdae4014c0ad2baf7be6b81a1cdb203fa514c1dfc445cc497b5942bab4c704a356f6a72586be5bca6fbc739fbdea024a7afaf9194989554a62ebef5a025c8598ed282cc14af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18799ba789f2c604943ec11202e33bd9aa28974b635b0ea5b1f2d6fad8cc8712f11bb00214006c37a9f201dafbb9e9b77e93fb6eaf5089d981cfc72953d673ed18baf4a2dd2649c6dddbf9e0bb0cf0d30e0b80f0a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h416d88f87d6bf2c6d7b1e55d74c4c13945c1132a19a201d7f016814e519806c463216059f3741688697ec961b6462edcc6daceed534e9eac5f5f1c5d107a9068bfeffddfa649d3d1784192dec4b03eabb548c1f71;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c109e9bcbc389b74646f45fea63db2966f21ae38ac2ada01ede581c3044f83f08eaf94f24ddc1586344dff700dee8b339f96b6b1104b2675a7d79705b2bda8670d2676b8f506c2ac9b0ade8aad7ddde15e829088;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25bccfe9c396af61e24600f5de45fcd18ec2618f0151fd7d142227149d67ba23c72add98a085735a9b3ae6de49bf351f6fcccc1f2ab0dbc60ec832770ad5a05bbce7504ad88f9f4554f4ac193d5e4a4f41a6c57c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd3a2189aa89aabeffbcbb9b97aab5945a550b24c23685d79f54764806423e72c08c7f275c5ff7db0680b2499d5b5c1000c71d0b11be98324affdc2ceeb8059e3a5594b6d8015cb9af69cce36b907e12a8685402e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa54488c21b60efce5455468fd522e80aabde1765dcb667843d1fddfc38de06866aa81ad121273bfd8b1cb42547b7a2dff38629eda5786f51776591f6690b826cd25a6123299e6db65ace79f2bbb9079ad7a35372;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h177c8a7ef0d94270aa3ee01e75b976e1842f8fdaa065f5ee0854d909de00d6af11a05c33be6fed7f14c77842b6b41cac1aa4d0f49277420c3c115c45a8770c61daae44458721da1f657e6d29b8464eb4d78ef16aa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15c4b3703d0396650eeae407c21e5ecb11fc12145bec91cc013ba4a510f48293ec70f9b2cb52afed541aba2c199ea7d1fd2857ad9acd2d7e1c30eb1e99fb66a02dcfadcd7933dc6a473a0ba53816e3227d94c2e9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5739050a5d315ae7133c0a07a7e149c6d81b133554cf685a6300c2e9ae9154d0b3779c3be1526a0fcaf321f7a6b7a1e8f23723ee819f42bdfee7099a5b85b8d086571a2c30ec4e2c1489f478384b2e25ceeedcbd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f137ac216ff98f6e87fda59463126c0384ef03d13d6b5ccceb4d4b244cf82e3e579c4a3b6c0195226fa6e3527ea83875adfa27ab2a7d4282233a2e1bd9c152da85c99ede1d9063fa4a77115e17430e4769143df8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd44ed293e08029574b2a1947e26d7036e729f2929292d6a5ad746378358f2d8cad3e8342ab5fd8c931c04276071f9c0ed1892e40b0ab261e681938e0035930e9a0d5fbc1c4815593f5e2b1e2839d32c13e542ad05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89c850d38fa1dc5ce02104ec7c03d5b142090ec543566eab265f29e1fd17fd8a50445998cc057de9324a6894d97a764336d85cad42a6d1e29d02c39039578e56ddb3fa77384a0dcbd79796b106c391678e5f00593;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd43d761aff7317a727c3b0b600c5a6ba3186791ee1b8f75bb52fe1cd25d14fdc462b76379c49a265279e240f35def513b15e8c9864367048551e52d9faa65478f0990aad367360d24f6aa9216456382cc5be48adf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dedde273576338565a59a44b7ac2aff12dcfeca181d687ffac1bfd198b3b97a5f9f75dc1938a98fce5e3e66eb15bfc681ec62fe6f8b8eca608472a216dc44bc9373f0a447056db8ad56ac10068ee86c6d80d69be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd75fe3a5357b28078f297af2bb4e22ca9d345a728b8960e1c9d043f7d237853ace4c01477b189534bb15ff975c45d86400abce0353ddd5fc2ad729fea5cce2a685730409f94ae3f375a3c085d6acd8f3bb11cc613;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17d176fc97c6a481260db659125b84489887b3b68d759b32645e0af63578617510baa74e25f09f99e61b5979432d555a8aa72af9e53ae2a6a811a5deacb1cd2e22c410a13d0bf9773f87aff67a77ccd994ae5aced;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h615fab80df968b45242338d0105a278c6fd6c7a7c058462b0ad4dfb1c1e191528a53d692994309054412db07ca4104ff7a8a2aa2686a73c9098b32aaae7af5767f0f253ac99203c5c765c930555f28d5ddf9c1e2c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2ce2eaea0f94a0e8d26cf86849879053d0374d009589757e76e60fa0e0ec5d1d76fd2df59eeb220b8a29bc56432675d82fff4d6bc7d104d2eec3ba6219a412ed71ac00ee441f6e97d5366f64684152c22b3d8d51;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62bf62da4fcb20b07c9eff65850718a57a9c75c52e46a9e7c69e1a6c17ffb06972eea9530940bf200f131f66e02741814ffbc90f9b85ecd1791efdfe2c64bd14e3fdc3a7007a226f7493755e0dc8c0b5262b59f96;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7dd3406cd5011665eb201ffae7fcfc4496c5a49fb570a3894d8880f4796fc50d27a7dc725a8b97bb11f420134429caca0593f8142b93c8a429090a7fff3f730c3f0e297fbd03be92464c337b08814380d9344b095;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e08d23e177196b95810d39cd9e16a1f531d977697fe61b0e152804f06f0aa5f295f1eece10707e7f899e9a8360a8e880e6c0dc124dcd792fc0c7ce9fdfe98b23658f7ec7180ae8c48f06264f7ea23bbf5566f5b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e28ed061e3432fe3bc0080ec8cbe67aa3abc04cd922dd82e231e37c5dc5f1ddbb74db2e7edce1686b4fcd1486c58cf9b6901bd4d80468e3bda4bff43397c830e7d5e692ff4b41471406d5af27722836df84281cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h837b29e39704694da57423ac6f81d2ae3665894b9e26b44226771ee3ea79c7440a2f720815ed38c150b0d042088d5587384298c80da77a4cbbc339598baee62f8f23c86f0be4c23ce542b6d3f1296e6fc6eea73b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c5047f0dd10f21da90d4c9ad7fa028d47f94364e61a1518c1c3bb9053579df5a99e5ed976d270aec07842734294a891d8b0019fa634e4621b55045f2a4856c38a160e7436e565413104a4cb21e3fc09202f9d3e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb70d33ba44051259dab01a75a395bf84fb58a8150ca468bc8e6403a2b2d9e222248c46f1029febd1b731d13ecec40ce1388e86feecf79c427cfe2652d868b6d6dc35c8b3ea4bfe5d22970252ac2617dcc5f6e257;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9449cc7aa40531a0f3ab8d68906ca3d27768cf4e57094fdb1768b0354f2fd88477c5a32acb9f2b4ad08c1067d978b1f6eac3e1ee723266128373b0be15d25ae1ba96aa530d7dd15779cee5dba26d36652d19bb9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfda78930d0c5767f9e18e5e3d5b15117f12d03b8ffe08fd722e6d578ebf5ecab3e185c7fb49eb4720b865274464fe9b68a66885d79b201a8e140d05b18dcd399cacbdd5c1787ce5c7f3a59cee46e6d405a56c0af0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfddeb59bf90d71719d31231321ed57ad52494abf6bba5c9f7b2ad538e48e9bbae9a312ed4e746cb8a01a08e6b62d5dc1b849dde4dc4e9552cad83cb3208331b082af15add5be9150040feb6e594e797cc3ccbc4af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbaecb1db814680aa12f05fa2c1041fdbce10f40fc9d30d628badf41c44b9eb6b5b63e7e787d395b6f921ef1daf7446f0bf0f49cfb20adf38f76991b39a52ff7b3e64bba114109df18242ef7ecbf2f0a9d2a4dd8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f9256ca239e15b8144caef307274ea279506715ebf6bf00e33b9a75584aac6a8991d88fa310381443823009f5015b79302e88e3db5e00e09d09b579f45174040c674ce3d0f67758be63a689bd584b390ac927d9a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94b5e398ec65f7ec23fa1623ea413b632bc6dce7f6732e0dacba5c13eb908eb6b4331a6abed38cf8358096402b7f01da77ca159e6039b9a7972bec131a10e55e3bf49697d578079db84b4c63f863d567a3c7de1e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d793fa227b1053034a93a3d1581971805cbd5062b93d387855af6705f27dd9069d95b9032cc69c82fe5e3f6b2a6079405dc60d1e53debfc31e7b30f2191bf3f37f6bcc5ba21ed0390aea420620d6ed54470ca5f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72b1093c2e7f0be71f2af1da87db16a9dff98edea7daf3e337450132d83a82b42fd9b959b25459a04a807482b0e085389524f748ada9a1a15a7b4b0078d34ebae72136f72136aa73a24e5a4ea6d6aa356c8f625fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51748db595e3f8606e83556f3cb1ca1600755cd48ecd6aadaa4e9e5949bc52c9f23baced1734a89e4768384c865208c823c3a8870458c715f59bd3866871cc8de309b55805f3172ebcff954a26c923b7fd6acc6be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he843be5592d063411cc2470df59c1ea5e2c660bb4ba105edb763833c65b49c47ac046d26eec0b781707e1acb16b3fdb86bfaedd992e23f796637ff4567c2b921d3f61ae8ec934310ae9fe5384936acc5a85070ceb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb00ed9a360fde0d11b02fffd22f20027f2e082c42691423e73dcb403f7060d75b51cfeff8a9940590b5f4e52dd3dfd4e4d63f1761de9ab21d244f9a7abb2a956f13a54e22fb86150a7da00aadc6df207b3a5c5938;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79b242fe3ebee88ff94aa52d99047f86c71db384fe919d1b626656969f44a1ede70d71558aa6f10173356a0397f6af99fdf1e9612873a7583323f82d002e317760cfe4b2c613d6ca15537ea15ac0b3c8f56e9f589;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb3d127d335919ae8226757315bb778bf2c1c647dd225b1f040d8b9527c797b35796ce96112f7afdf21a4e36f425c05e5206f0fec26c8528f87d862b183b4d3014acffbe82a487780df652fc3892611fd51ab03ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he8f4952d4b0e6a79feda40befaed1f1e0c84357f5c32a9ac11daef3cae1a78f5cf4b43c0da1be1ba433e845d73739ec99daf81b59588848bbe8a8bebe7d80351aebfe68de3746fbb7bbd43dbd30eb50de6b5d9e4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7617866a231629f3af566423b4bbd19d791d584dbd4b6028aa2a0303d3dfe17ee18f935dec83db32974ed58f6c7133cd0322c535c27c276cc79b7a1910b2a79c34fe20b7d3f99afdd24b726fda25ecede356c8224;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h130cbd105ed53a9745bd9071e6ae492f250e88694e48e2ad9b776a37ad1dac3b9cf6eb0a219e3889c94928d6fdb0bed10fff527aed6a059c75f92f21b4e36f1fec2107e8482d69fffa5512eefc6a600967e6e2e85;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc09c0b9abb1e3047ed777d741da4cb8768cfd63158a56bc991e7eb408c483e0173c47411dba0cef40d3e75aebf9f517c19c416a1db7f7764e236999ebf381ddf2434b89fae707ba520041c361c4f55977bcbd23c4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h165e65bb72b810b65c2e6c6fb6cca2cbf2f416618aa16fa93941936891f1fc53ab096338f32ea9cdf336d27424276e26a89d969d182ad8bc15d1300574ea45b5ea067eeb9b394ed943a9bbe1084b578be17244037;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h877ad6cd65daa191da60b488246810f4f1ef187e91cc76c55726c2ffa2f5972ded21d02760a59922e4bb69e6b84dbaafd832523150466561497784a411a4c0343b5670343bccccec5107848b8e88778f7d7e7df76;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf315c24c045ea1d65d88183472861a3e62c4880b7236b9d5198f5bb615023b76c1da6551e204b257484aba7ff3af55a09cda385560034b9e711ff9101ffabff59adb5833e82336f8b8dafaee2ac9294471d87e2c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha98c7915cfcce9a5d3152e1ae69f4ab2b33c9fcc42231b5c1aaba0132f4ad8edf88f8c8fa784d51e794aa87d1d862373eb7c084c78f786b880b26d157a3e10e2b9824cb8e90c951d35c35f0facb937e0692b3a241;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1756da1b8aa9279df519b694f193cd1c89126d079fdeae63bfbc3aa938de1863c05de499d263081968a2a88e9b07d6d47eee30ef4cdb0b0edb29b4bbb732ba49adb11fb3dd30c08e6f8f101ca2e2324924fdf3f4e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d435d567e73ee71ceb4166474cc6c07f4415418c2145e25a1fbb477e88b6720a3359fcea092718d5a62dff62f926a32a3661ea7da948e3b1d22372a4c1bc53fe9985d9a87f67d84d02a868f7e60811ae140d5fa3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd49b64c270c318730c535737ade115de0752100933c295a927a7e88ebbedf8fe0b00c74389fc92401dcd2f85f42ed93ea8fb78bdab9c8a20f5223c1d8a3039b23b94f875084c5222616fe0f5708595d0aae41c51e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14eb93a4fac0ff9dba7054df8c38d2a829e77363abafd8ffd884c092c9f24fe8a8f8d802138fc5b1bf99136cd75be98989ff6c3b4da1e4610b7449be66f2d6d3fd126bbff15f3555ad6c92ea3a1ec049cde326a38;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4ebbf98c6e690cfefa3b5b1767931a6b604fe511adc618a0f463062a3416d58d04058919ed224211f4ef316f4ae5639a722e5c8b4c1d7d8713806f21759996579f5a37161b8eb3fb09340183dbaf51a0c978ee7a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5316fda9a556480e654d1da37d48d2754dcb83b5919dbaafea8d248fabd32b99868191816aa78df0fc0ca7ef9dc08d2b27c354a5db881091958480f246c766616d430e1297a8521faa28274e45b6515f89b4d425a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ed4708e52a0bb22ea91079fd214546276848d753fa7e9649fda508cf08f5f61205a5be0cabfad467dba246861bd5e245db415cc7db787fba546aada3caa188de26ccc30212daf2059f8be185fdfe8e5eda17807b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49f8fe9f83bf2d71cb665710a3e997532bd207af4fdf05719a22cc03b1b802f65c62709f96cf0e22a24ee1161143d2630e12fbb5c03aef28e95193b74455fdd7763013f09bc759f0012992fc2681a74740a2a9d44;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a104b9d2abe26d93e752cebf71407e6369e828224dd17fc997e043bccc1b4610030f704c904ca010ddb463441ae8d2cc6c7bd6bcd175cf03ec9b4dd33242f9ed73bb909f465cf494731ac2639ef43354659d4cc4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1cc06bf59a5bedad63e15e6f278a602b26b698c74ad76a1a472900296c138a86f1beb72e18dec9b8d6be18278369a5f6ec6c7faaeac506a5feaa8c772add76dde0664a8277b8cad43fd6522e0e3044475791bb9a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b26063319e1b0e292977c6a75aba8d340da2e1bef446efd77b96b6321c9bd86862c4b90d4b666eedea7942c1905981773f86f9f34bb21717417426181f27b65ec7edb5ab89a5f1f2a7bab0bfded60a2c2ace35f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78dcd6a048dbf1005d942e8adcd6b944d3b35c5d22eb0be2c666d46275e929b5fc70e736725453370888771110159295dad55ce7618ab1d865b6e11bfe148a627cf46ba7a4b22ba365a0198a1eb6b4247d1641425;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57c2d190af172958fe51ff807278cb7855724e30066cba965fb511f803cd97f815f086cc28bb60621f60a32d90e4a983f91fc47b509f3c320a4319e951663eaa9735104c17da86a9af6976f1b969d604be187082d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb34b24793987363c2bc21035eaa22d05b7725c491e714c2c7fc21c52e7a9f35caabbe63063b941d2fff9c4363c4313ed78c7eeb26c37597466a76355439891e6b0abed89e380e3cf0d9ca5cc4b2b186f67f0cbcc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf89895b1b2401909b15c86e89dc6d7f5fb13996193c3c3f342bb20de47395c8e29854d64d85e6eaf51ab8a6c5b05c2e8461472283151c5180f9d59bc5daa06da6ba272095c126b96d15622078dee6c07c74340a96;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4ad336ea0dccbcc390b36d940348e71ed54aec5ab5cef1b12a29684d4eda9e44ae84ee55f3564f5ba0e3fb7d27496963306c1338441087cdb973c430a38feccbfd5a960a0c2ab69d1418440bf27fb542d7cd3b60;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b643b8cc56406e4dd0a918960c1ec66092000ac51ad89ca7f1bf5304319c0556772273c86b9b63fb8c9fb29c4ac5a832f4ae9249947316de42e7735c8ebebef3b4e4303d0675868ed7ada1a564eb9f1f772bdf22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9a41642bb0a0b73b9f2a0883cd870a8ea60c76ba1201402c3d1fa69abb88c7ea18c2e1554812f7672a65f761107889b32011a10beb6d7adf3ee944b0b9bbc283f6475b5ce85fa2c5a108ef5f2f4df27e256ca209;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4e507d15624f609e04207afe7112282e9b141db941a1ae20e93c7ee79b6086085a848cc48f531901fc1fb1e6bfd9df8bc62d2725c8470a5d59db24ef0e96c220ec39bfd40415379dbda67ad8223c87a955e481f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ad21e8437665ac17f0bb6fd6150de69f3ee322668d657373679ce321959e34cf8c2e451eebf17a41b7b7c6a8e9cb1a4f6b759c751d8c616e5ea2e24610c910eac28ab710e807d02edc07ca060ba0dbf365639c59;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc665f9ffd655b1e5001e7d50cec5ca87754600f9ae145333b7e644b57d0acc2992842c9c226b2cdd3591f09a738705408a7bdae878824a61c5dad847df279e653057e5051b8a57a6a6148d731936eb8a6e15693b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a045fc2d22d99828c755d65b8457f1ccb0775a53a73d9d3da746e72558a7d3987956ea73b429328b90b3a9becc1c49db1d24b2c76b3ef13f930ef06787e6a2582da7c4bad901b661ac0e61721b5592bf848672bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35b732681e426dc729323ef63f3ac24819b3385e59b20727abc3924709056c6f2ed99a15298ddfc71a42383f1491f90e9ad5da68086396e11e0c18992bcdce41478a1bd60d213f842c884c1525bee87d821e835e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbfe8a600ac28107bb49c6d31452e985d541986935b5bc8b6fc9a99df37b238d9a8a35964b44cf3b380725a4141759de8fda747bc0aedfe345c0d5ea89981eccf05ac0bfc388077c1b02322ef03471d7bc029dd69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h967580fd595b47b8fd74cb2712a20206d6be635a6d971c44b62a8f081c811df34c33fdbdc04249dbce019b29525897d24d6880b72b4da6475bc4352dc6c6a4d8b88ac984fdfe5b1cc187d5b321522b99a1dbc4545;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4744bfb244e12ce599df2437a574a2673d8d481d95ee265c91e7eb320d0ae6ddcd133c5d62071955152273114401cfdb335692373b2d6383a0b0a268238e53809f5ec971de7954a7fef19a85ea621b21083f36f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dbe7cb86602564343fe4e7e43d9b34ffac16c0c4480bcc032ec0c1de8d7fdfaebb80d2e57383cc3cbb878f9a3496b0d224bc5c8eda71927ccba87decdd36d8094309c8a61d0c09d6452559920afd0f22528cd982;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26421bc6b115f58b81bd4ef5b4360ee272dba752423bafc05beeda4ac381a452edfeefacbfb8f8d33fd6e2ccbef37202a42ad8a7ef2c4e60bb03a97ab2ca1522cf47bebb0dfe555cc264db370ffced865ce39d483;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d54c34495f8e42f2c5adf770b1b9de23e3da8ffa9345772e283c122561bfa25810db80968abfdf24e04690f705b8cb2b14084accada9f8f9daf81aff832d1884e4827d369b7489d42112041e5a1614003774837;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44efe67fe26d542a63b9e02e7b85eb1d4a94d61f10ec36468fd621ce062d6d0fe46cece37573bd8cecefd4865caf48a999c2fd7a1846c42366a7286f162eef0e5a480db361dd1323f4db5c52a237ca4891b54a02c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b43e43e524eca31ad761f9fcd4b44ca843b9b3819d49f793ef6702bfc7d38f9c0aa6fb7bd9c28356aec15ea0df00e409ff9172f4d48ac7ae148da12d3fe3c8d2fec0b03d5fd32e03bdd7206cc218523c314271e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h959351621e2a48a0886d9e29dde53f74ab3737c1d8baf9333abe6dd5bde805978cdb001fe56ca200ea57c151b737a4c2f4184a4e0540ccd9610946a634db112277843799987f07e0927663e5298fe84239fb0f3e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h640d59b7e1d22ec8a9b35442de2253aeae2f268db602a157fcf9ae9687bc318970358afd3620a7c2044de4a8145439c6cba534d4b7809640a0cab1bc0b1a4c0229680dbabb61094e71e2437f70e50b0e4f746447d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e1a62cf98c1546676cc917b784933184f8caac28a9cc667092fd0159a35a5fe54d73adbd925d1a6a06f2e6f9cf0d46d40fb6d07caeee486e446b17c9b4a4d2ac5496829cc3a9251554b44c557d9d105b34f89eec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he57bc312299065904aeb9209b15821d3bc147da8f9df956d99a96321265edc599ed71b38b671b7999dc6f9552e15e35f9082dcdafd4de555a3c3ab068e16976fc7b2f7cd5252de5a6c44fd79332b16165c521a191;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h935b28d1e987c2f1cc229410191d94a3836ce36b4893aa1da85e20d698fb29f87662c0c4e72a2b99297789974d7bb17b4feee0d7a5df1760391ec420909f7ccb9b470639dbfd66060b70a6e0d98166ce90098b7bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf42dd99925c16fac9f505e1cbbc9244af41428b641d696117402edc4ddfd0365dc7ac880c860d0ceecd29af01d08dc42ed8d791e07c9b957879c4723d706a4d23ce50fdacd17f246f769745557341fda3ba506ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b5a010c1efc891fa4920e85b9911b4ec1405357dc0a94a68bb2f783da2a3e0e07b51c2b36e1a63f8f5ea2a498784b49a248adf01f15f84ee8aab88cc026c83ac9ec5aeca709d28d9675b2f11406af7a219dcdfe5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h285ea6eee2b2e4c72bb5d61c650ab462e15db1d92eeab1007d9aa1652218aa2629877a5c21988d44039d6acd4c24ea0baaa2df382d5c421e2b860b2842e1a4e101f5f3c3318edccf772689d13663597d021cce036;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4804b1b79824952de487cdfd3efc3994a0ce548a263917e3f400daf061250d15df1691c985c8aa33f2a1298a41e512423eb9b2a5a3bbb12e66b1b5e684ac79e3fe071780a888408e5101cadc438a1a5b3088dbbef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hccef6b365f9b41052bd2ecfad32e7d3d281b743b52e43ce1baaf252be66c82b85b8951fde8fe54aab8af12a9b22eefac290f5d8dda200628c81030e20d96d10c155fca36203ce0559c45ceb75c3f94832b765d536;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8d4b221215818b51cb1b1e1a64c9391b751aacffbedaa0afd681f4974ec612a610520cd61406c970484a4f3b6f4dec8203afb12df4d28e307ea8ba978a4a69ab08ffd8addc2e164d15a968cfd4be4b460f4389e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ad5766cd6bb3a14452800963fec20fbd81aa89029ea0322b26404b2e27a8ac8238b7c0a23df943d98e0d42e63c742f601bb097091d5aa5eb2da9c9f11f02bbce6d3e64e0699d469a5c573de0e953f30a3979a16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4729002a292cb5585d65fbd06bc2992194f2278f44c4b9ae0c6b2ab122307b98ec4c28ac4fa948551f32a113aded08a260e1251ba28ab3879f067f709fa6586c9842577a14a517661e2c0b8eb2cbb35fb44cd264;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2def1f2f39f42aee3f8c5d610894dbf2257bcae80dbd5d9ec4769d84c753348b4c629b1480e6013ff7d4eac03ac7ff859773eafef7b551c3adf1febaad1d1046eca4a2a8cc43d647698955d78efd61ae82238f071;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfae32b07caec650cd352dc18c4c2416bd783c566b3fbc2ff08eca6c6785c46b2c7a08a8eafaaa6efb0949d2879875c86db4e2e66bcc899bfe211b4758c4ae4e1f8aeead5b9f499a45f2d6f3a497cb0d3a23e929;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66df6a0991452ee5d177c0636a45de12cfd43439f17e485596e5bc0dfa60f384b03f20d205ddd9220225c0da05cf67f279f25895177dc175a8e9f2b59286513f711e67b565f2a7e79c60b3b063c2901bba79f95c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cd00a3a27608e4996910b80f3718c3f4b7861ed3f9f1273a94a771b822a96fc59badf39d9621af41057689e408746db8ec94744cddec5063cbc5fafe6ecc7adfbed2a4e4bb365e28241c4596ccaa93606550edb7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5f1bf2c940b8a3f6abd63401bf38df3a0593516123fc2c698d801ca8669ceb6edb26f2c2fa1ce6e1da28347a4e1eecddedc31832d3bfbb75e20cc52c5745fb9c7eef2431e477090e5402361ee1cce5f6aed38b10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h230137ca811b3c678537e1fc6e3bd7f54822eb94c40f4a3cccc6ca1489867add244e635263d08caa7b9b7065d238bd7a7753eb14f8fd800adaac98b3ce12dbb9327e9ec7174678bc757824ff98d04251305d1dba4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2589adb6471bf1499b8d621aca27c01fe6f5096d23e282ce30ebf6f2955cd20f296cebc338bda43d0c15a4f2d072502f0691f4f71bf9f6aa9ad22fb85bad63c73932cd53a2d2e0f18e9d58149190911570ede8f72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h390f1d8db262e0887b7bf49c9f5282d0354b9a23497864af2dae575cdc4000c356e878f85130980b98d330e87cc29ab6fff26c23dfe140524c679f031a9b0db33075a01f3cde42e8490527a0678f8609b5c0f16ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h323a75a57362fb526a5e2b72cc354f993e924863067f84be4fba396dc4581eb40c80469e1050d7936b785bb5dea07cf4b0d37bfae2eb8e6ec6076e01d13cbb674d568b925f0cb7b772b4339c8357f9b69e0aee623;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8ac998176e6b8a9973c49d930470ae521854a69c655d9189453588686e994fa88ecabeea2bf61abcc6828eab09790dbf3ebaea36e6e9cbe838596eff4f54ef413e2fbef4e30dab6c99d80c7d2fb336899d5c747e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd43646259474794bca4a090dfb3d4a25c7989816c09f7adfb86ae75f100bc4387da324ac3296c006ac99d035b74a9ebf91de92891c289002db63f2887b796b26ecfecb269def1cb810cbd9a7ce3f35bbe28b78ac9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfaeccbb9bae5ab2a3285f43f5c76b5e2c56517597e5dc81832fe8aecc073fe87b9bf683cae7642b6c162c764ed4ed81d692cd7d0121e6d88aa74527ce387b4e8eeb1185bff2d4f5039d889d04b3225402724008cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45fd3a4551cfbb2fda348ce91ae266974cb440509f37b580c8c0ee75e1c0d8e9443f20b162cd036ac4ba912a73c99ed5c3289d357b52a459c2b97763bd3ea76de7feab9e302c11b48d232add06147a1e87ebe0d21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he119adbe5805b1546d7e2bc1890bad25f09749da39a80ac9a0af33ae7ab4085dee11c02b1bbb508bef0ad491df11a8a46c6f8e4a06fedd2f5a600863b2a190107b5aaf2800d1ea6ac1cb5e4615330162b848b1d85;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e258b0324bbff48ab7a63f340148a9c8d5f03a9dd1b2a5c41267a3813c5621a9187a7248c1e13623775275850feb38142adc1b7842840bb5535a4477c8c885aa20298a1327c6efd9c084281d21fe5bbb4fcbff9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4324ef5c82fef602a21db924bc0d57814d939e227d40e1e4a1a757a22cbadcf88f938657cb47b8636b03459babf5e6022cce40c1f535010bd584a9f116a32650570339e41bfdf693a53d84841a956b5a4363c17a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4443fe8699ad2ef0055912d618de103d9f85fae8307936fdb33710bfe0d565176516f4429f6e2bf4e05971718f48326d814f30036784ba78d801a876e5cc4de2f32a5382c59be1eed6a0137a061422029f3060e39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he94cc45301288ea85763846800f7ed17bdd0b7c8f7ed3b2bd0bb4ca2f27f9425759c1cc6766e1bc9f332fa4bdbf6a46beafd030fefc1b5ea4f6deb13b73505cd76e479f86028c873f38cbfbdb61984f196cd99078;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90d477a84252c3d35a593196cb0484e8b6affc3938fedad13f85dfd638b2b834ed1641fdf82c58138aa5e69c7f0a7aeeb33aa9d73ac9b0e1816e212dafd6d1163d44fd0ee8eeb26a77f6df43ea52e19125662f7f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56a0a1a1f280d6a931fdc3846f7538e8438b39d8792ff0c25eb32dbbadb29fdd55dee8d4c7dbf2bd3743ad5129defb0f19b38e7d56afa1429394a2f1fb23509410d29f732c66c85716c11b4494d67e3124f318ca2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfaaafeedbd63d435140e5c22bf237d17599caaef291f781cd09f3f9168828d5223f60a8277c0991f065b88da86a4fe5a2b8586dccc594bf16bc8af10ae8a356b3fc7ad71a74748c8fc97424e4c27fe7f1f4e62b48;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66b7b70081bd0ddc5975bccba6f1b21d276c2585c9566863b8b2070b56b9708a097d720206409d1a2d62e0477ad4e7f692361d69a25601edfbb7269466590f4f69bcb9fec2429a975bb34ab3fd2a849ef6970b68a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he107922d33251d5b692ce0c583a5c385e3cc3be963fe0ebfaf1d6965694b5cf2d77abe351aaf3f24b84a819fc2034a749c672975622e9867f5c65f055727f834fddf7b45a4bff175bc2149c9cff6c63a7709f8f2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59a939dbdc43eb03d73e39b4a92ecfc4436fc5a836296e56aa30cdbfcae342e71197032aeaefc4ea91a202183ed636382e4ef01aba247f3a3b5f45a2666d4c1b791eb4ee869b9b5af8a9fcb280c97977146dc6b16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3fbdd08ea61e76636788cc3adc4aa0a868157387788536d5abc89e2335773897c3bbcd736d5ee7b532bd88c7f110f3e500489bae17ff885981fa158399041b0d9374314add09d830eea53390949cd9373aaab277e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76d36114e6ca72a03c8a6abc063e564ec59395b3c3bec5ce7e304251fa5694345f8579e2e9132b187892ca74193442fb89364f3723eccac0d05cd50ec17c1d6c50ece9fbd6778d2cc1b07298fe31bdc37dc4be984;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb653877bc0f669b7db60972230b9ffe83fcafd665bbcf7839f02c138886e08816243ae1ddaf8c609a87ce6c73fa44b9d29904fdcaae5cf781a45f107696accbec9256eeb3209a2daf81553adc81f27d1cbcef1923;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36be75282c5ede44363317a6b0a5ed3bad732c9bbfe693ed7c92158be464228b8ddd37b4b107426636acbfa3bc98f2818ee2d2dcf8fa938129d7602fd68d1baccffab7a7809f8aaab0b52a07775437d5383f2b84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb397ef258d35aea964eeab9edc5abfea71011f040fce463b57264375b8dbc0a776ac695a8e9e0ae2a3db000fd7c7713a2cc9d77e853a6c539191d4a2c49a6cee7ae4ae1f742831f4b1cab099aab641bd61310e412;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0b3179ccc29d61fe55f584500db9b0676fc97d77f384a9ff8a678533b10ec31d0e39393936cdc2384b4841eb2aeb913495251483d1fb363c7020290a87f1fd79fe67fd5a283acb5c983a82f6edb16dfc48516ac2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd551a8d85e3b51daad43bfb8a8645c1a97a34fbd0b6e44700271987711a6ef09ccd1934a11b29b900eadc94738be46ba8d65e7df0c179952254d69a6c854ea7c6009a63a77842013d1d7743e772a6e66a9442c79b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0308cc01f35c97ca55c6227b1ac25cfab8a706edfd0069c289663263b8ca83c8c765ee6c6eb70712fbe1271ab5087cef5da0b440f1e89b7eae4baa0d225a7feafc37526c21eb2858d97d1a854d369806a69aeeb3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6dfc7db53b338690eb4adf949784c7d8c485504b1ac4eeabfc0bb32fc7f35e13e57a9e1774d591e66272529680b6efcdfd74be197b0e792c7102c13730cf3372e0f8dbdab91ac0e4089abea8a533fff5c6747588;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc955c0a88d76f6958491bc4abf4a107b39b5cdb2ec33dbd57d8e4d05bc117f82cf798796c1d69e8539b5364323dce3661bbdf602f5e65f0de8ab94b77eccaa4e402789fec50f0af4c75fe1d015f62b8d197b0f9dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h762f306054e8d8c67076aacd48fd00a423d0ebed0473625c7e1e94412d587f8dd0afb6ace826b6602b89b7e2476129467891271d32d385123984d002b339864a0b871a59cc3eb939e209b896617d223dcc2aaef33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h190aeca1c220c2954f35ae5e406e478b4caf43ae75f5eb4dfa72d0c36d9078b71d02431cc668770bc5ac96256135be208a0e8648396ad5e353b5d2aec7d2d8de1d44663f78cb42a04b63e7ec3b90ded5047f7aede;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e13115f903f26adb724262386bd4b750df27cd215bc764dd857284d3c177d02431e64daa6b9791b8448553f6cf4eb9efad6568f7d7feb194cdc865d8844bc020f85bcd093cc72de491ad7aba40834c01325ea560;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h338d7524ea51855799587524bf260d838a3a0a1999c34f32495b2397ac7625ef2f0f764b8d176a2bbe67cfb7414936bff546aa4dda3935b89c91f492de3a0f12554e9ff26320e6811ef50397f113ead9e471e22c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfad54c4523c9326044e10a087c2a74e13477f69831dc8612b04ea4708fef89b3990675d5e731322063af49cfd155051bf7d188a4c99104cdad92cac3fab56398f249baec58e0cacf9cd5082280568b6b6d8fd663f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c437560684376f8486d7c56f664cef9d22daccf18b441c471ee5fccd26f360e9c6883565d7fdfafffea2ce257490fc2a983cdf0d7bf6f4745b312facf2209de1669fb4f7348bd4e3b4d25da370061d47865f3a3e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6438c2731007a6ac1a7ec63ab29cce5c160a9af601dc259d035bb800911e448bb9f4236fabeeb2a86c187885c6c2a99b8cfec7fc8c36bab666de8d692d115094cb91f779379947be73f782e55c56992d6f5b67fd0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f1f0edc69fadab986f711de1575322fdfda1c0f8175aea4d5a0f4590bcb1257be1198a55bc4d9dc569f847b15c0da70dc0079f8172b6dab1f59fba18846f26d64158271feb54d90aa981f0d347b06eda5e9c2af4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1004b15e7944e8b4a6d334185d23493f921dbe92f0152d40010cc67f9ad4f0b0e7351ae9bec7e6377e072a0577a87af5957dd76602b187a7ad8441449aad5e949b0a45e8ec445b66ad5758255df2c585a78a709c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9cd41b899dd7ae460cbcc1f6d04a7e460d0fba6a124546198eb218475c1e4c64f7eb92b98258beb3fec6a8ad2c5a6e7bdfde485d5c2575a3d0e7e7202c02a7fc8e5e27e54181c430bf337a64e7598be6a16eb3423;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0f301f90566876be5ffaa5271bb1ddb168901c0e5935d28c05b4c597e09affd7d0b6a0902a8149fa573101a65690d7b80faf7ca1be3fecc436ebffa3ad237e5c7c9041e701af2c36bb9737d997582043422f97ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46c148da2fca6678b8138e44cceab9d4f08f1d59a428389e47329e7ea84ac975cfffccf4e0a467501329eba7f9ca6963f6839c67f2fd4cd09431fee1cec7a46f94054caba5a4fa9ec7bdaf7d24694012ba6e3786d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3676773a7b35790297c0841f918e1599edeea5b9a1f83151011c1d2a161af067ab84755f80fb8e70533b8848f830ad9e7983f94e90340ca420a4e57c37b17dbde62ee5b5f92aa1986350710e72871751ad5a5de2e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc55a513e9c1d113f30f66e600b96132b1a81464f407107c9d9740d600e3653db499c5febd67d8a9770cf681f9fc10173045d2799a6ef9ef873a43c308462f432d00f832af162f14b1875bbaed58eaf5a3fa01cb9e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6770e7b9fda444a3fc969eaf8beb2f40aab56a09b39671acd7074b18363c60ef373b1cbd5ad9909e5b5fdcd5100a6ed976f7a0c287dd504d60035808c3ce41a9862ef09a84dc6576547ec7409b08016251a31f452;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17d5eaeb02b826d74e94f09c0532f2671ddc6274a7fae8f5ba26e9a7c0984cd2152736fc2162850553d5c268f50b9f60be6edcab773754f5cb0ce6a372dc2d0a07dd8defdb8a1c7c70ab8bb13e128e710b3b0a7e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6df1a398fe7606228be3135142c0a826e4b88dd6fbc49dd1e0e0eecc5b29d4af0a77b766dedb997b2fd3e429f1c0f990d1dee4038c61fc7ac84b6573c2f6ab60b65ca29258223c25df6f86b3acbfb25141cfb4c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb0c3333e89d1f35066656d0a5e039690fb62a6cb0f3baa7a795a2f3ac305a50b3ec066fe4c2badeae03600c156aad4324e950baf0c4fc5c18902c5cce602626818ab76d169e15bb438818f2d907e1acd39905db8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41fa8eab637698de97f9644455494dbed23a38f9797e7b02b31d6fd7ced9f4df58e68a951ed2111cdce71ff23085c0266d654f70f4909ca64ed1b17dcac427ebdb7fa7c85f6d715bf2016353de8d144bccd6bad72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35352b9bc1b9d3bed011ded7b1d9fe35bf99d504cca2b72f6db1a205a5ef4d6ac5e07be943351f7a2a2dd8d66f636ffbbc08516d3ca35ece8ec539845d3b9b36b5acc7ed5fd7bcc29a0ad72abfddd15e2933908c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed7e11a67953ea1349748e1a27f6e489465940f154c6574526c3e31db560f2bb30551da06d1725e520be6ae534faebb741578f746b9c2a8f74ae10016119a8cbea7e9340745cb9b9009f66050ffa902b6d598378c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacfe26804c6e9da84fec4931f2064bfe4077ccedef3b547749f9f3240b778211fb683a47a231351d2ae6cab6940e676e0bb0d7d7b160f198708fabd61cc36132fe33f9d8a0acffa107a8cd309b6cfea46637178fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd78c15690f43da86eb7de2e3387430993f6bdf563a25623de95fb9f56d3771edd6372b83ed84516cf820c159a9c580782d8872bbdaeaa515ef6d72a4ea8709d670caf8e1a59c17ba9c3e2d7842d82e760bb8a42;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heac559afe6185fa57bdef6f75a42eb02cc206f4b060eb44228d01c9cebe6c38e214bcec7acd903a4a04c1045f4c3f15b6e86473787499b490535d5152beeaba217b5b5833282a3ec111932b77b07ce88b52379d34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a929c33515a03da3915a8cc0026325cc7b8951b189e075a4796a075fc79169661e4371612a565e9761c5c044d6b1cdf88649adab8c90611fdd4bfa1af1b5b648425a070d89f20e96011321e8481e838a6483e0d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75b296e9f6b879693fc1fd159676131d1f879e922b2fb3c136b7a648140c2923aa541e93ff6fadfe6e1f3dd51567d4e03042a3b3e1d45074f6811d042a4d52a779889b9f91fc1ae165e1ca942614ca9b18fca86ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc96e13adf62e581dfaf69149307fa2b2188115ac462809a8f36a1a0f31438b151e12554da0419619b643b7de0a233a39870f226a99273b7bb61c22a5612d4ccfd20de0c237d5375459bac1875de2ec1e1820cc03;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7aeadf336d46cc674fc714fa94a10696f4b2f85893a8124d7cb49ffee82d47807d9277ce1ff33eca32e4ecf21e19361ca030497ccad38f7fec13e16f65ee267ef93a72c327356c08bc2c3beae60139c4c1a61c27;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f6568b66ea38342e9ac2af0c52be5422247916a5e03ba4e44505ac4725dfe6eb546b9a197b2de8897ebecd31dfcb2a5f5b175b490aeda78cd83bf77a32bb24c1bd258c1f5162c9ca126d96a01359796de84e2162;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3119272cbc13fa1fcd92d8638156c07e5871cf290a2a2ea19d0c9d64b06cd738424303fde8248c4921418dd38de4e81088daae4923193de781d5cf23a751ee9d7b9a6bd89b42b32723f6de938412bf2ef0246be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93076a637bdcd86b70977465fdaf9ba71ae90c8bc574adf1798306109156163b1c6e95afeae35b88d24fece85d1f38bed673cfe221bc9cc7cbd5cf981d7359e5c2579b8b20b8c634c61071aaaafc79965904c98c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbeea22372f37802ff3c81a9a6b2bcd61ed31ef082c0b27ea199b6f13fcfef3c3ed8c83e0419ae61813adb0e4bf70c064e85a66ddb00597c9f17c847a258e0ec0c94fa98d6d065d52cb532e2ad573cd8cb88e7b049;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e7373caf4ce76b38802e9320c05de4d7f0a903b77a067ab99ab88c8e4763a2c775ca36b7a8af3e0a72f22b4feae6209fbc54accaa5a9438b93f33946f69596660f4652ebd1bd34653f949c84c05fb2e0b9890d24;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e00accfba20bd7a19bfbd6bb6441b3f611cbfacbaf80a1153462fc0c097872ae0b58231c2b9ce507ef601bfcc0eb553e778851d6c9823e95d14a323489c825dc211382b82510064fef1efcd26805eabdb9fae217;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a359e9555077b3a03765f174151832f4f520bb91cb418ee23e17ef2c19da052afe9518597ffae2ccdc6d9d6ada1f96529bfb48406446f119a765c19721144b766502ad38576ffb7ee299b266bc6d13908e514be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22a83511cbb7b13c1dbaa081132726c5d8a0c6e83138c246f0a29805a3ba1dd7bfd33936925a271db97b3c9452e28deaf170c645de675271a69777c75afdc54332ec2373b7de8baa2910752576ea29f8b55497fe0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89932444b382b44081b2558a3c1e54e8e8f8ca622f6c8a289bbe3479c80e95a061ba0e97064385e0eba6ff00d8b6caccb194a1ed28f723b79e5895b701d23079a32e92fef2c8be635d1f591f477136305b524f43f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90f6e78b3c25a9e036a82df2b6e34f52ce96d527665d1d4dbe843432f4756f486f909917a37fe7411f8d97aff409bfee906fbf1c073b2be82c60807e16bf89b8599dff09e8f30cb3072270f83006328b370a20eaf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc005520de1b8f050daec550567147901fa0a835a677910000998fbfd5bc45e82fc802cc47eb479e250c25c364898cac09524015f8ef58223c6bae4195067a22600ed46f48c004c1d2450bb8d4f5b9f0cd22f801b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2dce91108c862a1e27684d1f572fc74b181540d0178a5428ba2fa030d56b27034dff239dbbf897757d03b7772a34839f5f75da02435d06fb27578d6146a057e94c7c2b35addb62ea96e3ee3e34e2a2add9724f93;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9b9db4ac4f487bcb235c7518d7eac4b6bb5186e5ad0537254009d67ed83775abe9b25ddfb1933e843a4f9fcd9f63d709694027094e9e251323b0788b2debf84bc7572232806a103a99857bac54bbde6fc369f3cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac18698d043244a454926137136a799f5a551a0cc607033081a8d3209e138ce0a63083f3a061798995c284864554372a7f2ced80cf6223c611e086fc358f75a0acfcc550761fdead57fa255350bf18df7e58c0699;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e5e556a5a075c09a8cfa2c94f6b14375cb90e35259fcb6874f0c753d3ce75e059e43083cb52aa095137e21829962b4f7bfdfa226ebc49060bbbddf999b3252f2f047f8c4bc2d287827b41cd96285068c7f12c632;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc43d8628cc3013ae4acac79fefebfcfc792aad7cd0aaf063c8833430fb5bdf1bd0d528a97ab8be89afd38ef9501bae392d10fa552c3bae34b8fb92a79e0798fac9e687914b9edec3bf7d495b218480aa468eafef2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81d7b3e157b2528b6721842159496395d0f4bd64359ec153ea00912e8fd57d7a19e30069b13c5c3deb01a52c2f8c3e81d163e7f526a8dcf6fdd73826bf8582654d50b6a1d09923a72a2b2c575e74314beb103d46b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c3b61ccad11d426842c07ffed46636cbfab5bf14027bedbdcb6ddc8c3741d0e1ce1d068ff193ed213c47891ecb90a5e8eeaeebd053062e81b3649788f41ff38ae9c3f7adc472f9463943a3b6f12a46ce9420836f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6d927a3edb74aff493849bb6231d19d3a2182fed5b7488a448b9af90383e48b34663bfdaa9d5e479f252305b1ca34d4d119c7f72a816e513a2cc51f58e76663bbcd9893937d6b9b76894df176b292a7ab456d3f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf3a96234ab4685249fc1c59e1fa615b1c45c83b1d95b4b22f42a2e9fbda372d0cc233d39243ad6fa0d8bafc93d98e020eefe7ac32fdad77382ee401331a1f53d823e1f267f938249ce92c3fba2dd551fa497cb6f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ead9d677e07ee46a88b2717d85008d083ed4f146288589cc222d1927a2b6e8310a3f35e49f19112b1c0b47fe234e8c8baabee6b4916e9f597157dfedb5e8b245b384c67afc3a1a4c5bb38997fa32b2b401869a4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f8404c74c0bcd248a8f5c7a5f19d07b47b92df8696fb72b39ed2489cfc271547e4feea2052e9667d8a26843f192fd044e82710f78c6aed3f5409c8a312eeb8cdf844bfc8a862f2e1e1637d4d9707369900008eff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79f115133ce259b2e7c12690b4314bce89fb67edcaff0c3e01f0ed4e9eb0fdaaaf4b56b736e27396528895eb1c12e205575ca32feb8ca88af4aba0410064633735c297e91707f5c073818685a8cb391594de2ed9b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe3a04d6089766ffde110cc3f885436120f8f19fca575425c617097ecc9186c213bb81d7b84f2c7627e69c3d580079311253cc6f44efc1d5ae43f63b4c7559505aa24c3687dd3c2df5198a7c99ede327ceef953d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dc82774c58d97f9c4ada3cb620fe0df779e4f30435028d6888dbb4a78c0ffac200cde2d70c878c82c2dc399bee9a9bd45c1a765283b0cd6e2bca32b50df7944793ed0daccce734d1b0814e5dac4c0b732553f296;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2060755f19bc77e919b5b8e514c7874abef57e119506618abbbfeabc8e3b6ce5a6b10a6db37f4e002efb068a76e7afeda89b0eef93f660683cf3577afa9ac193e605d7a06ceaba3ee26bdc67f1b3888b59c411f6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72f2650a55f9e74348224f08c5dbe734e604be6388b3ea221a00a739478d1193ee0bcde0275f2cb6ca8411ebb97b416a171210b57c15165ffca06d83e123d199a40213cb9787adf582d02cb9765a786befcff5c59;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h169ee450608fd56cf120af6d8a45ffcd7b56af4202d7881ced2cdc1e189308df1fe466e90599cc5a562c41ba07b30769ad305d815c7f802e4dd805cc6eff426d5a58884a24edbd8651907f73acdd81ee99ca6fd8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac4b0c1d0242a693cd59f740cc4f8bc54404695e4d2ab266d42ace80fcce439a4dfe701a29101383104079e21878b8bd5be38b81714fff1a849f6f74305b141ed4b32e8e25d71fef60419ae43f9850fdd14608cb1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc444844091b0d2d9eb13bfa4e9286d12653706c3e66870f027d99b099c875160fe4fb7b685ad193978e2b24cba4f8b0768e0114b1cd064e81d333c146fc2767fead77f94136ddfbab9b1e8b978745f6dd5a91f123;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5792074c26706eede348262471e13fd5766ab8f9cec5e3261c3b43a47e6fc64be5a35b7cbf2d7573e8488928d198b4cb3cd59a3e886a75f603ed680012ad148bf138cbd54cefece0131ab1823558e26a2aa97f72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32c80cff9a72a1bbd33fb2dc45962c8433555a198287e09483c3a601e0ebed8f71f6d6d822ae92873e23173ba076a2bbe7c3c931f81da34d0c79eb132a6d09ef94a191f040cb40ec84a8e4a0b7465baa9f43b6404;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf772d8e5ef06f008635273866f78aa7f9fc69d30e8b8dc139dbcc459ba92b095b2f61e09682551dcf98f8e2d5e6a0e504451c9a3b6f226d1b32d528dd382f26725faee9d7d592d67d6ce3d5fdad3b8f2a96c15040;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c20d0370e88020f78221a0b3525ec1093246a22c446b763e0a98554e61a43379dc9f45c61a53b7bd5331f352f67430496a16b00c2d0ba7de34cbfc42dc00698a1d48ce13d95b65c4704bf68f35c5a4ba0c81c69c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b493e565f868a3196e9b152de09facdb14ab5c779945193f16899e371021f962ac4ee2780f187b35aca4905c482225eb69562874d6d35db8563971e9394d782919e6d38212c880a58032d3f46394a91577f27814;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2def23a5f0b509ed92c645e6dd8e0d9294a7699f3b6b1d02413634252749c9f5fc17567d52fc0ced2ee576e9ca9b9b98b43df2c6eeffbe170073eb15513cf39c69d8e0bdf2ab65d9c5d60eb8315b9104e439235f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77a9f248ea190ba4b921c569b462e3c15f5e8008252490f3ece489f51979c3c5904b30ec0027285a5c8a8e4edf632cd0ca0255e00f21a65531aa3456f0b7878c3ec72528376b4aac2fca7a9a92c6f4d92a5f19ca2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b45094cedf9e4532774e3d63161d7aa781dcb33fee4430bb80451b6b6ba9b7bc1bb8136d4c6cec327a9ab395314ade27001eb1d748dfc1d80c13f88c3bf7e1f8b339304aa3c074f272baa025009bcfd91b5af348;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1e633a7bf76e03b065401b9f5af1fb8c1fdb97aa21495c8f8656933b79bd9bcbfcb687cf10d7348dd360c15fe3c6c27b28d52c928569bcd99b091cfad7583187dec226622337ba3e4aead02d4d1588d1d512c28d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha99d392caddded543b5e62c9be894c3364afa8ccbe912ea4ff5da011c146e3f34ae8e7a5cf81b7450daea83b47dcf9a3ed715ca200490338118ec0f6f626aa4e42006894fdb52255b012dfe16f25e3ae5c04c57be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41e968e56e29312adfce19edb52e5fbb679f16254654565b74b8dc99b36ed451038f257d542a331f1c769ee0d68a6b907e93d6c2fe4c6f1290aa3152f4ec84bd03aecf4d8094931614a6ea5961155c18b2e3b2c40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbcb9e518e7af805e1e4b71e644af9536f9a630fe67b82df256202df3b1178482c4dcfb5cc9ef0a02664efc9ce07e8fe2caf334096482d2027c1a0fa1d97c9e7792352309c225b13126fbe50dbc7c53fc5eab2f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h964666bd2de52ac7d979f49c1962de7fab08f12144cc7440ba4e3c557c9f3c76ae8bedb409e3cbec3bfba8abbdd610885e3f5fedf9738f3f3c0feb3ecc2c2794fab91ad82e169e5e3edf29cd2f8a657df4de7208c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf989e39751b6fae03212161fc4a17a44f9ada96ebf7d060194e2e646051d142de15d6f07c00f825a500e09d8019e103c29d4b79b3132589d29959617b8af893b61ba861adc65001c674de777b54335498c41044e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h595ef6a0723ffabc089f5a0f90a7a789f266c00131be9b17c22360900bbc19361001dc6c88ac065c6f8b03d7f7b45d9a34a6bbabb368d0b21f0a0d8d5e40b8bf6ef9d822d05069f524b19d5cabffca29f3d102e39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ff63411ec249690425d60580b17c023ca8fe7c5b1ba7399993862c721744df633cffefee5f5984d59c41167549afc3ba80c4af42d2b1ee2e0c311cb2931104cb4eaafa1862793f599efc70c8fe6599349f659651;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77af3d6ec69ffc082e23ef21302ea3d96ae72a5ccbb99785c8a03dec5c53c6902081ee0fffdc78c409863b0b8091ba6e758d25a58d31cdbc1da2cd07e2cf5f57c2dca0b959f426de8eb169179c38cfdde13d203ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8de73aa0a4440ef2d49a9935674e49da2b1ae89a784e76631feb575eb645a1da9919a92d8c3f4437290010acdb9e1d67d8b00d871f0594e42ab656de0427d3f303d1b2a7c1d7db19867c2d14a3003d4b4b5290a10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1be1fbc06bbfa3b4a31fa0b04db6668ca10696075684df4717300616f8e9c778bc6e75c0c5d292bf47e6397951840990e2f9f83083e613f4bb122c79088745c3edee060c6b64d516f02a7e509083dc2c2977780d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ef6598cb94ea4857a5526ca87d3fc45a7b24398ddc46bd421ad248efa20f10f377b395990670867a550f79b5138cd3ac1d412b3a5e6a824d9d9062492f615df875f4e50c4558226a19f685c42f6989bddb5ad178;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hece460662cccceaa2986d948b69a8062245bfe3a6057a27a566550983ed068b7517ba5f29b1112410ba36b8a5fee393ce9577e92d94efd8773844daea4ca78af5de605996a7804ecc83889b35413a886e1a88197d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fb2ae1da1a9371f93e32a15a6964e3acd16efc05a17fa4c1c865ecf42de5aa6a3b33f64af6b70fc58f6673021d648b9ca23fb0af8345e48a76666c414f8ebf16997b54f4af3c03dd8423963968d79351a015446;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h325e7bccb3d5517df866478c59060625b981e0aff1a91fdb0e40819c3015bba24adae16f7a20a6edbc29ad11415162a8b10410e2d71f716afe385f21354c8019c6bf34dbfc15f16b8779f5c112fa36c0c17006f77;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcceafeb2695bd4452c53048e62d6a9584ceca2bc3d0e8303e0dc5bc8dec8ce77fe1c9958876e57ca9735bd475b41e96417478f31efa888296fa76b30e1c2dffcaf21cafa219d171210e6ad088ea4cbc69ef7b8921;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16a498a459f375ce9151cd648340c78c7c3db3c163888e9673d9b1f0c0759f671b2baad54e7f3eb67e29df698464e4596f45a9309ca10e093f0e72303eeda7cf90eaba0805200fa2f54b6babb83854de9bfba7964;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h756c60e3aed2bf3f85ace4bfbaa0ef4f708a425e04f3b48e5c1efc2c0d523e9422822cb076adc34c6158c1defca031af9de0dea17065ac9355450cc577324f7c75c727bc8734d783d9f3fc15903d9e0c37776b48c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5568adf61bbdb81a191e60f8020394d660f0f99a2088e54f997607919bb01ae9c6893151333cba47c4156c2ae76d360c7a8913bfe7be9a466056893af495417d94fad125b7afba6d499fc3945b1b6d27ccac354f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cf1419f0328e1212db1115b05c0223ca9085dfc39142fb889dc349100229f542715674c9427a66f8358fd590491cbcdef363a8e6c06c9927e68637dc210380573cafdc87a010b919e3b06440a72b272b5641de4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77f23554cd235b8fa4963fc63106962ad670a1a182b8c0c551b1afac5d269d889dc4cd00a06f8ac4b6acc6015506e8e34b3ef994609ddb145319c1729001d3b60368df869a0c3529a225865444b5ea58b0b496e48;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d2e1f72944f14f40299f871f60a4b66243449f63dbd8e849cb84b38f14583a68c3f2f707fc806a7561e2b360ca96b4c67891140d0dc33d3136b045763ae92a3982e12d75d36c0377267acbf88612eb8ebd45e6f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5627c4d47c1de9e8549e0c314e421ddf4cd9daba1eae35cc60a92bd0e81006d0c9f9a9ce9d454b043722a64048b6dbe6a8bc078047a0d1c3b5a37db5560e0209804f0a6c80744b3f1eaf16979573df86ec4bb2613;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ecb6f608638f2a68f8fd4c9c0742ea92cfb18916a5f9d5f6a089f350e221ba8ebc73ad72406c9b2078e12d5c455fc7ee0d7a58fc554d4c58d4d574907c0ed37994e01f701d9cc41993b88c95522b89085d3d7f09;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6613e2bbe62304302a2d8e1a1673289f8b68f3e07e7dd59529e2894b2664c1e0e7fc59b823f0e5155048ad557d4aed1baa85c970a3dcce2b0c39862393fa7227526b058fd01321d66e3b02f4c0b24ab85031a69bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf38a65b222d2b9e1735c613ad823544fc5d03d966807b845644769763438fd7dcb84189c19c661370861b2603a89f0b2fda5442849ac9143e9215efef75f762d5ca7a994828d73a9becc89dd5699fa952677dd50e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfea4c9f31ec07adb8851f852fa7746b4b7581ddeb673bcf76f9d1597d6d0a1150cb79b593624dd11ca693fdd33b640d8ea271e2428996457404d8278831bdd7689cb026c7f1c64ee02c55dfbf2cbcc4d774a4b39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha83b6b1f4abdf92389279500a099545ec4aed4db2cd9f4e4e433fa8dded457182ca722f766641e1c6bf89d6a4fd2c056dbd609aafb1a2f43cd450fcf3099441b89c0096f97f285efc82d07cec83724502c65732ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee143dd0c20656343d8de85c89ec8de0967f9c4051537f9699abfe6269b60a46024aa9737fa559dc8005868b6433c8affd06c8a543d97b9af2d406de1b0514813484bf6c7da70c49d8d6de3c75839974f351fa01f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb3818a2012b85baab953173b35266a19eff0b7b0ac852035401a9d9a1a7247becb7446b4661deae0256200b78171865b2e8df0323d8e82a763309da56d40de972a1019d4fc85908cc6f24455dd79e69d310b2761;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a7eaa2f7156b554129dc736bef9347c102eacd008f535175538e755d5a3eba9f58e0d915e1f91e73962f5ead1faacd0f7dca3d3202a848ee43832ef8779d6b1d2db542113599b185d22539e24aded3510a141d9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b78189a0ce079930552dee943ba7fd13652d54c960bb6320f6208fb638289274f40b0ccbc3dc9d41fd7614316196644fafecf792d6c1d034d8f8110479ec8f27d47640c521eb802b74947bb91a4830a8eca7f2d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86bb16bf3551ddca3bfae298c6074cc1ddcb3a57630613225a3559c106f851b2ef3e29e6b9b09411896efef7a7e1d405dc8bb8aaa31c5fae95a54efc32583809f3447dcbc636c0664d2f0e6eb113d2803f8b41a95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62b77a9d1be82671d7e73629537c3bb175f846dcb8ca1ebafaa0ba59cd2968738a587c751384a9ad883b42c24d8fb011b196859472af594d7abb0584a8b37fed11e8477b712840e91babace54fa9f220ad8c88e4e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78281364d0d705165a9f2e56cf43bf19b2eabc570ee45fd038036c808def2d709c93042c986842f85cafdd274e83f90b8794e6701c0c60f4c42a6457bc8167d3303abdabf96630e220442dc3609caa282e37a3031;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h598b9584e3654e545dd046a2b322bc2325ea86386f3de24a832d998e667eabdc47883a4822b81477d2c1cdba00be1c3282dd1ea4e1e543684617d836a7a59a7ff6a7987fdf8653147a1ca2261cb4b5759162bfd35;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb84b5d290c5733a76788acfd5baa1707e18b54a8de9010ad69db176b67d571b3324eb9e0babf4361e3e3b4bea27de03ca7e76940225e55244416c3285e9b93cb135fe45087f29183a3cc2b7cb21c19d6f8ce227da;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd0d0a1b5cd39e3132e74910ecf26402cd502ab277f0fc608a27c4f1fee3f8aab5a8f4aeb95a3faa2c2bec5b61113287db5d0103c0370e3abb651b70e646257c8e3a058c344bc747bb97052ef2114b679558a927e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1be2c111a573518432c0464d50880348b242eb7394bbc0bb5c364ad481e65b24fba315ec9f21367a641f61c75c54a7a25e753643795f8df19ece68c78b2574639518b9cd3ccc5f1cd1fd2984e0101997224e9ff31;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h285cc62978e76dad30bdf5669f49a873d8c462451453f34fd37d195d1d4e06eafa7371f66c255acf381e101d34fef226d0ccc8ea9ab843eb9821ce75fbc9bd58a16a111a9667306bcb625c444dfb8878fea883a5a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e7ef4ae55ac8f57c919d4cb9b1523566145f006752a8dbafdb8eb185c87c7c62505967fe42f66d8fa6371f82351885416650ab789a9aee3056352fad235e084449aa1186559ebbf8d980470c195fb80b83b5677a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b3665fababa6a4959be42216aa8a485acbf4ee42ecc0ace568720340681f737aac7a97e65660466c08a7bacffb355572d3e444e66eb6ae36c7ea80c2af87873f93a5f5d1a3e23129119097a2ea0aa155f8c0fdba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60c930367eba05e1f60fb595159f9fa5fd152ed162fa2f33d06d747d4bf39bb753181a9002b5781c12adc72e7a9da433cbcde14bc874214550890ce3bd03603f730d08b7424737555c0e95e7e8cb357c696917f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5b4c577b85e74be846d2b724f322896bbdad1e708872b27290796fe58aec7f8435b9bca41c68747238cb0a43e0472462c9071b196e4355bcc37efc7ce6c574e23ec563160956c96c93aa0735844c68fee4f8223d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd53dda67e42fff7818be5b15d1525aa8b5f4dd0466ecec9ccd42b0063e34ed1409807d141b5b831ad24b7ee8a7271aa4965aba01082209b4168bad344e289b6555bc8ffe9cbb993ce1d33bb664fc02e67a78175ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h682eb20372dd3f400e7fc0f9e529699d61b51eb3777b2f2d6fc8170346722be618a9d18d9dea4533e09750a12b4066b9e1340fd8302356a4dc8c05595343255873a4ef333a7dda98004ae98333cdd5f1e0663eaac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9281d0a6f04639958dc2d017b24d2fa018630fae54380a2e6c7dd71c0d1a05ef37c16f337ea924ae42cf82d0cb44a194357c74a5b0cbe343fca8a8904f287fce591d0bbdbd652a802fd49b946fe19f126242178f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0648977e22f4590397ba7c1d0ca92e282aff04180f687a07f18046e8d3c55667c28f31420f59315f10770cf74747662be464db2b5e11d6818b44e25a04294451a9761fea4d012791c38535b160279390e612bb92;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc866b470e30715d86e20b1948092a6310f72b4249a7689ddb61e58a101ec3a94eaf1654a64e7f3851fbe4145ba769d1f244dcb1f03a35e2f60e7545c7c1048188912fdd98e2eec05117fa11371064ed732dac2481;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h993bfec491de1fa240813c0827f7d7a7b1ede286c8cb367f955fe6ad00c255e8546c2eec956bb27b3df3bc8f03c1d8fb5344d6f812b2f94c46536a7ac1079062d2c073e2fda622774bb7a08b9910aad41779991aa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb152f807ba7291f963c1a2a7896b11c7c23a805dc37aaf35ffa17dfb6d9224f3bbed5ebf9975478664d572b279c4c3de3f379fcc0342c9585ac10fa2dcdd898cbba1c50b9cf485b38cb59edce1e5ae55da2f99ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd88300e60a0468e2852c9308a57f3a62479a094857c90fd19117bd0cc6b8ffe872990d99003d9f9f3b23632ed1b2a432705ba25b8ee9383438609a4e498b08070be73043185df84c5eb66145413b9ae848c84d359;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f94ccc299efc693d7cd1c7d3988a9db11d86b01882cbae0015621d251064e8998f87e0a14a7063e9e0faa97496526ba9f1af6ef39bc35775abc87df53f38d8294ff0b87b41800f086016c555a500c4669f7753;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b14cf1c6433f5b31fea9d15e53e786625b4e4a3852e33433aa5dd918bdbc2a1c91f5e45c640f019a0ba0096a6b4f635fe49cf065047fbf2e298f6d45bce1c06c9116170f4c7f7880d4b00810cedd6d51fea88f73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haaf7ac78b2f4311ebb71bba698d14a1406036ea122f6402ab4e54469bfa98db1041922ca575a2762fde92eb8e8b83fdf14daad979fd561bb4727bb63e1410d4e42dcc07ca83cf1e0ab95dc3e05143737f818d0a91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1a9a20236fd89c9e57224b04c60bbe36a9b912d69078d15c415c0e5a61f99c551cfba3c13032986a3a0027d2103b8b179cc293dd88303008b2e42273f20d9da7cd4bebf1f4bb8d15b4af95af0591d2bdb3e79bda;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5594b71524322d89e1f6278eceb6cf58a491bc7382563b450f5a2cf1eaebbac21c51863602ec956fd9ab986ec5ffcee1c60313c04208c268c34bf6f14ff690cbbd9067ab4e2fdf8b14bcf03e4d29c5ec13f2fef74;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fea8f6f98ee4b190320386070248ed80b9045d548313798c2cc1c08e49c5fb7055b69efdd55a478eff1f672234ad7b02d05665bf230e94e224849889029bd6429692fb49df0fd8f7a554903a05861d7d43926f06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb35ad138c2f639e0f84280e182cd66019b7b172efb6cd39d181471b008d41ebad9a9d303fc824c2da44ec875fcbd6d20c92bbfa1c542e1d48ca30df0d1f80465fdc83aa781d9f792d2d58124cd531ec78e300a1b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9b5c4cf349d450e9d6a45d6a40d04d8d118d3b598e5791e7402775007ec594f56082629b83cd0cbc9ce0f6f378f90246deb86a03cec92cffcec4163c907bb9bf269d5de9a4feb17d2529c7665b4ebb72f5bc509;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he55b932af5322753222ce65dd243372cca285aad0aaefad0ba61189a6256ce0feb18b411ed6d7a88de80f71aa80141bdc5d03fa4f65d727b0a9c715a33c4318c6f6d1444dd513a29823666785b767e3d41ced9c90;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c32b6601a8066ee2130a12fc5968666829af8b76a901e09a246cf384b48606117927e3903672d3ec4762bd666fb7c87d5582fb552936de9c5e4ff3bb06389b00fdc93ca3a2b5f6539622fe67a096846a0b34130d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7b4a631849514174e14106c5c64100c9e1e2892c118ffd1982b0e8060be9269e0354d515d353686b6dab7a76af9244233c8c47faf27e07f6c0ca177503dea4a5d7465688aeccb3299c9d9b9763cadc32b38d2a04;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcb2d399809ae7ddd1449826aefcb39d2cefac967caf95f56b091b3c974e9a2151d91a38c715e362db313e64c6827b5cd94ecf523126b936a37d066993695b680e9fbed08aabf055815c9eb28e898c7a0f2900c42;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88e9f4eeebfbb04d017bc20e593ffe559d73259d352ed8e3b24864ab1e92a511e3e905e3a2a8a8e01ab6dbbac2cf354d36f1b7623a81ef51207825692d2ce1089193fe902235808cbb0f34eceb6adfb8eba9a97ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59e97278abaf54a2f167b5a2ea9bda6740fc4dbe598d545a32678a233e9e5d940285ccc3b340d152a448cf50f1c8c3eaea71867adf1f4552a0928e692bc8b476fb77677344bcaadc8efa1fa2bbf68f740ef9981b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb748fda653466cf50fab67771fb7e3e26f7d0f419f57e6123e78445ff71b3aa8554ad881be31a3473c83ef71dbfd0a2b3bd9982c69279887f3e1e9ee6bb0bd12fad6faef8d45f60dae7b043b302bdcbcb5972615;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61eeac02f37356a3949680a25abec445837d025a0e090e49801d80a055d5eaf2020523e88bbedea516b8033732b02e72ec11210790f5f9b17fb44edb4c3c6974405ce2d0f6db66eadc82caebeb9ae164008757270;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd58901e08d97e2fa453640ff3f163fd311fcf8fe3710336186d29870752d103b1dbce45eda423c6892b7fe1f0371a849ec562ea68b7211eddcc612c766f2e076f29d5d188cfc937a36b703cef9d5d3d7cf786ee7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89a8debdf98be3095b52be5e23da75ce46f9aacfacceae429eeb3661b7dd9e279f7275f8e2b16c4834d0445218882b69ef34b3633a7278b406ec0621af42616ac7085a0ccee20ae423e1d9b58bd91c1c506db27ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87aaac19b9a141964e3bf36588605e7408608a5826537697108f33d3c64282bfa22bff667884d068066ffe204b732845b903f4f0d7c2af3cc96cf6e3a9fd0751b8a1cd99ffd7d899ed9940877b61f872802aa30cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h474962afd801d3698ba0af3286996d516e58f8e62d72afd91d37941214b998357ff7a896e83332e04710b2bd3cc34dcdeb7a65b972148b2d3a7a9cc9f6ce7ebe352339a63ccaaeda6021f651780ea58c86aa8fdcb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h231fbb11c526bddd1e1942ceab394d0378b4f10c23fb4691ebb490254a72924681b4cb6a69730801aeadbfd2e632b69be59254f67b7e59e3003c57285538de07c913d6e771e70a12186c5d850876a4259934476c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb154f430c7c44144a8a2b31e5c7a86aae20708455d7539805efd2e1437d2cf10c734b2435bca24166811ced82bb5ce72fd91dc56b5cd7ed70282f1a61f6ef7d3db190bb29115397169c6598710748759e1e7dd2a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37a81f9552029b8e83c73707993c2ecbede89c9c3746945e3a70ceb59032de160e7a7368f8ff53da1c511f0a7deafddfdc054352b24d1a40b24ae1c25b48afe3238dfe2797c140652785ef6a962f03222065c1bc8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h224f3c6f685d08d24f865934e7a4bdc8d00995c9f1a499589d5723f6035158a53027363a61f14ccc6a2054b89d04fa3db6f873173ee0f465142d20732a4b2a39b463691ff3f07bf35c8f5a1de1785fab7fbadb8b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc19b968d2780391487851b27fb7d82f2ae3abef7ceff0db97124400a080b1cbe720f44870f3aa15a0c357891a485708599a6d5a5b04eaa7913da46add4346bc257e323dcac78d7643bbaa0d755f4c78319484980e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h353bf2775277ea3730f89ddd9b8c78a48f866b309fbf310f3b46ca7b80e392138f2a91a5f5598d17d985f460bd7308c2ebd04e252f6ec27561d5dabb3fc3b7305fa53a584ae0b75f86e66bb12baa4759490755953;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6f0c44fb6db427bc46de8707166eaa51224f44c3b25fd05091efe3fd7d857d4253a0618699182e06481e1c2eb24edf4427191706d55438edd49b6ebd0c57983111f061650975c870cfd02046f47f6c6b42c70545;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0b40cbfbf8ac568c82d551b032fe396a46a3dfb08e8c9af5be06bfb91293cfdc4ba2432b576ea341700b894faa7180c3680bc1d18bb5942e5950a0380eadcfc37ac607000bc0aaa7d9b982053355b89d8fd5b7e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa22ba2e087334ac980534a14c4f027214aca88098f3050c7d37ae7dafd336c32698d1e1b7a9c0c7003b897b3c56eb795ea13829431e0b49d7dc40b5a80e3dcf629ce6660ac75f583fbce0ab89941f2bbb82cc62e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ff59987fd6366b193cb64c3de0f12a8d7fab86d0391a42ba7f3c43085871d3bb844f7f25819b4914ad5a3a5c7778aa43699027ed2a7f9d1e910c01521bbd0ec6d2b46190575e99c99f8f28ca7ba557ab8284a458;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb097e0d92cb594cb707978f8878990144bed233576368cc1a71c5dd3dcfc280e2c473e901674ee1f7348c953dd64706569e054fa7e459b44ef72b3e1b8c36e3d0bd15c741a5bc16a8a0c9f72cc7e84fb83f9dc43d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heace783f6ed113299d72c1024f19478966074d809eec620e1f3dcf6b2e40b7b2861c15b61ec02ba8535cb7b18608aee7d096fe7d015338f9b1121fdb21f945bf747681e79306943316e81a2522882f930c3c7dda5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb07f719ec6c4f604ac163ff57b9a997be5946d0ce2692c1a56c7e79e1a72d918cfb97a3f88523614110d32c30975677c5904442078c43ed65d4791b4cbe4cc04e1c0edd8780e1ddfb76285db8d64dfa56294900e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88d046ee6e578b0f6c9a04a5496c25bc364d44a4b64dcb876e2d6814a4260957358a82d17c09b7afa7fbaa3710b55ab7671ca7a74dbbac9a33c7ed1c22b6f5e1326cfb62e0b62acd4c1c6b66b03fc9f060216f344;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb89b96351736635b75cb8c938ef73f55e49a353956096031333d1c6758a625d3afd02fb845bf9483df188fe3a89bb2ec654a189da3d6f551ba34002f22ad883044084e9dd5df422afcee2d6854fe6cb42a73eefda;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ad2c760898e09b5f24140303f06523cb5747c3acbd5b772ee334e9780b4b70706ba525bb1c0a9353d91e82d757b16e42443acb04f73bfb5ce1aabdea0b391fc2845df10cc379759ba8dc23ff9a43d1230e611f89;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heec4716251ce39511440e1809ebfbe8d0e2a36aebcef5d593f970c2d71febbc2248cc17d6c30069d3e873068289b1c1b359cd6c10a1b9dce169e44baaaf15e440e379e7744fe212c889f042ac1dbac5e0026757e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60e91a9ffdda3ae22d9e801753c41dd8bdf6641d53f7e8b0261fd95f61c850c78286765d261bb6354dd3d1f7b25a7a6260fc87c2c4247586386650119efd15405e9767d0512d34b9f5a42083dd4578acfcf2f789e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc73c3c87211f96fb55bd2423c2c9357cccbf5fee079fcc004885efdd6577ff7b7a81b645e48762cf465d3a6c052938aeb0b5fe529f5d4f7e586cf273db602ae61d4564d9c8f3709e512e877fbe0f7a2b47a1dd94e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7baac3b2edecfa888d385cae6f367719d33fdeee5ee1a309910fe60d066293b3bd37d6966bafbd7011d0ba5812c49ba2fe23f9a5de3e9655306c52c0e5f388e9e874fc3ebc5b97268af3b9901ab2fac94786afc64;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b785d4486b78f64ea01973841c9a34fac90c850f7d94325ea886ba08a4d0695597d931966a73bfd92f750e3c7d47be144accb56a2d0beff7f5083cd939b334639091c35487ca333d60f43efb80a649856e3e53bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h884fed67fd44553c33a1996fcc9ee21b199d43cc8177bc0ddd0b27f365fc87a6599956d724485984736e415960c640690f08fde5e0cb1a3ad6dba8b11b0abc53a1293f46ba325d674d05cea8c9d89625b7373623c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd18ed24a63b898edc323a67f0cffab6c183143918c297680642ae5c954e7f4854fde8700c1108029aa52cdf40df2d53725a9e7a548ed33844afdfa13071557c8533630be19bf989612e953722515d4a79543c68a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25dc9e814d2a5c55e03986777c943f1c3cdc1eed889f050e39bb42b2d28df0862c3fc45a00bc8822aef316b61b77d1997ff38a7e84f1205c3dafcb9001daba72bd77c9888c1f560dbeb8a86233f19af6fe9735aa2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h787b3cb1d0b7c436147e79d543abd30aa5a14bad249f9d8766debd47f05f4f96a57bef991bf69eda9199bde0a99203e88c9819b9e8aea51a9c28385dadff0ada33a456f10b2151dc5e45835af2e5192ddefdefef2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ad84cf51ef1b97e37ca2872c93896633dcf0945440ec68a26299998cc8e38878b4b2872272002836b8d2f72faf739743e8eb661fdceb54fb28164840d549fd09cb898db961b4e87d99712239227839d2c3a24d5c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3fc15fb078b71ac03460d9967d1465a82115b9a793077892ca7708cbf476c01d955a803ba1445bacfe5ccddd2144a7bf0757c65ee702fc14112271e8e5394131a9d41291002964ab5901d03a30bba355cf0fb134e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bd369392d42eaf2d8e16892a61e9912169b8a52c39171370e55eea9548bbed68eb949e172af0d7a7b84b3743e827c6f1f0f57777624b80156fb221ffd3460636a2754aa8a1eefb3638582365944c8fed1c969b8e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h843021c9f17aa3ad3a89ecf47ffb84d8cbd52015e98412b1d3dfc21f3f18f5766e92c4ee859ba7e5fea950a7dbfa954bbf4205648b807b0492ba7561912862f9fd266fa61a16eae47a7c9c65c031328983994f206;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9b8601f67251b50ac51864f9d08728aae8d208f56ee652a1b5760988338e58cba55476e2e0fc74499bd5ca9305f0e277cee064b48194bbb73719dac637e907b22a32dbf5a779830429cb4ac1fc20b7af62f6b20e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1ab16f6abcb5dd33054f6801d4174668de93fb33c1f1214ecf24525a7e515d67c0f0b0ac7a0fb3cf3da0edca219ba5726733e2d5076fbbdff427333afe8fbb87e09399d0824e9cc860cd284371d9b4409331ddad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1b68a1da31cf224e67a80a60b7d7fdfa848bc55e3e66fde1c2a60e6326c73ffd78b2a57672967678436aeb4e91c1aee3fd4d4e0e371e4473c9ade0262320376274da504707f808b69f1250cb49f6fdbd57784299;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8575d5ae1bd36f721956ba0c4a07a8cd5d9ec550cc526b41e088c605dcf0cd5d2d82bf447e0b0f1ce9d4df34c183b47686c2bad26aaa84369bbf6670d3c97238e0741682f476a5e317e8a0d6a875127af97a0d1b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb55f3ff416cd41fb972b4c0cf47e3314f05140ce8a3143c883e23a9d5ac6db061a2134d67057659d5821bf325e077f7a449a853922112efffae527d97aaf478abfddc7f30684d264714b3e249b08acd8eec6579b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdabd326e62fa3aa20df3ca64115b1583a87b7d8230be2ceba54e96df34830376c220e22995413fb9834dca7d6cd92d4eabd005d3cda4c711bcc6916988247189dfe249c95c9334b47728cd25bc7332962d185babd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h511b3446b35375f0608104e14c74ad05bf149f712bf2021674f4e226116c922a9e3740edf91ea9af0bb948b0fdf23acdac6a1dd44850639dd9716241ccb8e4fd5981d9d6c0131222fdb40578c6d4e656dc624438b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e85f62cd93e3ab11fe2e27fac6f30caa7f62a90d7411dba63d4bdc51b9f9558632af19fad7b1ef277a7efd186f8d4709bc1dba2770a5a2e45f146309de3ce3f3110a34e0aef618005fb26563b8b2a18762417dea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'habbb7aed44c35cb0f24b40c490d2473be9e8a71b843d72e1a23fe3b2bfa683983a41ac96e5ef4a72cc6eb4e5a3541f995aa3ae10a88c1e83b1c7052fcdd440b8bc2ea060706d63a58d8793ad524fc8794d8262ba9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haca9650a0a749cc0d242aaa167fc8c574e16ee45a01707f1de35ccb58506ab44da24b13297501807a6ea625fe0f659381c19ad535fae5440cb20a0bf37f8220949be305a302f926d3e71e95b2bfc64ad204fdcc66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62b2b3d8b85af148123e9faf6efc403b49afd79268ba3eb910cf8a94b28a28f9c4b94518be3c6bd03d998d29001491e0c72dfb83fb30c4c5cfce7d50ca102668033a2dc37f353cbf9f42000fa321bca4e79089482;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa15dbe9f7bfda92455c3da3be4ffaabac9ed5fa6f5adb3ae51fccdcef18f3127c18b7b82d8fe1988f66c189b42c82c312cc2220e6e351dbe7b584c04abe7a3fedfbf72bf41e57e77f224d2af43a2e44651b83354;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb07ffdb4c73870105801315f8920f2da42618e79a2ab7fdca29b896cd76fb42f73a4121888595169f765a1fd69485724d94a46107021822640ff344d4da5621978e5d77ac549b01d6bb7a855adbc3e928cbc69491;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8753f384280c7a24260dd931d0d7a930d5ad9f33690cc5078f05dcf7537ccf3935cb2bed212c8f3ba6fab14a3e0f74d2673380abfa19b6c5fdf9a413b8e387275c26cb451276112b9262128386a1519f65381e2bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd09a9cacdc0276ffad132fb9980a992e50890d4bfcea54f3625f1afcbcccfbf9b0564f53f21a053802abf93663ce3f23c1845baa9fc4776b8e74c6f3c67363af6a5dd9573634d7aa8c812193f96dcafc4533a4aad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6db8a2f8437b22203814277886f099b94b81d44563afa48d7e4289cb1e1654a371534ae19be98231c766472f826cee63591113561b91b38bd010247c8189b4c8c51e04d2c1357ea0fb53e755d6aecd28b5c6df603;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53df0c08c638de35b51f50309b0963333e3f4c41ab10a24f83b5babcf5a5f56662361f566ce912ac123cd78450120802210bfd84c70ef2601ac4aeb372b31c7bf1e20e8114575c0eeeb0c9c08a6a78321b3e0e68f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cd3784a514da2aca48866841ef4c4d6b427ab846c544768f48f8a4b66259498f9d472ed909f62930dc92986c787a6dc3a1a564c94607a403e504419b3ef2791a7bf03be0a9bb16b11e364d97ce934d6117067932;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98d3404d8475565c917b2732d46427247841874e2e31321b385c9d13c449d64185d7b3d72f4ef9a7724a6fe975bd9ea56cb0d83853314770327825f7001fbf1a8a75dfe0242cc8f96a1808c6597189857bc09d9d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdbe8bea0f34b934121531db6198054f0bc351683745a5c47af9671a4d1dca8051b97ddfede9c1ce9685e552029399064ffc5ed8bc1c0c12e5a16a98b06e0af6f9b592bd4badab4b0a5db594f8511abcfbdf0141;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97f79e35d11afbbee2cdb1afe234b3ee72ec314aca6355e75baa63fe168c303e4de4ecedf9346e51a7d986d2d5e6e603daf1b0fe1095c654c8b96a034d279ca4a7958c0c43423d5f800a09d7ad59db1a5689d92c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15d020bd1df0c90b737cf2e9dfb75a5f49ec71d3e66c6b0389b8505062e6ef8fb51baa4b0de889929ac3eedc2c450d4f0e82ac0c31f1e314688fd2e258d5234757a2b211ef0f7709440546100bc8f26de324ee26c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7f5de5ae53214ed072aca2ccdf0bbe82bbe81b6d750df3c978dd8632b382139ded7058ea70b3f07eea0841150b2a940140126e0351e244fc25d3f30c26d0f2e3cab26d5532b07c5c98968d85892565405f9ca75b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d84f3c52c53f08356a1fd1ac7da922ec74bf5a4b9922de156fe9620460062a65b5917d110f17f8d2df2e3a3d9d4cdae411cd0b2c803518143ad1efe384b4a895142943c879d87670579d7997370e893b54298590;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85469b34e4d2ad40af74ebc124d9f4313889a0dbb40f693eb113b9882d023187e9d75f7a95084944851ec541cea14c07875eb5120af4c6ea1fb4a1421bfd7628cbb53a0c1f0add7517d8e2e1707ec707b7901605b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72900792a0520b6b941c171c0be0c967dac59802a6d3438eabae17e942ca5262a8a85036ede63efcec6a24c2737d339e8aead01786bdb5ab58bd50bf96bb8f98c2a1669d5650794600dee900e11ec1903b220b088;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d2f16541cf5e71d380898c81f6e8ba2ca61ea5703709f39881b16a155983fb6b853393a4568a5b6a7267393426d65eb5fc6299580ba3dca21ba95d52a2d7d8566db6b4ba356442148e7dec44fcb2d2db5e39a0b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9500b683da38500b0f53fabd04e1c4b273b67701a45a5e66e2e19dc87ce900bc470a8750d47752a22e44e4b957198ea4e25b6d7fe3d52c017011760755e4e8a03c5cbb2432b46643da47f118dd75249c1574d3b71;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dd11ca46b602633e4727f30a1abc5ff220a1ec1ea0740d80922a1f4d9b0e1b4476123006fc3a24ccb1583ba14ac7d437194dd433a8f63b9171bbbc813d2c36c349c9df915763109eb37b8361e449bd07fb10d395;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe489cbd0070051d15f077b13c280a73debc8eb0e6cf3d291e3018ee5a02f011ca7ccda58f7599c45d16dd222a7e65ceb60ec3d9eeb0e5b5a8fd4e4085698379e55b48525d59d3b46601b7b04e487e8221fb13699;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ac0042c78ff9969a997c62655abdec1413db5246978c9dd18189ed089909e9ea0b7f3544ef96ec3a1770418d116b7ca2627f54b1965d34975e7cc677d4067b25e0d6a56028f2c4809cbdc9650e6da0afc582b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5a7ccf577a17458ba74ec9aeef360ac45fd422a62d1847dc0569228aa7a3e13f283cb720380f143236212d2004948dae470887dc5da3b26d794d47d983c41932e2369bc05bb26c4510791ddaa66a83404f511efd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8c055baee48f09e73b564193631f4932186ef94756812ddfbf626c13286806017655f1df63685f0f379e7eb51485e1a5f0c9e0a8d2dfec29fae1ba18050a71cfb37f60b984f543934beae99546db6de2d8952cdd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d8996ed9526a8acaf2acd155f9879bd542c4cac65bc5ef97ce655f2dfc51bb5dc91781fea7f4bcb6b4c7e4ad0520f062e92c5bff5ca8bc7af05137186b135e2157ff1bde8cae5257db09a6c5fe7b2ed051178d84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h682b5a6cf6a48814fd026b21dde644dbac1e06a07259efc24eb7e3a99958a8f97a6ea6da8a2554043aec71ca43dd3050ae4e0fd4f5b181abb3df690148a49ba0d98465f67fb2d0f243c19924d6bbcb8d8b203131;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7deb9f0adfb8d4ad9cb1004bc8a638eb13c06fede709ac5ba97da3bafe0ba69d2704c154e198a5b785c85a30926ce6099fb633150982778b02e398870fde80339dfc0f63df66f52bac09338fb0e69b5d5a280c9d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7433fda0e1a0a27bb4e465e4f7020ffb688e5adab47ef0ec62642e0f610b787a6b5fc99d7f012f4aa767894acf21f8348687f7f045740f6d3384cafb1e9384dda91c253b290df8e8a0ed0b052cf2f58b81a58cdc1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6523efbf81eefe732210e01c98d4b5dc63684e95154429d6bd9eec94aa4d0a7d2fed3a46c0bcd1fc33c8fa378c2ba8b2bf395e10b74f85b59cfa661155e16c979d5beba06f49c431b312c242217d048bc8864255f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f3f333f2a1f3f45bc16fc07cbd3a8295aa4cf6ce8d489e775e42e25914728f5bf1120fb22b41fc1e07d012a19bd96b93f4b7d3a2064e7b2ec289d9956009384d8b6a8213fdefe64f9e41ab716bd0cde12a6fb0a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4210d2f3254a8fc0fe86650b378f2f2f580a25a7697dcb6c3c63d55a7a74ccf8ca8447e437704de2d1b421033d917431ec6c025c9f4b3d4abe67446062e7b34dae960d24128a95a45a79d45f24ee1e378e1c64a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ff03593e33864482914571f38bd09e4eaccb13ba1d300aef9d8cf9d62923e9faea96d8914e3254dbe59af21c39ae52db97496fff6ec75dcbc2ed12d95af848f61e55b64f59d9fcd51045002f37d2bf4ac7515d4f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc18c61d4af0a241b30ff0ea6803d76fc469681ccd57b69cf585606c02b716ae9a720adda261a5912ac4e2ed1dcace88443fee87de91aef9da47c8d53544a46f6e4b94b6bae68bc6ed247d8bd7c112b51cdc04dacf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9395cc8fde429357f5fd6d0df21587e86408d6c6d6ae9b7f179f3ef58dc8e0d383a80fb647f9cc75cffdef01d3822dd223abd7c2bf64e629db1d2fb8b0f98f5e16ed12d55dba116aac46e5b4b91949b141204d660;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h517aec015b71847a8dc5dc53dbbda1de3a6dc66f2de1bb100f0db628d6f336a8a089e2fbb72f5eb8353f8469f708c0619234beeb34085cbd542ca4877c2155f553c9aaf2af417bb012508512301ccf680e05724cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfce90d2072d7da2a53c66cd0e05a5c7b800eedfffde4afa6962e1517606ecb8ea0f50877e85d42a5e703fc0b745c51eb329ffbb60278e4ecde94ba0a2db207c3b0ae91d3e6b5fc2a2c338e4f8954e8a17fae17ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h845aa7845a3fd1fda2582025d8a000e517dbe9d0c54e537a8372fdc84b8b92cd357ffb2d712e31a2930c5b64cc865d9aaa3a2f4020a4a1a919e3e28a1f620cef33d2611f7540a123e0715fec49aa0004eb0ed2e66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffbf1f334a518514fea8609e4430d5a5718def01a3f18a40042a2d7f325ca12ceaf638452c623f9dc513a1c479415c36e71ad4ee226b0b1debd19f2126bada205fe5cf6f28794f234250b4de3b5c27f1ccb4915a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7fe1a554412e4128fb10593b5db40a93469fbe981d214741077428862304b6081aa90b0582bff2a1f28b1679045f2fa107d95460f778c387b97ab363740abfca31f56678d76e1b76d4c40b517d1b938bb230dc77;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ed4f677784e7ed9cbca533a1a2fd4d8590088c3aa4c910a3c4d7016b8f842690b55be4d447f446415f0f7dd89f8b02f4d35e83f03a1ed8f4aff289da98567e84f60ca18e4cb3670f92e48781b1f49840183fa304;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8c9b8d8a216ee719d533cab7f45e660c99caceea48e248ba9b0b02e32030ce3ffdbaaf0b366482542e039d0f48ff35451d6c226bdde50325d26f72c9df03d181d02ea9cc60c947e57c218b776e455e33ad37eabf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bf722d40cbc97882a1a087a540e14a238a7fbd1d85ec03e906b34e2ee96d7516702a6ab5e8af58d094c8eada24bd5eb286ead814b5f83b028b1eecfa6ffc8c4b8b01cf5c2c3b8cefff6f41acd84f60f7c7ca8451;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48e593cf5ee42870d005e18fecd7e656e5e2f33864ace64eb29e0c43fe3593cb03dc8d914895fdd3f8926ad7ed0eed46ba8d6a832fee11edebaab646b6f1b94004defde823bf62e12348f45326ce25c8213bcd6d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67fc8acdfe1651871a953a3931714e2f63f65b11e36373d52fab2a9188e77ce434e5471070d9c2b8b4392ed7a1b86b365526d2fbf17755f2a5d90153a72d3601f2aa34951d44e833f8978e8c4620139989a298418;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21a26c0e85d9c2fc9aa1ec32e4d7970fbf6a07706b3287df0e1a6e9fa8ce5f4e7733f2cc63921ecbed1be4a5d143341aa446fed665c38949570d0a24f4d0b8dd8a0d43a1a7b8deda2128ddf7b4bbe8a889e41817f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7732d318de1461590b11ffa8707d655d1084d38e1e6dc289b1495626c9e09f5691143ef0ca47c567916f6bc03ccabaf49b4604a8f6176cc82037984ea78d92f30b05176fa11ab3ddcbe7b15f3e377b06afb264eea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb14d57bf13888ee4979d9216d629afb9cba2ad219432f67613e1831f8b3882c0f4713d7bdcd867e7a1b66d2703c028fada7d3860a95fa0ac8207d69867f68457c669196401b24ce7d6772acdcf3bf62e36269fe4d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc36eea0946f4608dc8c5e1a044dd7c858491552c479fbd66b42767ec44e376e1b1a3983c679544cfec8115f3a9cbef9a7351754eee44bbd97a0f357f775cb1c94075c52756e9a93e598323ee8c24d3d19ac8ee825;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2fd92ce3f40785f42acc311f734e1847ad5f4c9628bf97040b3bc143954dc5ebef1ad364cd061c20276fd86b60077d1a61604b56a27eee0ac8bd59949dd03a2e5ac376cae9499ee34beeec223b2092a69cabd1cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h427f0f5e987480b50b70954de1a3f24c03b7995a1d388a53a253c294327b0a37e94a0903fc8fc8711c44fac2011538c0fa00fd15a615b76ffcc712bfaba654a9d638c5902ed4f77ab75eec6bc00d08bf075a2e966;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h393e9a9c5092beea2f25e3a55fc080c7a28868d1b5ed71b113ad05bfcf2dfb34e8a06fe96f74c391da34dfcf1d2fb2aaca15d8efeae9dd4a9d733a5e1e1e7773a33a966aa8e38775e6ea131cb41f9dd18aac97cc4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7673432e5afe6954932ab365c88af29b057354799ac1c061198a1490721ef5611027ceb47d9904e76c7a8ab5f3e0552c4c14535d500625d69e170dafa91debe291dbaca8b5a606682a798ddd18c3efedf446bf6fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h470f180ef2adb82124551d7476aacfb35246e30af7ac0e7bb7b92c8daf436c7ca0d8389f2abfd87c4d6a4b3835ed23d7492098534e6026b39bc14cf6aec8a5ea0746f031c2ee91c63f27263cee7cd18ffeefca275;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1980534feaeeb015cb3739cfc968c7ae02f27b1b1d8efd69c8df6152179900befb55c678f3519415039799fc5ddb43bfd6cf4ca28b5b3b4a19b4b7a553b0616e259484c54d496491a2e2c45a994385d3588bc25a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcb91a3a9fde38f61469bb6dc5a08f104746a8f426d33a5f66bdbf3b35464ae2ec6df2e23fbda3f8f8eb4f1835ceb700dbb8d1a08cc15001370957f87cb1bd80ee5e405c10205f29e6cc273c4e0fc0f33b023d442;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h363fb94de30e8aaa2d67256efb7646a25afe2d8d969127421633f55d1ebbcb72e3cd85e25ee188d16f394d666ffa56cc53a5044a66d0c7b1a2455b8f3fc8022850f451442e16fd7d20949fc004ddd3b33c5309d2c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b4d35f3c11c9a62ddc612edd08bc108c4d3349f20e2820d7b48764169dcfb366d1b4f7f42ad2f29a5b1e7d5f1c4730edbd23085f4cf046453dc2abbc08cfb15c182d81832daa159e605b5078cd9abf24e069bfd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf08b1ac8cea19a8d6e32914d2b9dfc4fc50fcde5ba200903b825091addbc413a33132611ff3164843ea565626ef5bf592d6935650484be88d1c657a34269fe197eb810b512d5a30fff73a9d8db49c651fcc9a07d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ad542e2c3781e7719ccbdeed66c7936b2f61c09d92c1c2c666a1144e668bb15ad3458e65a2cc2e661f2f58e39887386a387c3bceb34ea37fe9fc8bedd58cd307488904ff232cfea4ae8e8702c7065283c66f0b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h122fc523f0a3c915b2c22220f493279ec912a4934f326b227944da23041b2de3cdc28324379e09f0f6512d5310bc46118401cd25eef5ccb6472da07e1ea27580c5896b9a0b7819d874dd26eee4a9aae1733c42d72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6510d26238b11763862d8732912b2b7f4a90f17f48874bd797e2d278e2fc40f69ce2f5e3e7e027f5230c523a9c26239f280470cb18c3dbe3daabb525f50d3418ac8029f709542b5b0979b48d22a58572d2b6a5af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46be8668e16c6f40cde75e73eedaf35fed602905da48ac0527bf5d4420953a9e1c632206335995b4bd04d2ac17e7890f3f8a1dff75bfc7f0796e7c0dda7b536994c5696db80996e813a12c4d94d518ddb85fbfbd9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6931e23b29a9546653a06927c2054965f8443878167b7cd9ef5aad9385493edb56cc0f1f09d154fe3b4fea669183672f5e0ae40955f0aee2cdc713a906b19fe660e1f80039ea63204b81a347112d83da92eade00;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h629b222590a840677be04aa44094b1d87167fe95060dc25e060775b6ea465fb2b9acde57a007b5b51caa6437280f7c2ab7a893e7783bb370e0764c7b165248fd451632e82990e3c41ae7e40782d7e0d02ee89b790;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16baa2439877ed5284c60e96710e46b2815c45679e59d5849f8a9f78fb8cd71b271f484feba76f0ef80cc64e691baeca81c8d3ed61f6afd01b53948c2bba66f29ece1f9e6b180d27997be39a52ba07cd27baec317;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16a7a131e405828cf4768c989cb4a1f3bf0ee1d09cfa5c1cf30dc6ef08f77c0e89fb148fc347e77789ec2418b0b5d882731416020339ee6622d8e893b963650417f3747230a155eb6eb8ce48f8698d45a18a86f17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he23589a5ef089a700670488a73f78d74fb4944db6fbfdc219099868558ea63abf972e02104c49734fd47fa75fbb50f4a697215c3a1a369b5cabe46ae1455854734af0eb7b19218c36a07a5285d5ccb39e24c0b963;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81a52abcc6d2452c57a4020560ef472f6ce8feeb2d9527199e8b0d5b65730520425c03ca61521f1897dfaf5396cdeb233c672ec8627f7edea0255105298cea9d892a2c557e21048d1448e71816da93b9cdc7f6e72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb6fd6315aea46167d0081b8a983dbf613031769d6de957d8967fa96522fcaa3c41c70c7213d5861ec632d321f8561fc58a6a1c4e0132ce725be7af6269e4711ab9c43610e2d32c8942d0ca2dcdbd045466281913;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1127e189f8c9de66dfe98844b18098d839b797651fd3a3d538ed4cdfc7c1ea2b0f4bd7af415876a549e6a80f94f2c5b0425c08d1793467586196216e22b47519f4d58afbb6b4731fb1b22778a5a2b203a71c544b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacbfe2e163beb3b6f08f977e035326bd996653b17312f54bc157f0d393f86d2e20e856beaa7a74e25cf99c2dc8460928b3c1570f2a506331437e3cafcd80f14dd47c077e7f36c86dd2581b082385bacec7fe6afb2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32de8069b4f4f468e1e08373b967075673143f2dbf862df53a92f0b5f911e330495b76691af4bc4e1441f08aeae6e1714be43377e481cd7b3b134714ffef2cef6d7181c7d28edb4f61a9acfe6cfaed3033c41b415;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d2c9d16e708cd8b94b69fd1ad85b59b3de7dd0d4d01ce5085e48dc463ebb189f19c95bfa7627f94bc6a81c228fd8bffee4d7e063dc93b7b202ca607e35d4c5b89940b0b4e5f392a953707a0c355a07a5e353c60b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a074d419686102400e301f2dc35cc2003fe00bd1d887cd66d571748646595d96265789d44da30dbabad1ad4c392ba8e2632c11e914b48c926fccc314d87148eea2af991d4866f110ecca60b35c26ca6eff5cc77c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa67badbf19e87fe582ae7e6b72fd5630671d50551e0cf300fbe20bcaf5268cfd2932177c4af3e903e93dfd9ec354bbde9d448285875ae3c224c4a3c09336daea53cc739da7ad37b046a20e33eb92d21293ba2bd5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he753abf2dd85179024af96f14ee6be7621364aa3f3b170f69f315ced9a3029f7d41428661f72498dd9b7d3dd5e181053afa5d29877613916af12e1834be0d4ccbbc4c11d371bd6fd0a96305edf5d6f1b47a50572b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc35d124dc9e694fcd3d3a12c30485b9aee489b45e003103bcf718afe455bec737e430a9166343708adb3766a6a928a837bfaa0c0746f5491f14f740c2c55c53ebc0fe48a76a9c2123fd58b2ca733d9b939d4a764a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e01f62f1694cec62bff6830f13e5e668dea7d584176ea55a74090eb89f084c3663a6756fbc9db7f248fdebe74fb4ffe8192bb618b1bc84d593851ee9d5462750211aab2cb3b47ca7ad336fd6e9d86533270985bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfeb51c3ac942e02469d3e1fb935c303c64780a820d2d75f8d1bd065f93047423bef086c96d0a420f76813272efd9a8394c0197d1f9cac4bb631c20ea7dc48488712f9f9fe3f169da865809e29918dc3b989140665;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d281c8d4fe2cc3d81aefcb82c3a8796e7f2684524da185fcfbbf871d769bf0a9421327ea13603e89fc5df27ddaacc38150b853df35ef2fb13287a987252e8614d45ffa854fec86812fc0fec752afd72a091af8c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cace20eb065e0f6e6b7a940de7c877021776aac683e87d7866f2af7f87c8d958623a0b48484e25388e642bc1976a4d9aa028ceed267dbe5c1085cb4dd7a90c7d35d7f811aa3e21274bc17ee4cc6bc57ff8238544;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f394ae0c6cb07be0f2080a4e9a71c911f4051229fb9834c9a8210b688d8ac289f268bcdcb6a1237f773f0fb278e74f942b2f4085dd18452d9908c99b41b537430bf4fcdf4e796ec17063e5a01c961b5fc7dec00b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc30c86eb2ecc76162480fecbca032f0d2a3918204de7088d6809b87a97a0bf3c850a80614cfa4117b5a108dc38cd89e4d2aa772c6067570fe2a7ece0c1f6cc15aef5d0d42fd2bbd9d14ccabfaa58f446d526c3302;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3317a0bf71da2554f16ec5c6bb42141d16dfbf31c96927449b3c33c373680d14d2f6b88382ee89e2027a84828d47c841b6b3098b1ac65f87e785f3e923c7ed2076bd17f4157dfebac82733c9f97f944b6719660ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf05a35878b056ceabd0bb6aec018897ee13717f4b76fc1610275e5a8929bb052f0d5e45af27c8cba87b8bc849c7b417c227d136bf98ada0e02cadb197b7bc46d989a4f45f3d393d5d7e7288ac9a686ce265205a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15471fd36a5938e50eb8b95d59c67a7cf0608936deb5aee97d92e86805c7f607bdd811e4500e49d6bf785be48e65fd35e037df07629e05acd1ef34263821ed8ccd4655808f9923547de55921af75d923242f495d4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he996757eb19f1a734c20888c5e528353abd4dab349b7fc9657c0b3144223b7aaf026ffd8060bed17b2078fe49fdc4c5c7312b2cc0303d5db873b2bdb0110412650caf8677d31ae69fadadc668acce70e10ff7efe8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84715c20fc27e31b72a76ef2f1321fb6b6c3ae40ab68a9af9dc6894247c3e51e2fc16ca22177d9bbceeca0db9a85f2f7ecb4527123f63800c8d81f94877231311a6d5bc587a0a2c5c543b7ce248a42de303b6524c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7de183bf8114ec8ec1d69e0ff8f369fd59d9eeecc15332ac949706d69519e0e9fd36043d4eb2208b0704005c94472a2e8925a89dd4787d2707621a30e9c23e62ccffcdd32b0406b7f4640ca75cc3f1fccc2e4331;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7b123ba88517a7e74a2b202873f56f754966b31e250e3d08aebaf8cf2caace16965cb2f240a8a2454196b201ba937d56233afd0e61030184a3df61190f250478788b5a0246f21ad1ee50f32330dfada9c06e8438;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc63299648d9876516f36c1d24ab09b1cbe3251c6a1904a3b641c23849b8f4f1827719156393ede74ccb2921210c0fbd70b8062122e24e11a8f6f3bef8d605424623be07479b0fb309968b01861a266285bc3fb3a8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47ce66880014efec8ea7d15c9e8b33a08abea16cbb71e0a5afe0056d8f13f3abd7adb6c6d05a6702bdd5f646206aea2d7ad2367fa72cb7d079f1c1cd4c24d0bf800a000dc06db506db2d0cf5f804c15d7bfb8c00e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb275f6cfd6a79ca847c880becc483a028181f16646e9ea014f042250af815f74485b2982ac2a525419246f087e6ca6cbc6d0f3768f612093d18f3e95aaac4af9cb014940eae40556d0bfc9830750b4ea447a1195f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha67c98a658dff5ecc6eb2abe39ab1764697924db4e501bba6f43d5831169831c05695e0525b1ab4e61d1ddcbc83a1a0fb05f11857686ea1f7c6de5ed4d377d543d0e703c511901a9446073a2ae2f428840e895db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h185fcc9b20f2de17efe369166ece2fedbef4e27eafd3db7d9d230f8a3526d83b3c46dea0e2c56e5ddf8e59e05335c293e11df15f42869e0b128b79a4ea2a34946cb64e986fce3511e43d47069b6567d818a2cff7b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha369cd66880c4f622874e2fa9a3bd8684a7422ecceeceb0e033a125bf12c3f77193bedef0837cc21a92bb997c8f52b08e130bd1314988cc181a0c5a38da6c6f2c2aa0cbdbdf82071046803b474deade4adfec3596;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b9d286edcf38ded083f2d131a412f141a97dfa562252337bf2e9bad5efdd808af8e4d3bf219646ad4e63421ac11f9ea2166e6f4d0e7467610f22f43467b74ab443098a312cc6406a8674f557ecd5f712e6ccb903;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c7667bdef9983a861996571f4917a769f59ac32bcbec616e5eeab3b9bf4c29872a9b6ac276ee293c59a626f523d460d500da14b9e5f824f37439025629a85a23107870ff474137fc860d4ee895a3909c811947be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62d9ccf2c526564534ffa98adf3307e2e7642bbaa8d59663dd75255448e204859bd4d708624a60c8d72e876826e27d96f6bb6c565dab21abd20ba7bf1cbaffc15b875300edd88cb2a460f03a5f8181c827d08a148;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56305fc852d74d4d76a6714d1ba96b2fa3fd9dd2b9147b0258e1b095c56c33613049ad681cd78a342debb8d238ab80516e1dd4a2d35a1525d2e174dce9f3de013c47e45f9587eeeeed8ffcfeeff626c29fd0bb3b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9ce7b17553e5e214276e649d21c1ea957bdfd2b4d887267a9009f574727acfad3da58ff008739695ef9d4022d573d17a722d6a8172152527d31095e383b8d9630f1fadd2ad71a261f034a001299cfb2ea467aeaa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h600b6cd27568da990d4fa8143a6b454ddb702cda2b7606f65486817b9d8b35b4ef9793338b3871a2e9c451f05fbd8a7bfa6928ff57c3fef52d88a24a6cc9e0f2f80a3bf09f74efdffbcd631112c212bc78295ef10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb277c1b617eea3859db53152b71b269f0b6b900ef08f27c46b4160fed85c191272000aac5184267f572eca4188bb80b3428bca33c57277b45af4f2204a8d6e634c7fabeca38db4cde7172ef1aea200522abc7f54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e1fdf8b99fc7ecd555b9b5d007472e672f44f621f53312ae481fe303b12eff29531d09f9b31e21ebbada1c0cd24053e907f0e11e83cbaa659a16c0ccf4333b2756b88c93f161737b934af3a6c4ab24accdc29ac1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf92bc11c7ec9fc9cf024275ba3db17e473cfcc2039ce440eb4563e0724418f3d974fe5a59228eaabb44581f2681ec5acb1dfc64e840fcfd59f62b06e05c270ce1252ada6c7affde514b6e7ed0ba7f8521644ce104;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89792d9498db2910751c93545c8ff01c85849f2043dafa6c87d2fdb0b818b897bf5060b5423c20cf5ca0412039643d0075d26534fdfa0c28a7b7dbc3156064d69cfcd40fce2deb3a5580a0c751c8d75973c1c0387;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7459efe7bd807248c8f7a8030b1375c0c3de636bb3fa626a087cc376d0806bb156aa46a31d644a82e060e7e80cafcf59e6acc688951ad11bad85d0a36c6e7ec43b829e67fe214315ba21313a56a9df7877047f3e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd89731f4af134b5e8ab054f4085b46f17a4a102888e92da4495ec4f66a216451fcc18139ab7c3c32eebfb3722ca4e429dcdba7903b05e1308e6bc10d62025504c8db9cb3f9d1d1dea8496e7b8ac059dd0cf3d89cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h954f13f342b150885af37c49323674a9b1057a91c6ad493e4d7260682c86c352db18b83266fe3c6a6e0a32b33c38a331b45f4e5f3b47e2d53523d0069799756bdcb39b0198015aa22d707b1cc8e8cf31840b50a04;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ef7d13c0491f3e9af484eb323ea9fad9f7b11886a09d1466aedbb72fb5fbbc0cac93140c8d2a0d9f4bac18b9701dc9d901d93233d7058e27f709ffc9efb4c23b34a9c17d0204787e24356c338e9d5dc782036faa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7440b29bc52574b81b26be8e445189c75692bab9e6a96f71c5ee1d186cf10aa1ed725c6c451341493283b2b259f618f3c5e80e64fe25ae4efcdeafa3279a81eb1b6d5cbfcffbbf3d0525e56853c571301e46fdbd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64ebbda49a26c57d11327ae2066e1d5a9431e9e5cf6cb62a0386332fce738b2f4aea64e196e29bbac07203c589eb21b9377abf9313bb47d3435fa6fe7ac7490432ad95339d2524f303af753a2218301b092f7b8f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b587348d5b4485cc9daeb01061d74b0753da1aeb0d344c0d292bafa689740b8de00861717926532ad914e07b5a09df65a0af0f4a47d0f31aa8242b817f20b9272890dbcf5d3702d23eeab5e233bfc08aa2ab61bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95133feac67a23255698f7631e15fab0faef22d312fbef478bfd63c1670d6661495b877e94285116a6aab7b586fe08f3e69bdb096a9f98a7456786e1154bf23d43cfcf344e6ab23eb15f175ba9905f4e4e4bf4e33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he70226e890f2d6e857282d69ab572f6068d113bc660bb3902236107ea8cb6e47c88576268cd64b57e872f2fc88e7dfd774012da25f0cf4a425b6b8636b8ea68e6cc9c2e3324c69d5d58f74596541f69ea304ecdb3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h389c77060694f8c49052be155c155d200ebe5d3373acae239c1d2c4149d8ceb8d18ff32c4543a2e20443226ac1279aed5884e2ec0df3c6250317b5d5682965aa14e69f79ca7c83a436acd059304c9647fdb1efba1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc24dd89bb2bdbc9f58ee40550adafd645a544682858b8e4d7ff58979f8e53bcc0d13ff59e475d8ba46672b97f0faed05d93a18b45dcb7283ea6b084b692d4311774c639469bb388b2834a4559df7d7b0cc186b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67128088ea1a48b55b835614ddbe1b1014729319ee0aebcb07b557b4345b86de0b0ca4cf05055bc3bd3e3c4ac84835f4e8dbc9b03972685b5ef69fc7e9d6ebda153e1855b400b27151952aa66f5cc29747c82da8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7268c55162b91aeeb6fbe1464b0562d698936031ec6e493da7f8d656b92c4966659dafe434a2682d8dde6adadc23df2159456f3f5e11a98c134aa2e305a0db6678251521a2e42d4f43837aba51f08ab77bca91055;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf329959449c31875826d8bd829ee227da1d0e289a7dc9f6c968e9b3ddaafe02a31243775a61a2f107d0a89b8df731198073c3d7b776b6e15544064bb42518cca0c01d73a35dc535124e31b99ab6427bebd5c8482f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13fb24c45adfb45cc2c8f54bfb713e68d3340822cc42eb119f1bc6724243eede8917d790c82aff557f67b79177dfc54b2f2e6db48853827dcc2a0b2825015df2bd8d6492899cd030cef0a6eb43548390e09439e6c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8df6b98bb29867f17ae077961809b2eed606a641beea92b9eb3e12c0d75d4f26de20a8d49e6ab94641050434a01dbc2f16f021835f4d825a509904a587872015b6cabda60e0bedbc242a656774f66080aad7f6203;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb24c13b8b9b09c60f715ba80f3371bbb884aed5d9e4caf6601d2671c2ce59ea551962b8a42b690177e3e6626bd5863d81236f7da0b3952917fa53e1ed279b368516735c0dbe98de568166b4b6da9eb417253b54cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e9cbf630bd43a49111258f259506309d4de0075436f696528c8ea16ed2861bf2fbcfb07d5c4e5ef70182367e788082e9cc38661af0bedfc5783812f2ad88a4abec666dc9a75d631982690e74616e9b2affb8d3da;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2101b7e5753e587349213da4d337585dde458f1944d95c4546fd94808d44e075aab017244d7efb63776ff7e838ae7eea1754484027e249f1597ae9abd6b7f5df4a6024942ab2616bf75e2a34cf42bffa3719a2991;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cdd24cc194842b99dda959b9d9694ad7639d0e968e5d9fa17f19dd3b8e50c704e778629ca10783f71bbccf433aaf6dd2b2527c5528033368924cd1708fefad12ac3f53801a62402cbff9c168746ccf125f0afa89;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6d5ab53e2256bf838b0e586e4357936bad07a3e0fbff9568af0997225beb4a4a6bef0cd76b9008451c5c100c68e9a3fbe4ad5081e0334b0c709a7c7209c8d4df7579e2ccb67c056511e7abd8bc46c260b5e548ca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6dc6b4344cf621d8fda3737c374c47b898dd4c84e0131b1290c22ecb8839a70d1e00204b917ccf892d3b198d7038b5de3c816dc4977c930800b665864f1dd82022312b9dbfbee78f553448b638f2b8087af5a0e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha24ed20efdd113a674b7d6387a4083e19774349343bfb9430e352eded2b0f2ced2f937cc6c498a07295d97d38587f12a97e4aa30763b4e6fb460c1a08a13c72e11496c6e6df2f91ec4d6f5e33448b7639df37115;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h170502dd395760885d7808bd509c6b4873e93793c6d57145c87f525c42c31cbf410ff78748d6f9a851f0c42ebd16328f8868003ed006199ffe3903eaf847953de1bd98945f283b291cc96e0275361f964511b9378;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e01acda43165bbf0473be44b1ec0cf24be6c179963b3e13904f4dc8e19e124c3243cf523a1020ff5f0f241286d37c4eadc93eac05cb61ba56c63f9dfd9da924e8d2fc7aff5a3ae795bc7142c07368325aa4d5a75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4013252e0b246c49c7118557e2f41deb698582bffa5a6e4abb7ebb5bcefbce454e5914c99d61bfcd0fb7f8581abb8d0dd04b23ffc6ec1449eb87b5500678f920103ac0d151af777c74783f40541862e2c97ecb126;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4930347dafd6edc9d4ccf4569af948d3980c474705f91cef55e8ab6a7068188f0a3f9a0856e1f3f42e3fcb44d9e5ecb3274fa9a5f6a5d832b1ad23dbff0888e36604079b489d9b0e03e1c11d0c171cc88e021bf3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65c66145e99e363a095d9b689fc6a8e984d389a23ac64501a2dd81779732841536c8f24c522abd1f2fb2386e352837c91dd2b19dd5a0e994a9f7a49673b7348699ad61a630e89d1a52f2e4e6b7667a72993894142;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2fac544ed342c4bb938976b9353d8f159ad4e665878181b3e5efe943725e4fea435c37f312823f43151215b34acce57a3f864d53dcc52b24ac1382d1ac35082dba8283726ae96091a4d86ee25321cc473c40d202;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42561e130f005802130a74d9f1ad7580fa800afb3ed9d87a6dc08a43fbc24bfe7cfe433d749b4820e50ebceaa4b57eab50dd78c7278f0d0ed3b062d0dc3dec8f2571c682a4308bcac108a1bbef39049def46b7bf5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80686de9e9a725a363e266bc048d76f7eb96e4105fdea8d48cb57e60c242d8592f98fe81728fed0d4c6cc948099d9afed38d6c84ab20574a3f0c62e25761d29ad627f0c7b61ec4127cd9a1227523f1d3fe55fb015;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdd628177b9d0b499febdc160856a95819bb67267e39ea6b5012f992ab756488c2803645067686632e92681dd0785d8a818c14442ca08914e04b6d1a4ae62f4746d812a26c917ae99f3adc0e85902e5f209cc4bf7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d49c46fe0cbe257368ce9ca5e0eecdffc8529d9cb16afd4459af90033a6b691f420fbac1b22c3f44c15ef8bf4559d507dfbf66afaf0a99a99ab45868c923cda28ac119b04352617bb4f7c716333864c9f7a395b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5135e4909109eef1820b70930c0b217245d01369b29452a4c45af2e69d76aa752ca9d8b8eb9bacc388ff4d56dab38702220adbf2bc04e2cb3e72a6cf795b256e01caa6efc0f0b3ca0c6a4398f7709f02425d99dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he70b428e24e8f0671d9fe664bc5b5d62f3f9179b98d32b5d14ca822207d68ac53a2f6f0120eac8518a352014fc79649c1511018afc84a972a25897ee3faa0b641c2b22790aef13c6c3be13618f46641ebdf5a37ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0b8ed0578f8627018075e6639e0e66ef5d2fe789bebad356c267f3c811b7c2a80aeacc5c0fc3049d60f0eb9343c4c7f004723a410e2e7421c3a286cad27e792a97aeb74c74a355473ff23b4cdfef30f4820eb200;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfabb8c51e792cfbb1c4ed636b4fc0a84cc10c32b568d7b3c09005a01f92ed0dd1644cefd40de808f6d3be2c1db24a766d9d3c1307fb2b19db4cdc8c8386fa8902fa9063a25fbeb83509d10b3515041342b60ea26b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha67812931af071730d8ddb46cb4cb61635fcffa861b9e2b6a7794f0c208e601e2decfe29befabb425eaba0ef6b9044c8e5008437b011baaaa68daef1f3d9926f86959f35c270024760476d6f13000b5014f5ab5d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60767651adc8fb8be14833f020c9990f5dd97bd0e4bb61bae0ffe45c1b63950c6e7dc1459582b0c476b716350cdca319c45c4f6d2fa6e79369daaf99a0a9ab87ba3915042d23c2420b2e21e764c57de1c9977e802;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4550328bc5294d88cb23a093702d9128391ce1eb012fb6388b7b56c1afb24535360838e55b1fb5f081471c3b3718eb88b8d6c6021d0564cd2d38caaa2f5845085c1ca442248abd06593831d97155a692431cdeb2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h883eb8b42ffde604fdbca4ae0b24bffcf2315de8270346726891ecddc61212b3a1428d61595068dd97da0a01e98766eb28f9310b41a96ba999876b2b47fe5abc59134a24faeafd4ee412943bf32b849ef16fdcf1a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h442240ccfc44ff778cb3ffabd30774888a4117a48c6fe8bd2c0d790896ceb90851ba04987a1e85a2cd15788dc573450fd6f1da21ecea51ec10d0a3d5b2ee97c60b0d7f74a20d513007fd57a625cf21b9848c57241;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h456953d908b0861c4e41e088d894326f0cff84954427d9058b58fbb40a9fb839ebe75a2fcc89548439996692f7884e777098778b64f464d2f0be05acc8098ed89d28c6275a1388428a250aa832d38cd79a03a66ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90bb4ace45b4254d39c78515036ccfdf4017ea5d2cec88944b223cc1e2976a20994de73970789c4d7866020cc09028848a9a5408c9844587bce874586a7f617270aa548331ba1e3840758d765a1ffb079f6df0c35;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4156c952244ae7421c43ff179d3580d08f8067a0d570da19ff38bc5ec32c4bb1e20d0f7791b65903d3bc6f9434eda451be49d8660317c589c19f9410063488747501f8994a769dd6e9d93f7588621cb54951a9a2a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5c302aea9eafacb418ed99b8e2c29d7bb6610129e62a3f62edd6912c4e2e7202bfc64a51a2c32df56282db9ed1f467494e55323b7236b704726d2033ab16c6d2c3c581b24a86e6372615897bf88989f956b86c6c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72bf71af7fd43a285c10b24afa5cb7ed47cedce3a8b0e4006a50c2671459d98a38d1838b1575ec5b50d40323405cca65b9e0d9b304a3c7075c7d6c1d3e055f06c4b3e93bef3cdb0c0b4f1ff98beb3537df746589c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef8af4fe482057547c087cce18dbe2c35029ea35cbbe47d4e258d269a6a24330c1b30fa3156fea4b041b32f6c6c47c93ad3a7a6eae6ba015239c8454471e20799e7d54052e2069680fd5c298368362f491f6110c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bdf306f88d3dd9f37b1427cd2f474ab7a077f1ec2210f0e65b50a45c50255ee9622324688c5ac1c54bcfc5ce18e296d91e02fd77d9260aa94510488a0ef04f8f0555e88ee15c3c3d63266030c38f44ed30a592f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f7dc90e7db817e6fd1e2734d2546766a09aa1a8c44c620050b3312a75514d1dbea4a44c850e9a2b493d34998be2244a7944a39ec6a12799ebf8cc757b5798943f0ba2859d004f066203f4b8e3c2f2b128e8621a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e35db49544da44653beb2478cac2cd8d61c6762b87b070f3c66dda875ea203ae0e1501770cbc0b6f9816d326071bf91d3f3fb69ee8d982fc1c48890cb3eaf4c28c6bc2b975b28bae102b9016ac6398dca207832d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70123ba0902532898681eef0c48fb825820f9535ab7c19099304e0bc1fd37c8ac2b5031fe2a9da0cb7ca2cffa5d418e4272f1e768fdcfd29398273d95f03c39fbca06395405477582164b1020738d029dcd6b750f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4e85616cb3a4df1978d5f6be2724e5c63ca6f5feac531587bfcfbedab68962c4db9bec164227e5a11fca0b398e434df1886856b00467276f3d1e79611fd93f7cdece0b747de56ed2b010eb4276acdc99a4b26482;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2f916d11e5f4806de56eba41d67a0225a67722acba3258918d21927e9a6004427574ae1669e282a62c4edcbe96415d364320556ab49e97c4c75a88038c88eb1f25faf40705d12e1b031fbc8a8a4454df0b00cebd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd061c925cfd4157c9776a8b621d5745c2c8d2c8b580c2c3928d4ac54bdfebd4c901a105bc33860827812c0c723ad62171c72e3535ba5960601f39d145204892b251f9b0fb58b1f98d5fb32e19e4a9661313c1f0d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h988f81351a3150dbb578e73712ca991f92ed0558feb1f6e1dfba784a73410060a05cf40427bae06c313f5e1bb1470a9d474f654290bf526ac2ff89f7494f01e3be310ae25a3dfdc64f027efe05dfaec85cf1ae931;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54ca5326ef26f72c5e3db27a32fb67ef91c8ecab3e5aa33cdcfdab79039127de1530d29d41d085e2b2fabe952c739ed2c83c1ef3ad4fff7d3398df8fdf424076bb26bd38a9a4a4c65763de4d2743d9617f1c3cebf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40fb3f9bfdb08a3e2406f4ae0647061db961dde21316b96388adc8cde6c0cc538a82cfe83139355440bf466542c7411b42d6b5249dca31fabedcd73eaef5a12287ddf03b6d3cd0d9b3fbd0e3721253077e90292df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbb239803769f25dd25e3f987ff086ff367f510a25a87940e30bfc67a18325a0a9caedc7b483a9816fba6e18cbb2c89a97391cf19dffc89eb370982a17545f7f1be35e3049819c793c2d5266b4633b0931c95943f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h503a3467f9aa492263f64e8b5c785759eaf096b0271c2a86c3bbb7ca9a1cc4a83c49fad4c272044f93e8b964ab1ced6bd20f90e43083ffcd81362505974f21cba0f5c1a88095a0e4db844cec6b461bc31ee08a3a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5886a684b33098c83a5cc709e64c9911d5952167e00467e3117461cad07b2726661dc5fd127f6cac4c09d1af3d3f6a150a14029e59ca52d077dfc589a8e27eafb223621c35f48b711ce414231968fd07abb56ef73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c9b864bdad9b71d6885b80f87d287ea312a01b140a92ab1078aab9d749d5292b1488a83b2b484e474772b591994430da00f03575c1fd8472f72c776c424725498d8486138d16f12e7cfe2c0ac0784081cb21c855;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f18f5235c3236714fb3af9c72fc831df7d04a15e582614e5d58c72158c678f18ec31289c669ed0096e40c179f16ed1e97b6a9c9c640583aa25e31d5d6f96b271bee59cd6e147c574cb4cf28373db75c5657575a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde0344679ff779fc6bd66ec5f2338e897ab6ada653707ca0dee93a43cf59aa4020561aa7053f6f33613d661b3db17d68409f62175c70237ab036c16f0e9927d61525f7fe1004b93ada0926ea6f6d1d5d28433e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h177f791baf69238d76c4973544e0ae301d094a09e8ecf2bb99df9ef2caa9596c90df9fb61459a9e1de5cfe3eb8d6c5b8bb0a7019b03d8a0695e173d2adf8b40fda6ca0cc6f4042241c66efc85bb5ef1bfdcd996e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha12de278a07957c6d7ae952a8a8125050f4cbccf4c546573b51ca0c66bd87e160c29ab71a6b5f6be723eef6b20d0f72d528d1c106e8752652569e5d4dccdb8fe296222034305e8e4dfb171aefca48e5ccb8c24fb9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9d180481e37375664ce0052dbc68a8efa109bbd1ff515c95bc38324a6dcb41856642bb0027dca8f1c32b5ec06ebcf5c92a465e485a58e5343aba0a4bdd9b33f8ab274f063b3b945b9d6518f6de86c0989b099b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc58b9c6148c3631bec904e8078c978051c8382faa13a858fc6c574a820450ae3f779b7e27070dad6ef688e68121909f9c9c999509116e53973ce359c4aa56159017f7335f6f90f0286fccb3711a6dab1dd442457c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf38b96aea46bccfe4d6ef4dfb59265d649156311fd7cdca315b5d77441ebe73daede5fba590922644b5adfaa1b8ddfba21daafaed42fcf13e614c83c2f4357a88290f18b7cb69d39f3036c4e6abf97d5606b6a355;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h648ccb434d0fabb84d1e596468cf2bd2d5e0bb2a2c305ef3eb929d5f5f9e09f5aebe6bf3815eea642b0c394821e1720430222b3cb3426d04cc27e4da15174468739a2d83bf4a51e17d04edc4f3fa7fb808daaab0a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5812e98a6fa8e60b46a31c6f84f87efaeba3431e8f5ace78d4aefae9f4f24ebbd94dc1c0326e009d5ab05abedc3f5abeed1ea0e90692e699cb41126f30f247c28905c8fd767ad82c9ee13793ed5359e8b0339ce9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc37f73436c3f98da7938b66b8d1a70dc273eb7db9ab7ded8165aab4e8d2ac1740afc179ec249ea2dd64ca0ab472eb92c44fc010b3c8875bbb045721062c3db89dedfdd53d17077b318571b21e1c61a66de47e2a95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h649f5edcc27786ecc9664bf7b409a25e3de744a59fb430e624af4f3ea3dcf85d0f446f63890879f752ee0d04c9b1bca7d9e1cbc390c0026149e6cfaf97d4a280b137758ec0c8ec5f4abb45795e7bbafd57bfa9ecc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbdd0e5099c3095d117370cd7e217c3e1265d6c7616feaf986dad77cb043b0f81721dff737bfadfc5cf48d00c3f77ebeeb23be8fd23bc6cd9333116fe448e8dfcb2272497525370d087a86f2485f4530fbfe6aed7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h521055da031ed935b19293ea2b7f8e02f1d669b90ca443400e0b735eb0a15eb0834613a04f36039378f897da4c2db26db2816c785fe64c2f8d499a19591189f7fe0763e8bfbc62a4e6d17b5c0a8d4f041b1f8ff15;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20f4502bf1c5ec77dbfbae47624ab32ea1c12b475647528dfc215f8d2acca83d57290e91ed706b069f361b60b9fa386bf5a53e4192ddf9647e71f807a92e83f250c20444f72bff61f9d8855077a0a2700e82aae8b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5118b6f94b4145aace726f05d4d8ad92472084d18cbaf05e64d67592e8918559137bc47a4a1f099c310a437ecc546282009f3a9c60a455ea144374544ee7f03475afc7c97003a08ea77d60662a7c056b64332b37d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81a9e1facf9d1a2b12c19c3a38035c485b3bdc011f4f770ece7361525a4c98957c1ad00dd8af0f8df7e6f5b50c11c793bf5b448367a7321df3ecd92b4e6060b56b3e85a98dd1a3da0cd66c8eedc8d9577a4f0586c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5be9e48d8c3bd4a40fba7b17b311ff75c7247e6668fc9f92eef7c186ab3add73646e2775bea55db442b3a38e097c2239cf9529fdaf26418a70d2961ade94a90104f03532844f3d401422ee655464046c9db9d218;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9211d40240b6c34b55ee249741884191c51122e371874f4e5e04f970234ce8946c19082e5ba04f083e0d18746524c1f06a75082dcb4655f4a0ac7763119e0ba133f60905b5e6b524b3591ee65c974937686172fc7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9796f7e93d0eaf34ce8084de98161c9edebfe4564e933a22555187330266d49fc5377e1aeaf8e629d524b7a9e9a6220277bd4cfb13b32b70ae8355bc121479bc0f380d06da0fe60a347753c41c12e74fe7346177a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf511e9395b9b83a7e82a82d4128842bc42bfb3050627c8752799040a7b9d2adb4739dbcfe9f20087e61f5bd34f3dfd402d93b70bda3f2233e576fc3d9185a0a7cafccb6aa6e4db547246cf23604ae61b33b78d2bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h970ad9d0ded676c9a2714beb8b15a7eaae279f2e67aae409c149923bfb1e4068be17733d7dc9e79e9b86ef932cf22c4608f25f47492eed56a516fe5c54599c045b8538fef6efa5be57f192e791f423a48985f2a97;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c371804b9bfb9722475481bb7a66b77156bb04dd3ce50d9adbbb007066925118b1122abf9ec7f70e7e669799c09db125d30ea0e3187c0063ffd7895de840414d8ffd71d0ac66d9b01db5f80bd605ab36f6cd5871;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8502eecbdaabd1b1309dbc35810acdc4f19de7deee6fe8882f53b6381e048e2cf19ee334b767010dd45bb287d4a8608b063e7d57edb7ec5e89464101e3fe6495d97a061bb1f63f5f35abc2ffa8ec22f00c4a79e6f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2edf726dc7913c18a9ab75eefce9585d65837d4def037038b1f303769b10630110fb336c386fba661d38c2c5653015e250996711a0c96022c165b0e3ab8d3f544ab2ddc6a617ff75a5c1dc84bb32cb188600fd35f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4627ae078b7f667eb4d96e6202b049b28e1ed6d8459f21f361c6ff1062ca5c8abb68e3a4d329f8f2b2fb279f48581f56e6586daf15a9f31045e939e6ef6aeaf50511f9646f125d4715c6276d49163c1370e2b0e9a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9e6aaaa571932efe5bc562537f6b54461a073714a6aa04c6df8a91c6e0dd2ae455919b180d2a656732e998392eed4709b4c27eb802ae827926bdaa24578d62919d00a8e76d63e16421c4f818a6d13b140503474c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbb7cc7e287d0b3cefb544eef0fd9acd37d7ccfafd7486f2be4761e839ac42cd47be4ad0806b898c237bf20d9e12fcbeac8717fed9033ed261c8435d00278129560d621575c879c156c314cb86c5bfe1d9971d943;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he60e4d2ccdff7eea37eb919657769d0d0944d1759028337326857c19a8e98416d8b8f46895b486c2aa3600574a2239fcdbaabe3c8e9b78f493b6e5f23ac4594a73f3ec077e9dba8d6932020a0d0fa991e6774f3d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22fc9ec91c261e38f4eed00966e8e0939b6eef5c7f57ccabdfee399e3302bcba508a0bce7c9f9c494e5600fa8e742bf9a13f40bf14dd1862474620442690f51b454ed7e8ed6b18dea4722317130c6f6fe6528e5e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18a29ab99bd7243df6c691a06175a38aad8d1f2fc5e81d19711f5c8d1b0254dde78f1d67ef7eb2d6f8c4ca75397030a7271fbe03e932257d01a4f8e9f6fa09b2c8f73976b7936bf4de500b3bac48714841164c1f6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h844be631fc8ebf29ddbff78cbb843e958bdccef7a46d696d4e2efa2a6dfa38f924dda4d939d025259780d1648f6adb79bd4fc6103287d3b707b64411e544dfa0293cf7cadc019ec30ec7fbfc45d068bb628a6e7ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56fe91594384fadbaa3eee81911bbe59100c268e8631e637a5a3239f8be846a89cc13808d173c30d6d47dfc4cdd9463113e809f31d3c424d23038d278c79def6bec69dfff504b8798efbb75e4dbe23956b83d8650;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f27e12420b9cdcbabf74598fba387f9282440a2c23fd9cd779adb11365e07a288fe964a6f5d6a038a5cfadc65b4606739ba5180ce9db7f3c27312dc50bc6007f69c5b0bbefad3ceab4c841d2f0ba9760f5522549;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h352f4ce6ef0a4ba54c4587393cae2ced9c904a4acf8e1b87e1ce0c15fd58fc68cf7006def1aaf0e57bfbdd4120ba1b85804967ad5ca79cf84057c2d8caea9d9feb0fc07ea48833f2145ec6fa933cdb7f7faf54da8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50adf6a0795bbe841753001bedb96947fec04088cf2cbaeba37079cd056e386427be052874c235dcc1cf28581a06544fc21514fde4f620234cae0e7d12f26891f9cf1ffbc69c9a2753585fbbffc7d80639914c971;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44e84042a633ec5e1f87bfc64dfecdc290f0acfa08e66a28ad6cd0950b643fb32d7dcb056e664677272b023cee00d2b2642cee64d8c1bbafdac237c82736a2240d69da1950032799e9444f22c068674d0ed05bfdc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2af592b9a57e8277baafd0c0085e13c676b82308c752f0b3ec5564195d7b6a32b0f3d9e7b66f7dcdf4a37dfaee552c492dc4f9d0ab0afeb2629bf06c820f0da65318f7311cbbd355c784dab8572311e8f8a9338f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb3ea770b85b8506769ad6ee99b149f97822075a08d3c73c5fae9820eaf985862a1766802c1babf1a3c17e863239716a1dcd659731cb393a68d45edb62dcfc02778234f861fe9f5046b3c34c36e1ebbb9328c9db1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed2d786eaaaffcc754f36893c1dee2f596d5a08187f61332a9218a6f8ebf3bb69edc4deb564e8ca669fbc7eb83315e02fada28a84a79db2d50df30ab1def221f89eb731048939811f8aaab550aabee83a4b7ba5a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1251e499f95e3ed15a97de0f2eeb70f288879e0409ad786a3482ae73a3065173f2b37808868cdb400ff7d49a655c34e2b6712055565ac8448084ed7a3294bb7f46e3a948414c40d3c71f967b382cc767eff01fa29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60aaa70b29ff167fc772c98f4ba446122121325860931c62ffdcae74ffee14f42a04ec88f584837e961b4fbf5f7192f2ab8abc32b6d4c4802e39e2a20a3daafd352f9d460b58f3e0c1031790a83733698471bc564;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca98c655b313bfa66815f624e5f8aa7b53db5fd87cafd9e8547de713adc23d0e2c829f83598124d4087c6eadea3d6d87bbae9f1689d781ad08cf4e60ed48f3f7bb7ae004b6497eaf6b96d462338ba830e2c86cad5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h982c239a038ffd7e41aa72258c4d0937216402cee539236aaa0019c5b32b165b98f0226d2a49946d3961c7e3c30a450e9db8b2dc2ebe54a04d125afc4953688512b4d9d21d1c76000835857ea6a7e647d1f81fd77;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9528cb4f20313e6fa437a586d6bc7fa64acfa6f489576e8d6ea3ddff4c87137fbba7f3de448f20e89a462ca2f595ef1ef2beaaf622814fd108c2188202fe93766af5449273ed4f3fd37e0a6aecf9ec4945c2367a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf619027eff601bf1d518a0ee6b0ac16f09984014034961e0a01ee6efb782a652023a838a7d898728aff55860bb389f344ecdc853861485c5db20ba283f546e437208317ed724b27fdce36e8a86dbc69126b8dbb2a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf99ef79828fad59d6be3eaca2561d9eb0db5dd78a271752a657e431bb2ce245361a8eb716f368988a1531c57aef198f00c98078e528911de8ce4e2cc25f1582906358969514037628135b02df9f03e55b2f545663;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14fc69ab0cf0612fb698e412bfdf91388718d2cec3c86109d883692f66782a3d3a58133b4dc4a05f325567eb55ed37192652d159a572fc91f9d7abd967a1254063a61c1194b2bd0b5615b3618aceae7f566505d84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56eb227fa8d97fac8327d061d6c90d2edc8c6c16179efa16c4f7d818afe61411bba89d68bdf143a9ba1639252e5849648244a4fa31cb6a2f5809c943f270f9c40f570d0a87b7be9669c902512c8311bfdedd8696f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he515ed606800c11101001c5a21f7adf56ee2f1f0e3d1c40e0ceeb9d1f4955765794188ad7feef80182a687263643913e722dcf57d0d805f9af567f05fe1f081f82c9685ad1b8dc754c1998fa5eaa962032f927e5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14e6863b48672e58283a5e3eb0d8912147e6ded5c07abbc16484329534106995094009f9db981a18ae28ac4ba5ff3f5ec8d0bccb59638b16b8a0f790ac091cb970b3815101de67a2ee49d68567190172b7a851466;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0fa6ce71f2ac90a4c5a4e2fa916e44b53aa86c5b8b51ba983bce3a2fc15f683fe6e385fbeebf914cd622f0ca2c620b39963a8653f99a239e04612cabc12f10fdf33c37015692b3ad30ab3ce0d30fac1d94718c87;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83f13fccce4ffd4f9aaf1e8110c99131f4453f5568afa42acfba0a4bc986d6cb0195f237e501fe5fd65ca2a35d89af75f71d3681a57fa4beeedeca426089f4664601324aae73ba573a8ed8f2cd5aa3336b1ce2abc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd35810d381f2bef744782dd03d20c9adba2e5128cfba1b868f3f6a06980874d4f61028a53cfd7e55ef938b8b58c5c1c239627204131d3dc3dfa8d222defba31777764d94f730ec4d45e340ac0dc8514544aa090d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8719a0a756d677c5f0fbbced447034c524ac4d38f7ebee1a3288644ff702690beb88181f269f4eb858e1a829dd882e56bba0931c0e7d24e244aa7ac15173fa1ce7fb13b8f2cabcc2983823dbb9a2c13ca1e8e4ddf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ed77765f4d205db7ad0e8a3999385d2a6343f6e495bb15d8429ca213bfa472b8c578a8f72458cc847c08925a6852a7c35650f1b42e1dbbf4b86261d5d67395f935622a547c393f015c24bb82d9a8aba421fb2f25;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1471394e0942edd03651363e12b90a8fb38b4b55b8af30b06e152c9c257c2f7464a84b999ce3e2286cc934290be706793a5811b7cb30c5277898289c36a98f47c033cbe18df5dcf4f0e694d9f543eb8acacafd91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2959ac0e64ee3858acea927e346b604fa41028bbefc8bf0360977d52c7b0d3bb1a623905fc3f0b7b9d00bdce12fa169ff5437976f4380f248e1bfa42ddbde3344a9bd10324dee4cf91568ade691ff224bb9d9b72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c35946cd1f17cb49a68140d5aa65d58b90c68e6d4d8e1ce2114c29891bfa6ecf97350e49d82309c204436ee39363d64e98cfd6b15b752ee1d1a4e04c0ff4b87d0356553e36064114000f85d07f34b2b022fa680b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h130416f0400e967546c09ceb383ecba5b9a7706752a4e3997a66b32502c205f5b8ce647a7f1aaf5052b56bce672a301ceb031dd49ed4109bc2511cbe1cdfb0a164fd84f9cecc2eb3705c67759a3356d65c93946b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f73d641a89bbd5642b38a0f737414d3521980844e826d7137d6af477d011ae1c8e41b75b9cd38427c2c02d5b891785e9115f1a2e54628508cb9a982dc3689b313f1da5dac3f77ead049e72d2ec0606abefaca79;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba7f2742a9d04cc88c665838b175b42dd8b0a0f374b4daca47668dc15447996d67ffa41a4bfb332faa0e7521d1f53a5c482b6d53f8a7d9a463fcc46b3b1bff194420da31e419b8321d1a544fa1324faf915537911;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69537664dc6558b432b5fbeacd55662884d60711fdb890b365aac1bc8f07d95afc31a2bac7eaacb3d2a8132910f325b3f3b58172e20dcd64e88d8143d0dbadbd03dfc409237f552e3f376e7de44b99ab6bc121149;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h289eedd22ddc1c2cf36a36005e2ae4964da9c465d328ca4f19bdab20d820b69269220765d626f184f82cf3d32938311054acf526ac3d6fedb4a49ec362b04e8f885b94b882b08fa070a83839529d232e81f85af73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3c93bf9ed141135ae93479222d45857fd5eb4b87e19fddf79834ce763e491745d6e5e0904729accd256a7302733893645441b1b01f76e6b2dba6a091d14a022e9524eb27f8d6b69c62441b3cb2c19f5aae24a3d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85391418a25138075e33e60a8c2dc24a3efd5a2c6f19233e1e8623579c1817de2e805971ac7475fd913815476020a78aa63514063445517989042387175de9817ea30bd64a6260b3317878795122990e4b213335;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81c2e32d1a8ad9ab96bdd81515b2e61f02b05b9ce56bd31604a144d31db861e835886e963776c1a61d69dbb5132c8728af18910cebc5033df1ccac209895b5b4c8397db11b0d157cefebb569aee7095d952bfdce2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20ecace3a822da90f211e9c3e764c5b8974a1cc3e1a72c4071958d0d82e1c07395d90a17c06d113253e68a774ca4e2a8d9daca40da4a7b983774a7ab6ef2ce55662eb4a761edc6376329b651d236fe2e5febadb48;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3191bd5a6758deb45e46442248cc052bbfa9564ce54c8f6328630ea294bbba88580dc52b3e6cc9f568f5c5d57d46ceefe8ea6e3153d6cd1253eb15d12c3c3d4a2a327912a3e9380e9ae9c1db9174c1fceb87b71a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9440f2663d3efef364911d0c16a1f92dbab5d764c4167bb4409391e2748d11d911bcc15f46a604f7f12a9a87e394c3bdbb4ba9e775ca5897c6d46b8ac4f3e610070f62ca79db01f503e9c142fc9a387248de19ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14ae0827d6e633d360c51827eedee4a8972683251ceeef70f59e50d80a3cb351786daed53b75159eaf16bfe1e4bc2b2a314d8305d68171315a207a6c40d600681bc3cfdfa791f0cbe60c9a3b4651c91ebaaff29a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb199d4458d25be52be541821e4ddfaecae6debd36cbce390a379bdd397f24ff172ccad43cc88b7b83f304d0e66f839b81a24ea41ecf055cf2506a88990216f60c1a5b13b2890f434f2a37f59c961b6e55cb648b6d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he50acadeb7910bb888cfea3bf4a4ef0a2692d4523f7666faf89042f1fb64c754a877e5361064352f66fafbfa4bbd210450a1d6033f0746bda74981c58ab07f53037f33e1b31e4b139140f49e93180d5e4de4b15bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb82fcf25f2b313f449cc8612161394b60b7b7666ea0181ecda292caee4e609db5de203483a3600c736152838b4157ec3df6210ecc511e494cfa44740f5d108d4c008f88ef838ad114bd3c7a536aadae21d89c4ab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6542e47674cc00804913d311e16c264bc997280c361dff6f75d7021529f8532aeb668b93a8386bdc9ac77ffc23af017e3789baa4cec2165b4512c047173fb50d37f8d2e83c22b824df584f7e3a5513311fe3a4e47;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf053712a20d3292f99ba05b9e3d9381e39d7e3cff18176ce96bbb958582ae43f3db3e12ab1dd328987b6c33f2a51492cff26c2c58de1344ec8ebd8d692df50129a97c913bd985efdf374ec586cdf45e4bbb9f8222;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3b68e5e772555586c6ca7c96374f1d8e10403ae05c1dbeb3724c8378c56444876491a1a12cf8a457c74fe1b971a9ec09d8bb49fbe9fe427df99f8785331226ee379fd0bb6b82df19e50fd4cbc2109a1c5173b882;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he59731f2bd19104955869bdef7875a993ae3f480a4aa5422feb3ce3bc7409fe0d1ca790912aeb5b578dba1463fec1276489ac7b4cfaf5f283d74416bc472c11652b59182cc89f40bb3a9a3473a98a5e3934fa5db8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c7fdb3af6e2f6a8f7bdb61eca8ff2764a6b8f1c7b8817fcef572bbbd2532b389b6674ce3fd3408271aff0e785db65d2786a022c0c2bf07d740107d90597f4c773f84f02ae47e4bb897952e2ee52404d23408cef6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87d26ce5dcfe9cd3b4873843b5c59c0c45cd00e68ae4c7cb1534175c158df72d9e15d212a5d344063a011682d1f8dac4f76468c2007aa343b2ed7ce0c343981bbcaf971e728210cc565719061c1271aae120d103;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb33e83397c43070603bd8e673ace8fdd89de515bf2ff605a77dd9726189ba9fe15228a47c76bb61561a08a52ff4262940b1b78f47f42049790b9de79a8ebfd76a8d034c5223044e41f4f0de723c1b8f917db92142;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d1396dbca74590f16575179f66a66c8284aac51ba6b4de50c23652484dfee5847a7b69efacc13d47959098f9cc6a85137b4a3c2379321e649eb917023b3d6bdbef9e86def442c87db3ce6bd0f2fe37fdc3d94d54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbda24729fd68cb9c0e07ed28857e7c340f43a0ec9d39883da9f660a5de0faca9399a245c8b54b2ff9371d2bf0e859635f13087809d544e06586649cec3b1dae95d14e723a9290bab46a98c6feae020d0528fb874;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a27202ff40f15f4182542e26fd1668519a5041e7900c606ddd7bdb7f6def386e96e40495fabfd7bfda60b5b97e288f893d4016abc53a16294c9acafdefa2799f313b92081281d5aa80574b3d844fb9c922b921ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f06b052ec0316e5c0b187f0e2712ea91050708d74b9d613d607245c71338171b05268a4ae21813ab142dc186273996027fc1ca325603738dcd72ef14e3e1e33e080803d1bf18dcfb639f8622e8c07510b2c024e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b02a969cc35b055a7cbd1b206a1de747b19b2973208c5e3ba9ab5835dec1a6090fb27538786b07d7b622ebe6ec69360cd51038e2d989303f0fe6d8424b74849dc8161aa685fe018ea4fea3b5c1759a36d86a787d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3ec0a82308cf709254f14f52a68d34a2f9970be0560b15b3c25852b7b69bf6ad37b2f70827835ccbcaf14c17354e201f7cf7e7aa2a8bdc8bf81e1922ce11da87b02d77c10f00c87a1287f43e539dade8003dffa3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had4466373ce469988ba689bbe2eecc15688bc3218f96a2bfbbd6e767d26cd205ede7e4d7b3da0ed1c5473c6eeb578a2c6bc6a50248ad674d3af5d45b849c8883c0f7e3b5e1e92d9109f101d0c99523ce5093c3eff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11a65bab77f8d8773af16a1e40078e8618b4ca5978576195f363cafa2824e0aa45febede8ab63f41a2205df21119f90df27ab660f8e260b18e323a543660b3635cee874644a7814f281ba0cc133dc3e550111752a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbd23ff43c796b7bc531fe2bea9e7037b3e2c9a2ec1fd06eb799e39ef21304dd0ca92cbd554eceb746c3c1ed2151192e49efd4a58def5748953bf4f14831d5229f7433ecba7db45a90f9db6a5a481288a84ffbfaf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6282c39a7d5ed709414bcba3daa240dea7963bd802309be181f03f5072b2cb103af7a0678e2c59221c6553050bf425dc62ae2742900c7fbf8331b11b9d475363458142d7bb0e190b2b46cdd62e89a2c2d9f55783c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h200c543884d9e319e13fa8da898de6435e203e9c4ec858e09656702f3134ae80b33895de21edc49123eda17136eae717764f07bc6525162419240148d9a5719926acc3a7bc35300cbad982a1618a578f0d4c5c1bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31fe756347bcc14eec307bdc8ad210a7b1fa46bcd792860c0efd9bb365a3e85debddbbbfc5e54df901dad046ff2ee9394d99224cb52e675ccdd20b873aacb14b1bddbc5037ef6e04472011faaa3984660e0580932;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbaa79b18703c7bded319d58e8d8232b3dcaf5c6617dfcb83075c7430341af1a1bed4b5696d50f3f1e8512fc06673f6856daef792be92d05e33eda68256d77f1a36eaa9da1c01b57f6aaa752bad6bdfbf4d3967735;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87034666637773b1bc43e7a116fd50fa4195fe86cad286849185dbba637e7ea591af0fd4931132a292eccc56fa57a4f1adea6103fc60e520f7729d73bd1bcb27461ce26fafe37e8015be85b0b2eda909048252116;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3a28e779672927f47c10aef12354019e6459e70712f64b208793d235cd582e8597d2f462a51f39b78cdd2f85a73cc5824a00cb341d1e6ee1c8e2bec7d53e8d011170d72fd918963a93924fa78bdfec646c94885e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h652890d9428f3d60c4df391e5243befd5fe9e16e1db5dc15116e201833fb42a3233313708cb2365fa3fe5a2319c4e993a73fb72c402d18e8dd8b9f613cb78c91def74104cc4217a9ee7bf01024dbcd553c413f942;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce5e464659f7f1c0cd6cd83a24264a442f3b66cff9ddfda38c94d91eaec5bdc56857ad4ed628511630349989a368531deb73b70f53bd8dc51c82d33bc6fee509c99f19855d22cfd17bf20864b3fac9eb0a553b082;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e13ac41de842b36664ec53fcbb31ef7e7e3cde7a56d1e776066003f0b018db505a53e2adce3067f8821c9210827cac87279af0d9cd93e8ebdf5b75999a0ef0f12246e752061baf72dc22867e3f9d62fa526c4c41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9a5e30a65f732031da18f1c62316902cce223e8520d623c7dc6531071996da4f7c357600b81c2b20722e3cd2735c987e57892acb4d4a9367cc4315e8b8914a7cde962555996811d51b5c2858ee361817120522c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c75bba2c864910e971ce22f15dfa6f0f947733ebc659a233abf42206457434bb960ce5d1f6ecbccc1dfddffddc4bd92303e44122d2a9bc814eca3f1928337cdb043b451e2d1e95a8be9be22040e73b8ac490a7f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87a902e82bc5150848fac2f0ea3efebcbe3a6351e415e2852c867e8bb2687d7cde8fefc14fc714e9675dc5699327048b15d07c1629429c41f8f09ef9ad929439741f6005c9b6b75b1c4abd8ec8b4dc63aec118436;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbe659fd30d9464574dea6bf172f710c4a439a3d43c95d7c265ce36160b309741e9873e32929ba26007470f10875c93f3cd44dbf753098713b608f93d26f08aa2ead813a3107a5db0e7d34c78e4bce664812653e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f1ed74bb831261b895bc519d7eff0e8829e4f05d40d2e030adca370ea08421330be79a9d5806da0194f4de13afb88db740ac0e564a3f11de0273886e143f54fee2bcea9b9b6eeb4e1e358d3af332b6ea4242ef5c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9f7a9e387c3bae8ff932cc73b5bd0d7ae7577b9d06e57bb2d17641b9999d033b817907659936b0df095812e53fb17b6adb8f25f764284b6a8179c5a61bd4c022f28cbf0512fb06ef321295f50795139b5da79397;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3af3a4071f5c440052681bed4daffd722a039c92b57ab4d130890bca4522392a2acbaca64ce236875d7c808af6132ea6f43a698322059ec3a4a2e8af83163279c0592605a31dd2be0c7fd6cfb7a241897caa8dce9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha885e957684ebe190676e030253c69bdd9c44bfb9fce991d26651a86cb07c24c0d14317390c4ea24e84a3e961d83d71a8db40207f3ee6a7699f2602c7f31b82c37cf033425ce351bff594e236bde2c2de8577fa5e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b4a7a097e6fa0978bc8540fba764865feeface01fd10c3462a239db356fecc3b7bf36072b8e0d15738c265704c69ba1e34a26e5daade6ac31df62bff4bdab59d1a1a736727a3029f5cb91027c600a7ced9a1689;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dcd84b5558e73aef44e09cb219130a610a8d75d7ae39175f9a3965251d90f1dfb3cb052032d550c4b42f74c6583e1a96b300e224319942a610b341c1a0f2df460f495ad11c294ac618022a62d8e54f8d909610ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddfe9ebf91796e9e4ff8f052fad4f699ea1879d2401a18969423da9f0e690fa68e4808a0a67466d969e744d34bbf63698ef1dde506c011577fa2477b3bc273038261aaed51783ee7a227f52f9996e97c231285a86;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee092ca1e7c1ad0716fcb919e5860ce2a49ae2900612898ad98edf8011995b16e27f5d019ae70a76043af532ff8ce09688ee9deec54e65433a1a2c70ba3dcfcc22a961ae32f80f695cf99547c2e7f440a3aabe66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d92693bc694c7b6de7ea997e5db2fc8d61a6f47c5dfe5e63786164562ed8213f9e18e92539fbd0ed92725403286bb7077f80fe94d17307d5f718a631ebd1874836280550f2320f46dca2725fa07fe576c58b7abd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67749064695339623a229e1d1bc0c89a6c8527a7464deb9372cf23670ffabf58c388b9ae96805545b3a51a47959599a63ef546bc9b288dea05ca1594df9ec59549c28756886492baa271f0f4f7a3d070cf2009fb2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57bd9ea92452e1fec3b7e85ef69d9f3b3bcb6b1c8747b2b5995474c5485fbcfa94ff71d7405575b75c75933e3a3091c8ee9939dad3050bc67461f859eac5b1ae34c26fde88a02be8e4f0cfd9c37a75e24647446f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h912ffe40cd017ccfa661eb585a76eca4c21c71b422ee1f8b720af46df5f09799df38ecc7cd779b2dd71fe269027e9d6ff7647937556d9052ae1147228b100c2a7a06435fe575239cf65a32af515fe3f47bc808535;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2868e092f6138f4583bab5f0f069d89b7a2486eac1e41bd97ddd231391eba5073c49ccdb14c466b73c3f2b9482bcbc6feaea40067b0c81f344013967b2e06599d447ea18d650c63821ea6d3787d7d0b0800ed8df3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96f023e82ae5a053a7266634ee035849ff5e78dad2d112969d7daabda2ffeef1f6bc61aaf773a8e3005169e098ce122e588f0777e524a0c9c8e7792aa88377e7e29af2116f4ad8c09a97966871b02bd8f7ecef707;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cb7a450ef7e94f53ef97e2f5a3fe22c003f64ccfba1380b7ec2512834f99135363f227185676ee15fad219e594cfc4d73eee301f272e976dc1e9c5954031035b968b43db4c584c632af1e657204ca64d76acce0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h246908163557e4ae9ba50dc4c93b0ea3cdae4636187283e00d8dcbf136297b51bb9650286a5fa83dec2a825321eb57361f924e60db65608c38e9891af7fdc8d684c6f5cb16c1b561c7142ff8ff0c14dd34bb27d6f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f4064df8c01691c7654eeddfdca4f278fab60d8705795ccb53028982d06fdc61c9274396d6d57fd40a2e8a9a65906fe53d1af911dbd7eb4f2ceca3eb65dd1c20f62b28d438e801d79895a17cfb4f6da087c8afa7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h426e2f1b7713ab0ed50686a171b7ac86f4e271e1c4b20218298d38a20288a6efd075b77abea7286637a2dbdd540cf2db84f4f396db09a00bd6579ea300a606d028494841c15741e96324bf30b4616f40ee3342135;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25bbfede99cf364c0f8d61e30f3c57b302a9b6a3c41405825d36feb2798afff193d6f2222b68cc8830c8973809d96b0809d81da4956037d96e93cc0f15a6f77103d7f6a4587ec0fa2a2f33b8195065dafce03acbd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c6d8985dc83bf40739b4e93db2e3e378453271abf14a3c32c7ca8e3e9d1c2d07ee8e2a51245dda3aa204ea1d4458e496d35362342a04b162a16ea6d3a2d294ae83533d53cbe77635ea405c6f01ccae2177ca06e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8473860f68480951b31caf499abf2de4e1e7427131c9aa3e768459509d8d9f5489ab1ecc827c1b459c1ec6038c96fa1d1efc46e647126078ea59db23690c41d0fa292a2437726e93c15907eaffa0bb21c86d0a262;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd086a186b6b5237624c838b6e00d45ff85391ce6929664480ea289b5b321ad45ecdf670e9297fd3af9d57c4f7f48cbc9263fd429fb6c757e487e70281a929e05291ad18c5b1be2ba3e8a5db2f3a698c7182c3b0e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12e3336b2b30ba7d43961358ddce899795746850c1c6824e43c54c2c1593beb55608d957f592028caf59efc6bf215dfb37ec949b1f1c9e05b16f8d27e3d0879fd1874435bf4a017808eec2d4c8f48a8da360028f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9f80c77391af9bd4ac4c231b809031e572ddee1a9b7c4168c939901f9f67ef886413956afe6bb3faa4d13b840c3fa98c9374dcfc25c36fbffad86f7dd052641af222d2e77d8d65b295a0a53fd93e8cea4676cc13;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a140efda893b78be4709a5aad95ba2dd8f833ea8541008bb13ea94c17d6fdb4555ce34cec7f34e74f59ea10182c98d1d5168524accb29c38aba14dcc4ab730e1f38504b0f86eab166e896229898571023790e027;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dc3f5689929930753f124b2a79c0caf1a434307efa8f12feda6473f2ade6004b3ab0dfe707e0a28c1c7500797fb50c34fd730fd8b0eaa6899287f172366fc735b1c3283c6a9c8db39f76cf07e279522fd1666b0c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6677afd461ad6a4bb696c6b90b477f28108ce8cef15d0f89f87ac111cd9eca1d73f12fca7ad7a9ad613c745c0150f7c64acc705463f4d73ff90d0dc37c71e760ad67968a47439cb7f9588a36af2f1759f16df8c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27bedf7d78085a6baca0c7e55f323ed39cfcf7a71a2aa7668215e862da9a99860e782c6484d1b46fb3fbd59d570e92a2edfda9de357938749026c20e3deeef1655e7241bdbb3b6c1f39a7244f3de1c410b63becfc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f1da5497b3bb2a0e23cd516c804d2bc7cc27405850028014c56ac6105b54dcb6275b411fd1a2d3b9f7f9d6aa2b615c7a477a27708979e708ee886033e4467e4365d9121167421e227aa994c0ac433e76cdb33c65;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd25b9f87ed806322e07441d26c8b12942f4692818585361840a9a89cb521470a0aa3f0373c3684502a330dd7594abf1c6e836372a197880216eb27e753246d37157da0338a0faf222c7cedfea1237618021ffa5c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5d830fe11e234aeadc0ffbc36b140b672a511db834c4dacedcd47b354440dbfdc91d9d87ace6b2e8ff278f9794a450932b8186d5c55cb5cae4199773cc6778c581326e84c4dd8d1482e28cc6ba47e0fee66963be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfc127f60b198c08a573748c7fd0ca88b4d66a1add11d5ba23cbe5cd155a61c4d903b292d9911842a2a2f3d181d842548bcafbe164a9f2f0799ca19ec7833b69750a7b393bacf437a096fb4e449b5aa072177bf4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b6ecc01740c6de070cbac5303aa56ed5c7eddd2d24883f19ffb1c0aafccc6d3860f8621ed55926e64322b9b236ce1855bc8d6f278454b9d1dea50869c620647432726d9cb091035ddcb95d3aac3cda4e9f6d1e0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd40aa60e585e3f320575c3a8d06bb59760337f84b40a59cb4faa412abd390df16771b6ceacd035f5debf61fdb88281dfb30687afb35bb12f0b8d6507735a34b7b4f136c75feeb8687e522ca404c62f16393e6518d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa547235b9777cc2465ad7e6c1e617dcbf54d7131f2739942d2ae2185033ae95229c917ad4793d5805a108210206b798678c348ff3e1fbc8a6585a766105e8471b35976b3ebf647694d66e4416df91378f19aae97;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7175b75fa4e7cb3f52c1308ad9d63573167e669654a11eba99e595d754acd424b5577009d6339fc6ad0c7976e7fffd106243d9d7b1932866952e9cb472f478693a911e498c2b5d3dda217ff5a84770f34ab04bc1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h379cebde865e19fc3d30c3b8692998c1910c3d8cf57c9230439bb03999ce130a57b4a0411b527ea7bfcdbe42f54c70123939d0947cb5c5c98e4e774687f729b525f17cd523214a48ff1bfea87e0a38244ba7cd04e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb170bd9ee7710822ecec5fb36776f1036e8e83927d9ebc59bc4bd57fd2851d0ea07ecf8d639f939039ab562b8593dd010800dc532b4d838055ed8518583034cdd6980f4961638adfba0216f736d123daf2c099edd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7af4721b635a6338383f776fcf2410cbb7b8c079d0361f5ece12ffdac534533e47c157ebc21d7dea2ac68a3cc159ade71c6d7cc08787f2e29eb7adbdbafc677dadc3231446987be04b1cde13e4383847af428b6b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b9f6c1d0fdd17d3f1fcf27e4e184a466a302dc0e532d41d581aac560dfd8e3030179cf0a477441ca77909b984261143bfde9296a9cc27102fa9f64e2e0fcbebca8127c47797729b4a2627ea591bae1be8e058409;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4d3d5a8476d6e10cf3f073ed37b18c4459a72daa0555c4f474a7e6aeb67d5d7eea6c4b21bb38bf1d00dfe79e5d1d0e10fe974a0580f81bd927ddf5416cd6da3936c998edd6fa9239ce9792afda1a9a47807170a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8230242b66d0dd64ad9c0ded428b208d000f21e836c991a81aa6883688811df84543f5b49f07b87ba04ace6b139f986b07b392165874fcc101645e528fc52e8062a66cb7496282ecbe8f1ca238d2bdaea1b9d9b43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b3f32d4d32c393b122356b7b6db26b128b9db61a804e8f5b62f8d20efbb7a26680ac830483286e7e50ff0f6e230107d5733a032082f904f9a22391fb9c24c58b1fc814d3367e42cbf71331b9669585cec281c6a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h824141ed494a26d4c21c173c2b59b7750f9842bfb5a0e7ab7ce3eb9ee990edb8f6dd7f3d6907ace133842aada55ef9cd89fc848a279f028afaa9ae48314260b642286a8e22d0893fde226b7eb43c879f53bb158b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6eb99c5528cce35fd6a3291094f4b8d028c2158b372a8519c711b93d489cf0007921f3f1d4aa1d61bbce80bc25ce9ff96f589c88954cb7fef79ac78e20fb9e68ac08fe0a8f289d19ffb01582fa7fdf54dc4a194a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc68f6dee4c6e686b093175f36d533d8207b9869cd1ad10ac0e9c37f7d472d39803942406dd324835e22a701aadc375b1c1c5f3db884e625f6d876bb630d1f671334d290bd780799004e46bb52cb94a0deeb2ff81;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb05147477c4c3b39b7c0ae086ac91884c50ae65ddb3444dec35085ae8d9868f181c761e63cff8727b0cea996f7d3c1d14aa82913874e3ef5c867291b54a1d6b5862b0df87956d74df70284648a0aceedfb8924f6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf682914fdad42216cfeedfa17c4fbbab1b096403f2a2f80581487d4c66ee1b110892e0f9724316e78783445f46f5cf347016481cd3bbef362a241a4eac11f2739d2641deb132a8113b908afa81684f1f9bb94a8e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81180f0d5edcb2247687c635ccce719a95e4a08c0af53b2fdd1dae8eab023cd8ca2a474441426839b1055f83d6b0fac25e0151cffeb48de7b90363e4b4440de719366bd681103be05a8a864a35a5e4e0e1f3c11ae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83d60f812791fe18be442bd5be1a0cafbc253b39bd8c29a74816f0d98153e8b5b9f80515f9f7d433c604bdae1b47cad56cd0ef7e34afb83ab2c355c3664a251b1fe6ab9536e1c9b9d64a733e16d9e0e462d859d3e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcab38b55776f3a785a99bb29289d276c2266adb4197608f02df47aa764da0dc1cfafefa48824a9dd6e28c6360a21d48ddf85492c2a2d267562105595c01e6d9b1324bdf5ebe395f3b19b27c1af5450492cf41b078;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c32c3dc0bf9af6ec559d3845b22df4115a31a7f903b95941e82c1d09219638bcbb461b74d1c652588656f946e17eaa6e61ba64ba5608e43cff98e046b081d272995127b47d7bd7728d7cb423e4bdbff4c61aa2dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddf92c667d8ce9f0a96f16a7a0f8247ff9c07ba16487e858813aee5bf4fa449883a6832da453081b1c17411ca1d5b67a0c434ae39c7e8af8428c24f7ae8ec1febcfe56a2f58e5d2edd15186238db4e640d7d1614a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f4d901144ada970ffbf37581a7a85c95f7a50568e9984ef40191ff7a671ccff29327e5ae650307c08ba577ba50ea555c6194bef42712d8f5e3436e3f81d0bd8b207854bd7890cb181b3c8cf4e3794715e37cc4a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h563a7e38412d226567cad67e1a22b84a430a5750ba17aeb67adecfe5d190b57eb8cef9f6d1e7b3e38d537721d2f0cb10e69869c29bad83d36fc9edb24c2de3bec648aed42f0feb72c932e7170d9bbf146e8820f22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ad4597a6f08beff8339715cb9fc54ad1e5e938f10f866a9419e7ea81e78d6a9fe0c84627647f879f1f86ae575b2236e8f65b0d3a7bad1fda1db271a5cdf631369c07db7676f47ecfd8264544ff307d17c740ac6d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58e18fa557f1e2231dd0aa8cdd65c0221dedffac04b66d7e065111295a7a531544450b29dca5cdb9c40cc51d97e525fd75349eb13e7f07a2bc544b18aed35fcd88d8f0c195c2343158c594ddf6fc65c32977fd8be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb874af5b45f4b44ca7f270b2cc33c9c3fb34fdb24d63a27e36e908f2714c554ffbfc8ea370b996294f4333547358640bacca86e41b4667e09e6fc5e02d146f2d365a00138aa83b3c63ba01082fcc1615a32ffd60d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58302f57c6cb748475c8aa6d9fc97323d25baa976a533639233de1044701b49b53fad6146a427fe296553f550384c7e92a773e7d7b0cc0756298cb0c98381fc7149869d9e5d3c6a0952ec10469f7051dbcdc5ce69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h258c97dfd07ce827950fe4044ce7a9301d300a35ee4d911015c7a57c813f7720bbb91160e956df14754ed5767015c1eea57a62cd45349491bf320ad38914ef6434f4672aff5764ed6ae81d4e5588fff1ed85994af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43619719ed34bc05313052f71cfd27279f7a9e26b01db986320b58e3d6cb5a66e67debdb16d361263da34681d8889fb8411639cddd3ff4e08ce24f03d309b22a49165e8eb49196a3c1f3a4e8f52fc5b5ce0691866;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h429aa565c26a6485f690441cac5dc8689e6934e5d49a8961f31dbe0fc7d035671dea03a84e2ba174c1311bcbba0a0b4ac55577a9a69660101090dfa421c3dbfdbc0beaac6a5e5cec5a36dc31cde61306de9ba23af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha19cc96702fab176985a84af1f899664e9cb0dfbc866b00a5e5b7b5705b9b09fdc2ff84c7bd3352ced18237cbddf69734ad572df515ac4b1a94499ea1cccd9dfac6f338d937e90b5dc40662b64a3c84d1d6ea811e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1606ade977b7ded85efc82478a45509ae758820dd5138d63c67a6e733bc3d5aa6df36040a2b8a94df59e1cb93dc418c1e1309ed3192dfd5a38381a09275d65460cab52f5efb5547108e6a8a98f89091c9f5dd4b54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d56b8f1aa390ecbb90a1fcaa02f044d0f91eea6bdd1ebae7a0d089693394aec8c66724a5ed2a2c530a15cad9f375cdd2c3b08aca0d75579137f38a87801d0a0d8647fc6f10fe623fbbb0ff9523975f556ff84eb1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd6bdf22b5b4b50ad61e2409e570bc58d5cf494c9e22ff183b860c9b19d8d292780cb2ce57fb980a135a373f4813878245efcde2941af3876564b3e178b475a667f2461275156043b27df2699ed90c3ed5fa9d7ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2dccdd198c62caa01eb1b2cbd54c7770694a6234eba681f3d98c7904a1c8c2489e74c8be54fdbc502cbf06c758c55bd5f423734d2ed995303bfb43e3aec3e9841b39eed48062f3f70393bcc5007d3a48b04a3e77;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2afacd1308f0cfd098fc6bcf6f3ef40c70b94da6d545a17d11574f745c79193de8440c407acb32f667db8c5c14e500e7f5f8c397d0fbb209ab014c1a12e271fc51da936310c53b1ffae5ddccb58463878e6b9472;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce70333a0dbf4b31be81f8cf7709e9e60a565aed36c8d34c11e31c568d299c56c25a8250a515cdf5f68410786e430062373fd57b33f5dc043b39faa794332485cb3dcd0e951933f84cc85500e788fc945a8cb9fe2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h810b17e5bc1d7bbebebd7480ca71f2d702cf979f4111ab5dfb7679bf80ce4ce3f1d6c1dd9bc440467b139402e34f805f414436ed10b3c428718d21fcd7c5b54974ef17486675ed0f0b67331a155a1ec80638adc29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb02af81aa1e424e545c54529191bfc8cd2680c4a125b17ccbbac2fc367ab0bb6771a7db33a34b73f6a372f5f03ea40fa829b85efdccda030001bced81b66138a2827b1c4743755910c86cca1debc83f768d3b278d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41e3a7e6899cb6bd440ccba59e67e0e01298dbb3ef3ec0a11ff483aeccd4048b163fa3468ec13a66296111bfd0e799c7141ffd5e7fbe22acd69e524e7d6bc03a2c7d756c5e82ffbd2cf52869e5984bd28b79ed790;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5278a8f513374760dd2556d85f513a48c7ff533b4503317a050f674b5579eceebff9bcb0c294f60a4a2fd82d5562599f6e0c4947f16cf0d944c396fc10b90f0c38789502c33924eb70f28526d9d356c7689252bf5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h498c4455683fdac975783a6c8d80d512bd3f7b9645f71b11fb234cc7ea452e97e7fece3bb689a628ce91b8695c664794400ad86f23a249235ddeb125180c1d8baf1946165259bff4ce04b9a0b27deda5cdffe9633;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3479bfebdbd4e6109b153a5dc0b046d40aa13a66d6b3ba190481ca5699a0deba405d5b57d3398c4506a2e6a724ba816389ae96f09bca40f2b0982f92ab3c3ffd8a75864a1a638db9cfd0838c88a82a29bcd7a2af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc09f9bc6e038a5830dddfc5911435a42ef4fa8d7be251ed6b5924804b877d7d3c6fd42ba9bcb7b86681f3e060bea7c647f35f25522f000e82e98abe5508f0862ea04b59be2e6cb4417aadee722b5366025ed5723c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14278230c28cdd2586eecb89162c18f923798bf3e08ccede8d9913c986f8586f3d0f8d8f8bb4dd475e73e854b1a54be7b538afd5104e86644629b74cebb9f0bfdb40cf2ab12724789e83fb6d845529ad58621e33d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf92bb9927af79d8a181548770f6d6d21c66fb77c2b7e168608304eee27cfc3c4bb767ba8669da1af579cba4b039dd5112907a32e6a0bf9f5701acd17f8f01ab2ca8fa10a246fab6d71f8f3e32201421b6e68660ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24c2589e2293594db09ac7e9aba0ed11592cd7a25620cdd4e4c9e7472b32ba735825961616ad1faf53f9901a6215ab2abc64d4788e427eefa5759f6f41d777079510bbd28b2043d3deb968d6bd387f977a2541978;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8332a1839f9aa6bef2abfc1f6d4f02a8cc64b1ef2a3c2876b76a7050777d08ec82770cfca100a9539d1c491843a356c0a0565db4ba639370bdf36206ea040e6da19d3af0800e5391d4fe5eb91490b447e74beedc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70e677dc1da267aaf62463d969603a140239621d7c297d2fbb181cc9bb621cf1aeb36ba693e634e8b99896cfb39133a8ba7aab26ad07fc3bbe937b76f9067039ba94d336e05cc7f8efe309e6843727a15af9ea57f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24029cd926a0d4d12cf55f45fe004bb2ca688c29ea0318f24a238bda5673a255568e8758aa632bfafc3e0bd3a680d1a71b9c03902c7592a911bfa0616502fe1fb29dac27a5a5883823ff745fe9419e83f31d5a69c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b5868d3ce22c0b1e0f309a76fa7769bf92f6274477fdd01b0790395efd6682b3a131729411ca3e7488db84443699cefb98b273109a4f940c3e86d41b9e654f7729d0500c6007c9d7797cad9a78118df746f03777;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h299f8ba3c725856621ba5d131de4b6234aed1febfda76443bfa5404f26a954194c337ce2a8dfba1f53dd3cbcbc47e26d627fdfe106c6c9583ac0bfc194bb21e3fe1901e8683c077431829c40d7a38cfb03febae9f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haceef06b0bf7e9bfe1f3954f7776263ed53a2e2b31ac375da32da4447db4e71a1395fce826d1b2df95215e640da3e1257e922ba70da5a548c789b5c841953f748d48cdc787634aedf28497b9a5dd668edb604bdc3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6af312853d5a604b2f964d137852d16d76ecca2fceb342454ec6b4d81ec8dcdea5bb342f9150875e1616ac4bdedc10668631da27d8620de84275554af33fcc048d74d8ab8dead4e135081b85ae176f858796afbf9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9242192ca5d020e2cd879a104935e36befa0ca43a4ff7d36d5467f814d512468b88447f19aab322228ce83abbf5f1b7f1581c1eb97eccda10eba001d7b84e43b200aff597386c39c5c3d5c18101ce828c80bf5787;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cac52519b7236716e89fe2c64d5e1ccc2759574f9363016c3fe436ae8fefb5202d77444df467c70d4c3c0fd6aa85778eb49195779321f36dc28366bd51a418394b2803c9a79e7b25c3e59163d5787087b1febfaf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h464677c28f7bd19285de0119ce0d55b745535deedcab5ca228eec5e71746ae65b54780fdae447c46c60f2c9277713c987840bffdba5b2cb37f1b6d527adc38f80fa395d443ae4d1c3ca97391f1fc5c3d184a29a98;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2ca2fefa9acbd733c3be6a659959149df76f8edc2abec8df554b26b35cffabf7359bece717f194cfc5e814adfd5f70238aeadbf1a3361ca67cf8355e504734eaf1f2bf3f42a64fc118fb94ca3c464e3d687e133;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec50f5ebfa9c401f6366112c6bb8240e1ac45d65ef5e1050bf3ee2bb133dbf929ec2f0ab5c4debc580c42bbe5a507e6c5d17b5c5775562f96e0f3f8a3f95eb366fc34d18243116d5087a8a679bdf257903a3f23fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h156ed7458015af7c98c565bcf31a84593c443358d4e16b53367cb5f7b63fbf43a4a66867379745789aa2b8101f43f8a0571f0488affc952b47d5543fe03840c283431bb5fe6723e2c259fea13a4a79d7ecbb6750e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf20fb452125e35645513d0441c1d2ac2e433c16aaa3278aafff59a21e97f155045090f5339536f7e5c259727c0621da4cc2447440a59a6d47643124dcb83d67f303057c15ce2cbcd7c0be5d791bc6accbd9910db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7a07dc71702e2aa27bdcd449e05690c5b5277375767724f5ebd4d30403221397c1729729cfcc8fc42baeeaaec31e35c9a21976dd0a0fd24e0c54aa8b75fcea89ef6224337972780166b5ca2173ff02abfedc9be9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24c1ccbe505fd02af3d479952725f42376df42f3d153de95b36ba36b94dcc2424f57d3ad72ce098f6f129c1c423b04b059285e3474aa3bbcefcbf28cfe00e48ef7b18e781c46ca16bd8daac1cb2e6e5a24f5c5866;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8a91e1aa5c8400c75f6d1105167c94440c6531262ea7a5885e2e7d3d8a478826e589fe822fa467f290dec8e55b6292f93c6808d1291c792684ed03adf40cecc74b61b9cd399056e353dc6b565f0b9baa377ce1d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51b29c2e182ca64a07daf4ed0b343db4d4e8ce49360f49dad49ed5df60abfff4f442a9e0e927b0d6fda923a8d6abaff8fa0a627c84363c03dd054c88e5e3da9f80717d23f6051190b3195c55f9caf449104b9d60e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60da5218ec3284c661cdb2382387f19db3dad02747fcecec7018a3a3cd9e7f8ca6540d546af82ccc091ab0025880355abad58fb557b3808cdc8b6eb84574d6a42ccbb85785e1b877cf769a47ea7b8e3874208eda2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2b247a60a261bea7a837a89e60d6db12efd586dcf12ff6904f53b17cd90c95818d3f76adf16cdfea4232d98bdc07f4a34688e304ac0ee25f342d2645cd958a9cbddb3a81ae5c9a18cae994570c4672b6e1e96f32;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6e86917c67ef9a3f68771ab08c1052f2547f5cd89209bcabb5fdb32406802db8bd4fa2b5c212db13b09e60b5584a955f474ec2a746a82974777a738c54e4d728e0464a006cc3a374a843ac9c035c2383004d37df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56cc81da03e59967344fd8883d9c8bfd68d77aed7ff481dc99dc2a086b33179097b6f8939b5ceac0d8f3766903781b5d5e62ee189807f39a6cf4b07aae43d9ffe7036c0d8345573362a0c103554e85499b1f39e43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99784cd5b9ccc207f4783b2b2ac7a98d9c61015d5c62a117edf5497c451a6c5af3cbef6352b079f44ed73ee4c332c5df8c760d5032e1d1e45305a7083af5839a5799ab59c798ec89df06c35290474670026fbaa97;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc280856c7cb8a8ef0e778b6414f5c8c643fce99b858f0c5494d7393bb56a7a4210c06c5fa8e02475623133532cf563d209def46cdcb07a48eabe190ddf908fdd613ed4e5747e06966ea5e0978f61090d20e62a39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h245dfbdf9d2c751922e9b06341080cc5453deeeb49e4288d83c622db25d4a74ec54cd4af35260f5cc86897de3769398b364f9156be878b5fc6b9c6b672f1a6e484a6253a394f5de1717d8831ce8c1737c1bc4fb8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5d951671e9e51cb2448e473313babc8e55f2156dd041236e2ce997bff085b4794d8b538a23332035350da591c4884dfec40376ce356a76b096c904ab11fc5687a72ff4211bc43e2c6eb3bc1af49143d732e63925;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h889580505dd07c30d60d1a044b8de0a46b1b8448aee7ef2d91d70e9bccd05d5239ffa5b0660196b4191cf0b0265edc078c3e938dfcc7d2b2a43f5bde8dc36d44a4b28ef3fc4fa55f39533adebb360a11d79b3ca86;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48dc4719359d0266d8fa929964066e840a4672820fa4a94a71b476476fd761d3b3ee0f8c912f7303736aae383bc1847b7408a07798eb840ce290e58b2aac07e420176e1cd22a61ae3c5244c1bbc1b887821c76a5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde75bd6becc5a949f5a2fc2d06a4d0a3fc2ab6b2b05da524c8a8e3ef58d301bacffc60687ab9fa07c688ed1d1e65e542dbf215500e62d88c7f41d31f8cc5d30956c07b42e43be213a9c016565dcf4f88c6982db6f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2da76cb24d306447b28d6ae1f2da3f48b72a846fdd87eda20ce4ef897962205724aff25c50cb13f97dd532410956f6f34ff8072d8626169cb78b96f43d0ba7afb52b0a5a667e2952caa67fe83485097aa41127155;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62844185b4c1a68c69d2cbcdd01352a7f52b991b5547b98a15d5aeb84043fbd743365ba6b43bfef68050aa9c18bd9b52e762d34141ac8fcb54b564f9fc826bbae065a300b8056c95fa23c6a0d6a73f9c2b08ccb8e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h518fb04303e28ccf8c3cf35e8518e1fea70d44fcd1250fb2fc292b1f6c3c0b69fe2b54336a455b3f8c2a61bcd9a28e81f28dcb3384120ac8e95c1b44a96aa95da5af3c78de9a6e419826ade357aa9584fff2fbc68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfee702a77af704b8bda4b3cbe419fe151024c6d845a7763dc5e215d62026b9db9c10a6ef081f7c671db9de6e6df627419aaf348a4d6024c126d20cd3336a976c19a63400e265f1e9ab3b6961af1f17adfae69d73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85de7e78f858bf70b7a01bb6bf4f6539920933d611fdfb242f7a317775fdbcd10dbe410701c5553d49835eb8eec28fe5cf6594035cfeb07e3e8b3e8ef249e54749cc407805887aa459d48e14098adb5123b56b7cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce32e4fa4ef860dc4e6fd67f9daee3ae8d310748f80909eacb88d3dd590305695a2e2d38e77ce9c2d6fde1808d940b0b63bf56b2860a60c41617d47648bed2b2bb8504a4fcd7b97a68866949e69a0e23b072a5fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66e4177d4558dddb4e697848e7a5f9bbc2d8e4d55b4fee9118d1cc5c6c07cf092853f6c2c5bb901d8970220dfcaf18f8fadda2b0e1d4f9ef00c9fb3a438183ea89fdb85747492dd3f1acf36659553beb437d73bfc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63fc7402bdcf7b4f7f028b4e831a73a8afdd6053f3e6a4112092990c26b22cee5f9f402b1d44a30d0f0cbfbcd6d909efe4a393179eda4aad1002d1a23bd70d5144e7f5b1346ac6d01598bd3cf14f30f0b032f3c9a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb46dae219b1890b4c2d3d034692a38886c9ac5d10c5b2e98d8ae2fea1f6a92f0dd0bd25950e35c79c78a4d58a4c1ca963c24231574abc5d07ecd158fd425a3404502241f66eeb6d72953b34dca9671eeff7eab27;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h613cccb82663c4a0a12ddf5d6b7bc6ef905862469e0fef980099710fc3ac940c4b50c4a582e1f57c13c933f5919ee4f0f05688a09d6c41c5a3c95e2782bac9db9317e3c22d25ee5434846ceee9b1cf9722db3dcb8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40e74d22f375ec1d3042e8082684ecbb541d8c2b0f1f52ed23d50bca0d5014d5d5d79444b989724e6abbeab98cbcdd03543f1ec8c36cbfd3856ef556b8dfcb05d54d5319eec252cdbe75a573b8f403ab7e8becbf6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c976c00889fced67d5576b7d47fbc86010b36b6f4c17ddfcff537fb36bf10da1e4ede856fee09806691ab8df3a12c1cf238cbbfac2d48f2e40d8ae5d8839d85babcb562ecf27a5323485e29d730653e2f4ce728c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5152d1a0d8cb3ad39ef8eb4801b94fc0760568a41cd03fe43bc6122377abaa445da3c6415e6b6f8444f2e1fe2377b488feff3e59542d80c1e3fbb00eabf0b1823645a58eeca441d1ab9ba3764b4f7fb20b0b9673e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd852d21476416f842b86663cd6003d33474e3e90e586936ec87e5be65ab75782d4e241c078e0c5fe831a900c6a3da35781bde9d0372c39d8675a322e9ab12d81e9b7199c85d95c6535a4a63af079775a2d3afa43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h435e41f63c43cc4ce851ebccd5b6feb02399ecf79982a0345d94c866860a2927f75d3b54f0ee9b9e62a7bc3e1b1f3799263de957856cc724caec44bb784db41f39106b1091bb9fc2bc4abd36afffe223ef9504fbf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf54eb74331d1c283d38be348c78b03ec65c4467b9b5a2c1d14d52f43bd6736f40d550b26cba72f6c37c773319951ea09c3c9cf76f7450bd1e47d1927435a5ecb941b3cb8ed5b145e1742c4e6eea7b04303cb5c22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcf83dd098bc9e1ebdc49d778c3a59f9b83f1a60992c5287d17a0761a751ab792d74428e76df37fa549d622ad5fd5c38d76737de0905cea298e48f40beb932b50b9486bffe5d95f372e99b3c2cfc8b5985b88941e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha85531835691db905ecc0f10a65ba53796fa666a55a91fe8dadc4bd73dda9c628faf83442a34e863ecd8264dac396a78c89e91e220be803178a8eb37e1fdbc73f10040a8d254bd8a6ca67997f76a86a0215584539;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1a5afc0d59cc54ba6fe13ddada66fdbd55770796e3b53f8f707dc63fc0a8e55a33f60e64bc77e9b1718382c5d22cc2f2b6a190b5cea8779a3749fbbf38d4409f6cd823f87bd4a8c93dd7545f84d13e847f1e54da;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbac233dfd5fdc4a52e5bd7a0e71bb4ed5872284c6aaa130ae77efed593ec419b7681d6b495a65eda8e97bf0b81c44b2d3d3875310b0a0c374d2a0aeca8173c78c275cde61dda2153fe1a74f17904db32cab50d9a8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79f8cac6c688172bce7f5e353a439032ed018dcfb60ee04957ca5e47ef526ed974c17e7ac1114e77eed6d2856d2a1939b7adc36ac4e443a330a1d2e5ddaeb7075735f9986f48d4f8987bb7735c9b8434e332b8304;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h756fa66c91d818a6be090b0fd58cae53ba35e60d6ed1f496b778462cdc24adafd9e49e70c6c44de73db423c928ac078ff926757a16099ab47ceee0987c9f43206c78c7100bf4d4b60b627d9a0d6d9af746a9ccf16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93ba3a5864c09c87942761b2d5b09555251b4f73e32259ae46c356b7f34c9230a831a6b1b04918dd8b3a658d31ede0d135d35e1b27f8d8593d3d6ab5ab3f27de320aebfd71d03b63bbb744ed326c223924e1cffe6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ea2fff54519e9acbd2d5d716629988c3fc8070b7a1b1865ab6345d43ee511e707f19ba010ddda999c7d912e54abcd8fd7d4c32795c24be5ef33c0855f2b517bf683bdf2a92094eddddea53138bbe9ab10e304d93;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e51afe6bab5c2899fcb92b7a2029d80f000da3fb4e62d40976aec46a87c41d5b2a6b9e410365014fba49e23ddcfe5e8b61654b62f1fa0e5d1e05ade6a86977a305ca6759b558bd2113b9659f906d184bc3ac8957;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdeca648e346449833498efe03754ec147a9863306b6859acc973ffb3a97e8dba8ae29724b7961bb8144b9e304abc2d4d4f0590c9e01c00c71d48826735b2c39fbeadb568a945ac97ed8764e3979cf5c33bef6b98f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab45262daf419ef9aae537d22e4869399a58c47541f50832cf2ed458019144d101482dd0b25778a3f5e9268da623b2d4dd229bf1c2735a5cff0a46b216bfa9528319d03f9536acef0e3d7138628b5ba3322e241c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21cc5cc86144a6699fb04ebf6d6528c705417eacc85b9fb4587a9af4213d2778b79ea9a1ee8d5ae3158653adb7c15eb5de50e63ef7c893db158496b6eff2d8301b2a08b5bbaf1e7c27c9913a4baf40b71e15e73a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9838b304752812d56368e52d479946aae3dd839f872e73511d0fbc4b459c80f6095789e7a58a5f254c8ab2f9466f667561b072ce088324357228539a245c51bc1ca11a6ef0595fc728361ca1fcb6c7985fb041dc7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfc9c9ff7eb3e5a1f7d166f974090fc639cc93323e15d33651d456b0a7389dff916ec6953eba4293117289e7b68693e96050d875c39c4826aa4e32ce37b147ea166f672b05452f72720d805e32fe71a297152af02;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11b2753190070e72cc64c5987d8e28f7347222cebaede180d847e39e45575a6d63d496f17a26a35e13f26bec030279c67a32a7c447f7225917b5eb1cc244feab15d24a2131e3fb3add30900a1045f02cb97b0dd9d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4760d9810d62bc5b3c910d87c03124b045b5baf71ff0d1e1826c388f8dda7d0f9f3f8be02fd02477bda3d592efd5ec657a34b7a7e5db6e5a05aa2e39b39934d8c054d84fa4003c1a4e25299313c0b3b88e6a8e90;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd660c9740f4e188a38898bb8f694c3f049e2b146ef059fc0bb908cc09620106ddb44775c00b6fec1a5f4d1a7db61cfea6243c0464463617dccd38b010b780bcb443a80229b7e2712773f14d6fcc3c71d049496e5f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf72b7ae2f2eddb7280abd831b652f64f92975c7c2c3d33ca0177887ac660eacc812ce2cf10f049e46c347507d3bd9024f4ce102f8338b2ebf3af13a5f4f5fe9e26befcd9050916c9786a873e9c2ebb79dc7d9b243;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he83af4e326766ee2e5ff9002eb887c4bb4788e293cf54e9e1a17d9b49ac58b033e535a442ae3c3892233ffbdfa1df16696fd7a3f9dc6541281325c016d0746a65362980113f9dbb1d66d7bddc2367f9cd49f5383b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7833de9d7437d4897b936c14f318c9aaec2675ae08b350587c6f7b3699e7c9c1b11f26f7ca0da2a2ea14f5948fb505556f47b54f52d4e8a3dddb205d404b816b506425141bc6dd678f01a2b5a98b52353a2549176;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd90666300cb0b91d32009cb49353ea1a691a9f918afbd0dfcdf9ea036d10c105ee026d9db47ba73f817d3c7029e8b8601a07339c2a3ee6aabf0227be5909f358caaca6bc7169de8d61927a6c6ae90c78e82c0a31c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9369a868698023c8496b39da70f61aa150259d1ce97fbd8baaade59df995f2247d77dc45e37119691807eb2c3b6147039316b187de06f178dc40dd4de8a34f5b94abf137b5423bb503cd0a3bcd45331fea79fe653;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79ec26fe1fb4182f898717cb0b90b82443626940de1da524a53ec95851b2bbc6fe863c672c83797bae88dde6d87be3c53f5334b8422c144851bd23c9e50bc785e0d62045dd45c837d62358260e8519fb390d4fb67;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba0dad8bae5848d878f17633d1a130401bd8d676f5acb16fab708a8faede257062d7bdbf74ddb25f37502c78e427f81e46e8f8ede7ffda76919dd62700f046edc9bad5f9a7aec00255b8d775aa1f89d54ece9c5af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58329507b808a53ec5ed7a07c07fc6d3a44605fa6077f88074db80bec4635c11e6f690323dd28c57dad144aa2a612c077695511b9c1d4b618b48ceeced8bc9971c8109cfd51b99ef049f80b77f9899e4ceb89e25;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4046c0f5f5c6926d84066abd9b0a94ae7e0432fac81f5919456e5a87ccd13c8744ce62c07bc541768a4444c61cfba7d45f0442206bcf44f0d79bcbf9f1679ac8524b6b5a0c46345c0e498e4d28d1a605d3ca6050e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde2399313e49dad11620bb5a0892f8e3289dfc4566d0acaec0ca3791272c31f5ce766825a0839017bef8dec3a38ad0d7e450b728b67efdabe50fb2081ed64e13d050a801faf2e01d544f5cb2240ba656a4e047e32;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6ba7a859f5a6d1fea44da1edc1925a1e4071ffe2be2faf34d540842bc7d59f47e5687074ec3d387d7bd00d468cbe9fc72fa54c19bb8f7ebfea55eb974daeda28e176650efff1372b47b9974d25bbaa2d0d8c40c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45fabeb2af8c381120767d8e6148f4bac276f8092494b897b0120b22ab77c4e98fcfbe0499a1534ad3287436f657e0fe8553eca58f172083cdd5af3a03513c3de7caa05c148c66c437c9993d55f8ef0013e6c6a16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf04dfe7ced916896210119d3a84dab19ffdf6dbbc4cf81bb061290043a53a5d377aaa926236c86ced5ef45df96f634ed0e9c22db8149e7f05dcf494a27a25999c38bc4196aadfff0697565bf5ae326ea2136c465f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5e6750a0040b3dac974bf6e5c5b3fe93b6eb115aa162839d6b5686f7e1af097cbc96a96b007cb42d793a47a19039fc0305a47d15bce468a9a1ca4b8e3a778a54e305234b0f1f43afefa2ed344840f8a8d3bf9f6d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32e73f2e4367b7fbd76a752e5640a559bff011da615b2ac0eacbbb74836d48bf2343b1c44c72ac525f749cf020da91bdff4fbd557053389b46c21f4ac6190df111d0a57f13ab3641ac55d010bda5b855d9ff56467;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57be62a019ae4023b8fefe845a4849129a68b1bb529fa3028ef2da10c546c30613e2ac621b8c9d6ba2f62f32610d196ddd3b01f1bed14328b19687f97f64e697784870d820fd8d479f2922389b8afdb1194c2f6c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c724007dfd0f9b1b3cf65c60acc634917ef7c6b0b413186f9e83e679e986b57b6cbba64b4078fb707090eafc8ae60a79d3b1a6b1e44a7e03a53a98b4d04dd8ae8130aab8b0d992ac23474355f3f76db2c0250a29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb531c4b010510b8d1221326906eb60d0e76a0fcdd0ca77656dfa8614a9f5b178a82a0f473c56cbe1aea4910a554ac9797ff31bdbe3a0fb60dcc9465ab9cde655c037d12e7f9b2bf7c55e170aae940fb8c44d16513;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haca03a4f26ec9f20331ec13e799c3a75ddb0178d4b0c3970991edad61f3d48640d53243586951970490d3aac96b71a1262ad61eb3da41a70b5f2f9c0f070dc8aadcd948a704d0099fe960f9a7afdb13511d2eb438;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7626c140a5c0720329a730b13612c9366b54ae23c63d20efc7abb94b38b5656934704964d03d2545e764f401780e4c6c175ae7566778a8773fffa41ea039ebd1d1ae89a3c7d1d3821b1b0c887ef81a68740cd435b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8376a9bf29d7f269b79e5a958069fd5bd25632f2b87663cdeaffce46bf152a546c1dd5406071f86ccc98980d3ea793dad60f6ec0463f01e6f9fbb2852c34076c2b1e12bbc4b552687d4f7cbddec465a70ce205b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h975f8e6539839ac4b90d53fc2e08f173e5c13a871fe00699325f3ffc9cfcd74a2036f7636b332b767325d2b2aae93f6e6804955a0a3adb694eb73e41237c5f3e602e8fd1b81c280786d2dfed5081047b5fec51f37;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff7a909cf2a09ca3cced0e60a06ef8a58c9290760a9de4831a12465a14f92320b5bd168c344c84d481ba80235ee2dd090db1975995b55e37230e8b087ad1653d2e593b5bf0b72d042163fbe5c2adb85a64a3c1cc8;
        #1
        $finish();
    end
endmodule
