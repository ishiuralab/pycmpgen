module testbench();
    reg [26:0] src0;
    reg [26:0] src1;
    reg [26:0] src2;
    reg [26:0] src3;
    reg [26:0] src4;
    reg [26:0] src5;
    reg [26:0] src6;
    reg [26:0] src7;
    reg [26:0] src8;
    reg [26:0] src9;
    reg [26:0] src10;
    reg [26:0] src11;
    reg [26:0] src12;
    reg [26:0] src13;
    reg [26:0] src14;
    reg [26:0] src15;
    reg [26:0] src16;
    reg [26:0] src17;
    reg [26:0] src18;
    reg [26:0] src19;
    reg [26:0] src20;
    reg [26:0] src21;
    reg [26:0] src22;
    reg [26:0] src23;
    reg [26:0] src24;
    reg [26:0] src25;
    reg [26:0] src26;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [31:0] srcsum;
    wire [31:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ef9a9439064bd75149ce85b10cc8c0ccb16b3e3e3122ff9cc4614719be3c842a2e958e99b07ec846be6bb7eb7966b1f0adc629a87f8591d3a1396e29472062706cc32f113ae13800a6b92fde9e5097c1d8bce8a9b3dd856fac536;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69b4df9e4837b6f165e594d1fe751cd1fc0ef4643d8ecfd8742c93737cba7cbcf6e0496ebf9f02979b84453c9874748515acdc3a95ffcc0614f3c729bb81b78496e13ed218a3d669711744cb39481406f2afc64e1bfaab0a0cefab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115f571a0d7e67e695928f336d7df26ff7135ce93dce7ad4ba1856e0bb66d043ba58efd12be1de3fd5becf1d9d0ae2aa8135c4b2c41a34708ca718670d5a7edaafd62e47a13e164f1f1e3386f322a27f4f4d11fbdd845f62b902bb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ce5e88d58485c8eba869b558d2936b72156d8778bc4aad3d78c72b61a2d82fe8a8db2f4aced459d9f908fd478cfdec40ee3c0b29c257e7062b3974b9501df58fb323c68d229aeabed5dc765212113e92a3d726b9e4cf48d4985b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1c6362a5fc2ece088d762e496d8c8531892bab41a6c8c4a3ec908d4eece4ff1a9e1dda1b410ce510b34ef10d8145663b768cc8b86b1a7dfac44aa643fad1b811ebb5a81601bf53b6d2af0f64ade08bee9cc6ef8b994301d134236;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72ccc0a255f396f7a67f04bc62568ac2687894282ac60c1b75690b74df9ba27f8a0a865d27bdc7ee6148dd607372d8a9e136e8fd48515804d9b01c74055efc5d540d5e89a35cf7e839e0d59b9c068a33337dce8201ae23d5a6d7cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2295f12c8e7ed47c3f68c34ed42e2cbd2c12e34a6603491361bfc6ebf3f7207f448527e46d32c97e3a57a913925743ba9fa0fe2f50bffe4be3a46aed8e494456c671c173be36c87acf0670ff7214d6eeecc10314c961f51017e225;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he83ed6d798c0b2aa9df001e1eac2e806b143f167523c34644b75d58d62d582abbb871a4632e7cf2cf0506ac013e604144cf7c4212bab14ab1ab3626e01c45204dcbd5c801a83d1c5b77e382b603e040188b889d415b1fb07899c87;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a99c98b1da4ebe72696e757f6827df2fd58c7bf60dc66f95400fd5467dcfdb6da4086767100cf1b5543ba8c68e6f0cacfc6be74c5c1dd5a407e83a19f8387147937110dcae73edc979d1161f5f5ab1d60388be22c4547769ebcfcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h703bb9d6b6eb31c702fe42e28da430e63ddc9f39b34694123d7b80ec723d00cf6456f628f43c801a55319815f78c6d32bb9252a4b63ddbf77f57c3ce798344ab5c3e9b05b0687db2a3f7bb28e5b3f1ffca26574bbc0d80e19a0d53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5f62f164d61a5e6f35e2994be25829cfb86f9c56d811f74147239a19dbf8372a7c08ed08b89bc034724d50a487a0b6a2a9e90f86c006514cb8d66556c5a51e288d1d725483aa9a0ca0d6befd40d81fc4ff838ef887d694e4cfd23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fd0fb91328fea9cb6e2b913944e854aa1158b8ad920475d7791bb7c2a7612adb5be8d7ad8da2ac808e18b213aaaacab652a5abf54815268548286c263a19e5aa7647a0820926ddf2cbae4f27bc09f40f6f47fad29840b48a2e4f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcfc6990a2ea002a1890ea52829f745569bcc86898702970998166dd4c7574e89242ebdea4f30c6af608a0d9aa5ababe0dca7897f6abdb5754b32dd7dc0fbe03f7f7687d0dfb81e6fff961d6ffde5a79f56b36bffde64f233bff35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18dec90afc2fec74c15580129638d332505ad6d13eb98bdf0d5432ee6dc46f3068c1f598dfed9c31e03f6baaee557a130a5b10bc2370fcecc169a16c02c6b7099b60087ac050509960c2e6adf79297ea7e122c22d95515dcda50b72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a22886be9ee51f1b9f6168c1918a9d3a211063c9b43d7e33dc2a54a86aeb9ab6871e3e3c3e154a16ddb51697e64d7ad8c3605655fbad97e44f7a8deafecde8480c3b662178591c80f37f5d3c18fedbeefc42882e241a4415f8684;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e18ee88e8364bec40619b11bf654e7e40ca245b808d23589ac20d448035e98c50052bd06c5975409668bd83a514827f36a404ea7987bfea8b6e506afd474858ae2eef643f5582bca67472b983ddb2d1a05a99af3837c75d504b302;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec4168a225b817a0bd328678ed8bf16d219218ef145fbe492a7ae309ca85a2e8ebd57e83973cd312237b26b188799bcac91f44c64779c3e461be026272e1a3b23e4148a807826a611f5516f895e6e041811cbee36ff21448ca26ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha7774ea80e10031eb5a3c019d1579da0956ff500acec682063ead0b133d6fd6c5608b9a18a5f1b760f0698b44efa96639fb0205f7650ae04f8ff69ed61ae9e1e12f4f65ac17d704209df5eb0b8b14502fd23e25f4c7d7996be33d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e1741dbaadaf66238abda1a0a88b8ae80e9b50d605b1f7827cad05645457a46d245112bd824c68d8d2326f27215e34e6dac7bcc3c3e8b6d8a9ff64614c36102ea131d7b564bf9e36d9ba1356b3168b3818e70cd689cee7b270ddd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121c478155455e487a2aba5987114086951770ec0eb5a43a09e470d23d152883d577ff1d4a81b8d9968ac432ae90ce378aad80750bdbb84d0fe2745f807db45258ca81f16e312c9c70db06f3c705806285f516697500fad9e1ec492;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14755d3796a728f8508cb814e93c099de6335f5304a224303327a003838ac2a5b8a8d0156fe0c18105dc5c9385b5306eebd739b4d293c9220ccd63d2968076a57adcb41c84afd03ebd1f8be1d700de2c0343cf810d354052a10ada9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h186802ced2bab09ad6e6957b4dad3ae6a7ffcdb17532c4ac8699e901b77836b712a64e6154a3cd8288794b23b0fb4bd4f97ca8c46b48d85e4c493cda13076f8c833e505742384b9fed7a2ac11f7d8c3a6b5f894fb004184dbce1e63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1816fe80937315b05af67e1249889fb41cbce7125e966ac6ddb2beaff108247fb24d8805d5c2fa68977ab77da8c68b49a0e995c78d1c5fd2fe1203dc87b437e98b86ceefd687ebbaabb1369e3eaa66505b6ca894dc428514b2fad35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h563676b327f4c16165b57c20af276722e4536d1478b912b0d0c1b0479fb114880636ede22e7a258a24d01c5a5972f3dbb9d92627fa63a6b33eec112c26c19dad02e519d6a7ce8e627f044e1ae5b403c02367b4499a2cdf60d09c1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d4f7a155042eb8c9c9274c20d4da6bec4483dc409a9051743d0d1ab37c50db4ba695f81df12ed445264795994d48ffffac6b028840e1c332f6929fbbf61cb1002415b208982ecc5f6c69c3b31479837bcbdb729b30ae9ee6c5e50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd9c8b0a255baeb833dd4b45790126a8ded55156eaf84cf1c9c9b5bbcbf8e7665635a77b8c49c5d7202939542e67108362df55108ce93f2c820483b1f57a247144d5168e8ee3aae6c857a3513896b7d554ac35062274c316ac18ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e144d7e761f0cc7dfd3b05aa98c12710d79fb21d5502d7d8e15c310ac54bac7e884e7614cfc6e3beda768b25b066a82d6093ecbd48181ff995db5ecf1b038b51900f48ad31e8e62e60b1992acd41dcaf3b548367ab4166b5f940;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c2ea1941fcacad768824a348767552fad9b71f853b43f20ad3c34387db01243259bfeeeb398c7adaa5862637fef88f1c6d8cfb07b73e097857e3b1008d95811c51f5fb60db1216b70f8b22ca072505d612df85dd7ccfd119ad15d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2da2d110c1bfcc4b73102eb01b4fcdd07a7d5e76ace8198c4e6af119e1b9ab862ff189139cc7668ca22b23595e9f5a9f6956b9ff6f7ec86055e979d3bdbb31f23be59c350fc3184291c34ce4b228cc3e861599837d98e7a882c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a913f1c1e36223dc1fae42ff148d85dc94e129b210ef037e9f0316c30bee0164851130aab47d254938f1e54bc7e97c6edb695197748635fae5a460fe2e920e6f49f9772527bb8e8f98206f5249ae9ebd236ca25877db00ddeef38d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h621f12fdb657f38db2de3a25a31227e24065a53df831dc2db7e3ac3c81d36235e3ad322d9ab78d6d8cc79b032aef9fd64affd0d8070c5b5e7e61a24ee1b0d2842ccf0f2af2e387f9345eb0130c1ffa3d28007aba9b4b11fcf3bce3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde5b1c7214ec2adda2109ea933bb7401e291b8c22ced00731b9f2d3b84866088513c47d6f2a87a66cf311d9bb3da3ad41cc96621f565bf83c22a71ea126e159ffe24ef301f1c5783025404a7456fdc11b6f5e27b0f67bb5dd356b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc67ab08aa63c38a3062bd9e34d9a6bd1942d386d0775ebdd16046c9092aed21b4f4ad29e49014bb05ce740bada77640a2e934cb7cf3617ddc04107bc96e6106d52e2aafeae89c0f0d01052b2f0c923d3efe71f45d922acc396932;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa54789690dbd1106bd3802ab34e71d749209121bd09adc8033e1803ad6bca03a04da3deaa0e9a565f98c45dd68ec211ae0c64583c6bbd0e896520154111f063ce4b3d81de4c2643e698567f7458c89b2e7642db1f3508183df500;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd040f65d04b3f3cca503c1920281af16c902cd1d2c8cd365b498dd676f889c55896fa09e6a2fe7cb0b35634a062fbf67bd815ddac51fb52c47a668d7ee767ea31c110b9962625c365bd5ddc7d3a29b93150019f51d93d5403774b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f982fa525c12ca2bf92d80746e76bed4f7041a1d47a7817950bfcfa80ca99c7ea11984b48efe562e0500ea9041956607819c27a33c02eaa049b59a142b7c3ec457ece7fd57f5e5508e7bdb02879e5b13c20754df3eedffe060792;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49ad76f19c3c2bac58ab2cd34f51f7e98cfa8d4a66e3fc8e00ca13591b67ae2c64d1bb23b9b74915f5814c4ff8fa8d0291d4237a67d7bbfc6f9cb00a142023f5cdb9ac51dcebbd18102085085dba461e5ea0943ec7a2a0ce1ba980;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbe75a977e00353af50449d1ab74d0136e7aa75bf1626f667562ca9ece6b43d985f60bf194e07f071c93fc8505d7e81106e5193b74db90b714bc6901b25bedcfa242d3632fb167be46d7adc983383ca7575d76bcbb94e0981f8a189;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a523f005c292cb3481c5f0848632047f15922b2a7b5d6b2758ccdc7579d084e7895e33a5dc72000ff20bc0321affa4c200e91255aca3576bebb8950c9bde82df6d317fe502408cacbf5a20c0b636fd47178f15d094224e9326b95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e0927a7cefe35ae1e1b04339f4573810de1fe7f39c5a8b216069ebfd99de9619c30d4f25f8647eeedb430f237903cff687d9c4544d7f6dd608badd5fc976156fbb05c2157a06aeeeb499d96099e2f1add909503aaea105d37a12d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14805fc65998d3dd4347ea8c84c01f299898cd24c90ad97e0c5fb63b7baea54dc9f10260646cf1fabb85f9bf26e1deb128519c475a62ace93770f2e3746cd2c82654b6f1c7ba38304ca255e74ff2c654e9e9a3a09869dc3c9b2c15d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1088a5f437bb424d933fd7897d2517a9c52afa7130cf6a576859012a282cb6cf2ed0a4f5b18e82a4cbb44a753166ba2a92f2c5478228035800c816311fc4d756edf9cf8d8929bb6f671f489858ea674624abed23cfb979b4f4a1cb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1df05a8371b3801fd83d491b36d450c6133fa2f8fb8359408d6f9e4c481935369a4385f92ee3adf832b9dedc418653a95527b12f77013d2c5e97046f4354c38b22fa01624f61fe08df8b31e96a694b47c95d381e0e206772ee6b81f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb23fd91291c379fd9fe2a1936bfdece0ce7ee824f16b8434e9d630cc66151371c723e262e360aaa0e8685e84012d4c1a371a7de777f73afec76ba48e14ba8242d2bb1043a06ab7406887d02bbaaf97c7486d5185432deb750e2568;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8444f0c6b3944c795445a542c3bedb37ec68cdf421203ed388cf1a182c98349b96ffbb16543972d187d79bc90aa21528703d04070bd3fe0e2689c055ba272af78ae5bc64a1fb663e78a9f71fd29fa9637f1407b387d9ee8ad143bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f9a929f6201d407c15622ec7231cd5205f4b9a4cd72934e96154e42461f70316b462f11c8c13793aae206bd6a76532c3b90573ccaacecfdc5d51f55b1f84f0adc146eb8dc417c782db257d60d800a26cb1c380f3507520429e5ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb8b4e4fabb259027dbc22719ff5a4df7878918e138d38731c66e432aabafe23f0ec3ec318f7dad3e4427d3efd50605816cdf267f525ef853aa09910371c6b25eb702e59e290e690598f274603dfa84d2f2729e6e026da0110d4208;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7d8b7b002f65be550bfcd45be14a7a9fa9974f007f47af8d06d359696430c8f11aa4a0f6f4e6abaf3eb8334c1ed076dfb27b179bf181ddd07fbb3fb84a1ce8c4e7f96dd90bd43beaed0f8ad9540cc25a04b19fc7ea00e583416d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e29105c6906195dbee265d9f47b463060455785a061dc2f35445bfe62f6cc4a8502ee4b723c1708d8f8c0db84d3ca45471a3b641411fd1a33aee20818cf8785720cfe7fe6a635512ce1c288f0422d83c418d000c716f1561aa91a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93ccd730caf80c66c468e6d80adde02cda9df0142a206ae5500d4e1107f83ee4f6d6107807a28cd9931d7081d8b845cb22a432b9c9e9af8555d91785ad26deba4455ebc6ec9dec5b3fec10b98e36c06f89e465eb3a65ee056d8d50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7122f68fa0ed2f8ca54cb5b381f8a9ae16b51e9da7b81a9d15a5496c648169703f9d0fe6925d0d1e14aa814f0d17901ae05bc082c6b6d080c4cd776c48adfdfcceaee1d8ec70673af2ec84518614b21022a62e6814f34c56bc6d54;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c59b9dcf705e824ff0ce8bb5fd859b2f0f256fe43fb66aba7204315ab89ab61d6384b836d83083247da9def9d70a31b0e790eb26d5f733d57285f09c2da70cb703e4e6651f0e64c4468c230cf005ceb9d7a6524afdfb965ea68d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a5009958d58d3416e91f8b4fa5e9f71d3275694defa8dc00b3d2f226a57f7371168854d15ead4181dd148c801a7ea280c36409f35a815b7e87f03a48afa318712330cb62262dda2bf3d3a1ba296f1070abd9ec8d06c8d430dffe4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115692dadc1eb8775bd983324bd6b43af6be2e438adb9e25c080c1984e7ce1f8c4aee06af20cbb54b2bb132a7d0fc2d3e60315577c85b3a2947780b3268d6a9302eb0912961ff098e814dba9881dd3590df1a7b8656ea7612a12fdf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ac338f24616c1264e657c2c729370e55b0eebd25512370c354d76eeb9dec3b1679d2443e7b62e2dc9ce134e5f43ee39eb8212c370f3d16f335d281f3bb701cc58581de7511172a1eabb025f60214971b9668559d5ccfe41796b01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5e41e84f1dd1cea4a1389213e554bbf0d27b0155bb02a4811bf06678405a3a1ce661cb7810796a2eca9b47f6178f536b9b4dd44fffe1da9c70289b937426307415787ab3ef546fec3b839912f36a4ef506cee9f59a820e1efb18c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h124795e09d3b4f611ff1560ab7395150a66d4e0d5e670dd3e4995a74b6ae3df123be683d4f638bfdee0e746a67e1a8dc1c54d9f15e85ab3656b84f6d1010c218e7c7b7ff181d4e9763d56f9d6c9ddfa78cd6040abc0aff238a78b66;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86388a456159120c8244822906a0d2d47059a59f1b1324fbe9ab7b69afc4a31202e15a101c31df2e7d8e9aea2b6bfec67833efc02b1992515b86b28fa9dfd7e8cad30cd3080d21f63821e99c5fa8a49cf3f20d53d0c18d6b9ab91e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e79646af65f224f9de896d5ee3f9bb4aeeaf1c5edf2479dceb90043a2889d8f2f7562066fe300173ebe99b38d3c122a565aaedb87fb919f6a524fdf74e3eb93b8e525d58483f64df6854670daefdb4033b7fd4a5edc544dd0cc96;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c5ac53ad8f8037ebf0f8d24258e1fa735c859f92291580b3d513cf84c03e16b843980e738c225ee637c416a01c81a43375abb5c321cf7f4230c4c307d36d593a7da021f8990de3f33d449b0c0f5e28c0a38283b581982050cdf93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda465e29a4dc8b995767fc9819573a39bf53d30217c837e1215221476dd2d005f3064079e06fe75a939de9927b6e45203b1deca07564d8d2311124d72dbdc00957ceb51fcb1ba79c10a5abb98509c392bdf90510614ec2e7e1b461;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c497869d9d02ce69d46aca76c95f7633af797451871e477adf1b63028fb293ef736b8a3ce75bbf1e1c855d059a8b3b36feb0005b67f151de8605cf6f0e05d95a1f6a459245f1670345baa0b53477fbf38cac03622f58e13b894b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb42944a647dda3fda193b26148e7a4c919166cfc9afa6a0de5fd3908d6a005824d54867913ff8edb0028b47002e035133a52d4b1e3267f68ecfd56b5ef9ea2a434c71688ad4cc459795ba7828ae2fcc3d17657ef65846954bf5103;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e9cfd1d6b1ff9d4dd24627bd48541fa5fa5b4edc8beb1bb6c464d1636649e61cea3f8fa5cb1c3bea36d4714b71caf965506e8cddeafd11d03edcf48a7c097085bdd807f6404085f14b82a7dd81f9d237e475eae39e86494d1ec597;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f0fdc3b758b72a38e394d82980ed298510069535a6fc755be9dd02ab756e8ccb7155b31e72f64a04b8bc6e0e65b79d2811ec6ca843fba9e1d876083dc24787e51e0b479912f0439eac0ff248c51285f8eed28b3fc476265974d986;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f21fa0e0bfafde2c3a0871ce90134ba18d378f94061e1c053f44d0520480d955f8e1abe8a3f1aa9d4a95f4f23f2c56a89b373333dc353a8f3b7dc8a10b24bf3036f1c144a4bb84ab84fd96a0e3daa280e30a239f3829ad09f008f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16629668b51de4edeb830ba2c8afe50af45a0034d8a7839feb573c2532b33f2142919453e2104d24dd15d62f5a8371332e8bdfc1dd7adf9fa888535c519c29dfe4bbeaea62f6dd1f29d42ccda1017f40f637542471a3ecd169a49a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90d8c18965a0992725c5c888e0facadfc0eafd9d1208e5b09f13df223a95de2753575391fcd02139aee763828e98f7d790a2ac66da41d57bb6affebf7ba1075e5b68a2852066f79322cdfa52adde8e7a08b1dc3f0d06ec8edddb53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d508e90f0160590953659eccd606cdeb28023bd861e95fc61948667d46eb3516e93383be26b67948a6a28abc6d3f3dc4cc73db8236cdc3ddc66ad4fb1929e6c17e3ceaf1cd33612636c9ad4202f6c1e00a4e68109d29194be82c85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed16097e6a0cb8cfe6c201820fd11465cfa0a9d8b9c115b8b13be3620d7cc7da9f0b052ec554af1037da335a72b730191b6b0cf79d67d2bad54d6cc5aadea00590fd1f683d2097a9625d5bb73f841c9bbaa1362d6d9bcff0cd0679;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8663b9d7f380d0536df7d5cc871c1d5bba905daeaa727fad79f7989e929b007a2ce873e2751f6811a21de616e36f296a7289dca79d5ea9e9725a5bdeafe627f168fc663068329c23279e3edef42fd7e444b4cbe97707dbb16c8526;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f692ac65da83251654a6090f8b60af6bc31c91c54deb62fb10fc3dfd8a8807b45399927f0f830361f9984c35b094666c972a631b42112bb38947e81919e932cedb1e04dee50eee985083a638a78dd8d2c1bac6ce3da7cd4e4a2b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16713deb6070ef48d1b3c113bc4d3fec03b9177038dc9e823ef2cb8ab80529927377e1a1b09e23c32d5b21b0ea0f59ddc75996b768db3908dd69bf744a9c8b5b1d201012ecb51f40ccc07b66019e3b48f5f2daa7fd413623d2c9116;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hea3270ca14ce3477a526d3fd58f9932251416889504b4f6e67fca2eed63c36b159d5aa8767779d3f2bb01aeed9621af8578c7603519a968f701f3f329b71f6535b9f4322c3a2838a4ee39373c5c35bdf19481ae917acc741f80dcf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff19ea40e2f0cf99dffba11d08edc573270972d636457e328df693b9a4d43be626afef55c1daf50cef676858a21f6bb5ba346ef671b319ea47732926b0644e95feafc5be453dd028db0577d7e29bc4177e664602aeaa386b51a838;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdcd1a3961162225909b69d660685d17def5661c64e2329fbb1a48fb1234ad6252c4b303c221557c36595689ff6c19e8b35c6ee644e63b5b755862017e501cd2c21b82e8a4c23d506f5cfc25c480fbc674df01789da810b3e4259cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5caa10e135e78dbcac04b4990bf4697eb165795177a652ab4c53e55978eaf45083d2b5b9bdc6f850a9e0fb5e96ebad24ab04de5ad82ae2400dad08834d6e000ac7efebb05f5b681d67bfd4f000ba4d1042f3a5075db60cd3d6dca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b52eedc27ed24b91bd7f596048008ad5a6244fcc1978b6b0af016430356ff23ccd40786847c0a6671c2d3d52ff83767508c3841246d1a447136916b400d860fd2debe639f02e9225c47feb1ad1f4e738b768c1e178de216ccd2d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136383d24048e39b625e5c7efd918b70126caf269f5d17059be76648522ce178682c6ce754014038c4a41adf799c9b5fc5887a989657e0d9bf81a7c08b9775b5e149ff170f3aa21926919491ef761483d682630a5a33a2f42953e93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3403a1ea19033dba3758637d3012efa033a13e300e53a78051fd3cd2c31ac212fc93649f1c7ace430c1df5c96cf3b2e144ab8fe16ada7e0e250a25bc0af2f0233faf54bffbb03b72754328abf9b8ef97cac98dcab986db0a65eec8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed134e2e70ff2fc30965e1f4502bf72f673d42224c80a79a8bbd8ac349d47c0e23af27562aab3587718e6f5ab70205d6b5999112a6395d76111d6011e2c7e46a62c7668d4fc476528ab919fc4b9f12762568d595b5901a1eb2d282;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ccea3fd78da742732d02fbf492822c3fbbdaa19680ef825c1a48e85fafc57a7583975d8ada45fabbc1a76f148a5f44f26ccd0d11e1e3e6432018781af65a8906b838bbef366130b3fb58e5092a85fae1157998bd2167babaab33b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd059ac692c19b7d60a2c2c2b09bcbf338c785d099a28c07d788f036d24619e71108cec19db6d22976bda2ae8909e77815a2465d8be093d46b4e2aed9d5aeb5d5a6a9c89ff7888d13384b460d43febf21d404400cd02660a21cd3c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0be86e4bcb124e5d0615312331d8c2be5fb7788a1dae08ea9aa0af7aebb1672ec72a59096434d0941b8951bf20b3d504d04cfdc1e3f0f74471e2f901ab42cf40e32da839e975cb3ed1ab44350d577270c0f7e7ea2193a5b2b9468;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0cec4bbb6213a6190158aa6c6115f27eab7fadfe60ea149ca11d367f790b688e59cd417cb5602157f85318338cd1ff5231ec1563979eff75b8c8cb1a7c6a96f554d405d7d08ddafc0087b3a799d1c10ffcf73200c04cc1ee1dd98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h120a7e0a5745ce61cb8fc69f310deec5c0909dff89e71efc06c22cec8d74bdf055af97c58e2a836394d5118e9b314f61cd43d0c3dfd17a07337daabebf86c1b418705224f47a275489526c6d24ce78f6ca3f69093910bf0fc0ffd46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d49a53b6706a5711cb44d62a7b1a98928c0d61c20d2c4ee85c053520e77be11756c2f46f9f5401203199e3d3518cc8ad54f59071b0b9559c295648e64090bdf138ea19be37a34b2dc13e0b69c677696d737d5fac09e37ff8a726e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d0432fe8904fa50b3c2647d396efbdb10c8dd91db060737d5892341ef3d13586ef368ce4c19b3764f35d4e9bc7ce76a5ab5eaf238cfb21fa9ab157d6558ef1cf0ec738429355b360129380ab5f559d8592d84d1a9a6d04f212790;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3dd186a16ae82eb960b5a29439356d76eae6ff1b1f7b4087c1302e30abc703d00386ad54db52cdb891b41ded54c69182fe52706a426c2a4707917a6f347661f1f551a74adcd36afc5bec83434ce7773997e8941cad531fc5dc5b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a50093c6f218cd30181abf34d491bac88d7363b85ed6d169efa0155214ca8cc22eb786ea8bfd2c5b3b3cb133aeaca4d89e22b829fa41a54590fd9491b9b0c90baa9568996ecfd420aa92b2ced0a8483a08f3d16dbe7c5086e7a66;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfbf302fa26952d8d79f5c9ac56018c7f63088e89c4ec1e00074db69d50b9b120a25b08357994615a757191ac2e98b492444548590d936793d8a9bde64d05df4016edc4867070be1db95daa2dc23a21024cf5b005d8b986bc8cda40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1896f569b77784b8621f4bc60d687f9015bfb6ab4416e0a1641e934940d8023b8d3d4722744b52ffa06bc61bd3c692c9d5841a2f5ed43acec8ff2dd41a686f788f4f9b8f59f00706ca4010d8e06e727fd01d68563c672fbaffa1f2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hac7b74fff2101a60abb5abe5cf702d9dd1d96d818c7aed257ddf512d03f15515261b81e4f41770dd65905070bce2105daada8e3a18a1a62348bfe2306936de8b63cb0b08b441767bd4b6413417cc3ab5cd241cfa3b7007eb19d6a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20b3a43b6b603556422f6e00ae5b71c06e8c0b393eec3148b542cc8ab13e02cddbb463451e7fe997545e32d79a63d66956875cda7b797f0e397eb05c636189daa380f10337b7c0e6d68bfc0d07decc6a2f02efed31a39742c3af6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126020876d2b7c00fff969586d7bada6507f993f22cfd53058115dc5c360230d2a5870c36209ef626fa98c30b3bf49fc5a4eca4095160727ad97beaaad001638553aba45f3398e664490f017136b8436d4d6f2ffe2ba7941d73c749;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h117ff61e23ab364d020bc0f15b29bfbf6ae5383390fdabbdce63797840a93742a832d19933872d92f33c4b66c07f30bcf68416d90bb5191759c22ab73808377335743d87381ead8c8bb42578289f04991ea3a8ac4b17fe9527ae199;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h625861b2e4a4c88ed98512d144a5cb80af6aa785d9afc58383e48817d6d3c9847dfda18e96e4231b10b0ccc4c19beb9e412d1fb263c8754e08eb9c4dfe2a362463d776c017a74253e9780d7fa557ad7ac9a1dd65440ab2d574a18a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fa66fdf447dedf930f82d9c4f094437da5c26be6b51868e94bf237ca2350b4a76541f041d2713bf3ede16fe3f083bbe90d825b64278b8ee92875ab4200dfb64a0c8a14dffc6b2fb669f533ffc28e2dc78b9a4ce01a01f87ec4314;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0b1aaedd0c353fc6e30699b493f790d0ae60f78114bb6dfed626d726bfcfb9f7a544982afa5a39523ac3f032c25fbb158eed7e54848af3052250361e986f36fb9b1d234c1bebf9f3dc0a82047f3e0c1ce74ed741a7306a611a875;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ff80bd6245d29d72caadec0525a238576afb71c9f01844472fc887b39272a8e65f41f4d89b237f35d64a654859eb5d1b1f39c97aea8780d87c86b519d00fa1b77e71e04b01d3bd2f47c6e36574939212a02c6335886a70102ba7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab542022013f5198ce9c531e6dc00c63567bc224e18d6e4e88fc58939d9ab2b95fe5a32ba6ad98f3d5cddd473c3bc554427cdd37a87becbab7f7d44b967efab873ce8b8b55be4eb4079c0ad903bb738402ab012e2c1746ac950849;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h978c41328bbfeb099bfa724d3f0f9f296f2da9a4fe54ce2f8776a387018def145a70522e468ab0480480b4d1ebccc4116d2a8ac43696703f0d8459ec7cd4999794d611ccf4b2fe263274c16ea5d841534dc005930fa8695c212cf0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ccbbdc02b3c2c10ee6e900b348cb99862851bbdd1651febbaf7cd593cfdf83351d80f21816f69104283b7a2c1c99c26e4e7c96816c80ce465f6ed02763f08b7170742eaa788de22e39013ad110ffcbbb2ea23dc573389d0e07266;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc49c870b43f5b28087b3d3a415124afc985d9d740a18879bc8a066ab141299809b8abc3d332c6027b03e72e2e4459414093d28f9c4dd86a2ec8fad05a93dd19f607b10f7da686634996950634ecc952f36cc3ae8b45172f1d7440b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a6cd728fb31122ee67d3a7b61e65833abb2ffb75b2b1097d96eb1ba04d3cc0115898b0d367ba3b132525db1bbf6ce02cd6f45411ad4820da67c91ca508965d13de41059b3471429813a16dff487c59432d26b639c03703ec0dd01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h141350179a53a68c0918147bd087829c0d4aa2d9eaa81a40ba03d4bffe6e3ae3c30cad9916fc7b4ba2f470e6858d996f3e0fdbecb14f78dbe2706ba36fc3c404ddd1931d082f62b9db64e014814165cca5aa8f57e04998917cba64f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h77daff736d41ab95c3b7af24557d3b27510426d8f5b7934b150e86c93efc2e0c8f89fcd7c506e28c453c251abec6d91d3e86a42eaf84f0ddf2fbe183222672577164e7f9ea3aa08f3bb44c085b17020fef8a33a15c5439a45fa318;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193c0ebdb2a6deac39ef3a38bd37b68b8512fcd8aef2fe4d31ed772bf0b6a62a24a38da005bbd8a82ef4fd0a5e0787302afce3bfd2200f0d8d093096aebca0ebab6b6052e127fd165292941df410c85f5fc456330fd6c311d4d1b94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6685f0a5d5f0fe9276b1b18daade58605b632383252a50f7be4b17db5623cce63b947e3ae463da6c387e95be32bd5d1e4d2bcee5026b413ba54a34e50141008301bfc47fed19cf72880e7dbe4d4d47c88f858405e427bc4e953d4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107000380b02ed2f53278e590616ab540f93427976a5d23ceb257cbe48cbaeb62d06b15e41b642384a266349e7d5245460edfcc0317cc55f8368068e93af8fe4609765ed4c4f0361e11afbf47be863eb8bef50a1cb1743cdfb9ba24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f17537e38c957faabb9cd5ab122b3ccee5ee46776484b22f0c76abe6388e5ce696719322e856d852837355b80b0bb39a70797f977e7f17bce5504eb3d55e041fca9af7c92bd4deca53b2d47d43faacbca86c9478a2870eeb4baf80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24f8679b7078f6a27c2be3967a04b79a2076d50c672a37536400f6b6a9d6c2a5a241ea855d022ee199186061c732ba22a625c9b8e3529c599b67af0643058df7466f65d5af3a0fa9589fa2ce1c61409a599a75fb93bee37e713899;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1755ac8d90ebdeb43d9497baa6089bd48e051b3f2148142c5c48249fa14cc278507b22c5c2f79b988b62dfeb363fb1d90925980e622584a383166ce0e6ceac7fd8a1680a774f35cc7575b9c63bb7afdf41456445672ee65eeadf684;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h642a3132cea505fe54203e36b97f3ddae6e241212e399dd188d5d59012742926975f50961e50e3d338694595542fa41d89027b0ccafa8ae5adc91020fd2732f8c0b1cd1815aa704309c316b7d7ab7cadd020cbfd3d94b65515ec0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4787a8c1d8bf1336ac93ca3b3b0d53548e047a7cba4c3eb449d7be11d976c965060a2cb65cf8f0d8e0835c971fff334e1bff386df68ef9f192600a6f4673ffe4fa1b62b93058e267de3f80d48da88424e5346e0c22b768dc92b978;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2b1eb41c7d050c40d8a151c6aae7501405f50485d1e8d2fa39fa69d5872fc49782038cc3be271ff37db97b139c2e7a028488f63bf395129a32805b1ebf5a66e66e28616daf52a022cd3ac4a78dd68e24c87a630babe9ed1d210cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1557500124304e74f7de76ce85b26f33a24d29fb0136233a364f1af3bb561a42a176f96577db499ab1c4d20aa9c09c2823bfbd69bfef4c39e9f46f5194c6f86cb2484d220fcbc205c0599fefb9e95273aa53ad2f546887fa74d471;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e8e07e78d6c17a1f92cccb838f8646a199b91b97c18b385d1abf7865cd2f89d4931c8d20a3ded62c9be5ce9cbcdcdd0e63c9674b07889dcdd38a4a7d09e43e59cec48401d33e316dd9fc9b0b9852e242d1bb2c6af39b4a38179e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha70b8c33eff3e9614d0f6dd72916af5d160012c669714197ae529e08582ba7510be70e43228cc466455189dc3ed2972a701cf6b9ca896d15a8dbc6688829d6451096f4ad92c1dcf20f7223af358387e75ea42cc2ec079341feabc3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13050b85d648511e8eaa0a2a1da130e38eae6b787b0536762b4679e6a23619cb58f6483b5ff47a39e3cfc42692eedef227d5ff721953f7f3fde098e45a25dfca699fbf1e7b052462e4b152ba6429a8bde1977550224a1ce605dddf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ecf9b522933177a47e5881763ba5e48548e7f3d7b978b4e328edcd990646237d8e7477e82b5a97e6f0f03d32bbbc69f8342b66877a456f5bb96be1499025a50dd326045b376590ee8f049a74a9a48baf6fce678e51918f7415307b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a5e05884791d7ddaebc297443c12c8767006c53357475b8d1e99e22c4d78d8e44bfa00415a0ae5a691abf5905978c3355713bea759121ade7265674fa4955a6831bd3b0faa5b9060cd40141bc1262926e0451eb1663eb5768124a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb2dcbb8f4e4f2da9fd3fe836bf038fa18b5b606f0fef8a8947a0d0477787b0a32fd2402d0f2d23db3bf3b620373858a5e13ba1e4c513ee8381b3165b74ca980d4bc29f89172825a223056eac598952802e7b27f3b7f4f5f21b659;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c943f223e3ca3e346327ea38183ee674a35dda2d3ffc8f2de0b95b59d8f4687775687b2083961c01f5cae0b6eee265edcba05ce0ab525d9edf0d9b6ac945d156be9884f9d42bfaa869c07d018b56ffd07649bf6d3fc47b2d07925;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34b3582064dca1527eee846ca12255571024241759db0a3c5d64dcd9e1f7790393346fa8054f7bd84e3964ca853f89e2f19673f236ce0b276d63bb94c4983107eff14c2bb64974d65125ec9dd92259ca6ea16a09667c6d7ff7ce41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31fca271f5cdccc338511a2f7b66b04b49483b2dedb6d8cf2256732bb7a569975560f734c79582f81f89a79df6fd971c7a43f44ae20d5d336776dfe6fa5b8cb5774b862c1fa8e99d696c8ba84bb3fe564c61e3c99fa8e7a758e096;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9a9a333155fcd74513f199f02c58a7421b38e116df920a29b9ebbf7dd77013cd44e5a20019a50b1a239234dda0ef42d558ecd0914f48b6ad761494f25e4ca647c0c6900b883b72f3f3dfcfa886ac816b0b31dbbe6f2a7dcd95f2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h645c85a76363b86676c1fcfa1e4db0e0a0cdb900669c7cb998395268a279d610d9767753eb0f68e8b3f0cfbd491f688feae2bd7545036be363464b53ff7e4158776fe8c5b6f1d436fc519c90d789cae00767c3bcf78bccdabc80ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c40e3701d568178ecbc701544ff5847139af9b984c57a5f175c01772451f1fcca77c5fb1a3e260e8d8e39a4014612d0419f2e34a362bb4f5523ae02a5e5af7c0560d4cea72818645a25b1f484872bf40dfbc1cc9ca04d8e6fcd009;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbf0095bf2bd3ddaf9c70a650c028ce4c42859275baedacb0137d85f77dcdbeb97230c82855ad49e5a6ff27f8fc85def0fb49aa55ed5a70248a7911abe6accd6acb61cc8dcdc3a1231b6dbfa8202ade70abfb24cd8cf41283e861b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h60d9cf49a08ec6cfea202a4cdeffb896031af0f28cd4dc02b185cbc5ee8dbe4302cf2ef3cdcafb588056b022f9915bbfdc156222662e54d1ba60cb866f5aed514e32db2e9759f55f7d028a95fa4fd23b0f3c0733947c4046dbd002;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h163d452acea31200a9ea3bbabd33d43fb2b17b276d4caf16b5ba467921b784bbdc5ee13e7fbcc1affd0870ed6de3248d999d4da03463a4ba197f92ddd7a1da30d181dd9081a7be1ef148bca82a766a05110e356ecf5e62d86936eea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b017a90ea224fecedf64582a177a5b784c5db9b277aa19c0fda7109e6f76898a3ac7e70703a0077890b786b03ec9e9914f546838073c8446fe010a66fbd5cfd404287adb44b13b30a213fd88ef034ea1b151a8c3001ce0b25bacb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8fc0d70c3b900fb2507684042e0f3d50b356d33f0dc7b98e37a4c7030cfb01b6211e3fbd2831738158f39c90abe8b9c85c08c8f6ad2555742a1d21c1d9fe45cade43623f508c758fa13bcd563ee8ddac050d151c92b1c92705951;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f39408bbd647390de07d78c287d03f2250a7f4b9cb86d687a226c095ed65ff8bc2f0d75530569a0a51af9e26f059606ddfcbcc9e708850a509ef429d302ee1a497fb1cf3629e1a371a6af95b6b3f1b4e7fca81a1fa9d9bad821b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d1559aca98137fa2ef59275191e3a2dc86cf3677cf9fb2bdff475923bb086a18a7880943192812cb6fef0cd94bc4bf7a26ee570e395734a7788b9384604f472e93a6748ec5f5f0471b3745cf42bccc0ba0392061bc4925e4e2b167;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25221fa45677461e0246f5275a1c41bbb5b9a5421995ef171341cd8b825d4eb9afb6cf3a7dac4bd40f1fd33964e7706f21aadb0ca7a0695c92051d7e3c2a851b3de8db051b47c29ec696169464819a3ec185838ce6a89070231578;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18201f03c25fbf8bab44331ddc4efb08447bef7e845c19fcee6483fdcdc73e8205494c148a85c0122b17bc9ee6a3a9d076a4510c319cb863181c49222a9f96884e1308058f0d0e221da260575d610f6b60802722145fa290f0a62db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc3ac81b1875ac934e7b42bf06b17b45a8813fe329fbcd64c2ca7f7cffaada13d8276eb4d0ab75a7e1671c200e967f3f5c7c07d393672bc9286564b3a86b2e898814d37e13c91e22e0803e652c3ba47c0092048aac7db534d58703;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1449d3daa846a86781e4f5d852fa881576a9950aa7a3084bde0286b9000b1588926d95c5f74edb004a05a9cdf6d559c351559fed792f30d45bdd2343bb7957e4654ba35e109e637e95d5ec1e446a6911db0185efd12333369f5aace;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9552d1ccaf9844dca30ea46805eef5433dca9e1308cdc49741a07045484d0716ff34fa01539901e45601e34e75169423f8c93873901002846fe7bd917a76cb78c7783428d208b95dce94c0a718d31a159a285b83de4acb3555ee09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cef4740e0d52ffd33ef63505e79b99af11ce11da6ff94bbba46df26dc540f20e565ac3280f0ac11db766817e55b157aacdb101f13f4bf74468f4870819eb64bdb919710b8731df313ecff131bf2c6d4d6fcc0fee1674c2b9a6ed8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1d4868f9589dd6c03b69c44d29707475b463a9e5139f959147c4845bbb3d9eae68f1b21e15a71dc9ad55d30f5939ea6137f79f87f6d43d2e1c005f00c01d3a0191d58c2620cb234a0712af909ff40712f03a774b0710d10de4683;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12576a8b005a952bddfe240be28087582be070b18ad9f5806a0a99378f0cb8e31597279cd32f5caba3b11ddbe375e9b8fb6a59c70fc8e956c8dd731f93cec6d5424cd91e2df601c29fa23b5af9640168bd60b241b9e854a8872622;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6f8dcd518a75f2254c56ad5393bf527ebaa4911d6adeac4d748960443ec114407c4465cb9ec99cc0d4e4f19b1cd49c8df7150a75915ddbfb65c86b16bdbf083572fedc7244e1142fb0f842947d80db1982a4b3f893c3c8a3d0dcb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122cde74f4fc7be85fcaf7743e3a32eab595e19a973c0e78cf7c008dd1fb31ad7e3f6931e908dafd689b3b466d61d374e731522bd196a0c8992cfaebdc95fd18c4f9ecb9b00092ab875ee9b2424288055bba965bc367f777c35d95b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbaace38e7b4d30ceb95009f37c4c56ab52d50bfb2199255b11a711209c4e0f5e5fe8abaae2425aba367a494397d1e7985f0bbf5e409f6d3689de63f86a43cca37285955096d3e9aa5ab5619af1b97019c33f3ca7aea5d42b9a9492;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0d225bf67d9ba232cd1db1d09e2834e68c751492380c6d9745a23e255f2f11966951eba769f026aab146ad410716c7d5c575ad0c5161e122333260e24e60a674807d68f44b8b51f46e14eb9e17da583af9ef4bd017a4a597f8110;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd478fb428ed4295a22f12356b9fc1e80fcb5ca7593fe3ad48070ea83dd3a06a4cfabf01864ba1afda3848cd34e4468d5df3c6a020eed5bea78864cbce207b3aa309324cc19df077a1bf32794357ac9abb56a1cda2eabde18b6533;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169f1b5cef9ee423982484eb8fca411a4c80db2457afba42d35a417f1666e3516799e391ed992be73449794bee60268befd24fb1cda6cb36618c8886d5a33858765f7be9a60209974e0319323553f77d8390f4a80562ded111f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86a84f45f7ab75f3f5c98f40543eda1fa1e3628650e6de1dc11485ec8344f2894a2af60eb25458fefef5d75cfdca19068da2ba5b0f077a4228fdadb24456c70653a156e7c802e0c829dc2e345490f56ca7fa5683f9d48d0d8f1ae6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d1bfb606873cf7489908538aafb94588cb122748609f74957980438016e6046264766c5bf9dd074c342028a1db99fa1a3238c785851e8fe930036e4f63bd689eb736c548948669cc7a3e989fd1e1e8de8ac6a2733397bc397182c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5784c7cd532f61686de7711ca674211c3e7eceab7e68bb7b5fdc44ccf4a0f2b9bc86173834a8daad46dc67084d3d86fcca5c6bc2deedaf709377dfb94665bd0b111147252d13b09809df8cb9d8fe054e67b32640cfd9ca9c1c5eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f937fc871d28e136684f76bc4ef87fac73c76b46a7287fd0efd782d0fd5ab71322647d9e99b64fba593427de4ef507d25f815e3c08ec01e73895313230184f83a07a03534913cd3e61ea18c410bc49a2d8c2e50c49f9e08be168b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ddaafbe41c023ad89a7677e602f6414356a8237d7f6da95e81cdbf5d715d465386cb98c7cfa0b42bae14537ad3cfe8bf4f92bb4878c2a9afc2cf4f6c2094c67a16a3f671837c6b03dc7e0cab8f0d9130c9dfa13065339b9f9f0c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdbc8a7ed065897d323ffcbf492a4c0945378fbb362e5ff19cc11eabaa5ea1bb5d49e2e4634b1ecf687a3cfb1a489f48ff5df5a4492dd85ee776c79353d4787d052f203bdebe27aaf33583965fc9da4060f54905a5655917ab24750;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72f83cb325a42510351c9bac4ff4a64aed1da4b991429212a9c9910f80e617f933a26478bc957e79adc74272ffb98428448a3c157cceedbcccebd5c5b4adf6df09e3656b0f5406284135efde9110900a8f86d8404486cb8b5d9a68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfcb41c1050a62c96941ae763a8db776a7ae3805f206f67386e3e2e0d99a795b8e611beebdde49b9da0f05ab901e48947a0c042d3d6bb0fb8ea8a19cc73332ff6085ca8c0ceb35c22a15b0a22df9ccf3bc855af791b343fdba1e36b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed6e738e483a7e48f507b11413477375d359157dab786afc5aea1eaf135b068673d1e7c58925c5ead0d2c39d161843fc3ebb3d2c5ea590502014d67042569e0d8d11364e09655f44518300bc615d4f49b7d00eda40c3595fac13d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fc7fd95e002bc76f477f74e0e832a5238fdc7935b4817a2acb3e48db35253068508f28ad182f614803f3ce461edb15afaee8436610a70a9d461176071e9bc95947f9babc5db4bd41646eff3bedf82c7c5ad0d43abbce9b10440b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160a5dc081fb8b2dc8fc3b6cd7d77c8d5f4584593308ff629544dbd42c3cbcf1c4796a7ed355977f20dc9f6561d76b26eb50f13cae8013362701b180770212fdb2a92c1078fe4836d49d3b8ec1a6977d3c92ff09450cf27a14fd3f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173105fa05d9153a4bde632c2a1a43f93ace0e7d29044930d2a0bd51f54a01c99306a0324f80aabb6edd5159303e9e00603ff8a28f8c9d491021b57b075e3791b66041485a602c5f8e2f00bca71ab4eb75eb9b0fe2aed436bf19315;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f13fab0f47d5eff89c91374df237d14e9cd4e7bebbb40eda1fac0e3b25afdbd3a02412ca27f708c855a893a3418fa436a00721bce867221516ab1446168e086f7739eac856f7d4e23e85a87afff64e6366fbc65610d8b11c9a9671;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa3e197db044ac86c7206b3d2eb7bcdb37d382efe42d418f5d14f77f574c3da22df1143c34fb003f9f50badf9fda5a2230f907b644657d51cb04f63c69f5468266d8a628a87e6613c6589c659cf3fe967bc9ab90fe00c2b8e8367b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h503d7b2534c2b5b6c2366e21ee69b2412c695fa4b7b933429cd8955a00ad293ef2110276a00c4d886069d33fd31a9f4f59411348b40b175bb0050840ddf4a8f759d8d6273104e998211d9572c1a4f7bbf60e73cfb298e5f28f79aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15fe94ea61d566125c7920ba14e886304928538773c1797fce6efd56017ed9046103fd4362ba740892ec17b49ca08f7573b0b52c308cba41205b1160421be52454a09521bea616f2a2a7341aff141fe92b1bb6de832ee4c7bb29bf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc98a4fb1bf0e3500e71ff4a880399c1115d388af334fb5f67be128d9f7728e887ec48b9212191e6ac0db27ca83e6c61658df44d5208765a4b86ebbba027d003b506d9719b14b84ba3fe9342eefef7504addc21491b4bc9c856fc05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h149eaeed392b6f7bf5b698a137bcf74f16673bb5b70c5bbe917c8e1ba89d85fd73adbf5ccb2bcb8c1761c1b75cb58342142932187eb7e2feca32512ceb5fb320ad601fdeadf86a5ac84b6b5c4966b6c7577007486482945fdc11a15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9e7925aa8303e102c22b656deb101c41d507ad9c676d1ecadb7b3a73a0a71ddde5eab7c5cf11f6ed40d2dbe3a42cc608a08068e6c56e719edcc3d7911142655e0192d2af99bc7f1a8b595a9784601dd776e6cf82c053074308505;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6fe7fa7d93223e667df89bc8d1e5873c04f9cabcfe65997a579e551bffe7458b8cd6c744e857552a709aeeba1a607315acb14ac78b3737d357f71dffd174236c115a664307ecbef57d6117878f7090e40f8aed002f607cf5520d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h795d8d1f49462e9c9beef493048007840ab310d59cdb67faf1b247d55be01330cf30e630ec84e86290d506326d6d2e83fce0aeeb7410a1fe4db3241493d5264eccba1dcf4afc53a9d1c0e3b3794504efce852935c88ec4dccec12b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he37119e9b08b1ab4a1ab331a99cb53366f21e3d22f7e7874a6577357a13db972082c67870ad5b25acc9cd2f9e728a68cfafb944c342ff47c2da6b7d704c7d9ecae5c747ea14e3e94f1f2a2026b3cd179457bf6ef75e6007fc98d1c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h73797d4ac97ecf3e8c3684173f9b87f648d8b1c74eb1398fd0aea91a2f3faebf0b2664da31f1eeffbe3de9dd5ca25e3cb17714dc9a4172e306648f2a7cb28376240255522022fb4e7db7c5336fa110cc1c056cdc551d81ce88c799;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8ee096ed77c08f67b3d052fcd1f4dca859aa6a37a18286a241a680175e678e4c7d99c75f07f975fec3a5e4a1128009135422427cb57a1675e2e22d7fb8c47a36758cb67fd80f0cb2e4aff972e396551508823f0d3d4f1851654a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142240261d12e678a802a36e6185bfdac24c2972af28929de6e34d92e9a5067bb91a91c42b132f744856629b72efb64b8341f264a221fa15d32996ffdf00a8b8861a5e430dc09afa01529e6ae96f3a8d3a7f1a47bb83fe0099392b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15eeadaf8b22dae67bfb8a17698dca49d537ee56a6547429f3f62bd448121b2897af5d4a1ebff72e0be3d276ead077278d9f58dcc8f254edc03ea6e24d82e8ef098210995ac41e4cbc5f6bcd4eb974e516d33f84e82c8555774f1a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b8d20bb398b1b930ed51b6ec306b66df79935399ab2fa741160f7ac882bd90da3b99e188e266b64408bbe3fd3803aab1109ece6b6ea618bed28897e8769c37a598a255dc0dcd23c5a8bbb882183c28cb82b6657566f979629de88c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd06a9531806ad8cf6f145404429b01c337098ba616569ba11dde9126e17ac6dde8a4650e1a6cfbe07b5748a669459a958a7144fa56e8f9873738e3385114af74f6650f772e5eb5b8f0b8ecfe3cbf353ab98f218b367a41654b600a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e78daa943f61bea06c51e90fe3c38f1b829002ed7d36bd418feb328b68aeb467915fa4d229f49f4e6e1817edf6254d118329b4c4b9f5ea41dae43784b6095c976b42bb529b5279e8a915fa3faf78ebfa22b310ebe823032dcefb24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e1bb4b3802e9b275edcf3da40ce6afdfbe091b755f030281fb277d141d2ab1791f82407da662acab1e6135e5f76bdec6c4c69042a002d4293776278b404ba7933931463131d3da8d6b8f4c7274fc0aaaf206994a66f3ca4f2e1db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1833fd5d470f76462b473b35c91a38839a59ed8c76a76f39a8596b9977aa2bdf7a0e3b2d0b966b17a491fd6533a5134f145f2747b95e7ea1087c6ce1b9fa5d4333044b8c92790d0f64d39881f4e837c9e6777ed2d0cc1909e09bdae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba01b6c4b8d9cfdb3983f56b38e29d68df1f27e827f0b7eb2aad8268ac39d797cf886aa2879e602e74b7af944c5786d3828562258090e1d34d696b9a2313c7734ca5a3d9bd28e62d6357ac0e7926fff3313b4b92730231218e6c64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d7c4b6fa76262e5297b98b8a99510dfd6dcb3b1b46abd76341573d7c7eeecae413a3b1698c2480292a1381c2e168604a4129b63273d2d0e55040f5ab737016091f381c586fcfa6700909c7319695347ba07d0b51c3ae700f038b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4cd4fe4c5076aa476576c86cecb1519627702e4c9256d7f6d24a65ed24081ccf72ad38f9e9d079c7a28a57223d761512bfb46882f0dd81e7778c3a22e0495a5d4806c699e97107541606cc388e7c880e989d62f6386942b963adf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc33fd7cea9df984fafdae5d3e85b0894de4fc5cd06985b257b9ed17d5fe2002a1ca2dbd14dfb72c23608e595e4aafa243037dfc08232d48620e7cb04de6e5bb827d8ae45cf0a0fce4aa0538a3097468b8db3db5eb4e5bca05b0669;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e22fd5020bd3bddd25f9de687825c4a13c7f024bcf487962e123767e10fee4bc5fdd143445f2284392c808c1d3fb95b6a4fe95841e8f4c5f6c36b8ce5d0be342fdb54dfa0d5e905be6d133866935073b3bad9f1e27e12b43673588;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd6366af78f8bf3112688a680e03e3d6b04294f20d07d6a6400d3916105ebdca320ac4b03df642e9b074654bf79d987cc6e4cd5c2094822767bf2e0286ebbd3159f406dcf362c324cd0ca903825995b394de61784a33bee35ebc68f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12585f714c6f200e3a4ecbcd6b68ac22b0fe67de6e9b818bbacf7a1aa3fbdb49c783bb8adae04b72d8c8124eae5a2ed8bf3a84a1e7bcd74670dd89440eaeef79248f6ed3f3259e79f1ea1f05e52b8b2a39bc6d1fb8d7fe6326124ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2de073df88df4b93c02b4521200a56174668771f732c1052fc09706b8f647ea8a6b018c418f45056535d89e5388dbec7b5cfcb3f4b1bbe8532945ea0d7843a1309b5f6caf0579d07bc79d963876ded12c7e57e45808d5622fe492a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h110dfe9e5fc80703dd36aa278831dfa7aea0cb1cf0c934da29d4c101f0413fe9bd1cf6ab394f40f7b655a933855c176b92083177b6e596fcff3db28209705716949cbc0446fce2b7f977ed18e6630cd90d6843c9a05fb0371cef7ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14337dd8fc7e859bb9f68cf13bfec53cbdb992be773c5ec6249773f1f08bded41409d12a17b4a5227dcd388a4f71b6e8dd6182156efe9e701d6d3d5cf506ad9b9637d9e2569ab9b058d49e8a02f589f1b1a94058b0b8d5aad0d4c7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hacf4576b6c098559964001a78b652fbedde91f9002cbfaae9dff393994aea0cca01408aba5be53e8260d2061d5d69fedb83d86b52253c91d3bfe4cdb5c6d8e249c7bbaba08d077b5e9be64779e7d9761d33736ddcd9037728a02fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3101e0b74c5a63d286ed625857f10a74c04fef763c267041ba3c3b6271044d1ad8cbc58376abcefa45cf230ebdeab3204e23b0c004457601bba7b0ed3bd4a82000c1909396b0a3ceb049670d838d1ac5c3f1914d96ea06dbd7f034;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc4c4d9d40e4a3c879d3ec31eb2fd579c9bcd9412fcc2a9aeab7ecb821f7238250d2838d11aeb0b28ad59504843176158bca1daf3251a8b1d5e3aeba4bd98008e703befcd73d11a96ee50c914eba9e71f605c74ef20c47acd3ed7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b808f4bdf35f381bf4f3958c6b5d1325f6161df926d57c2e3dc345a4cb1e6d61235ca8d636daf29e8755ad6339d821dea9c27fe06a1b64e6209a31b3bc33b5ecf210a4dd57e1bcafc5a88cee3eadf01632ab338a209202490748a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c67735f25943624e85da72c261bd4b7ff1e1e3b67b2d6ca6a0e12a1e86cb0c8fa894c78b5d258737b9d40ecb2ea9e98b97aac6c59b2ddf37bcda3957ee15d442501f565762e56dd1a015dad671f1fc7a66a8c5b499f99021fc5ca3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8efef01dc550936a63bb6a97df58203196fc1d42f44f6eeeeb4d05a83d72be0bbe79b7bdafaa2d8bd92d84c25a97982b3e80919674d90193043767cb051a7bf4eb0db3c66b030b0eea59eecb53266cf18f03e928429372c834e1c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1816f76a33e99a5525a5a6a8ec872509fde044c4e6e6b3e282de61a8b6f1852406b60f086d2b6f8430b09c9b4b5b305c8a758abdd644fe80474528bfa4c766249e87759243468a981a4e2fd20cd5eb55573257e791079f6eac12126;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1900eb1ce374945ad1f916ebbb8e22de46be765d3ea39974cc85bd114b384c4852f20dc5eaa319ca53e14f8019504e0daebdf3ec566fb74237cd81481cd4134036662bd3839c4d1cc6af6008a60b53d2647f77317ed401a9ad0b624;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d20c7da9bf6a8e90486cf5ccb6c1bd3473e733bd301b886933f122670c5576aa9d2f5e50a24c9b075580594bb36ac7289859affee943e657d739c681b3502e63ea7ccce2200702aec851ecb1fad7172a392aed724f4cd8f19b94b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3045611a53edf16a5de3670bc315411ccc43ebca58d164e375771d64df6331b0db045baab7d05daa328ac0788557ad950d9f8b3c83fa33569874d65971186e0bf21fd824c04c4596c2c1d663931e019b1757e4920c00518e2ebfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0bda7194d65c5c0987b69b77f4007f90d66455d262ba13d18ac3e78b65f7892db28f041702567f1de3b6cad03531672a6cbc7b3e55bd4f0f4f6eafc6983046b89d9c110be49aab46ebf31bdb05ec4ea42db9de0b1ffd9aec38d9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1baab41132957d0bac374f7359689af0e2a26656df0ce122d55a6ceba1ac7d2c0db695c50d7efe7118da6517f94580d70d7240ad6312ab5243c9810d5938630247027e32c2e204682e83593d856c2a3666463856c22d914eba7ba94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a13f098e4a590b2a9b68844343c122069a8537a7288f09105780ffa606c5be6a80e1d161c04eae29d2567741ceaa4f7c12547e3da8608421c1501a6089b1eaaa85f001719a8bdad04906b5cc555d0ba69b239859a95b8a699bfa1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e077652253b93fd556858fdb7ffe2f29f9c9afba04aea71621bd60d1561893a6b1e2de32d2683725d9afdbde6e16610d8e5e028c2b430fed1bd3147519111ada18e28e5a1c3264b5061eb01668abb64b955660d6278335a8cf5ac0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107d4824bf4a8dd06953cb44f3d25371fd62f087b96fc5dfb7b29127606d725cfa68196c01626d89048ca23f014b12de8ea19d5d55727ea101833326df0cab7b32e35c1c8a6ac0c8520e1955c9957aba8632df3963987cce88e26f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c43530750a44ea5ad4411c156ce3eddeffdab6d603331dd012e758f7ca9c3b0d951520cf0fe60d01f9e0d1b43089e4fb59bf24ffdc91c7e002efbd8551ea24dca3443088c333726022f3e09ff4b3cb876d4c111a52ff06cdd1d71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h175b72c7c7059e9f94a60dbdb3957cb975dee34ab344f16107358a07a8afce61de8304557342fab61584a9f2fa366eecf31116a73991d06c0f7675c36cb6e2b4120825f2aa6fec8b2a8bbf2587f98aeeadca543349382a4efaf8e35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1010033e7c2a4183eaad04cb02c3d511f8986446cbaaff6e2f40405fb2f2439c19cd19b8c607f9830b5b349df5c62bbd96cc3a2c59d931d2940bfa6b278db1e367c7ff37619583a6053273dd37102f2693ae062dd8c90371c752e74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f078fb9c510381e5c74604c12f54b4196a49882bc7ddc5535fd3f07d3cf5c31ec39cc669ec8c64fbc64ad375e3fed6608f8b982ad6c92fa4d387ba972388c120e3be9594e79fe3a572534cbcf4b0923c9ba275a6355eddcc77bc89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98bf20ecfa84cddf211784f99b5853a887bbcb987cdccab32e6f51f3aa8d8a86ee83d5fa50a9b5cbd9c39d6c7654229b5613f36a148c5ef7bd236c99223ced641ded2fa00609b12a314a48154172d0f2026c604805e42ca2437be9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1952c5bbdb4a71c68901bd47452367f5cc1a13f27011fc3b7dee3c7705d759c899b753767475160f4ec0ade50d72db4793781118a57b93b201510cd861a861bec62af773ea5f8307a1724cb8e238c2175e10062feaf6863cbb70991;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h119c666e66678f9c6c049e8758e2657d01ffb272d01e8d3d7cc9626ddadbcd387dd979de57a40712e4d9fcda2f7f36b028e6bbefb9dce7b97389e7c63ad42b02e53fe49f0b67e25ae72ff70c1436c06ef6fc79fd566e934def490e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80d02d43b77b97469d62eeebeba6bf56e72da318a96edc66d8494178b55e17d8e4e053bec331ba97f9ac8a2a9d1123acbebc529bb234fb249a9bb771e7811b8d5033aa04fb589825125d80191c7ad0c14da3dd96e15ceebaa73816;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e61f696f73ad22b9002e5577106283d4807eaca81557e026347608450c52c4ee73e54ed6029bcf507403986863bd072a62b9b20229a0b1a3f1483d39829688efa0e6eb0932d82c4c937b8fa874f79f4dbc047eadf7e0041d49680;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he704f689ab8061890bb347be0194c25c6455ecbe2c1f8a5f15d5c62594e9899bcecf8fb99650f5138c411884f183c8693759016bf8c97f672614f6bf1985c2a7c679adf592a23afe60975604543c90310da1a2fdaab57c30275726;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda46642c03807688f018c85b17177e591ce8b8070cbbe9f08353b1d20b6394d0421e71c3946a43f02f0752d31cb86a579eadd7cf782ff16efaf99f2b5cd81ae5e0f90f976b96fb4163d185a78f7976d19473b392ba0544591f0a43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7217def6a9ca031bba89fe8055c9e304581b6a7ab5ebbefaede1e53af3e49364a3d2b21cab47a7a97e2742849595a82db3bbdbbe8894ed0288339c0cbbf894fc33c67697fb6aedf83fa19c89c6d2103d5cd0f901b890003fe0741a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he29b6b707afebed0ecbd2d39bf39486fe4b0180aa5cd5dac8332e9e2a5342f4e07968c2ab5e72beccf5332d93650dc38d0b42ca9b3c0f592a396c8a93d9e6b6478cf7fcb469eb6a27c9957038bc5485a04535dc3434ce31ede7648;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27f80aee06deddbb290788c1185c4e4e6c49fe205e21c023b51653966bf353ae005e138c34322f0d6d79004aebafbba8dd1c885a7e2499f74937205aceefc5680996ca66ecfced77e5ffacafb855f746ecc9eb62755a6cfe44a942;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f1a7974137750943f7175e749dcc468eeb6eb922c877ba1ac7293df8772be4cedeae23f2c70ef402cd75519af929f01acc9396e211f876c8cfe30ccafd0081eb161a6192ae53403a8b417546cdbe96a04d6cdc08fa3eb89f18236;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a921c23794158d7a3d3fca7cbe70b998e0f3e8c7da9ba656480dfd257df9f8216f883bcb20dde15bc786bd97a4cc5b7e09fa11eaa68168224005a1e0e02d69ec9793b3215c7fcbfb989a100752e49723362e36acfe9a04a7fb9a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e6a6fb0323e6d51a2f1c0400ef6b59589a5b367480b062c589bf8bb4be39ca2d6d593a9102e1caff2895b8e05d439dc968cb86c7274a35699151f19097f01640f610fd96431187f8bc49abc751596bec617b1f83472b33cf93bba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1931d6ff3b2745b627a2e5b50132fa1ce306dd7b71c5ef594fcebb212f3731116eb099db911d25eab0fb7d2b5874a0129dff446cbd40bbc47f732686229b7efd9b881e4f1c389e2f833b24e0960900c44798b053131b1984d7c32c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h341849d95e5b2414f05e7feca45691e59453c9da614c626460ff117b53cb855e76ad7be5e1c04ef6a68b702de6d4a9e157d3c7506ab6d88b65d1acb8d5cb8f7f13e87d7a58fd9f9c7768f7288bce9044d3e5ff0ab0a3d2ab2c47c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1debf9c271af1faf7dd0e2274d7907298400f091f7d93ead9a489be87e768e099de19ba4780e7055699745fd3b660884c8ab5956fd21accae3f4c97bd3f821485ab6fb4b3e908f4ea3824dc57331e3375601ee887d8fb8314ac79f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14f8e6ce094bb7fc127e4c4b3067fc0685a8bbb702473511facf81bc03c59fbc13a52f53acb7c08daebb21d4a0a903f7e6e92eb143fe9191e80dd87d392fbd6b9638a8d8378309fada1e9e92a958144226f9af6f5bc630f91f8caf6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c7fcc0efb7610c10b4b3ec4d1c4d1285398a52692b6e45c42997f30c37639d437cefafed422cf8c3f0b42cafd2d4bfc3669fdda3c3410ba1ce3d594d43ef3fbc6a624ce91e3fbb10f02baf9f121a699b1cc26e696f1110794f87e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a4b72b2dde3524cf3cf6c3aba36dd5f77fad198ca6110e6347effe8a5f7d843558c4333413f87c6bc8e171b0637a59edff5e0746147f8506881b594091a0d564e434c14e28c474d63d2cb652d38b4b509df3d7cc8ca36b1f842f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7301bbcca56f85c1bb1d76c307dea4785dfe1025a2095453c761dc0e6dc1849c806308a494eb8a1f0cc7812f4af7461f015b6aa307595b3ac09d1b3496f8d3b10e114453bdf7ebf7147c8f3cb7868f63118c39976c7b887588302d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h96998a934d778d2ff66b078e9bc5766e371808202c7ae6b45baba027c3a3b78214e3f9c27fa3aa6a9cdd21f81da070a7cce5d318f039a8e1ce12763b2b4f5da2038fb9d865da96de968d92b9cf8103af28f9bcf017d3f8beef43ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab804669eeecbc1b78427f89b3d54633de8e924ad7f7ad29077109d8999527e5ccabd2453b1eb631b647798b90806f7833409c085771e9663b1c228fbe31e38bd40961a219f3ff963799f7e6bb46bde3c9ea4ff2c31e0b8c1c1382;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11af77bd4e781619258c575c077302ac238fc9d14a058190d11f956a78a62749de82b5e1778e969a64f7425a08b637d43fa58f6d8ac951138e246ee0544d865d28b627f0939d343f1aae86e366650928e8231975c930e9167646d0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1826fde536b46a594b9280ee3287788b014d9bd4d97a915f40935ce8d0d9f94f4ffe13b5e51e8219fba07ca22af7980d0cfeef9252dc1fe3010f706cc28e69ee80d5e9cc987a037ded87a5812148d86ba86378438b8b148e9402d2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d62ecef6e28a2db777a8b9345989c3c8d07a10abef9bdc695fdd8c2830f14306187f87d1aaad3d466f2322a3f3901df2d09544b134ed440ea3175b77b08e2026f3c88816c9c99b6285b6ae74a3b5ed7a6539ca2b9207dff48897be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h425da023aa0a92658fe0e9c602b6438fa29d2dc2871f527e95970aa1236991833924f400363a506ae72afd41beaebc5dc4f8dace2de22952e796f1b7bd7b70e7543758f7e6ecd5ba62676af458edec4e576a945f7e60a727c23b91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a6c1e550a2bedb29455c35fa05deceaf66f6b4f1f5cf5e0a35f01af3d836f382132ed70bc2fa6d9ee1a08d88aa1ba96aab066d94ed780090dc6680acdba025b7e7342aba7f2a183209f8aad4237e984b110d68ba90b0587d339d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5f5907fd4e4a004fc4f69c767d93c5124a1215fa62f116bf0b51fca162a45aabc72b642f499a4945161905d381f50e1d3d87486bdf667a0e9dbe9c2b6eb0b1e47b5e4e31385fd4ac048a1dc0120ea885c07a9d1de65c5092d320ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d5a7c9726942b323bcd99359ff32eb87eb727928bcf1d468cb55f6b95a4e18d61dda000c2c688ee6dee72a77cd31a76bb14ed240a8dbcce865d7e6e52e007a58dc7768a987babd6580114b7c780122c5445f747d69d91ab54a51;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18aef095f3da2a92ee0c7418e6deb6517d527586675fc93e7f81219ae5c1d2724138984ad9fda7ca29eb0b656e6473cd6a59b78c399ed6e4f48c91fe3984694850b69552b2b4a7e6d0bbd4a3b9a3940b36dfa31b5f67a2b759b8821;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa493f616f591882ff612305585ce4a41ad89581b4180a5a207f34f9e7087b64f32066ef3f86cab22d92a91936d295ac048fd4813b1e836b60fe6ba60f16f87e50ad4ec4b877da0b5bc0736a8c5f12f3c765a240173c6af364354d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1974855725b691872523137fb199c40589c18d520656c8b6d654a2102f959de7121fac31d11846b6ec984afa7210dbf3aeb007cc9b421a6e172dc2486061838aab095b6ce6e2abdbc668eb8ec5fa068307f2f7cc1676df74641645f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153f2aff081b4982687e2280475ec9bc2826775aa4ea42a93b048651e1bab1a51c6ba6f0b2cae5894f4ff62fb4d707ab4515bbd809330e4c5474f6e21847451b69f5b58f1608aaff8cb95b08ff9c4f09c7d0b79609502fa54cdc007;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h563dd04b94d742768c4e318bd49fa9c0b727c7902905cee51784831fb63074b561099f7d1e8a0f6410bdd5a70c1ac580ac35bdd0974697ee7a673acb3a2715718df96f7037e81ec868ecca5fa7c2ae2c356265f49d9cd16b215ca3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179c0aaffb938cda20f0c101e40b254ab31eaa9dcbb9d809f3d5e3ff85e67626f5263f99a5b59f3aced79e629879d3360ecc8c7332f7862f1e98572529d33e31d3ddfe5242449049da041910d9b4d186402212029d7228fc9777972;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc2c7bb54272bba0860ddaee4867e9fcaf8ff21c6c853f03b399826cd9f9946c657e78da5a50782073f364ac995144c7cb8fd71d83f84ded00f937415621551b381e313a4ff5f4d9d71044422e28075c2af189ff1f914d5689757;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1109720b3e701afe05991a9f9917e7b7b51a974380327d51efa75786a4d6b41779bbc2c8194611705597003f4bc5cef7da714a3deb639a2c6f2fd454a25032fc353b150cd4218289497edac4f266ecf76660eb93c8e1a6d1a8ce58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h397ccc485a0de55111c24ca08084cb0acabdca0ecd2251f74b8c3f1915f0659b9365559fad77b3aeebef89b674990f61b43742d208d492b5d9c1d9f814518a91f92fbba910976c553d48e7508fda6eb84a94a6815f559fd059765a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a5d7de7225cdf0696f537b198324f4d1e4c936656b903f29cf9be5e466d8aa6e0608a10491e5186113f0c08076b7561693848431b01cf051844a696d5ec14dc3564bf80c0a558fb08c9e633b4515d6bf16f2f222f7304e8b52795;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca7728383105f546d0a51ce30e37624c960c227e7d6c73301f3fb671901664e082f1a2832b55c6de4d25761943efea6e970d2015e8017962e1d941d81a253818f2d425604e2fadae3291581fad94285b23be4b94febe1aff177ccb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2a685ba73dcc1cb0b99cf162d14bb8960d5f6ab8a5d3b316daa1ac9ce23ca91ffa1eb39b8117ecfc84b60eac83a695dc25381da371f903a43d05ede61644a40d3bc4d41f8d0e8bfb04480353591e8af2a47fb3a1435015a110399;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1542077c7da4f4a2d608f2458b9e3188780db016fcca96bb63ef8acf430d00430c307fc5e04fe489e50c361dd30324d511d60d46737bbc928d86d0758837a9bc1de35996b544eb2e84bf138497b6317d13112ea222193660dfd250e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ead180502e1b519480670dde44cbad94acbffc2f49ea2c8855f03ab73dd50101ee65411600f26c5c04f13477c83fa1788bc577b484badad4c2d258b9d8fcbe6cd21352e0b42b7aee85a7de3b4a62d0fd4810ef041b28c13373b50b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbf96b70db14e38c00f4b471949c860e6517a31f63e8ae09a686d602cab485828bf38baca85e4e81b0d2c91971accfbb539c3f8108302afdf33ae8c53a48c075c843f73665605f276d6db0bf713a6e8e8c5e14b29f64fd1f694f5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h145dd48a6c7f055400148db11114e791e9a8daacefa27d6855b5f157c13c6cdeeedfb3682c866cd7864415b92cb4370955655d34148fc99631e31133aa6ef6ce2f1eeb0eab5c29c5993268968b5a2ddd5f8ceaf2e1195b35bb39a63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5839eb57acba2a029cfcb12a4f25a1820b89a2403bd32228276a6f595865467e3662d9006ce16eea5cd5092180edc16bbabb4f8b8c995ff9c287661edcff272e0321a2ed4197ac1fb411d13772b87b0f59365c43ebc176125815c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c72b6a694a53b6cfe71700292092d66cf11d61672f1af48084cac26c6796590ea10bbcc966f4509f95e7709763c4fe39205d49d9305aa81ea234ff5d319da44bd94441e98af62490f550eaaf96bf28453ebd46952478a14b0f59c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dfcc25c61f345901fd400c460ff147852db072f7cd40fbb074c4d776faabcb9520d9a1f622fa805c230c34fee29bd0f7e9de5ebec129a563f70d71bb42e7aa2d6d825b53c1f7c69d22ba05a5daa1230fcf868797e1c25ec70837f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3498e9032f7a1025b98536ac35759f6db9ab031ec7d1fddbfef3f0ea8673a7b99bbb8fe0af0abcd4eb2fa6ffc1a79cbeb320fc22cd8169c4e8b3c87d46307fa811c162960052fa0368b498b007d4493c1506a845f4043774227e4c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a64814ee9d2e6a24af6110ab395c7153749c3e6e10c843a65df303baaa739fda7e136f236eef852196df9e5b010ab2e42f65694b36881427b5cf78b55c8fd88bbf64c17c275d64faca487b89a30b7d279846606cbed67ca923092;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h82a4c65e97082e951951c60bd8d3bc3efdcaa38b0db1aea7cd81ae53d2afad9685e7230472fd6334a63cc1bfc7af302c6bea8e65eddb86163d9a3f800f7fce8fe9e9b8e7f8698e1158b44a5a7a6a3082fee7a9941335092fa24427;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152cff0dd20ae5c8e6a749adb4a5fa0e819633f25c11a94614af59584aea406acc0faf7f6ca174734dbc1eea3075cd6ae600f5a17ee2ea4aff5a4f10da2fe0f7962f70763175c2412e959ba0c10ad573268bcb4184a63756a05d7f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h201600df2205d6f80a07ac8b0d438535eadb219d8fab94f421b5d56ec4e220e6f7ebf13a77daa4a49dde926baadb8ea2116035e5538ef8090bb63ab23600d479742ada580341540051f20e2b16aa8bd4a534c34bf82b63dc607d23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5be4ca084cdf27c50eaf0d2d862bbd519c9adabcdcfa6e6ba4f2e7fb044318d187dabe15251ed9f1077ec5001274cf90fc992e7fad57f3587b2959cd2836bf6b146aee633b4670c1c4692a8d89cb6917a4ea9338caffcc4d3416f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157523be0ba37cbadd1cfd8fcd3c19f488d88eb3bec4c45b3f9a63b81baee2a302fca3d514d306ac802110997e5079467cd5d03cf4c8857392bd5ae92cebfc83e609877138b2bdae91d5678149aebd36b38f48f9d60c17524a7a838;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9aba7529d78cf8ccfa96bd5878e6ea4c363198a2f30162fe9ddde878109cccb97cc5f465f2f06ac705d9177e6b19c33fa1b4c7be0e7e836542715fc3fde18d7e91a1156fee24412546130b30b25ae399996f6ff9d3871b486b2962;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a002e9870da230d39feba36685f0c80e17c9897c9ce97737788809e2a07a78911609cca9c0b2fd9b335707f52c6bbcfaa03f22ca04326515f4ef5e45d5b01f0f8820af4c5ab059eabd06af9e40f1ad6429a3833329e1909058023c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1919ff758182f07fba3edc358c2f0903cad0e358afe5b86eabb7d9e34fbb3758442a15470e30778afcbbb65475fd031f986d80505340e022988786ecf4a2b179c2960278474e0b7de1b3e61532616b59b364b73fa1edf249e2e20ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3fa2ea5406eeaf2b32294386c03ec93fb7caa6f6a26bff87fc94768f0f54b5adde55afd8ce7490cbcd910777f57d8ee8d1414355366bdb0adcd02bd1039dea4827a59c51a196baa7360406a8336a2f16ed80f8db2d82e289ea845d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9694bdd1d4c7c903c2a155345267799e3030ade732fa356c6d5892c29f31b614f23935ecdb46043be514e3740950e372b01e7cf25aec7d1aff846684abf3571a2c686d908fe80f01209bc98f20072a70e0d89144675caec32beebe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b638f2c6d195d6db223254a2e9aaf0dcfbadadfe9ca12e18311b96862162da09231408fe6b860e745f51e90d94dc63593521929f09e5845a250de96df533acbd8ca3fa7c28525eab80e63a248cade6e375b4ebc3985dab05e597c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2feb263c2cf67e0325df084e13982a7425f8aeef54d2de73c7f00b91530a84b28190c578f727f34fad2479b62efd484380caa77acc40ad2e993e737454d89ed0b49cc3a5529027038a382d2529fb4b08fc7c8c0ff20bc231181476;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc19c61ccb303b88827c380589d2d3f4527d0c4732d81e8c51a58930033824070ccab0623c2696dbc6e39d3355e4c1592e6bf169aa939c6a3fa2b456bc966bdf5e77cf2712b4c785c99b987f76324fcde6cf09139175f70e6e88985;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a304be8eee684ce14f12d54b323a0fcb5cc50cc8b6ab0037074ac345afc016dc694279e101427be836464d8fcaad2da9fa9170a160102ebd4dac78a624d5f30191f84b8b95e19b2e1ef4c615ff3217006610a151b3621881a1ec53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h44eb64237cdbb51cf75fa88a192763d161161c8589eba0db0952e457c4d37ae7ebeb1728dd857fd6952b35da752adf7ef0481078df2feaf2abc4ade437d936bfb63ac985cf433b645c8368255d72026172992c961c2c554414efc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b75b7e79f3b9f2751221857c6b0aca97fe899368ad5a54b08347bf754f29daacf2946dd1102032f45f8c3c08f05ce77d83fb25584a594fdf713cbe18c484aab2b1764e1d6e063e49df167283e63aa3f18ab96e86f6212f04c933b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a46d53ffc45ab428ebeb874069d7932ed326e362d4641f81f14549c6976a5edc5a7a902a244e05fd918fcc07a354064be1bfc481a3f3cefac8290f5a5cc2055505d08059d49cd352e29653d12dc6f3e622e17a279faf88d637e1a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f36027f4057da76c2e919ec87c7b0ccfb171f20fae0e83badbf2ba60d215bf79773da6a1c87e9d616dd26eb254bf3bd85b9ca690d54d7a4b6d113b6fc175273b55c955a0841876c358d2961e31c1f7a1b27745401b07f3f6782aa7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a9765158b4dcc251e574025735a7c420e8299f22a124515e0cf92c44a94f5cad60a06e24ff9a4b8cde2a1a99ffdbe925d045c7aa5e64f7d9751e21422cbaddd311ded95e53af0eb3be4799f79f3775dda64722b180e8f194e7be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf45bf4b1b0d9db09470651e7d1426e728184f40fb1fb8787f312c919e89c6eb4b2018691d12d2fdffefd13b7474be7a32af05c6c9eabb6ad1838f4e9460495f138b021ea0a4bcd9769148f243b10cb9d086ccb57d4183168cb32a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1768005a56d452a4e58ba7b8e540ea827deb0c016575ebad3537d1b025db55b8062a3f8944241e5ad4653ca19c1972a3eec586fd24ab327e4c75d06137e8464337192d3f456dd32e0a88fc3d2a6de9de10b4e9d821fa8ef84ae5088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbecfe5126160afc9f818599d7dfa02e5ce0bfd9ece5c2cf3ff701e6df8337b77a3c576eeaf3442f3ec1def54a80e4a4474ed2948092075cce839f1b4ab98e2f80b6952a4fad48721549d79053db873a0547b18a37c64a2604efe81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19089bbc48c6058240b644062d533d70a9c76cc92629f8c6608bb9cd4028507831aa423d37ac32b3921e3e2e515bf425aa44023c402fa023b299397fb38ae215dd0a6f2a412d55c7a3ecf05e99916fd22311fa8a4ea8a0dbb287da8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha52db64cff86a0c1a68c67a50b26ed6da0ae07d9681da9c5028489e255e83875d36c3f9483203fcc0243a0e6ebd86ad68749a0e2c59b37af6fbe82f94b977427d76d5d1f5bfa515fa983a112d0c274a3b10f612be2dd024b18bf52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ddf944cd01ecc2c05069ae945597a821229bd87e9afa68ccaba18eecd6f52eff79c442aa50dfe3d204e25a851efa277ea4077b4a3b2b8d43d1b7ecff07b6bf80903564c71cf19daf74bf95873b358d79d89b2bed0614be025b0dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9de93fa50e2f51e27d6f6f61c24a4d2edfb9cd84ee0cceaaa9c3b96452fca20e7c43e2292afafbb814820500ed8565fda461c983da7aa879b64dbd2713e37163a7dc0bfdc1b4d03dbfbbdce3942f5974ac2bae3f9d6c1d2de24fe0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6b03ef7fa3def13e5bbc1006dd27a7d15e539963f5aadafd4d46416bb4d5bdb244691408724d4d3f2d094ac1fab978453db774b0ed0a0a0315f0848c80e2b545769f9202aa0510b44fa0d796a92364c821dac7dba5780d06a3d60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb8ff28fb361449ae688c38711c35a7307f38a283cd2e4cc0cf2f25ea86456edcd0cc9526601f6bd4a895bbd49ad3c067702f5a576acbaebb6628c28fc73ef1aa3dd9cd7e76294d68a3c4190e873eeeb1b9e487628e327964fb4cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12bea06fff9bc2172ce18756831956de1ae019c1b4a8c5dbc0f78500509b0a2e0709bfa23f8d6af15c81192142d6d740aed151258cfb9a31b20fab4461405323c0054ef27e273b9580886de93e867de61c3e8dc1006826d3947a73c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hecffd71ff899564bfac77b738af934868688a05f37107b626ec39781ad50c4fbc5bb6656a698f5b301042cd0368ca6adbf01e05b64225739a1e79eff58ec1f8be8df7c8c81aff144c1f63c2ca719751d276585be486b81b06fe680;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf34864fae98ba962b26a611c12ef22167734ad9a0ff3c45deb449af54b0d7e007fc5a176341b9a371c4706f0935c3a9ce73e1f83a2363ba988ea3fe0cb6690c6d91d7caf36c066c18017fc9d2394943ba4318284959612052edf79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5dad97c7ba85bf0f8b3d6ce7ba9b56afee627c9967c147c073450036de56d96507dbc77cd5cfb32ad0c4df70b7bca3a780e542c18d2a2fbd8433028943bd13b625de0ba903212dad707a37e850aa2fe0c3f27c695cedefac73654;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe5fe3fff4985f6af7abc00fba4a4b6cd67b8b9583e250f848db9ae04f7c3e8e4362719ef1aca50f0c4e2548075e0ea2462c27f6f31ea8b5e4a26a583c3ec3f20f50ab0ec105a00d3d29bdf5e149801211af69082201e66e96a762;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e671c936d4cf0cb331b93b4fcf775a16826455de99b5ee38e0911d5c51cad74061a4632cc4179e6f2262e61493ff10ecf85c71eee0336888fe85e6c9e593eccedc1847f16d9f86034c2ab9965086723b7145c611ec4f35fb59809;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20bb6a32422574654c102e58178935c77e7a8702cd957ac46aa79ec347f41e4b8b82cfb07436cf63b8ca714ad62cb9f5ca2f68dd7085ca274a956f2e9646acd980cf71ee9153af9a8f0137793cebf35da6fbc8ff99fb14c5767a46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129e4ee17f741994d679ec230cdc9649000b82a5482c82ef63c5806db38d14a85555918c54ce5da9d1373d14cbbde77f4f04ca703e1b21b09101c7436a569f258c1a90355f2c559aece2539c43940d1dc3a6923f3a10895e322399f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4484acba344dc9a51a32d06f30c95d82a8f05154941e616ae208534913187e81211b8ec9ba67ef7acefebca511ef0f63176e7706c77e792acf2625af728586f4d5111f182978f7a2dd1206fa64b4c375d3bf36f1f062a02d2a07bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1cfd888373a8a0bd25bbbd42dc47ac58f087f604d1ecb09bc45e5aa4eddf2fd262890a4f67eda95e541a98ba9f88cb2880a9da24f7cfe8ab3d6021889ea5d94f62c5350cf5e3d50f176a389f5ab11d8ddcf47c9763c2235436208;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e29c7b1f74e181f213413159d47dc4e9748e1238859cd294ac67373602f6c2f0d06b241c74e3e4eac76bf029169b5e3f7becf51385e691bce10a73ba199a457a3a37493a806d992e8fe30768139610d571918ccf4afcbddbe35a79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd8f831f69874edf6e7c429ecd7d88ca6ce2cd1abe392127827d37b391d83f84d762be28f2c349370e49938a84881f809eb91d35b9328960cf6f73b921331ff6cb6ce743d940ff6de3b2fa8c2e8cf6263789158229007a435b70db7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a40b86b0e68942cba4b2c737267503292b74c443b78cad42f99be7f90729780dc1310c39a381778fdb804b7a97d002e6a60ec32a6e1b031c6c5978592b52ebb31741189e70f7bda7200db52a19430f4907d55064dcf39f0a6a523a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51d088eda09b2a99abc46c008570183aab57e96dcec73c23f7a87d6d85a1e3ba9338d95a8f56ca1880af5586871feb23278220403070dd33a8a3b3226954ee68b28c6888b45b50e2d00a58f69fffbfd0459b4d19033e0ba0bcd20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed693668ac33b29cb9a54307ed47a790fb255a5957152ea19fda27f5c8e60bef8e5befe4f6d18dcfb9207c627bc39fc3b4a1204f0182f65d561933f7f5b91f12b42e2a17d50926a05875b5e1043e884b45af90d8a53afd07374e9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h419aa853fb81af3896ae77dd236c74d4cecb249cdd3eb7fe84a89d4f5bcf2e25ac3ff975770365a206f54a4f05efc7020eb22d6587a14c446988466ee6525afd6de9800265e915a11144bd5cd8ea3b2d733fe775444bfd05837960;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ff81791d93d0beda69b3d30f07ad10ac48e27e2ace1933a879b32bb1e99386ca60c8a478ff00c5a393752835fc3be09ca32d90dd924c2a948acbc4a6ca93c0e99dac36ccc86f3fcb949112222db14038df1a77bb9cb62581722b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c3a6ed49124eaba5bd2368b33d429f3618e601c4f189c59b6aeae52b149c790818a5fddfaf105290ffa1b8b810086ee1cb620685ef796390e0c2ec0d51359b43ceb87a487ea7e4200623e8d46dcfc5908182f446d5c3813e5151d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h101c866bfcad85806ff49abeab3b033f26cf815bdcaa7804d8626931b0b7211b32c36ce3cfc7fa2b0c4bf319726cbe4e6385bac4ff9d2651433ca95fa3702cefc65ce0f57945f64f412af5bfb532d2f7359bf415d9aa19878d234a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h295be3e64d701ad83ef5d490d703e9a6076c6bfe09d75d2e18746114855c6bbf4ffc7887873f45bf3c55e8505588a7ab7cc621e0bd32b8251c4ddff882feb55a31c9497984aab2a8d53a1dce74bc07ef320b60278e56cb924ae01b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168b94181fdefc244e589f7461b0b21da9308ab2ad5306ad7696229676a9d3913ea75264c5fe96cfc6059620f00df716b3e96a1631d6d08cb1af3001d046adc16fa0c409ae2288db594b513afc306aa29f54ed478ef892c2dffdbb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10c26387844b8b4bb5e09a09564293fe73961649e3e95727debb4e6e0262912237ea93e9fbab09f5a04b4d04a02233a199daeca926e6946835988df6982f9a6b051493ca21204162c720346ea9ea4f4783d97fd469d92bef72d8bfa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111dc78eda8db4536f356806281e7ef7b6433a8a3378c4f6a40c8987c72f27aac7450f51a9e5d3202a6f8c299b8fb78bddb6b58898906cbd8d5d84bc0eba0ab163c3ad623dd947c20c2c755fb8e85c31c5d3d4c5a687a75efb9d522;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e9021fde7e99438dbd17da5f3272c7c613c76a243068c4c6c6210b899cc8c06e3b9c3a2444b654e33d976633662a9fc5c259551bd793b65817b0373b15a116cfca1d0032b334d65216e055d5853b4df3e9aaf8d4800d1bb5e8597;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190076ba2f8cabaabaa8b99c96033f93ab8f4c8755afb5600b9f373d7fa7470250fbc2461a38e0f0e580016768a07b192b5dd3d7dc66e3913c978cce9134ec0a741cd459bf3de690858bafe8cacdd4894dd865c8b6c1b6e3081edc1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5716637815b6524ef53347ae053e4fdf3e0490bb23fbb7467e8433260755393ced683b9b7b8297fa04f69cf875804412aa25d0bc0e278febb20c59110817090db13d28498d39fa3b3362d6e68834fff79054ce41b5bc97bad2761c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6202aa338fa6644faabc8625440fb4b40b45a1f1ee2557a1e9a2f7a6811ad073a1355bd8ddf5efed9db9a9112d00aaad3b7e1036877a9ea5fa64c37db90e00bff92e07c3a4007d02b3f0ebe7ba34f8482defd66cfe325d29ace3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19973e5b928651ceb6e1ee3ebcb046e17d28aabe3ad3d810bd5ec2552fe66622a758cdfa4a9031e6190a1dfb8e403212d83fe3f5aeccde429d01cc7b47d6db89fc0538335383d95689b7abd98e18ba85d65ea76ffb398ba8c962b62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d557927169187419455d91642077f9e3295c49853cbcace816c87864fa0b2b4b44ae68d6b698b6f02ba5f7160c8ef9ca786656616796fa79565663744570379a7890a682049a69e0933fefd0f0db114b636fa7f10cc229c563792;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14f63e01677b7bea8257bfdf076029e238f03c747f7743b643e29a86ada6dc11a6dd89beeb190788c217b2060e2284495c3ada47efae6cf992cfd9297314ef59a9831ffbf6340c204140e28d52c62b426a62255bab5f3ab104aee73;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf7a01738bae1f5155253bfa016d197c9b2e991fe7f176e23ac7bfba2f42293d18361501ff1d601fd5811736505c1475fa5408d2f0e15edaf41ee98093407828fcc325108a0401719f315a755238086d4ec138f1968abdece412d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf45b9bdecd66f7b24c07e0c50ba1e893411f80863c5032e085cbde2a38a45703d1ad7ab5c572ec2727e919d05a3d085cc3608fdab4dd1805202d1a42084ad3c8b5228a3af8f4853370a8601da9b9b9db0bbab495b0d5257a53088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa45a5c8a225b04c2aba0e0358c2fb8e4199a2447edb5bec1a7407876c872799a031427080f45600a40bf6614b94befcb0b1d7b4282a522a7d721e3ede51e80824e61142ba9e000b192749f22d05a3a257a35f661f95d67913c832;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e506904bcac8e4d24394adde1f9e118fce93af421d9945a934b3956c973647e05cf5b5644e9c44b15f9a126895159df439bb4821c180e89e3000e496e17b43ba1e7be54e0e957eca1e84625c584d8b2980936f8c1430c11f5aa8e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h914e14d2696def214068cb0034de2735ebaffbecb19d8d469bcf628a54c7940c87d6e13bb726af9c34af87ae44e115195b07f9e2677a26a0c2cf22874b395407f99f1bb76875d82204704dedcb2b8fa9d644e47e6927814efa4e93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af85a09a18370ec9ab55e65effb70cdc285ba5473e4f33ac798923f177e3cb85fd4deb40b07325a1f699b880948c71de855d7e2e2fa9eb03f1f13f58fa1605e3e55575144c0411ba133c078d88fcfaa97b625946f2b15d502a0645;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14616b54b1709a0ce18b1e9306d0b22460332f2da6568bad1dfa0660f64b3d670245f27f90bcc41356033c2179ce156820cdfa854d049da233a514fd59bb640084b0d3fe0b04ded894a95ee314657fc8c126906acb760b57ff899c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a51de1970735e7a9b66acf0e833b372eaf983d827f9c178c443497b5f25467518e7aba0c9c8c886c2cf765a6bc20dd618f6e22856c618776e88ab2073854451025daea02e481ee24d39b2fce71a52d9bb4d307c2de77d042f26da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1162a1bac3704863c6be040f52ecf91d32644c7060aa755683eb8724f98f1579bf4d89c01a6cb88caa14d10121f8d3a9d3d4fffe7cbf24d6cf202cdbd19639ae188bb4bc91616424c3e921ff19451e98c4d1de3ad82698204c5eafc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11cc569f42405deefa9e6c971bce49c7ba4cccda6ceac28ffb6b3577bcc918ccedb6e7bfbc457f4a1b184e86b5f814819f9fcb370cdb19b5e8014da17ac765cd9b7dbbbecc3c2afc9e47546aa93918d89b24394d3bd4c6d3d1a22c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e091310dd97fb594db6d27910aa5e1c89fd1b4e4b5bc73b3c07f3296a72da352f7206d36ab769181e0f428a45c67df87275a64b2d89c5fe07da22a8bb9b90563a5fb28ecfcb3c3282e91eba1ca17592330df3366543399d35ce458;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e9bc7443ee4ea464305997930f222ddc12b35a0dc20da2035c2be10cd0547ca59ae5b7946355b4665bd5d6b280ad4cd69c5c5cc0c49e6c7215848dfd724ada3c03756cbdc652fed57298517409588b95b746192bf2f334304ef3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc681b2878137a6819008783f96766b5e1c8a665b9cfd204de995f8c15131c3c4c97d7ecabcb1d8277b1b729ae7659df8cab44c5d1de379f005718782d2f805a0efbfd2785be63475ed8a932d7f4b8fedc3c94215320100a359b98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aac980292f136371e52e778cd15c27b3704eb938dc11070f0d5caa5478f22a11df1a3c600e204cf69f22c2dbbc6ef3198c305966ce9ec81bbfd33fbcbba3df8de87c4fd8c72e76f2cf23e5b433a66dc69c0fcd206bf853f5d7911e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16bfc12fb307b3f4820ec57ee187d7d5acdd918a180923b5c68b8455f6876da441422b17d31da34cc8909e9916fa379185260e0dbd4c44cf7db0132ba85a19e09a32f71eec1a40d63b71df57fbf39e451f8d02205bf7744f32acef8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e71888d1bc1bbaae586beb70dd0e5c2557941930128f53c06c0ff6ffe3b0ecd72721179cd582198d1eeb08fdc3cf9cd64b7bef2f7e5c2a6128f5ad1a74e070f3de613587183305f0e469b40547b96d1fb91bde9be2aae055d5551;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee826395ce2ce3d5e379c9a1479df1ae44f917afe77f2739697f2dfa97580fa495715353499d91b8820a46113683d9a736e77238dabe4e1865c647cdbb9e9bc3ff80bffc2406ab6ae6a673725dc491a675167bb0690329061cf7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127f74665de7965927b6c127f2a9fee45b9a34b87e05b8f90a08b538a61822fe57eb4d42294e8294c449c913d41c431f442aa1aa8524976b10e4a51b8e7b67136e1a45aefaa53b759b9651a1c71ead269a0bb0b4b1dbfeafdb420f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha21170720ba9aa78fb8185473e4b68d89857d2ea676a15b5965132447a7eee2f1a106e239cbfcc9542889d824f1174914f7896c414bc6fdeaaacf6d81393e78ec090211c783ceb5145b0916bd0a41ebdd97c43bd79fcb47c3a8d7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h604760b23d0a11e4f0eab2a903a815577f02fb8e8e9f78fe5433f955881d45896ef2a5b8ca2404674d79771661a573e981c15f8bfe7a4199915457be28cd3e5de94f397bfd71fba4ab0505d79ecf79a3f70eecdd13613556104b49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc136ac630465e629898eb839d577c9d2df652130896d033fb492e7716ae20b64d1a9236760014442b3586ee972ca9521dd661124d9ce379e328ddc09b52c97fcbffa0c00cd0982039a2de3c4655527145d666208a1d5c4162b635;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1612ec3d53991b3214cfd18b48bf33f44847869643ccce4b711ea371fad6ac515fce443237b8ecbf58742fdf5283fd17016bb6f536220d779054a06b18528e23a54f33f0d6354948d8ef5df724b4f5e20f5e038d07762e750238044;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h165f32614294190cb32cac402be19b3f23f490f5492f91135fc855439e7b8f2a379e3eb1647c2ec7133c356eaae718462583336dfbd0513b455d03fdb568b88441eda11f5bff0bd1968539d94ddbd0d4c9f05e6921ab7563aebdb04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h52ed7887a3bc386152c598148149bf4b1773d054c359f9986ed92e853b2112eadb3801e1bcb3dc10dbb81e57e7de0e53b023d351ee798d1ccdfe4c4d3439a719bb4815656bde7b09c45a60faf3a6c7706c03e88a5bb64728a36c4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10544fba3acaedd34fa37a34dcaa548b0fd9f83b40170c1611ea0c8759bd65a9c2b93d3f63cebfce16380a9ae1840e6968e98f5cd0e460680e999d9f73794f308eaf64abfc5b45704081e38e69eb42d94de9d7c195dba5a9d57aeb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c75ea56606d3c9f6e4ef82610fe57affebb0b6429f05a053d4b6144da9b222eea0f44ebf25955fcff54f558373be0ebe90b7fcd1f94142ae66ed17a4844eb9733adc5d2a879a5db1b4347f5679c6bd5323d955c64deefaa412ee63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc9cc8d43282d46fb60a3766749afdfd3c6152ee2521b5577fccbdc4528bd4fa8b4c773c67f9a3a5e97a0bf307d09e78da789c8f439674d2a7bc7270c2f08e50793caaa1da499f9b57a5e5a38898afa91623bf1c6e27c3e0cee1962;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12aa964361c6a41ee4dd7e023c31d224e38d81023e84a86323956d0f99909ba766975f5527b0a5b9beb5a260ee912a2c33634b3efdfa582644515abd9017e1d5a891cded55292bfdb28bfb4a810505971753e061f117a5fe90f573;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h81f7569d988020343eb1264e3a817de07e2374edb9e09c22cbb92161d9af11caefbbc3eef26e9596a074f0152b3c66fe7423a50d288a1742087e96d09ac5aa6ab204a1abf3bf80e62096baba7d5718b57256c5c5a860d05b36e245;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb37e5fd1a051635c55e9c4613b21783ac3ba17daf1dc83279007e7ea13937cf76dcd1d9e32e7321dc5f8be0488fa667393a322b22075615fa6fb11307a80c0988556fd7b51e528ab70a2db13b951ff9e2cdc16e7b1c30b60db8522;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47bed1fdf6a2533bf690c17ea5db42278a8b04cec5c3ae0cf31a5c04bd68a17a4ccb08ea81d8694b9c82e48454f73409a7c94afb5d0beccec6b1ee8455e0a8cb68e0fbfccd9e83c753ac76932928807ecf33fd889a553f685610fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c298a0a04bf777f133b636e463e316dfc83180c101f703e8a9d75cc2c886f5b86d16528e6d7002cc2a7edad259b9d61c25053106db10c7491137c5e6e245ee5b24b4cac1e90dd3dd454d68f2e3b2510ee6ee314001451b42d6c2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172a7521ee85992e4b9f6443961503347bb532c73706f3ddb7ee0f8cdbc287f81d9513c06ab2cbaa4ed0c78ebec9f601372af768357a9dd58dc648f9b17427a090d0f818d285a634709a35fef65b1998bcba9fbdb162b405fa51b69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116f182094299a4b6f968db98e4b09e70b5756816f6f5241c60de9261e37a8b955a7bbf4cdb9b1e55728d14d50eb0028c73c85a74140449fa117489912396e946207778e6c0b99d9b561e5be77f0a850aedcbe3a5391515d66264dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e4110fff659dd4af38021117523fa5a9a7d71f772d5df4f34f4b01dafebb3f6876854d8150b1d099fa9f3fb1536534d7eab3c1d9e23ca2bb56e261a9a485acf1b28f92ba9e2dd8b5746f96d454600647723fab6f74221bb756cf6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h783a05202e180a444d4ac34a3835396077fb45b71cf78ee95df13da1d252b272603130a84d27a469eed6e954914ba7243d47d2c30daccc353c5046074d14af638b65d0d73820758baf31d3bd06257964cf1ad22254d7dbacd05bbc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6337e7618feee49ea3ea9c6fc6b4cc8a5005907ac6c6ec48ebd96edc2fcd80c6b31d28a76f4ee2e48497d73b893011de9efc89aaf90504ea0e8420dfc121a71a017fd3fb487acdcfe06a2b4bb51f3805a14688939965c8b5349302;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3d95faeecce36fbbe94b0c1658a6719b5e55dbbbe095af812e344bd7bc647cba221ce4b6853c561d8a44e79e7cecc430602a924fc38fddba1c64256a9fa26644d87263a44d3ecae620a2a274f7a79c6e6062a8db1702f1cf937166;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h530bd50057194f9be46451f2d8329f0d238bd169a39fd8fbd7a4bbc7c70c1d87ded350ca604295b82a58f1729a69e513aa6f398e2c08397f59d37be5b1cebd8ef373d35b4907856c0477e72754c7ac897246cf145e9958f2f85711;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h175c3793c0f3ffb923d96c4103d7d366825f4e7b81ec14d48e4fbb28277c9fa004d282857bd4a6bce98011c9f1eec99fb2387e1617cff9d454baab58858eb6f4143a2a9ab2868443b90f9b4241938364fc966f6f1c99419d30ad37b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h45966f8a59bb35a3515e5d7f805515274f259bd7caea6b9b1a4b5cb501ee1f8ad6a92946759f5141c02a40046de539454e0f2d74ffdb6d75509e6a6e63598a787f421360d0c07017febb0483765b67b62fa607c8e214d2f0bcb3e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ecfc0c8c9173a9d41c7be51d34d620b21a7d7b3bf39d5166344ef44eeb79cba481ec40c69cfbbd505d5cc85410b49a60344e9575ede40151ca9df96f80d77ac8e9e11ad1ecbb688be69abf43655e75fbfdaf64ac46c7b3e8af693;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15220b94a05eb081c56a20f743f5288198658a02025b996b8ac16a7e3bac4e3e5d6a2640ff235dbbccfaff9f7550d813c57f6abab3211e2e998b3b14ffce9d989cd96f01f3bb6d4467e1f5173e22993ed540d0bd3e7882e9174984f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff3442a4c648bcbae1cc0643577e7ce4b186eb9c3e4848311f3bc65ca172f8cc8a97d3966aee11f01bc4916810076ea5eba9005bd7748c4c4303a54e5d9a4e0e18e26c8b4361707dc670aae326d08ee6c4f2a32ff6f1ae5ba7384b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd1a49f393a4f959cf7b06714d079f443546eafc417fa7dec7f95702b1d8aca806ad3c0ea82db39758f3a0543bd986eb07176bcf1908a171372b94efcf92cc314642f458c5a68a7aa0c63bedaffb9f25ebab0c6a5e6c39395bfdfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h674dd84c373eee68173a37fc53276fbacf30172d18b5b4735e4a0b97b47e3378235d87cddc62971feacc2c224347333fe081df082320cd506015242d0c7bff2c864188218afc7c91d42310fa5d903208105c04f275d91485b5b63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb5d20d657318f2c9852ada6fd704b4fd9d6fed9f3910ec95daf29ee05c05c43248c7ea2027d39fcb525eaf99d0ab00ca4cb8035c1aaabee24eebbe4970e365e67b4daed348d84092d947ca4fcdc92b559e88bc358f3f7e1139645;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146e412dc5a5a9fd7fedebfbdf0bd7a88e002bd06ccdc59602060bbeb49a807d436d8b6070cdee6c47869308e40306e26f1bbdd28d65bef2af6e0d8180696e997fdf65f167c942ce3bc7265190f182d640404f0b1b5762e3a841cde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe02d3b71254300b7e441603c57d4c30ad178abed9eb08910a772090cdef04ce30533fbfa3d9547cc3127659e98ef72c7a60768b1f57690de97ea3b8105afd30d7ca20eefe59bd95d6e0d9f95bfb7e63112ab7b5f1f0d6b97bf1a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f3b361c219a328d03fda40e8cf4092b7c3205f98a405892bc5314b460a089a5c4478431822cc32a54c5a25889bea36a10d225e11438540b74835d518702cc60a5e22fe24a528dc296b39fa14afab96858d96f4e7c49db62e9a097;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1adcf3e45a9ba18c09b2dd62f18b3734b04f60c49b18d0e8ea4229b23c70b24a1d5fe94efd5e9f3a02a23c3dbb04e7c46f89b2dbe4297b846bcb547208c04b2fc9df6f8fc412a881fae3fe83236d9ac43992c63439544bb77e5b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ec11ee734712ad9133e7b6c3f0eabe3ba421e684b3d5180b4f9d118a060c6d870f556ccb354a98527b891eb5c81bb1dbc141e53e2037ca16c82a265d242eb85e7e48fb9be0f00bbb51a6118c14ae96a2e6058861485afcbf9a0b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105bbf720c0328a0236fd52a76a4d682cf8f69fdeef926b77e0568d7b426cd4ae932c6a1584cf4f65a2ab6567a34c1483c0895b844844c97689047f553a0fbfafed572ec8c352a601c286c7587824f5660b589f916d80e3f087d3a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h175ba559e4075725ebc300837c2ab1e996c41c7d060c9c4b46f184eb50ffab24a7232720bc453648174a3c002d212ad20476d419bc9e2ccec30d3d895c160aa55c5429c7ba65dae8b3db5ece9c996b3033388e0d6ea951ff1da4dfb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185e78888f6d6db327a5e57c00a54559c92353e5542bca7edb311a60999bbb727f7a51f7a5b11cee8f06cccc44155a799a2124cbf84334fe1836a73115e485b6c302b713e661770a168f161e5128184be06ad126922fa180b1f50a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1886da70130be92479930e335910d1e3218012001c12c37cbe1d945887bc9cd1b2a9039bef151f522d6daafb7b40b33aafa8b80df509172adcf0d889cfab74ec02038cb067b359fa32b1f5b883c30a91887fe7254ca0a3e158b9f70;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8065360feda792196c4d51d858197a1a5f92bce766fd25af232b11e66c65482bba2bc439776b0f2e2af75fe1b6a2215c0ac22021a2f94b9e5aa7097a822c1c6c50a446311a46091c5ecc7e2dcf38d0d68353f805322841e84c387;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a72c05444fc0d6d2ecaa30b722a572803495df1e60d0f6616f7b6e8f87382110580f0e82b25b296d1bd0f9caf0012c08c980ab7a0d82621449d2f850d33e6557bbf1a66a9bb609f5d65baaa29fdaba45c6c242712ee128772888e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefbe3b1f76d2c223b6adc9ffe4e79dc789f03ff63667cd7e802f9c2fd90af6cace8685dbcc8c0d0ed06d180d4971d80faa7466607cb1821c19b47e80dd0e4324bdfe833ec001bb4ce7340490497a2f4295a4a25d72e4980fdcb401;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a63d3b10f50d0ea739bcfa0a89a6e84c17a3ec2a718cf88cbcd1c83b52b99e1a631b9e7bca62d0b33086ff7a5f77793b6c39f48da65114b4ab5dcbe1f5fe92deca81894144000ee492c1382b8b58caff3fe4b6f878ae1e61b6cd5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9b8a0b2989803e1da90636a21f94427dc99558202a992ac09f603eab44bbe23a06d3b76235e6699d499711edcc2a4bb5180451c4cc3db11e83e7c495d1b79978e9a1c4f6a9d777455d57feef453077382df51d5032fd3b514f4ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195cdfc6fc6cf38b6a66f460658ef81fec72d26afefe2fd4d4d9c0abbc25fe5a1313c8ba6b72f27b95149dd2ef0b89e4487a5788363ea3e54235ba1527ae3aab6a7d9c339ab272ccb76d292b939f894f0d69ddca2536bfd157d9853;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca62672176e73a3b9a54f3046d071e1e526af91fdd791a1f7f51f74e29ba0639a29ee28a4ec90b5ee8bc7faeee48a9f40cebfd4d2571e50c9b56c355274e0535a6144199143367336980542486f0d768d8865793582fdba62b1374;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b5c0ab31e9df9cc104ae4c375476e38c47f85be48e3de215663a5c77376420f5499067496bf33a8d930dfd6cc51929bf350c7dfa159f5325249f0ffedf15c6840f3c7a92b527ef4b806645a710c892f814a6dd488efe7ab201b18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c33eb4f8c630facfc0f663164f57d234ef11b94315f5522e9b37b13240f671ed41cafd8edc1ac47e5f3d7ed5496015a217354e93120bc8ce1ddf71aee7ec9f13e0128de83d357e3717c5449407930c3179a15b5d0745d7db46626;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c10132a754fa4a632c295cd77afa842230348fa281703f0d0ce5c388bac38b89eb8344d592579bf0a5bf504c408c63b8a0576934d3750e6ca1a5aed9f0eaa3e3c1d80ff373fa5e1c019f2c5eca44030c9acd950cea255e8ccbdb5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f257247a503e2b8d89a1bdb31480045b26f146ff9399e403e92b64761e5c33c388340bae7eb25d864450adb36dbe5c2a75ee536d4ac2c72fb57875ac1c680ca151fe208633463846dfc4f130325d2ea5906bb1c3a81c3f67a67552;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1240659d9dbf8363a333efb833135dc8e93971a4756d757d9ebfe675ef1990dd2f38accc52b4df72355dd0d7ba4504d1e162e6bcb4f1904d3f093ccae9fc9f54e8ae978d1383732e4452c04be7de595e9432f5ba51f5530e5976579;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0db1e95612cfce40f77751bb1113c4c9b3338f8c796bacb9576c58ba2f85544e3d5ad5b9fc62bb121fe6a48aaf07ca8828ac62f358326fe96f6ccfbcc89872fa45200c66405a32573d9af702e7b8741be68eafb7cef12df641c42;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ef4a6c623f61be95ea879486d922dcd111ffaded0fd0c84a13b11757b5daf097e2f65bcd8fa1f833ad9804d52e47a152ab800a8345eb8bef2e2ddbb557a7a8bbb9851dc3bd401fd16e4f14a3ca9b80fcb12e27a7941a41b477c1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d80046629b1f82433e88e2991fc38cc79bd630994182e615cde49d751a2a5b56448f3283f0f3c63aa9051466a60f587d6af4d4c0e93ae27a152e688f7b7d7e8fc630a1d0a2c0134300812001ff736737820242e233e9d46c7b710f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4369a6de699bfdd3891a6182c1ea0fe4a1bfb61e98556e8433c867ea3a67a97ec31aaba5e7f03341514936cf6bd02f09d82b2bae171591ddb9f57b82ab11192e0b0b6c7056eb82449e20e4a9597866a71787813b1552d261e6da8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc3025c4bbcf6a08ff69beee072e5aaa2c09ef590c25ffd114765264a30b537dc8b6b76cbcbad29007cad67ee19a0dd82f69470ea919716c0ed6bbb0ba6d7d3cde2af17f1a31b66ef18a23515333429548a4a4d54655b3c8aa3b2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf38ef2974d6a3a6379a0b93dd43c77192ad24a6169ada3884d07f14dad240548aa284fafe14c5007738c97bb0f645c4a57b7a2be7232c8e387b1b45b05b8a81594e716511f13ba895b0c8536075b390c5b02c172bd169f2d0af1b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6db41016490a55cf0b243b258209257c0fe2e4289086ad36d5a266690efaa79029781c0ec4a155ccb60e416e6e330f48b421bf16009569c055b6efc653ea0a3fe0d8d55eab044a4ff6003f7e633b924f7d5ecaa5deee434898845;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h131724e8a0f2586636dce8ce40c895d860162fbb2d1faea22327b116dac6345b2ff0d28d0fa0b348e3921ce3cfa0fabd5d2b2e494b04c017db5a6e6101fda1e5a6923efffac7b24cf046d7eec9116984700282b6e63b5dfa0da2603;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185dccbcbc594dd9e9bc0f46abcf174f45acf14be871f1327b41674f37c45aea0aee5ce03ffd94b1f1dd06680b2a04178916d856e0d2ed11006ae9ef9f8793aecf2e26b8904042915f281f48fb42fd08c4a936f9c2dbdb86ba01a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3aae5e59ade0688bb72e94283526b7330cd886773046b405a0655c10e6fccaaa485119d60a28fa65f64e5b4b51e1517adee7289edf555784d24480b3f2486b2156d0d81634dc0638e57608bae9e91880390cbe0871938035e243e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h181ebe55172bf2c65ed8994f166c9fcffc07e14e0a976de97b4f2e647948b3a044f19432d52f3ed4a3ef7314f3dcd49559b258dcfc989c5c4ce4579575b96eb113a8a3e18e5838df195b7eb3671c4e738f3c66b7039f504d38bb01e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hadad0e6728364ad32e9d6e8f3cf9ff76b27eb8cc7c062fdbfaeade0b5bebd7f902d6475b21ceaaa6135c84376bab8d5ab77e0acec2751a73059642eb7dfccd1e6c380ea85e3ab555902ed8045a67e94360a43c641425762a7830fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8de54b689e922643f5aa81f38356a17286dec7ea86f2f57e674766b24a14fef0d38154e232330540758c75ef96bdd79809ab50388ed75d54bf0564c68ed1a97de4a63dd08c6e69d7ca2791f871a9f785d1a338578fab61ba905c02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bddf54f9e3c4129ccb882634724740b15f902290418f4c550674cde7b6d7a378565ebe6460bf1dd4eabfac903bd33bbe63071eeecc4fd70a67afae07d10f0538af26d9e763c8353694fabda99181ca4141a2d4b782dd9f332c5054;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2753bb5036ea2b1ab1c74619d90400d555676f4355bfce787cf23d20eebf43bcd914a82982ea6908b18134d683a6beeca18f4fdcc4c33bd0a2694a12f22ccde2c75a35059f82d6f3132e3a5c340a7a1eb8d21c958b3a16b03a6f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1932c8f82d0b485abbea97dd35df7b744eb994b61ef32d864a743dc9e628de8dd77325e576b50df81387e8298b15a10eb0c37765ec6c5a36d8b387c6729594191933c30d943f019bc8dbd6be61a7da2d6cdac2a8be673230a5b899;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7a1a095da1da03d3ea1c78c7929e3bf9759175287456faebb370b1649410f2c5984cadb67f916146f28492c89ca62188cd28fed372327e739c242a20409aa946726d7bbb949db25eaa71995af6bd67b2e9dbd924c6bcf1443ae40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129f7b99ed7a536f9b3704d311054ebfb63a1e6d7acfea62ea71684db8a1bad02ee9c38ab1f7d7235887125953584ea035186f36cb97f6647ccc97b6dcf447ed4f6fda89501229522e4a39c11e76cf18543342263868b064d5baace;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6626d28cba11e4a6b5310bca9bc254a9e5322be2fff2c8daab36932b0b951833cd1ca8a6398bed0d297ef40ac24d16ac9db93b7e4d03efa078705dcf9f39be7a668bf7cfe700484f22c8643aca2e0d349afe7fe7542a8e46467f0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157a9464c592508cc590e215a1f7f8f09af3d07e6b1e96c2b9082815de21d5e3d21f89907c82773da73ce238f9ee1887d975829cf2ac4b7d049fad95f650738e7a6bd7fb77ddfd7cc5aa8ed4671601e6d3c0867b987fd066f6c0772;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16cdb0c5a2a7e2537b7cb221d7f5a595a8654b16216379a5d3ab04b9d174b05d1a71d608e3d33ce3993ee7c73f4b4cf8fb8497d7a11c644319dbac5fde7edc3a62a925a0d12149d408b5a57c0bc6a06966377fa227ceb0bd6f8cbde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90c3d675e367326f2538e914d4fa4c78c6176f58f329d07fcd61fc49fa06834bc0a596a52b0bb88d311ddff152c0153f40148bc1ce709c14fd68e4b04b163506a36e98c4d5998f0cc134a68356bea4ae1114dd42d149b65d09280e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b645c10444dda47a72070cc2ea6c4937baf40e317b62f5de0b6c58f1acae47af9b5dae4b2afe487ab2c337955ab78349ba8ee0aabdf5ca681e1e32d7d98bc3a3ed0f54d7860731ffd83693abb76f5516acb04429b4bbc1736fb728;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5428260630164e38ab5e36e6f7677081316f46036daad1d34ba6479c28782991f34307149132b7d9a06867667c89b0925817ef2c304b5fb2f9f8df18c23aca6d71b1c82334b10d0c351a0d8091777a0490017f70f973b7ffcaacd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef2e2b4494f155b8252eb3a79ef94cc74febc580b3780f27a1783c610af3491f77913325f820dbae19717c93027177dbb9191ee1eea93e0c8c17502bf7774a37c46fbaa348111df13da97135ad3af46b4ada6be696f6ced27a89d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5755fe0737c1e21c587c3848a6ae023f0c7070ff560a30ebab548d981af228b1f2ab4be30b66fdb243facc91488e8207ae1b2040413734be22d369ab1d4c3dce6591d5dca0b6db4a8e0696c0f5297dfdf48f3f1201773e55bd073;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b587064e15842a4b675610d267230943fa3a930f62947cb75830d7f38854a0c6c9645498a1c38147977e81a3aa15765abd9b2b90b25739a55a61fb8a62780d5c0237cb0b4f9078513e2ac7e19e0d9e4c3acdafe7a5ef16540fe8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2620b3f74c182065fd4b7d7fa063f766a07cb71ba9391e9b5a50642c409c91d2e461766706b23513ba443cade107b91e5b4d9aa65602c53606758866678ac486173cc4da36a326a39375a93d6d9404c799134cf2b710853c6ec39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4212d4160152f776a6efa81f4b6102f2ce98f5af37850bcc75544cf0f1457eadb6de97dc1887caf4dfa97fcbc4a0053d0bd25c112996070cf6710d122fb00a4857f6bd5d3437a2594228d5fa5230e8481a908be06c31f820575238;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9f34a53513ce42b59f5baa8e94574f06fd660a73a2e6b2cf9f10759ae5edfee791d4f95faa8e1c416d517dec97af5c83c18b95f475b3ce8a615749202ea01905d8ed2bcea987ac5c8b1351d41f770e698823576f75eed0a7629c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h963ae16c979c8503e0649ff65f5537fc31520710c2ddeb13e0bd805d0e3eec7b483d89ef7b17347af40481b572f85e06e9a4a7be6a1695162fe3f4f573fea17d2524d2fd67cd0fe287bc6cf60e1442d6d4bf53dd3244eeb094c1ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc6a8f9e66cf341e8f41cd11404d22e47c971471cd81506fe42e2fdedf4c1b4629f184e8ced914579b95a082773f42a9a249a79e840c49077a019dc80122ed30858bf40d0c8b7c98e1a39a397daef03e9cc8964de10b77926f94c12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h161b8143f7e3f09d3ddfc0e78af4c49069c610135d4fcf6599c5dacdd1fa3670cad1e7b166eec43371ad0890e290e1c6494cea090e95d5bd1d2efdf9627e76aa0e2d642da7d0f2c702ceaf0f74e26e73449d293d4d968896f2f6b91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb13c7135e0e086b9460a4cb455f203b537554c2247d922a21a72265a7f5ee6392824437a058b828ac04f65c0d023b89abdf2015135230dba73d7d229bb48b50cb27e0bd13a936f1c53a7e4adb90974347a5755fd2a48804b3c6e0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1245f9e6c7f8ac246e71924ccece0167e2e41bde0aa510353f1903bf40daa4adb95520277da5728d6760b4137671369f0a2e5cac3c39d07afec2e7cb1ea12fe3beee313679530ce7bc463e418a9285ec82e19c6cfd8871cb15b4ad4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfbaedcc92cce1a3df6c1624479b4e960c9a8933db09a0a9af60eec82f46261a4b8880b39a6f02b63208b5908f255e2d06b1ddb9d2ca88cb328df3449a619dd84ff5ae927303af190dd93c6805dd48c6b98578c1c79cf6749dfe0a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he34bb59e9c573caae1038cd7f6d5ebbc0c6faa01bd8b4b51489c1bef47decd2783090e3917cdc4a14161de3fd469ceed93fc868cc4e2653c8e91817f0cf7294003faaf645913fb9fb9f90174fd3505095a7ef2011837a8a785387f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23c5b1d3ad2bd37966ae7557696c5d87c9ddbbab7c9b5f06fbffd6c3bbd5319c96a6cc3e3b902ca8a2e5f7ab402a20a1cf7a79e8da7e2cf9117f51b1de49e50b2f80f89781e3a1c4f578b376d3e1f363c1be008081955fdf3ce2a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab469792dcc47ba1514cc0eb6aade5140e38f1e852565683a1780ba22a3efc595235ac2d62cae4ad63ed6a1c445c9904b036b33b546af6e395a768a4ead35f1c4bf28677447afaf1fd1d4eed3cf6140ac2e58ab14de75a18dfd1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h120821c321aadb63f3a599dcb08dd601b6ebd413f8328077e699b2db95b16c75e23f4d6fecfe13af9c4c48829c733bd32ea275a423c2b97248791a46b936e67d8112c09b15488b793f2450c239021cc5d06e40dc32ea703b51f8c0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d2cd73ab5bc1115f0502e2f764baa9cdf0a6648724799d54d16b83358014a9badc0d71bd68301ddc12979d495e9acf5eca99dd18eb5d847f8c5e0a101cb1c9782431a40fc115f39646476206ba186b886caea7b0a1b18542c9438;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb8fa77735b9a858d0c41316808b2f47003289343b974e5760869b05f603918015f2ea01ca5d4eaea791d20d255886e730073d0c2847a67c7d02d261a5d2a18a955b5aef193debf90ac65c75ae68f018e430d888201d6a5119a8bd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2a3d0b06bba07f8c23cd48d7c96aed7cbeb7adc45bc8525838d7709b041bf0acf5e74f41ed6f4c5592382495d8b126c7a615650e04d9e04fa02d0aa36a845609ec5000abb9aa31b2a2b7b85fe1ec963218825c8de1812541a58016;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6aeb1876a99edf2dfd32351a05ba93802094aaafaee0414aa6eb25e54d156319d41570ecdf7e194cc82adad9167b944ed77b8b3cf4bed66b7dfc90a077a15549d9a812e539bdf072d3881fcfa70528e22e643aef5c87a4e293db0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h140bed81900770dc18b2937afa84ed26bcf7c6453b2d526a4b3dabe76c6dac65c4212f37d46ee332a8f6cf36f8f898fef700b6f54e1f73cf08717db159d07256979b8896fdf228ec6b38bbbe2a0e3b35f6f3b5e862c528c23ff70bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2073c2d4a87ce68e3891f47ee6fdfb9c6fbb78163625aa622b77bd4f5f7a9a170160853a5bfc5cbc3463df6faadba26275116b2d98660aa4b4353ad3ed5d2b6c5a9904e44250bb7212c2ac67f55f23b64689ec78fb1bad93b957a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b365ef5a3cf77d1cfaba06296a987bc7aab72dedc3a8cab52a3779f79fba1962ee9c9592fbbb6b9512d839600e309bf080f967ee31132a188a72c6d628a7c431ca032906a2424a294819b97f48a1f59fde3e9c0a0209b008d93df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173ed5648f3a99e8a6cdc46c7755be89a1b6f16f90c10b1d7fd1208a2199284680580712423dcf63d15127f03fb44ed81309d680aec8e2b361c5c8a4efb58edb3b7160b228637da66631bb223223f1a9d65d4a6925a9bb18e26f19d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1927679ac9d0e9e27ca2b14039fa7b0be70f9380e3341bc037ff71a198d88e105337724766af055d6becb3bd1d98d245a6d8ff22bd8bb14c036cf764b6d38bf7059975f7f13819719abd510a4de3b894571a6a2c6e6b1ebb40ef7eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d9b2cc4f1e2c6f40a5ab1acfd14e403fc325704d5350fd8b1469eba2450fe40b96dcc9cad0a0a1ba9e362aa5198b0a05584e63eda1c5d42221fc2a081fe20a389d2a6b1765f2cbaf48a610f89eeee4d5d2bd1391d1b22c84836a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d8aa70be488f1fb7423487e3f461e7cbb1af65b5a06e738a8d1581f11542f0a38845d733ec0304717781373ade65664b4d0d96bc2b9668a2646821db59dafdef6292bc764cb949141cc8042947ef463068c9d5b4816b9ce8a03415;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f730c5cd8190a04c3f1cdc8c1f960ef3f043a91a2d46d8bcae47d2f96d1b19cc77ed650c4fae99f75ef25b3a287f2cee5226fe7a71c5c9d04e67669d68cb013370ed0f54cefcb10e42f94c4fe496f0a4df9fcaf5b9232203f8eb5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f746ba450fc118d9d6164d9583377d06a2aef6995911412cb02e76f75aea4514399293ce473ddc66c136ab85172c812a0976743fd9459b24f39f6816f3343e4fcf71e1f73d0de561dbcb5dcec8d78672f92fd7f89a8d7b95703fe6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f60cb505172590a70155517becf872f7db70b94bdcfa932ad673c6c07539bbb6c30c7915c4d584bec5866f1549df71800955b0434d6a5406cbeff08780495e508fd71b2d698c0037817c782b426f5af8ed00fb9168f679d08d043;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e2c8ade2d2af078fdabf70368c0ec5b2e06cb4cdcdf94c0c31d74f211e8bc8599fdcc93d4849f6a57837d7b23e466fb60fbfb4403055722170e5a02948fc5a1854d9edba1862b6b527c599ff55c377f2f404a469f88118a647f75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb8ab360aad249be45bc281707879393f3a95eecb46f12c1c5285896283b9ec6d45a339ff32fb78841184c2003d22fc1033614ec3168c160c0f889d01ee1687ffefd741f1ce5bef718f237c1396618f76388f05029975ebcf1873b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19311b4a49524a84afc8b71afa2fb9888c31795e8c0d53e0ff2fb6a59b41f6d8d7518417c41e09c0c637e1144aa9e2981ae32b277a76f3cb4ceb10277fb97fe8dc1d00cf3db35995741f50c1d7030fe1c1b9941e73edfdab5cd6510;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hac29bf13a3b394de702d10f7731f8cf527c998cc7e649c992df099737ac16569be2fdbd44551b4772cacb53b6d3f922c6015990270eddb3ca136303d36b204eb5c015d604c4ddfad9d31512d2522a83982c003069e717efe33778d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b1ac7a889527d4a73599065d6ca87cd48b162fce384ded1db2125bad77d6dabcac77e9057f5dba5dd3a74d9eea12462eefd730dd40811ee5649988406c07b66cc9012469db51f100b4ae1033e52c29368867a328da4d1509b47847;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe63245e9e26d7bd03a37dacb88191103be74bdfe2488275328596ca8ac8f3616db8c7d6db87648c8d706b6745091cf9b00a496e91fe396a0ed6b0d5483133dd791f88850e301cfdc95391928e8c400bdb427cd7032b323dfa27eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d44fb7d43d02b316ab8e15d4b7c13fda85134fb324c09031e954867610eda3646cfbcae1bb6ca4353c7adce43de982951f9845bc4df7e32d7b591eeb2d3eb26dd71e0098800be74942076df3d54271aaaf2426cc1aae33c5250cb5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51712f52bf6deda0355445676d8663edd71faf7e9c8121025c5a4b06da17d9ba9fbf41746b13bf22c576e083f23d39a671672ef4b72ad379d5a09de1d242222ec150008fb6413d8872437ff4ee43244a0e399e7a0fa970414e13e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4ac5449d5d8b977f98a274d2ae349af1a4707a831a4d90f035a05480d6dfd53d5110e45ee1c33b7edc6fc49ef042daf489b441db2f4302a8af03e01a1a342306e1d781f686199572b108526f5b2c8474d265f9e22ac27cd687666;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h390f451fb86e991a8041b6ccef7451e5e282e0f93000d8713f0636afd37d154c0c49d7c6402c6b63b627c561f39d6a519497638cf3944ee455cc95aea7aa6a6763bbd68cfd079579fe865d09c7715060cb537146f73903148a0be4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h165b7460cac2c7f6e6f8cf1e89b7cea7490ff457521f6264273e1f9e6aa80d09eb3cee358e3ef4aada0fa922605f86513cdba7d17d45d21e75f24a8c2ca627ad6fdd663d1486f2a0cb2e12338837de1f5490653c95530d5f3b62e6d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36d7f66fe9e952524186ca66a5a924e7ab068593d3a2fc5e7406ab69f85d8b8d3d9bcdfc6c9225d6b1a03817e7dd20402015ce434496c1575668d057afcbcc23ba9e452e1b1f3d2fb6904f8bae80fc79e7883dd65dba6418a90c9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f440aaca1109a86feff5b2ad36e0e0c263df16821c37938793dbe9b268c05598f888e55cf976aad3eea3210f50d0b2db5c80a4ca2e0f4057909822a596fe892f1a975665dcf4c7f1ed9ba7c30d39b1535bbc1c48d3b78f6001aad1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18761c6720861e7ecd574fb873cef6bd8b1d15213dade4e3aae70f31c61abe7aa801b836fd3ebdcd1c681e788224d173540d8f859a90f9beb42c7979de4c5b3069fce247652cee5e9b1e6762ac493651d32627abef9ee18f87a11e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4b94e5e9f018886feeaa47c22a07ac302d5560b6c87076bde21fba103f548334d4516a3c7835e14ceb7cd78fbb6699d11ed69e88f80fec47877ef9e24d2a267eab98f62bfaea823395cfaec9a8e767af20943e5fcbdd91fad0bea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa49fb4e02937cb6bdb45149a0adb5b49eeb0c3ebd626649bc8827cb9a594eb4fa1378a3b3835c7a2e5d31689c4452a43b45809399e51fff0d637b8df9884f7786395f7bebffa85ececd1386581c6f40acd0b504ddd472f907f433;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177b3aefe2e8fc0c5253a3c7beff486ff80dfc67aa0e9161bbbf5ef07e8759387a9c6a29db45eec30a1f52fda5731d3f3be81e87f1447d9175857c24ee69605e1b8fbd6806217ba7b297dd58a31e016726e488c47546f59c40f8057;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7fd17d65b4fb93e093dbda5450455c10924aefd8a498ea3e02b446d185049a04ca5e044fc174c1467f7143fb5f35ae3c4b1f491d7d30c4f87438992e90f7f272b67463a8ea6e795ec462605937008a0b01105c384dc3a7497f35f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137311aa258ba1759f1e14282331682fe09e48a9e4ade7e602bc3423c9464a1a497f2d8058c65cd59ca95ea497478aee4a0a0ba21f09229662aa54c67f103f04a7ee033cf5fbaa052bc914aef211c84e1a4e3b6512dbd75442e87cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35644bf8ecec25a27d0ef81c3ef0660603e542634e6bb709d324ea71b3173680e4c987fd993593535344d3bad0b8730fe64a6efa3f61da8f9cd216a85ca3e120011e607f2fd0fdec0bd8fe7c478647a864eeb75e07ce5fc12e0c9d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10be38ecbbe0dfefd8827992b988f403fb63e542c09d503845d4e0d340f4d1cbda319e29327837339c251972efb20d56d5b44e10c6ce378c52cb2e3b70ce178de33ea1eeda980def3cf91c6842243f0549ede8c5c4a55ffb2a2a749;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2e15ace0b40588cdeca833047dc1c937678371d9e3922b1cf70f8864d39a15e9741e57ca2c9310928526671a306da2e46b4f35232f6b6215035e152680ff3680b0f9922fd2021ff4076c6471ace20d5abd85094fcb59969fe0bb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5326d0817fbcbb65197aa567dd08f5690f2a7b2312a10a517dd33076c7deae4100646cb0f824bb5d18d0516a954a8de26da217ec38a2cff4e563ec6826df079ba54eded40513ad990f306d5c000b56d91cce6ab96dcdb815b878dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc0695e7de0728954ca8a852b12495504b003ffedaf67a6d8fffcf0bb58eec1fb90bd8b724e3ff7de6afa342c8e429fba3bc0ab64fe5c74cb611bbe6241079f42f9afba549708613e341aea4f167a50107425b10d043813f9523dee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d196b1de2fed321c872afeaadbf2888b20e57ac0ac6da1bb1549d86cde02ce27074b3f3054810da1b3f082f81e7af514cc48c0de91298a1d2ccfb5e634bf7a00648900c7e1e4d5a18e06b0b3c9dfc61f49c76e6aa99e4cbd3aa7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb7083a0afc599f5bd2967f1c707570d24556e7448ec92970f1384d59882286ae6fa0d11ef2c953679612fb528144a252203593e011c35e917e3ec310136e78d0dc961920fe52978ce4e09f3a8211abef8f2aaf26cabc40945911e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176687cf6152c4e2a0785021e62423b10f92d8b0b25ae5d1708e46571b8274bcb181734bf10ecf14af9b4ec55e920127f77ecbc4da22be47ada5bb3542257be3f923446b617a05063b63823075a6c84359c73bb90bfa5ce0226c03f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f28d63d3e4841c5ae728d1aad551f9cec6d5a07eee95d2584aa118becedd1a516ef8b7aff5240a31e58b33d940f98658926aa7b6e89150a461644534de3390c94f9d6128732e9fff9a15319d6bd44a2b08a928e465b1891226da86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ade5d1856d554983719e6aa78c3085a74f1f3e966b415728a4414be405ced841fbb223a25777bb2b8f307c47367b9570a9d3d4a1b66c1a0a0716df29d88766fd6861d5155b113b7b6614f0b10f3d6d0e1a852c0df1d542273499e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9f675a74ccd66496a8f7c9232a6775214000c6c7e2528a86335b9014089b0c67600477934cb58ea396e56e7d8f166ce50b94d9e458c17f33c867145fbfa926f42120893e7389032aa5922b4e2deed8ae728e5f6ed3bebbaaff021;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1627900889aefadc48d65d934054303026d517d1aa0b5192e3419c12671126263ba25c4830985c3f52ce36d21bd7463ca9ec285f06139fc5163566c48fd7fe5cbb4228e84c3162efd7f3394c561e10a103b8e041dc34572ca5da22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h559c5af2bd16422df014d04b213e96284a3a731a7e7fe057e638c6d75ac29d26f25d6f25083fac2a674bb5970a4a937709d95a764fb3ce6288280ef7ac05401721f7a344671e0ed35880df35af87562a7c75ab24d1b6df822af074;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h323c6bf8a75275eb174a574e1f879ca7d6e9ac0c99d8d1950cfd3351e8f1dd01d1383bb51504f3c8b99f5f55c1e4b82446a9c004feb4f7d097ff756045e4d2124b12b7481fc09ad5118d8fdbcf802f1ff3cbf6b4ca9137848d2e9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb9d00ee1a74d20f5d66fd2c34ba05329785a38155041e300d8bbd887c40bf086dd19c4e5833682cd817420ff37aa30751d63a4bdd24f332572d2250cc58cc0841deb87219b6f82140d8f319ec34a109bf649db4e3535137980c55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcaaa0d109834698688b96cb6f3a22f308db43d4f54befd2a35f67e369f042124325c4927b05aa2f6e9022ac1bcd5bf35e5cc5c17b4d657b82347133e4b02b337c9f3aa0bd5bd47bff1067088c132d29b2ffef885f314b09a660dd4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he27c9ce149ea1f13a0889e0c3e2609d7455b17eac77e5e6a7f92e253a99b8c103f004c281207d4d24134453acb112962a823a50ba056b9cc5f7bbda67aac08cc4278591da7c8d26f062fe2b21b1bca2fd7f7481b9de3cca836d981;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heeccb1f6f3292f57ec4e610ea302864c6e00ede0b24299e6e1f0f95045acf64c9372cb1c0d56ba80efe4d46cfce7ea9a9b7ecdf3c5d05ab5a2f478f716c00846d255a8d4758cb59806f14895000d0ab6cc47498ce642682dec89b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h781973709e183de7f350d8808d242f32b9186d9220c38073a5fcdc23ba273800181668ab664b5576c1d03121d505444d3ac7858e156753363fd881bc1b1d28b14c5d30f38aa56e2ddb3e7d35e197fb20fd267fd283b71ddf285c7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce0f897afa2530afaadb1ed8f40ee87a8df98f9d43edd61d74523b066f6e8af1ea55f7be9f5c7cda67ce463fec16ce439eafb68d1a3dba21345f9596654101df6bf9c34819f2a63c86fd42b75bc2a821eae393dd21dbd2c82d5a99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121e73495264d38e5441818cce454243c8ce0f06dfb590d6162be1a35f43ca9e65426c2fa60137831f0fdcd7310f1dd2b8ba3b5d48a0ac90d62024be27b5fbe9deda43c176e6338baeb68a5a91efb1b8d8687ea3ab2dbc9ce36a3b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10dc9e37a8c8508e9226c15ba4f31c255cf63f5126ac6403c6430de59029ed30b8c38e2e9b67d857d3b6fd5dcb62541ef1dbd2519da7cc5ca650d1db5e37fe0246c2386a588724cca1cfe49082a8abb7384fe4bd11c142bbaed940a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f7ba42a83c16ae2b6b1553c94555f3c3ef399c2e1ae982efd8fd002e4ea1ecbae6e75df6deb0f738d228475790eb2b3dedebf709bfadde04fcc8bd207a33f1f5753aba470d33dd8f486b2cf33b7dc830ab27580cb08fce713293b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188faef4fc316284f2e8b42fd3966574456e6a94adf14ccc681baf7483abfbb149c4a5f2946e6cb2fa93891d5fe6eda7b2486422e7e5047e2fd3c04f2e89521012bbf8e06502487b98b03f15625dc04d379d1cb941eed7515bc5495;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89da2cdacf6d45ad85d86da68d486827b4f1bff6193522b0ec8bb46b4278f005d71e8697f5fe05a8a7e611b40e41d2d73404b7618c302c31a4a06cedcdbb87192efc1fc325c546744993967fdd78eae8a1729e5c9a107843c885be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b0e15cca27e5acfa2ba1beadf899753ac6388c8734ed72bf3130710bddbbf1da4e99c79a318bc6917ed72dbd7db22e9f8bf87b41ea5209554859b9ddc6118beee54c4785538d9b46e33867ab45d9b8f27961c58992b00a66fa137;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d98ae8a6fc15a4ba022c7e3f72690e3ee445532370da9c8e254b3d6c9b038572f00ff19e4d163caaa1a36cb6fa7eb87d244213a15d7c2ad3f3f5e7916b7afa600b5d31d3d0d9c0e2b706cfb7b2f5efaebda73667df960b3d24110;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b427d81f04d6614998d7780e48130c0bb15f386e467c91556c07716039ab5f5cb93e804381e7786297772d132927b8409aca7c8bd0192e58cfed8b7bfaa31bda81243fd22267016e45f45bedfd79674711563b6b70492539789bd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9977e27893cdefe54f5302ce3f72b7d285b512bcf498fd9770b58b6127471ea43ba97677ecf511e35ecd47d8247d65bf4bc28001910fbb9b542146d578a29ee72319ca27f327a579a5503fe5b4d8dce36579ebe11dad1813bb110;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2a29201ae73e75fb474dd451678317b6e0962f50e764b58ff0658b8769e94d4485783dacfbf06e72fa9330efb1d2e3e7ff2ff2e24bbef603341dd899cc502143a1bcc61e74e3bd3f2678603c035ca8d38fc9d58943ef14a6282b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf2b025ae5b908790e4406c16af35b2b4289de4105b43c66618d3624121e32448b3fe4cf2fac111e01d28b4e7a3d75ca358ff407fb4a4ac319888723c12064a2a9bed50e60471075d3545ca93e0ddf4c4701e6c4302a5b50684984;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7eb6ddfaf24a1be5c6b0452f619f692ab1a704710a9c392634367b33aa313d1085c602184bf42763a047c2d631bbd81d4037c9b4bb8e8830290fecd8f598f9b8745bee117e9af3ae8baa75d2d97dd2e3e4ff79cbee3b7d3ccacb5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1513a7d8eca15c6889cf004d94b38ac6cf74f3a6947d76c8913f1a4f9658711956c8a26a123744f936637451b9ecb6f0b30253d040240034091a45ef934f6b9cb1b3683710d1716033cba6434be99110495684da5486caade68c5ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5fa95c0ce256f010e3e8b3045b3aa7fa0cd6b2aac75f0af6dcbf7acfbfbfa7fa911bd75b6247b8eea1e0b6b951ff344abf84652744097688ac844753b0dad34467599de92400eebab1abd0edd3a7f0869cd3662e9e56aa19dabd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbcca1716131e30e72e0e1be4b8992814218b0c888a32aa9a3fd492fa00635961ce80057da416fc4e6b23b0f94031649ae4708a2d3929f6ed6731ec62e14ea7f5e3c36032545cce14967fb41b7bac486e28cdb5f0c71a85877a4b19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd99e462dee432f513e1a7bada5fe0011b95bd56594312fbc4621cd14d16065289c014ca374f3b7e571f592770bb4729795f5cc94c792827ac7808cabeda9cf2ee05c461cbf9458c1e824019b0b771ce5eaa2b74cf78721704ad586;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3bcc179673846db80b2aeba60be28bbc3692e7758b2d8e646bc5599e2ef5c9bfb2b61f5515e369c915ea38b320e26484311d4a9319450fae03884cfb8c76ef030cd150ce3bb7847b8950b79fea38d82aef996c4547a52a54b3eada;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a6bf305d88d99d1a2b264c08b0e46fb6a6c39163d84af5346f0adfc91e56221299eb3f6023155a0b53305f7b0ab5b707c56fd90bdc732f308de607c6b5d8e5777454a775f7c05bf10999c3e782829477e44586841d51ff840a084;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d276af8481c8120c7190a262826529db0c0edcf68674bf329259c4398eb6622b695c02f6f3355f56fc074f1f9358ca308df1081bdde3e4f111b8498203bfb0c33c369e2a44c858b278ce14af8919b5f70837c6b445f27972291a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ade1304fc9567934232b682cc2d81c1b950760edebad4b49540044f4d83e5acf3a378cd98e827ddd009aca19db19677c6000b6efd912ce0e0bc4764ba0ec513b0c62508449c8af2775b49e51afdb7f047344b1dd5d08663f0b4e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188aacebec47f3e846b8527463d4a9ae6e18a1b4e1761228b95fc431a9f573f9a09a83b69cbe458b719f4fa170de11589df27514038afd6c8e2f97e76104db4cc630865dbf26ec93aa5c906d6e112e8f4db3bfe5640ccfeaf98aa64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34447753deaba8ff01f2c38d2ffadb00818798e494513c4979e00dea723ae019576fffa0a10acc22ee917675ba0cdf24e6521f2777daceef39e15c8bd39d361b81b75cebbb60769330817085c812ab69b09a2a3dc5c04dbcc4f6d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1105b903c76755f74333763de9a1a8fd382b52b5cc983824d970d649b57253360e7616d03b6b553124cf9263fc25f0692521385a68cb75115984824f178bc4d46dd3392270f795c522a9d2b101c10257cd16c5cf5d40a9f24b6abf1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3274ca75b068ecfae0f025ffd6c1ea6de104be4673bae0ba2ec45e61fbdf9dfed707783a0924d4197868f73cb24e95dddc54d9d53a3b84adaa5179daddcb3c12d992464fcc018adfb8689deff8b449826098eb01feaa55e2a208ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133351cb3ee273e5a4c298d909280f9b63125a49882ab958567a6506b44da99493c38d6f087a2340ace3fa3e4aebe96941a84f83d5e8250450367d68cfb4b6dd6616ed9ff534c401506ab7f8dd3c6360aef10034855792018db2c5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129ded747281b7248bb9e331e7850875aada3a977892613cda3f85e4b44629807cee43391c1898467d66edd30105dc31af1266df3826152fb150d44a61e8bf6ad9bd71141c61ddd05daf4e84c541adc9d24ae73e5f28db76b790297;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10deeb1ebd3c59109d4e7315508ecfb375534af4aae467fde04081456b70e7bd16bdcffdcd2ade6061274a6e4399dacecfbf1dd1a0091bb5d02436a3f61f77f76de52dac82a9daf758927b18184870dd935f81bf5423b5414e78634;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2805bdb36491070f14596b6e853a78404285c2a405ce953f714b014d5e5b4fce64c7fdd71d7647e7ba6e0e67b0c38d0cb65855f4430efdaaf7a21ff9ca09e74ef02869ced67f0ac18a7ebc36e9b4b9e5fbc91fd98599b7160f873;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5f39c947397320f778774933a4103b475d140d9177334e2520c7dc6bbf7c375e4aa861f0ce6b0216346b5ab21bcf6a2057300526c3d488589b47012bb9f9916b4d6f656c4f7098c9061ba11efe19d4725161b9e240fd91234b69a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h774d66b8716fda482c0886ea284712ebf7fac82b970960530aeed74db354c4d30eb0aea402719a4594da3b2a0b32514ce52a1f7cdc66c87f1337f09811d57cbc20fed61e56c1855da12931ac095a29a4afe6b7cec70d7cc13e7d9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c144459d9acd2a22f673d8585628275c3a28b1d2fa7c6492d244255f717d063371fa37d1d739474f06448f448ae240e486190acdef6f9bbdc384e0418fa6ca1091138652c79b927fe311ce2a19b15c23c19e56dd2b7d316f4c21e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h837d5062d4d173406a13de29d7a56ea542348ee09c2a640b422b47c1070cd12b4b2c1fdef2041e80fbb8b6343be8cad716717e3f364053ecf9eb8e4af4a46a73fcd4ac4c1c98507bf416e89ff2b100507995649d0b3e0bdc29bb6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15abacfe9785dff5a57439f60e6da673e88b8ede39713d3346bcb282a6ae28b251ecf4ba1b17983d8eb9c914730e35bbcf5de18cfca978ee8f6482a44b0f1f8b9ce6ed1051a04deedb342d20ab9100d8ee278263766e79b2527463e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb4d0d92d2da6652b9b8eb87c784ff13a6d1fcd2101b489b40572fe9df2fbf88c351a01330c63401c6670dbe04c491dd82d68a07736ff9206efe82517efe2c37c8461f391a06e82f1ef33999481f632e4adf82c480c388365803c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33f46e7582cfb02f1b9f88ea61f8356fa7f313a4c0361931d50f0432143f5d8e58297b750f0b0cb3d6f1f1acd1c26cfd7e28162272f795229fde6d2168ef4bae444c6191b2890d655cd7b5a381485eb1ada892b6a7b7986e919908;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7cf90059ad0ca55703e9a926b97f89cebbe5d18b180114d64b2fb37a6dd2488a815c9bbe7b4da815f53be201ee25486fd97e80eaa21d58c42e2efe130352d235253e1b99c12758f55f95af69c986dcf9bdefebb33d793c775f3491;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bcfa03e5ebe72c4a6033061a96532dd6b8c87ededeb7a96f5b9f3e867fc0a372d348cbbbc145327ae5f22859d28cfae8cefae7041d1e64674b3ce8e6b03e25a3299f7a6a615c327979ca761376e6b5c210f396917f5b94e26b21b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f56cd5b4b1138158ce4195c3d66e575d9d554f1ce5831fd4a37f83c3569c2ef65d18a6323dea95c5398eed42c6263c1f3abfbeddd25d9832f4d9e553827bb90f86bb3011dc831fbba0674e7865683323b787d9db868b144a1365c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13db05eda70e80c96428373c9e6ac93e25bb95d42a466e85d94b683bb827cad7fffa6c116b19239e549111ea8d4475e22d52b0c1d57f3869105ebe658155caaa5f21809c3d33ee89621a4d03775b93854c959d6d87beb589fd694ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb926f83471c741f724ed9ea707d1f19d547d6e03514e71255bc1c3599528e75755f9ffb671d1b4bf042eae9b70a6354ba50a761ee9eaae6c84332e4fc388cfbea022ab31a5ba3e94669b11803243c8b11fade33ed43a69422b96e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11790ffa85f96215490cfd604799dd5f08b116e31e499ed259f5b6b9e9f1258a64075e3160036308b2ba0c992c662a4883db48875ba169a9c42c9b62c00c0d2d5d29c2f3ccbfa2c8cfea75fa3235c9b903df7221537726f8bc67a6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b500e6443d2c53b81ce5fdb1f644fd49efdd79ba5f8ba13770f16c2bae8bc750011016fe09a72ab9b1d10a82871fca613ccbd4aceb02341f7b223ef1b57bd282eb90841926b41eeb86fd153c6f2b8be7146b0baa123803e9acb102;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1c3500fc18975a233a509cd028ed0c27d9049d009c9819fd719629752fb24a6e1a118ddeedd166e2468152e18ea37a3f306f56a5b272cac88c1e6340028baef37d126e723fa88f9c562523a525e191ed207df49e4b24bbe22f3c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5174afcfe8997278c6426a1818ff8d9aaa4473a242ead71fbf891c6c8d57dd4f94ef9b6a3f9e7371464bf57c024cfbfeb3e17db39f34f102cb4f2828ed39fbdab9786f784d5937334c88051949b8262ef827fb5e5f5df47443343b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70d2a1f167037e97c001c3ea7c1f8ba64142db94fbf0f3a6516629f6f6c9c1bfe6045bb76ab949973028fa6b10069ef2a8811323892aba9f6fa9ea7f53d40f0a08d8f025746c88ca71db6ea25154ae86337d10ef9fb7ecfdbe831b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146f6163f09bc69d64f6e8ca24ccfe7ed77e740fb5da18907895f9e15c2006ba70df6d2a3cdf57269a276d892cb639df1e9c053c7fe1d8dc420387b003aa98dc2d59320f829b287600cbd6f32b8256d36c7af7d05528c8ddc3ec2fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4359311390085059b8d22cdc3514b5f6b655bddac62b852af3ca2d2a0770784ec3f7fb10dbab390c12851c06b420e812f83e424f13774b4b3d08ca368041f6cd33e3b5d4827544edc92b78900978364813173cece74647652d3c25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a6adfd4a245e8ee7bc14f1b3e47523a3f7c63576c9c80b4f02a759278d1ff8ba69a90516aaa346d31adf14fe874282d7a0e6328033ccb0ae3353a0a34f34d0a253e9a195cc6048adf6685f17bc3464be9b99cb561810ae553ab6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c253af86e156840256e143d6893c560e4eceaaa6f441b683ad2bd3444b5cd4ae9f14d91deda86feee346c162e27dc7a60e96383e2b25370dc515ab68329025f64706c62bb49b60b07b731be4fa1ff137e359bb66b4476264e1b26c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d266da6d77d9d0c0cf09deb9fa6c137be707497a896f8112f29e6e37de22b644cb718eee0e7d3c229581e0fcdc2b22cca4667351309d10755593fb26c351f18d0dcf8ee45cc1f40c66eebb9cf3e14bfdd41d5cd97c6aa51932231;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e73ff7c65ca24ecf3431c3aad636477c8b658da65431657fc61e3e1d5ae347f50acb8136668929abe0787c549d02432fb6c7c44ecbd38163d31c49d4ad8df11aae5874be4fef9d996b5ab4e594c3f29c1a7c24c99c375fbff7915c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c2117c6fd816560fbf801558a488864be6dfb1995cc040c906ee65849373005e96fa143baa9bac0ebcf71ad35054d1da46ee5b648b175ae5806fa77ce43509d3d84ff65b17f972b6c39bb2dc0ec84dc029a0367b51643639ebf250;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136d51015d6d8437cc9bbbc997869a71c054890aa90bc9424547f7e1222561f5ffa0d864e36d6cd521b194846edf54a738bba3978440b7fb6af0f7e82875e8663c2a02ee00c270b89eac1c243130c724b37a20f7cacd25ace545909;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a221887b0b31109b37e37d695e89a8178d28bf04aa5abb0cce839a5f6fd3f0607d5ebd9af1f933f6234d1545e80d989df8adbee7bf909263800303e3f9fbdecb586d869d50453d41a36db0437ba3f4084db3585daab844cb89baec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13246b100194de409f475ed891441941acd06b59768c49bd5974aa333f00bcefe6f152d3311524e5e00e0fdd78a25b0fd6ad21cdc24ad8bb1178116f1bc955b35c8c738979c8219d30c7d4652f49a82deccdb4001d0190848d57855;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d1b709d6bcfdde1ecae77e5f231ff5682b9645a953b8038e4de45627c8b12c85e438e8ae2bc76db95a100484a280a41bb6609c6bc1e424f348b3ef8e1acbea1004f7b0f67a8452555c551404b2ba620394aa7e4d58cd30c1e1b5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cd83de59bdc7173849f2b68fbf6987f416e0dd781382e0b4c8c68b151e6092a43bc6f87b64aeacd5c8c1b12c26910a5aeee824418a550636935a9f082290692475fbc136e78eed0f3917211ef44fdd770f1038dffb204e9f28ba1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1560eb594e6d0849511fffba8d92356d5f9bfcfbac1a4dc32e1159ce6f810a20a6097f52d9f303696595abf7620253e90af5b9d561b0f2cf15f5c846db77a058652e45fb20bcc0dbb98c9781038778d02f3d2ffb011fc63af565b68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c474908454332f103530fc81296075d1d5100201ad12673d41a78de916bc82175cd3e65c09703c3a8298494d325e5a3b39abdc2ff3abdd964d2768abd0cc8977738f7cc08b186c0413e89a19bb4b3ef4057f89cbbec948ccb0882;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h489ca6864072ebad14481128d6c7767d68db5411e3128f04e86cf5c068f5442464b17258f57285c158e718012247dd4dd4c4b7d0d83d3e98b69cc4e2ee869c9f276c0ec0d9cc2f8a01d163a5a919b469d17cb4b86e69f7ee014d67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17121313680d61703deeba910d92e4aed326072dff41c1d682be899f245a60deb041d4b0ed7d8df4649dd77b29f36fcc557093de8edc7d7f9ddf61c521fd26be362ab82f5bf69b49a92f7db553ba10556a128cad5d6c6b53328f75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a567f28716c1fa60a9210af46f592fa4fd183c5cf70904ed302121c767563723eea208ca37a6ff87d83b29ba9a2c1038571be3b7558c8f03cb72f31a85e3b3918e00ae763b9b766073b4412466643038709b25976fb449f9e57ae1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab3b1c1632f34f67560f779c79bd2c9ef6a7809d374e413ea7c7179edf37d74edf4ab968880ec68589c9249d48d5351cd46b697efd478733caf6879695b3d2bb590cb517925c135bfa042e35e9e157fd85ccb36460db2cba4efd56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125ea76114c26318f2800128e7e83ef2051ec97713b7d1a458ec61a9a9f19b1ec2669503368826ec4241afa5efa369fb7c71d0896f23400d134864370a84fe2052621679abb2511ab8d18e5eda7c797e1bb0cdecb3e024e0900c6a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c7a75ede87bb8cf1a6a4c7288f00ada0f792dca4553efa0c9f2074fb9456a3a830fe2545c37a7943e26055f41e2ec926bffcf37fbb7e4304176a72e07d5c5d3f9267d93bd49e837d729339d91874d41866cd2aba997b2f3c7d106;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10efb7824ee5cdd598c229e4ab382a835bf5b1ad7d10db7c29a7db9aa12ea2a1ce67a1c6ff85e39caad9e39d2461008643d5248b832bfd4f30cc398f566ef90e454f92c484dd1db497e7f53c8c5747ffa572adfacd1a613be408eb5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a54a8911cb3c8c530bd16eef8b970472a5686a825e898ff8019896f2eb5a605e1c1cb591a891e74575bdd944b3654f0d55edcb6232d52c55d1a94920304095a5804bd3ed38a6247b5c5b258038e6d0b0def9902d65ca1dcc27e5b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf1fb7f12ce0383c0175edc5f24b219286bfaa8ee1bcca9994b2e99671291f42b53471d62ad1d54c86a2cc60ac35eeef065caefb729869da53c140172774094e82ecfe1ffabe2f07b534b9a2066fd722aae846706a4ce6f0e60f72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153779c9c3abca4e596c87e4d9f85c3b2b610fea9c9ffec3e525109962f48a489f3c2c5d7a93224399cf96c4de55d6fb6391d3e296224a7e611da5f9f4fa7b204f1969170c3c9bdc569ab5ddc9a480d9063d2e8007a853bea29b95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6195b5e8806f09a9b0ba4269a9e6dc255623ee5b326c0becc511e838887c15d0c8cd0b801ba2f3f912f8a38bd9afb970400e9050d8239ef690245e0855cc407217776c2d7fdb931a10a85b78203dced9dd8cddcf608fba74bc4adb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2226eaea3335b70e93c163c7c5ed318821eaec4e6b5c2bfc4e885a19389c08fc82e7d1f995044223e43fefb6eeb1206c47fda4e217635e286f473dd2b2aece5889507ec8fdd983cf642e50c8539ee70f2ae08164d0eef1f87a3a52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h48f80edecfe12e05fcad548d16344818839dbb43337c0702d0b44c894548c300017192a18ba8dd5abe31865de39c379d0e23b88eee1ecf02fdee2b2e20263d6c6b0b2adcf7b8830a4e93ed584324e16ad4d70875ef32a9c56cbe5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he10b4009767d17f3e6ddc37dce8393fdc4c1ecb98fb314590e6695cf75c2441dd64d4261c16b1340c0d98312f16e333e341b8c9282584add2972c1abbe8ae107c6ba2f05577bce193c412980d96bbaa07db3f455534f5ee8bfcee7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d542a0182d79e60dedfb199f357ba64619a2bc9dd4e48b2c71047cf8900e4c3b42a4399b7ffc7e7edce0be6ccca848c663431bd7950fe348fdbd1d1006934eca69187c08e81696b607e355ce33904bf134c8e871785c1d44443aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47ecf5502fc68ae6b8a2c88bfbec5850b82f631fc10f4090fcb14666d607e847e046e6cd697d81aae64784efdbb263f4f09e5b51d2956b6888859f3659c116be06427def49fd6979bea2d174e2f72d662b747a46340a88ca404bd4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3098c2b4d05958b1dfa4d202da823e05a3f5c88a54562c58d1721598d47492a49dbfd56d5294532e5b9785dd95059c4629a2d9e330dbe46990b6b122da3826f9de15376c787febfad0467021f8c7f5709126809dff622fbf3549bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb82716588b2fa5617f3c72cfd368f4f79008725d5ffd13c9c678fd9c7d769eafe7e7f83383c3fdd7f8d5b4a20509ac9523bd3d3338019717a55b45b95950d5416d021cd47085798e537adf2caa3a1ab28abd5529c88de83b0f9800;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e8f7e376918c64e65709d1b67e056fa76676780d38dfd670c0a40ed9d60c8ae8e46152614be92f8b1b6cf4d721296d12b57d8d75f694dc48fca192c3f35f02d4778f22884eef2dc1d0d7a925329c2551f5382a2799abc446afea7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50f53b011e9830d5847e55a4521d2ad09982c318b43c275c8560b645ac1c2352b9976e2dedf2a019f6a88472b3801358f43271885d8312aefdba8ad9f386783a4988413e6ef505bf1db74069d35ddb11d012094e02191f20bb12c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h109d751d3412d9662c83ec5816d51de6bcd90120b724a436d92f849fc06155e6cca498be33a2220dac8a560cb3de63927430bae60cb0418a093941a618ce8e61f0a08bb1e4e64494fce0500d561c6ef0638ee5721f7047ef3bede7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7edb3c8c701e60ba84c5833ddd1a7d9d3660b2d1fb25481ff50ac08527cd2dce9f393df80441539f8237b1f140ab2c4f484e49dd5c46c568ced2311866723e728988ad0d66c8dd21ed535fa86f27974ddb7f4e476723dccef0ae5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c96e5df5e04f663607bd9a14e0bc69e766ce806cc5493925f3515f9d217f7560dbcb15e654d823caf2ae59e196ae0f13ad5dbefa49f8bca361b03d75201478f1f10513c3f797664715d530e050a134ae00b83b44a5657c8cceaf11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e40be11fe858df301f605bb07788aa52da3e811cf927c799beee6023b937731eb1c8d6e80eb10521d24e0a2736c3dec45e8d4064c2ec78794e228211a9929b34e32dd6f622c2954c92c41d3b365c8b0b69f5c5331b80331703f4ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179061e3217520c8310e1f20fc13bc7076affd131d703c172a9219493915f9e23ec9c6cb4103bbd15cf16862141c82a4a0bec5a4956327f2a9dc74969c7412b8b0043b3fae7fffd5d868cfb9ed79746d03c3d9b399a502dc9e0536d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7567a5126b334d036ac0bdbae9f58245b5fc56369625252aee479a1f0c64f7c4e57874252a9e3db18cf4eff69964b280d8c60f114863cec760cf4c95c79d344d67f43305a59b4706e1b19ef40712906b77c8a98d45921653297160;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1abc252f6270fc4cd06310d579aeed9d607327da1ea9de9355fed52bf66d0d2e03c69d2b54d75111a824648329986e68d6274a83c9f6d2de57bc98786fbfb70252b25f9bca91efcbc40bfb5616d531e9f55d32d9db04eabb306862e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aabecd663495189176f6c552f141b2153023409456f1459f1d30f392b61332bb152d241da1088897502a7dd23986d74e5ddda36de9f89d102cf000b086bcf9a0d3959db481daa3fd4c3e720910b279cd6ef2453e66c7dac0fa00bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1228103ea0c554c0489e1e6c0c75858bd5862febca1836757eb0152611b1417ecb7faebc45261272c98033745bde47ae7f157fbf4eb20396813f368c15c1a2378f00a7e66bed989660a4c2abcc056ebf31624b5101205edf0fa9186;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e04ab33de1bcb3f4c2f627e3afe8844212bf35f86077ecf15321a5fed9b064b9d888030592495f06a47aa223c200632fd0c1847ff0631bec7d95bcf1e00e39e18cc01e4893112450c6256976939897336eef010dc3e38b4111d0cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbef24fba321307b2345935388e98e88b6a6404263f73ff44cb495b802d5f59638c280196543013c3e38b18f4bb76327697b7b4422e0c184f7a4b99e31b4fe35e3ec54e75dc29a744e470d9b3cdd18075026b8fca6ebab342edb33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b2bf85fee3587cfa69a74d53c20b719300a34bd3bbd1c168fab68a81dc252b83267251d3dd0bc5d10cfbf89ef3c75db9d213a8ef4b4020e3504813a4ea7a3887f77107d9f350e4d4163635fbfb98c232198b28b2f2f306bbf0f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41438ecb3082a05ea06966abbe5e3d78a2bd20c92a51203ffb48a0a8485cbf1ce334c144e9019aaa6e53ba3f816b9303fc69924bfa2071551041f89fb0a0361dfea4b8eca04035722048df7032749892a3234485696058f458913f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h77eca232fbb44442c5f8d0834129dd81e48e04eecc8e9b8cded2c3d522dc893d8e2e4899223ace04a8881df6322c76dcd36948660350154dd5051aa31bb94599bac7c99041ac370a34ea2ccf0630db20c71663e084edb788341b24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8984414cb23480e8f0c3f4165b64c0d9aeaa4d76e90c46b9c7c8fcdac2c0529c8e15277ccf170b32ee8417ce26f25c9c870c78933905ee58e19f073bfffc9c51bfbe1cfc1ffe52e377ac7afbd155dcc9dde800f6054b77b8b7e932;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2bc0812ecf303e3444b9a30d1bc403e1c18b5e781a5359161bc2b21203d09a1716658bc780f8636fb634ab8505a2a8f8211265060209b612e51df7879867b418d08e65ba4e9716f208d6a69aa23ac8ee99e70229250c8ea56f5baf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbcb161814ac148c01bc348eb6f39af9ba1e56cb68cffdd9e1f86108bc644efe18568be1d46738c8be70cc593dd955b8f8ecaaab0e2b7387f55b9318d10f2a1ba7c5d6d14073f2a83220640fb9ffe404cd0a1509e282e99f3c96376;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff2c8640b0ac8f6747ba1472d19914c373bfa00d336cc2b81fc6ab5de6c85980701bb6cfb9f1834e19b20f6b8c8e3ff8f4c70f0ca64e4d612e3c38517b8e265409949b7fa4018401669929fd88ff24a7f388507d1eff0e0e6586ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f21b38fedfcbf8011f4bfa39f9609d40cc0a84bc463f82607132790d15676ee89b33e7e861936a60fe18cf7a5f1fd3ee815323ebea1b66601d404004273b3a480c93ad35a58c9716905cfa56384ece45f06145c4d26663d088e10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b6aef4d020a0c1ae872892d75c06cdafc19bcdb0547c9d913b4ca8ba54aa1b8ae7af81bdb48a3edcdc480100224f7da624933987c344bd76ad73f7804ca748c2b7fdb9878b90f207071f3b76a886435c4f83f5c35bbea1f1b25cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b5b6d10e9ab12cd8b2aeba111a59d236517ba200f1f763726c58a7cfee21295789bee860ab2246bd0f56d48faadefdb4dab5d4346a88a13b2405f33740909d076d6b576dfffa5e45f8f90006866d052a9fb136775754fbc8292a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5ff8cc42158ee8ccf7208ac7a5fcf12be0e3be9be9a73a9918df7086c52d578378f2c0a0adb9f4f8be323e3d2f733cbc39c29908b968e4dfd57bdd36702b98a58413ba42340f0a363a46044f2fd09296dbddbbba14aa7bc49a5f25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5ec3bdcc24dc3cc9b8693f0213bae852c932a5b94f1c916b2625d999fc752a688cd25163e3ce4b9390937e63cb6a3f59ed35e596cb6ceb5a90d49486e86ce773e906a99f86a1a1bfbe5f787e6f41d583776fe4287be189c107ad67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd65dbde022a8d73e38c3916af868e4138ab86c6fe0f4b8e2cae2ba68ac075142d4d749fd64f2650de55325358de7c022a4dd2f08727db80f0caf7892998eafea01107fbf392a7e4ca6e3be8a921c5552702b49faa5c7c1279db527;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ac4976fe4efd8565085865c78ab9a6dfe0ce79fe593463080e8f165e855b58bbae4e1e759ed70877ae413539802eae7e4e9c6f3e6dba93b0d46acde49a79e0f499dddf1385d5254f365453f53ffb6efda470671a965e043f0240d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33a95d77add033fdb8f1e9e75f9874df9c268692da6755c28665026ef51668ee92a86863047a66d57b0889c5ae39f2e6d65313f64b8b049e37f2cf59c0b96d64e366758fd1ff77049497f3b273d74c1592fd7af2a01623dda8bafa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121f9aa3d0302c47c1520b8eb6e2d32b626b8f4d4695b35c2761cb92f3aae03b619f06d74664ccc1d7ea565f54f1c5227bb1941b635a7333be58c071a6386a57f43342b107d12374b828ef607d3b8808b234efa265ca6792826cf21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8af2d43ba5f348fb4e386215dc2cc75737f440f3d2cc0be56a16e46f6767fb9acfc7cb6ddfcbe0915fe7e190ee10124ad715a1f356b73f18068e290fa9497dd2985dd2abf390f175fa3bbe11777ac2299f22dd5362597e3369485f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he88be420b00857dabffd7a3c7192a0caf0e2b9ee5b46595619d0ba114e4e72da4ba49e7fea4749b883f5635e41bfd58b4a79bed94e0eee9ae1d654212c3277ce46cc59202ccb0b17dd406533f7bb831be74332f61cbcb6b9136cf1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160bca597ba9ae0d0ae0b8e8de9b8f2a2bf8fa47631b2000d1d5350b74c51376b1bc7cae349a4fb6ea5fff633ea6b65467b1609cbe448ecdc9b043d6c8de6a617854017ff6b16e1e6468e7d4faee44dea95a25cf0d200b0615f9804;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd6374dc30d9446005b588ce96cf0068fde4ca3765aa08ad80b2eca0f46b4728cab03b644e49be1f88fa4e5901310fd05a26e446388da7f9d6d0e213464132172fdf576e344aca706574e9545e2cc82ece0953bd98ba64df74f9c92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1159c80077b0b9da4164fb84b7b49ee3e7256f9575ee8f59653946cfd655f3edb9f6b44c58516ed1d58d89578d37e7bf94b411eebf9ef2e03fc78aaebbf0a80f344b9a5acb1aa37a3bec607e800567b34a625c5d0983cd8f14e0dc8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116c61909886418453dc0921dc3f1ba8ec3a7961572bdee5bd59e42f4487d63c872d2a7f12e69619eb8f4b01811e2685cedf89682c2692c27e976cbef45dabaf436b176b2f844ff99eca093aaefbb2bb39d52f703db87c4e529d841;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143a68d80e19d8e05d7aa589f545c4eb1001afaf62bb6160035a18b515762ad619daac4370822ec42d947b21721c4a6e6389d9ef6945fa22ef21b57cb2c0c173f5ebb56f86a8c3ee69079a8755f4ba2827bc21e7b631a33e48bd817;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e963cd6df04c57c6b58c14ec112220f2405b7360ae0f6e9f8b5511d6f8118dd494f71a35f9207fe6b6304b5719ce5334de147bf83d0d7c9b77f00ae243e584520856784b81d30fdeb96c5f3f504c3bf03b2d636fb590d7cf98cdb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd3c293e4e0cd285b261f9edddfafeaabd6114ce557b4ee109c39c8b9813ebb1ec9bb31a35185973ea698afef9e9817c1fcc2015cc08a8a1eefd5f58cf442c080c18b9a12eb8fe312ca757fadfad7cddbeef12f52525904f96fd5fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h401ad2fd30f22f34706b08ba304cfa8b421464a5cf9710c608f893ea0e069474cc72d90bb62e9c1a11f4edc38da8db14a9ae64d76c7002d9796b7be10e572c6f6c95d8347aa6c3716435c207bb0fd96e2babf3c9d2457ee803b2e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174969122615b8dd0a0ba8477358d04fe68422c3629af776e209a3957b9020ea50dc8574346785a063de5ceed05e842ae364283468b599414350861717392b1d55da3dcbabe857580b3aa0f21600b23393222a16bbf648d66460c99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb511fdbd846e8765b0ce5e86bda72505f7456132040f5ab7e74127d013c36e341de27ae54920010ef7acd0f169501fa47f83b16e20ed80e2d978a1b6ccf10d347b6c9fd792947b473f932763cfde5a9e447b15836cdb1f0d2b77e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd017567026a1eda8eb73ad57661773608ddbdefe434ad8e61344a79bbd6c66cb2512f7d05085c23601c66725850500a49bfe7b6418a350736332dbdccb40653489f4c2060189505788011659914b07ee8024d70c96df4da1acc9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d5134e1496d335bc65248740219815c4df298200c01b7dc2ac1aa0fe2dc50d34e560f2b6c657e318bf195dda07ad2b46a2d6fd66f721e197d9d2b8e3459a02eb5465a694e3f80ae7fcad9eb18213c13bbdd62508d155d1e29f2269;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1021b7f3305d5fe45fb74f2731b0b3fe000b0850bc72cc2f3556df279848836058fa24109aa441eda4e66019d3b3fb7489e88a78be096c3489e24c1403959e0c46a731a03e39aa2e85cbc53e18cd0fe6bb76aa3170ac92b6f6f1b7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b2208ba1d48f417bc7da3bc43cb740c5e284bad9c78c52ad72450ab01c9e2f44c20e150fea0abc4f4ead7bfd8a8f646032e99c7a24f9d6e605d6cb5b5bd0ca1fbad2df1bfc995ed1fa5475e0d7616cd33d728c84b5ab0d53527dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdae8638c3e62adc6b1e13ca197a7632952de77f4a12c308535d81ca36accaa1b2e9f81d0526b94d466c4e300198902b2d14835b4277b60c4ea5962349d80ee0a7cf79aefff4e81473e9a48b29c0dbe9f4ccccb1ea1edca166f1064;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1446bdf7855492fc677559f43d50dde228a54c150846a6dbd44e72022e4fd47e79a6375485192f9aa6d5a6a84f38963be59ca6463a3d1d644995ce095a284e216c055f33c8454d97de0cf1dfbe6dc1d45eb44a11eba77ed944cd451;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116e148b02056e63f4d3a1630ccd963da35004d2ee154a3068f8edb6b7c321c918d1a8a1e97f077d91e7b2e778ce49f8ec66e6db6d28e05a2bbed0a052630a3fd92f6d86d192e92c0b487f655876cf92037f9862df1aa9ac8c645e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160223177c13e9c2c2a4f6901ad0ce53baffae61218e067ba6d147ed21b6cf295267ce8d413e350f1156e9182edca5d69ef8301cc2c50166f75f4c1cd5f68ebc5e1f3e225433d3de1c7befac1eb22a8f5db749f9be673e4fcea8854;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13295bd546faf9b254487a9b82cb02626b315f688ac3eb3e2a532d8d902dce1c048d9033fe26a0a732cbc36a74cd3bbf5c5a22bab6d8055016fbda0d4025a42ca5b5055f384c311b12d9421f4722d9e9eab9014e5c8184896cec143;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95b5a2ac17089b8db5b311d1348b3e5dfcb559d34dfcfcf3de85184cf3e7b1feb7674ea8792f2da5187c852313414601f93d7d804cefd4c58a9b06550a0f7a0b5db85fd5682e3a09deb1253573e775fba9e8f7503fd5b3979a6e86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h864f895b4b304be1dfbf8ee8b2f0f805e720816b438c9e245dcadefe8f7c11778e799a1f1842297c4f4a65347a7ef3ea5421e52503cd37119551f371074f512a3cac7f88e34fcc92aeeba6c290ea9cce664d81530ee6eb3fb4f7a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f022da6a9562384a71507a8c4532c89f64a25ec31ac9579757f5447a3513cafc2c47cf5e5f5a4565f0470cde3b46bcf22b3f61c150988ec0e83c40e748a8414b178013a9001c8f933d461e71971cbae43da09e9a29e1f9bc654708;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha616716c87a2645e07cca1087f52f8bccf923b374ba7197fb94571dd9b212c8c144ce50fbd334029c96f166a8026a8f6f473e9209fd2410eef6e3e6d9aedecc242b9e4d34c8253e7936ccf9fd5f731de46c128c8dfb262ff94d5ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8510db1e8e135194de442f83aa4aa77e514ae162fc95c90a1c5c08774b604379fde67e34e586f8730e17861d72b3b47e8ef551305d4d7cbbd20e57c04f77dee3fb04f720908b0b0c521d69334ce0f0c3029e55e059c1dea151d8c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h607961377b7b144025a848776d4940f0f136fc721b9954f1548d0593be786455eac0e1d7ee5b5218cde4e6150fe23df5aa98ac76a8b2fd69287ce10aad717648b375772e9bb2bd583fc2c46e59dacba49b31081ade7752f012bbad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1717ef19ff4e33f6646d03b48979d7451687b06fc472b94f8a16d998b7ef97b729bdc87c47b0d9a2c7d690eb83df314acab676b45d02581fc4cf7fe9143b69638b687d0726760bdf8556c449777f328ffffbc82e98034f32a79660f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5a5145e00074fe3f1c0a60639853a43a8f7202ef727e6079d52229fa7382b55808fe708f184804a523c66290a18e65631a7d9f438b50f6e409c34f74bff0fb49b6e3a52d3e5659605df3617b40860feecfa1fade191c8e055f69a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he85001aad89498883488edb739104f3955f8fae581c297e08a8ecb3c86f5ec66bd2002040c075bf1aacae1cc7a49a0b1427ff8c8854968b632ead714a755f64de2a1ebc2dbc94657686f7b4847c95f683154c2a67eaca91b7a875e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12db11b6331e2c61c7273669f1dff6125a89ca456d41694cbb06e6dc01b8b96645108e0131a2227358ad17cd6e2737b5ec9479c705cf3b9159d30c7e48a58ff8e13c5184736556a4f93e1956ddf5ea6a94e9962fb015c96f796d944;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64513787fa4ffd31211f26797f9ca78d0be6f506b3bb72b397ae7d897284311fc89970dd1f82efedb1d3db7add9cea9f32776b86cc38ff666329a6254d22031c7a7a2af05096df3c346d3fe3924a4b9ad3f281844051e36692a3f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8050a74f5f250491f820b79515b26b039e1a619398784e2d8dc95782958a52a06a09689fcfa2a913394c9813145353d84acba89a4c8bda5fb4fd807eda5b0bcdceac04d6bbc3d31e93bd0ffbe961a05a71c45ea708c635681b9d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h154241282ba000545fcdf10e388dc22d2cba2766fcfa52e7f79cf162ecdda1547f98ad845fdade1bfeff5a1b079e93c9a9a68e3daea57b9cd15d60726923c936f1cd086d6aff44ae9170983ab3a09d3523f5beb80dfd497bec0e267;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hebd3049aef732deee27656d93e7ae6b91dd17a5f054df4162bbcd4c7c04a67a8205308bfd3b7348322b0501e24205e8ae39d22251e010ca4c147fe0b7f07413dc038be7b112379b4ec57e13a16b08e8ffecfa18105a8da75ed70a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1546f5771c0d257c6ea370a276b2d8e29076268a36bc784bed5dd8071626add0760d775c93d3b1285807405c7a4d682815d75cd56f4fd5b1988de21cdeb4df3fe4ba85651747ffaa8d0171cccd53e8a9374fbdf31d1ca5155e01af9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h903d34e1731cc0212a686e30d41510ed38f669a23275baf440196fee13970b0b2db61b4d570f92d41f9a3e10a1174dc52d8a7e05fcec3ee9297da95cb21334fa021a85fa191e9991fe3a33a9ad3f01f2227dfbd5e2d0f08799f097;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffd6ec61190c4f0557258cdcc15c5d2c7026c2db05e9c03a6fe11699b66c9989dde008572efd27d8919cf8449832ba9e8d2e03d6f7212ffa56da45750bc3fe5a52445ea991f094bb9582bc73a623df8024b60608a9dc9f3280bd6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68707f8944d0ed613d0777b1abb7f162353cbb399e5ed7bd44b971a6e1ddcf56d24f353d0670335bda64cfe629df646cdada3d8b737a2f690be33a34b46fcec79c265ee9601ddf566a5a681f410b5b2a6919aa2bdbaedef76ae297;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h772eee7d26add0c3a44b60355a6d23396b95b850f26acfbd4342bf83b58f515525af38acaec507f6687ce6dadf5c16a2be4a24959e687815c9d655d52f7c837a1c1aac1695314ef2e34b25b8801a08d4d6924c211f370f2f51f491;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd07eb853829b843515a0bb154f2e45c7ec07773bad656b9ee7998f427ce2237ad5ae1c1aaa4cb60eb2b329b02da4777418fec6b65871bd2c3b7c5340370b9bed6b2b2bfbf2cdb4adf4dfe8bc955e2946eab549e8291a3597926fa1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fbb2c1e78485bc1cbd5169ee1540154316ed51c04cac8d5846612912e980a401f723773624f13ba554b791911b5effc8feb6da4a65b88f9707b12364a53635ad8bc198e5f90551da783797985e7acf6d8a27c8b1227d24177087b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb2a0fe7ce0047b9219b96f29ace95f37214873cbe523207fb5816c629d6ffd2b2ea4067e06b1a4d066923a46bc7c580c358cdd2f4349a87429f8263f25f4ed3ef67b5de65df5479c64bc5932a599740590215bdebcd6320ffbd7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b5f745e0ee7be21d206af4aa6e764678654a4bf850df1114c15e5ace84387076b869a2cdf705dd666a2a52b7cdba45a0ac842fc672354703d73053735b724c78b077380b47d3b1ecdebbd9c104efb4bad456878e0808afca9568b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1291111528cf65bdc89bee795ee4129e78383207bc8e8da7ed44632451b98b15b0628b84f49284271d597e58143921c21f92d24deba24ff03a98b8df71fdd2bbae407c7f5325ee1915a21393ef2e21ab3720125b143f74792677c2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18cfdee31635b9c413fc225480e54894a35bf4aa92a7d7e8a0198de45fbdf7d3afaaf8c39ec114a51789c4fcb0fd2489b605bc434ea2f526fb851bcc6aadb9136653f119efe0d8b4221dc07841179c493ff98dedc8441f2b48a3aed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba2df3a6685223bea69af20a9a1294b7c31e8fd6e5d3c6109b1c58a420183867b2f13e30a6003efbb32d79b408e4d052f2acec3633f077ec8f77d13b229520570fdfa8d8d66053b7aad00efa278a52d8b80088e1333609acec7fae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8397634ab1b43e3994adb3902265390bb4ed73ec9a560d9f082a69f1b76d7532d3d9b7412c59bbe70a9e2683466c99541552fdc270be9299e4e70e24666f339e696e01104c376129fbe15f47f52d39ea18186456d1078b12134e14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148865656cd0fdb0a18dde3e45c5c54dfa1c402abeed64b765a7eb825965e4594d7878f8eadfe92ecd235fb8abe0e321491af041eb1b8d189384d1752efa3183fbe67dfbfb2691a457b8900eb1035ce932841b526f3568aea2565e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f01e1f986babf53bad13d6955136d1d98248c46fef287f8b96bfb766d5e94b55e89c520a8358f1466dcb49a1b0d791abe296ba87a6aea903d945a121e8c646316448d79b8aea7d14ff5dc327d17c577d3c6448501ce7e231f6b784;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bef69d7689e8bac945f41a5eb2f4b1220603231fa8ad8b9d9bc825a4d1adda43b0fedd367ef1ea56c3b5b7a3a7bd3e85706dc3703a7350b696a749a258535dc365ce15f9490bc584a2a8bc9f3e0083efb9067f76101e89310f5683;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf65f5fc049d11e2cc558c45fc1c2aaf62f9268a631739c66a4bec43e42cd0156b37568bbb6e8af16eafac7e414496d650049b6c5fc9deea3bc5bdf8433e54fde519cfbef82bc0d14e2b1d109c60248170c14259d8ef98ac0bd4bbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142019624250289dccbcb84cf13ef3fc6ecc0620b1978999c31f8510f2e0da13daeaed3ab936069b7974d7d8856899a4c3120228b702674fadd1209d2e9d3406767cd16ba9b6a715ed237c4b3f9edfd23519f3082acaee33320ae9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b02d8fb9fa4eb39046b2236620119b975f935ac504e227dadfc954934b5e588d114a40c6511c540f623d427eb5c604cda96365c1e2ac2a7d7f9f335e804b5e1671b1572901024a0a4ce7e8b74d05a1c2be1161bb9c3b2aab3c2ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d139f449d2f8326d0ed5fc1a97162d7a951936c2caf37405448de5c367a97357588358f924596fafdc2ab567bae5ba6a2398f73ad43a8832f9fd030f27d1954af9f4672d40f7efb68c161b70cef985700aead5f60edff14ea2f815;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b71dd1975ddbeb740c5a76723243f9dd98424e81688871e121664d9ed0807ab4ab4cbde8534442066f7ed29c5bf837d9086c59d050a72b8280e9e0a78fcc1d7d4db60593d0d6f74ff1821be42980cdc939824a75c9cc5f8daf3f6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e19a059840adfff8081dfd37ec7dd9853eae45c6011c8ea032d9687f462f6c3dadce6105913376a82db89d65f4c338fa327535c22b650a9aaba811e0cfb9ca2ee13c0dfba04172e684a63b159b0610853808095b002110f9c148eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h77b0aa66c10b187d7e124d0d7d343bce26d9173e027c9be133b2dbf1147d872e8318fa7f1697a176382729f2917f97a2ef601fe598ade01f1dd8503f9a8dc91a13b56a3aecb2059ec28392c046ad03f0e49d83fdff5118e18efeb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4e842f38fda08a29e2765f9d7522c0182de9a011031bf06754df523f1fc5f2524a0f50eeff02c75ebf2facf89720634c4851465fd1f62518e9c0c13f76607244833250a081c29fd52d101186d9335cd4cc590dc65c4646d6c333e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc1a1a51829f701a1bbd774b45d27dc9001d1035c9c6d2049684b7aaa9a8bdf4769de170452e247122653ee5c6c0b9bf8c26601393ce47c80ea4808344a32a4826d12fa99336f507accf390209af57907e46f7264568528d5a3edd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2d8e24c664b3d2098a2816b30329ad109c9f9fabcc6fe50659cd62c981575908a660bfeba8ea987375cf4624f0afebb0a4d6f5194eb128fde5bec0ea6bb9d6d02323ea4fab6caa227a7d266f3978eafd89e43c4eb61b71985443a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ab191c9e052a2003580edd90f9a801ff13db82bc5ffdfacf34ff6f83ad7d2f3d603874ec3b8f3f8ffc020336d408810dbab60dcf4b42f5fed243ec2ea91c2d5777d885667bfbcf67c9e1aaf1a9ad0843710efa5ff944c04a4298e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8fdb160c1ea2be8892a361679eda0dd6d301e81291e8ca6a687e53014d7b05e5d01c8b0766e306ef4cb2c15355fc26d84756ce0db325bd36ea5b9263de9b3359855ba6f35e7a3e96b510dcaee9f5a44ac7aa45cdc300d7f664e5de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19618f1b20e1e794a9d57932ca271f1feeeab0a9c4c66ce518d8548c3746b6beeb5475af33ecc12989281fecc6e81bebf8a16d88ef8bfb47355a01db94b7234ab870d0288a8e66eff9571e4b1feac9affaa81cbfd70259ce8932163;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5c3f693d0679baa86e4f34dab62d898733f4815b4baeee8b8025cc1a19d33905dc25b246f654761832c71cbdcc943e22dbe84d58ddd4b2c4533cb7c848db2909bb546c1f9944dd997f0a59f82bfaa4470d67fd59a217f5c1d3ca5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d39fd9524f42e638bb5af72c04c1800c50c8270599f8dcf1857981ba926149036d1465e1bc6aae02c1e2ffabce07caf17e760e7dfd337f16a7ceb61a138971d6d995211929ac441e05b3aa49764f16dac4ed38deaa11be911f8af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9fa7a41aa02c3459bc4ea9ec5b643ec58bde301dd0b92816853d740a812f7aaecc38aa9e39692be3c1fa0a874f03a1c3cfc0ff68f4060d0cb043a45fa91f7cc02147d6d88af581fa13c96f404140f7a3d7825a398d7ffa243d3bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e68c053582171f87980a4e64eff29efec021720286677555b06ddd5feb355158964b10ce2a9bf16683b8fd7ed906264468e984868b9228dc07acc7ca9963c255419e5bf99b1e9514a4324619ee71ce81ba14a944f48a2a3ac9c45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h319719acbb3c58fc012819ecb0bb7b1066d3464f4d87c634fbbe5d7691a887f912cd43674d2b2d58251a5d722981c00a4b360c15732df2e87acf9ee7b163feb53f303d0d00b951bdc5a4e668c040a5f3cb7fa5256aadd54d5ade14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f543d02ca952845cd83577b5df4990328a877cb95a2e3221533506aec295ffe25e0729c5baaa39d0243a21f4efe8ddf9239d17ff64ad3e9e6ef98b4d83c0a2508704b4c6c93008848bb169afd73bbe3ce3239c6652ac6f16e8858;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5e09135fecea03c8053c4a1bc5382db2d6b9efe3c6434cad91b88d7594ebc453e25b1e46208a851a7405f98ae41f6b4d5a22e71c7b15237cab1423b89466fa7689c8b204452a90780144bd07a544618995b46eb30332652c7f831;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6eb5c7476079aa61dbd2b287e69ee1b788d4d4b4e8bb149c3ed14edd16bda9fc00b04a4213638a33016fd336acb472ddedc074b7fa137e2097889c9b777380ff13fe74d081ca031c83b8ced4baf1ce3a35edcbadfef1caa4e2800;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a8a10fc7e9457924ebc7cdd14aa9f67bbfd9813bf22749216c9acb7594ed3fe941fc24f0d790d25a22d030d96c8ba128a7ddd4b54d6f565c3ac29b1b347b35aeb6dfda6e68bda3b265dafe9f212662f47ffc5bdade94f49cbc669;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h722d194bdc75e195b36a716e7453f2326f4da1241a540c6a912270332121b5f33368f165be77f12edbf2f7a6b7cd13542a3951fde1b2bbecaaedddfbc298f09b6f4e33cea2921336f5700873f6cebc02ea92d87fd15dbbde52b0ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7e217d2a70967ee2aaa48dd4bd96c67aa0df70e4085ae8fea98e7705329e8bd8affa0aa1dec0feb6b9f9425668827e0a82ff0ea492dee32f785e9221669f58f28c44526f2c89c6293a05d2e89dfdc88d4e52feedf3f51a470850d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5fde01644669efddf2d1627b51ffafbf3f18b60bb2eefd8f662a388d00a89c98cc000aeb5115aa4294e2a56ab10034dea71eecc3640b59587724c935e0d7e90a391e959bddf8805ef5f5fdc37f0135b74e46eecc257dd1a2f6271;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13691483c69255df370e3ea068f4263ed1dcb8a68a4b91ac81d3f15f3a951caa800befd59074f983939a03d258354cd2c1cff6bba8003afd3eeaa3acaf054276da979a17024bcd7c85d89b6fae61ffa18a8f19e3333485c9f226152;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ed8f6f0ea67f7ad3a85dfb955ecb60aaf8e4c3278ecc75d7855a8ff077a212aa836231f81442958d64f6b216638175f9b8479801f89d36c85eaf30bd91cd942f6a1bcd92750fad9dece3dc0ae321c99367d9b3a7dfc5cae6a75b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfcc70cdbefc0cd1ce40b3353c9f1feecb9fa6bbb38f41b476e5c3a9f05e8fb70e44e22e061c95b2e848cf419bd4d0c478c56a9d1c6971c9ccab58817be1176a05e88c1c460d395f42d0f8f047bb2f910d56472c794adfb46f3f269;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f2ed3102a07baa8d4b5a4b56ff356c79bf7f224ba192885b95439fc34dc9698192cc93bdef7cb71c9ad8b8743c108b85d5113de893bea9fd56fe72243557d9017d045e3e2ff3c83f473efe2fc9c1ddc308b889aa0bfadfec9c31d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf48f093581e9527ff447080ecb1f889f98fb888c693adaadbdd614f52cd594b888e93b4c0056bc7a88dd6d2de7e17c9628bf5408e2498224704ed75cc99e884e49d4aa673f933bfc4e5b25ec62facb5ac091895633eed19b3fd6c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hebdf00db6c9efca206f5b6b30800b22808fea8b11473be8bc7a6bbfb7a6538659e9d94eae3cfa9bbf94c34984785fa96b57a2229a7676f2f5f889f40098eecc5b31c46df5d1d9572af6f3bc15f4338f2ef95afca512fc04da0a46c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ec9515f8b84b7e6dea7426b9f2bb0ee05b89ecfcc7e3d34a7d318d28aab1591663f2ba2057d12a367af032f7aad2bbe2a0ca456e4bd780f206340e32ecb34dcac072b47ad8f1ec900d7a1a782d38afebf75ea4328ab3befaf1fbe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aac1c70711a6250ba28be198b13138f4da76586de1ec6b7df82dc286c5c78bb53348a8654a57e0ba7e9c3370971ea60aed78ba04c65ae95d5827502c4b1c980997f2df799367d6d863dfa43c023b188886361610fdbd6bbdc6598a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h175e33d8a8e4fba3d361d34e17f0c4e0af38b012aea826168252e5b401bc4003536c697e114889b8dc2af0627860db1ecb71fab974f30dc23dfa9208b5595ad4df2a9ef923e25acc03187412684119520c5e4a881e200ffcbe64df9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5f8f8647847b550bfe7248ae8b69309c06b84cb1738aa9b6cd11688b82e4fa13ef0d47f8f57e625ea46328587753b50a91e36af9d7c7ea76ec4c8f144f998541dcf93986dd4189e2806312331cff51668640cdd8ad86ecd227f5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ae5e108b7d7c788dcac677e6d3e021e9802f40bf85619bfc2f6f614f19521ac94392810a13eebfce9e5e81ec4d6520f1a5125f352897930a4028529f8f2bb5cf3cdb772b55b6b070ac2b080165b23ad26140226ed453214275eb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd436b933801e9b2500ed187758740d42690976135e467148ba9ff49a11465396850d89668adb7f74bba3053e5421ffc8c002d35335adf875915992c4624014003f9cb81aa105f77ee6dffde6e4eeb6e66ec98abaf85d8db773fdf1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7c6f83ce5cdef57472c18ecac7921c64780f07167722955bac7b5eeb3b1688b228f17f02d43874fd76a343d9d6d6b96a66db79c1c8cdb77508489f5357baa38b8592fd0feb015f8611bb0923cc0c5d39ea15be4e1bda04e8eaf29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c998bb59b7ef172994615267e0d2df6805a7e0ddf5cc4357ce4a157733b56bdbba45956221ec58ffe496c455d97a4f3ece35e63a15672f109dd738fafef460e0a5840b64b56dac56ff3611472339745e04f68d3d29afd114c1b3a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7056c31ba37ab3961b29d52eb03c2e44021e560bea15805bf1870d25d002364bede3e374a221462375dc5b536f534dd3a775d4658ec35d7e465f112a3a5e4757248fc5c6db3b0bb6df86f3de5930f7dbe147a809ffd56af988cc49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d878915aa73cef22c517ab4133232823f240eff3e3b1155ec70ef3311b366f3532ee5a9cca1c068069e34737a21ae88e565b32404a4299559b5602e25419419b06fa773150aca99fb9617765eca4a34467de44c20723176f425e32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1805b00d3853b7f062a9f26b3a221574786eab58d3630b2df1a624e4524e8af2c7a62e26254f04e49e2073e798fd0019329212abeeefec55de63cb81341f5735f1d8626781fae84ea3e0c10cb8818ba9681240ca84602b549fdcdfb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h73b2aa4203ba9d281988537f6db31fb2e3f44c43011c04805c23f3721f9c78d2180b03059717d29a8652e754fbfb8c7d91c061624596e6262e81a7dfd66d09822533154f7ef053c03609a852d36e7735c97ecf10b2c0502408b8b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e2f57221ac4614e91d1da8b0c05a12fa08865859e421e50438e9aae7379f51dc4580ea1b1c0f04def545805c9a1dcfa4d043348991688d653a6a61857349319ef318b15509455133abcc17660c9a03e6492a1dcaf1847c72eef2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17d66113f9975d285f61955aa0f0d416f6b28e58f217a5258b001207609f8723fe9bef97027d581b3b354fdb0a0107a47e69bfe8452f2b0362482d0a9d62809b2482f46e50c0ddff67c64e4ee2011d63bc2553b4e32c6753bc43539;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5bf42bbe8dceb5c1bdfcff6b42cd2453344bee157847016bb14ae1baf5b5d7f6e64bb9e439ad960d3cd8ce3eae8f34451c0a3a0abbb81fcf219c478cf18f7923df6e5fc05edb8ac8f2494ecc4cb62be60cf5e1437a5a5aa12028b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13cb4f0ca8bcccf8e33707429d5d47aebba2f8f41edddfaa35308b622e3a774f79464c3186dda9dfd6ec5a4bc855b1be1297b8fe2998bb65626e43728ed9d1cabacadc98000fb34062300aa89cf34d709d5ce497bf8f3c1f836e9fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e945f9a0d5fbb96e92129ad761c926c5d2a1a74fc6acd691e55b8ba3751569219373d2d2d287b23c3a6a7fcf84d4d9e113d9c10c08af3eae0b2849085598657a8efa65755ceba7a4c1c2cdf08b2da810ba6853b8d108fa7a7c4d36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f0e6af1a87c21b5b262334bfcdeb267e91e12e05ec66aef5db5349d570c2ffb139b8e21823933730ec8baa1a61e83d698bb84cfad0d5586f86ad9d66d7023344c4b1f4434889a720cc66fdecd7599ccf406387d4084c60e06cab1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41563f944739f528af7e01ccc78120876903b9d4ed1e76aadf7464c4b1d55c421f5e85bd3e36049ce19dfe1eb4f83e0bb7c4df66b376e4254b25c621118f18cd6b424b81dd6a2e907ed3390ba59aaa8f428a31eadf02db61b978c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe7499214c80290c50f5d60d83aef6f7e08264a5992fbf1888b1e8efbffc70c3163687bb01c8e9052ab6116a3bf67e76eec17d21c3c8ab2aa3e7dd44e3dae34b5d2565451a1b085b96b8230cf60ad5593349e49343f506ec7d58cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h267d37db4d7421b0eb392a0447e1dc6e3540baddff07f161c8401098edb81c6143f1ef2f714f1b1e43df8abc2c5bd19272f4033b83ec29caef4cae8c4c59bc912ad12974db7f2fa4310e15a4c361eead2ae9b4b1c832f679e17a62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a5ff01b7d8ed43ef59783e219b3c436a3754dfbeec306c390eb7d9958e0b44bd081e785ab757b1a4f0695b480ecd5cca8e89b2bbf4ad22cd2cecf12eed296e8f351b94c1a169f81e57f5b0573d0ee779e17d206d15655ae00085f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed5a4f5a0546274852917ddeb00f942acbe200ee419d9a25e264344366e11e2c2d8180c63ee89a4095349aaa7db024f462537f203f983f13f373f5f7a31418a7492f9adb20ae661e06de9251da11774f155172c79d54d320d5799b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4880e7d350e93766579f1af49bd6ef30db10d485d1fa6fe80e20e2da803cd29741fe0cfc11414edb01617e3094f2814a37457fab7485289065ae311b743aba2251a2eefad188059fdf842ea5b185ee0f319203beb0dd22c10ccde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h178d4d2c37a050e5d2bc141cf162334b6c1ba1d86a5256d7ea1ed6a4f97fa93502b9beccdf57995625e95cdac597af626873e4a15bbfe35a6627d7178695f135deb750756ad7c419e12443cf7194e06460281c4662e218112603af3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15475da680ddf01d23f4611d0b7853700265af0712a1782230854c3667da1cf3498ff739d842c4d5a99fbdedf54c1d7b2cbbe023c2d18ce1f627a7ab198c75592c677db401273a57fbbfb467a84c74014650bc9d38b2ce9dfbfd1fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db64f0d6fd2d194dc27313a9b201c6e3f335a28327d00f2bb6828fcc21c130c121f6fda1f4f3acd9c33715f3452bd2f97f275c63929e08dacba718b9cab5c645ee495a94adf070b276ee738e45ebcf88ef8daceaa5e281c20a68cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18fa7129eda714002004c9e8740eefb3f4bc735cb36b97cc1a6475ceb22705ab1c3e17db3b547c4fbddd0b6f3ec4ab894597a4121092dd2cda8c01ced757e3dd26c8c9ae9251e7f36ff5e4e93034c97a49a0fd44a1113c89dbdc3d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11347c3dd9bfa18c7ac99100f74e000a6f796a5ad9c730a563316ba61023acd64f6b2786ba3da8ed3173c9dcd39309a69a1b237845928009718cfd756081cb7291be3113037aec3d474a3b53500ad841e803130e8bbdb2bd310de86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2fcbbdcb2f14a8b18170eec257108e2e21968d34ab4e20443adaaca0a34accf4dd628953fa9145109da31b291ad6f8ff931a7c3b4a66db61eff0fcfaac70e1d44c24003c201c6761330e9cc3c5406366d7b545bee66c5dc8842047;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17baaaf2c54ee5608534df088a1cc9f6b1ca3922d00cd7fec236d00e3698632eed6c190d80eeb407b150d7dc6ed66e3859c431daf62ca1ef549725b42f03364f5e713524e395a707ea722afe1b478526071451c24a5294055512da6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd3c980b70f9fc4f0c53708f93988cb917ec2d51ac8c0de01f938751bc405b258d11cd6d9257453550a6dd0b483ca71810a70694164a011bf9fcfbd2fa6d3041a8ae6ad899d1a70b5f9711ef48af86893bf345cdeaf86b6bdaad466;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e7956ad1c41a6cab7669ef6c4415692ae7586b4c832304fd59c1ecfb4007db03dbc5b439b9c966c0166c37895bd2c47822254c73fb8f1c1da4b6f2f04a140b32d3dba689266c0aed93fdd6104faf38f0067e6770a7b72e823d640;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3fe6f1b1e04bacc45e3daa98ea50e7b757cfc175738a6200a17c48aecd7814bf8683a3005040202062a6c6d57069c61067cd8b60b00cbe8a96e56ea88574673224e25883dcce9af7931efb270d3b3509ea89a0f4ee0e2877400975;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a1c38523d4bf99b6b0d71a41d1be2f7cdd42f40dd479a6e799d3557d4608a0623455f397ebbfa1e4e8b9fe8262cafcb92c1baadc0ff597addb70a978110830b05cd32769be9f5843da59cb5a4e38e2e34a306ea25d24d2984ba94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de659c6b4a411d968fd4c261ea65acfcc8b6a51e652de718d04b8641c43ae563da15edca7ae77adeed163deb15fdd5a28bd06bc4545fe74787b3cf88de30bde7792698e5ae9f1746fb36ddae0fe7234107c21ffbbe0b7a3524e99d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfdd877c7ab1c6d8fc697a2086232d09c6ce87c3df52694e8186c48679d740b06156df7e69e65da50320fa08bf9199457d8f09ae87b5b6d034ce97ab10aa4bbe679f99fd9c51daae555537bc5452c2c46ba2e954f57b2d549526ee0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h863b282edef4d2395781ad55cb59f6946a9b764ea216963c7ea259bfaff105e9dda99628400f95c92bc18ac9a81c6bdd5e0aaecd81447b580539e272341f95c8ac38ea7033a6be8b3e45dfdc9c86da23112838c89c0f80dbbaa29d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130cfb423d5e1d84d41db3ea47b4a7ad421d14fb62120fc9a3702df51872ba1b028a91d3c177884313150c9a9a9a5a9d6f151b3475f90f09ee3d22b2db05d65b8ec1a5810d8421656abb15c7e2d20fc79d0fa8f9f400912b09f6e4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179584d3fc2e69df00b7e50add62c4f434328696c4083704bc9ab31b4f5732fcd38565a80b375d4c02c91f7fdb88f8c0c09d5147ea3706737abaaf79b2c1b969a41051872959108676cb538049d5db58bd5e6d529f47b36c74cb96b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf3dbc1262f3ee32db6ec12d75d54096d339a0599aca67e1dd95db3bc926f23d8dab9559a9dca51c18f8b9ae298998050671cfe0571effa8bf52f9fa24e18300a204f6b4e80bba2adda93527f26c0cffe6ff09ecdaed39ff4ff907;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187355b0f42f2a8cce52296fa5c5139a496bef1fbafdf8c99b5aa1017e875dec6f75ea678ee722af76bf6a1d0b1f83c18d8829ad6f67de18e7765e614dec8506a7e173977810be5653de1c413125f09e3cb2e6622a5c1cd3330c088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d76989a110f2476b7427564eeb58494fdd70ab5a00577e52b6368a7079272533d02e6016372beee3dc54932a9ee8479ac21ae864fc76211751bc7a3a859935a7b85fd0ae1b9d956db07d903c68e5d1b6fee5ddc74405f72db7ad68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143673492f3ffaf059810ec4e8455b7f0a037e4ffa8473535c3a0f6425cd815109c3ece89b59ec88dcf46e0ec9b6afe503faa2a7b85da2a1168ccd03754353f081c74c431cb63aa654afffb8ac4b047c787500ad61c6f74362b5411;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98308b7f040db488039f99732d4b124b3a7505a8801bde78c34393ae4d8c41b3c9d4fb638203b9c777adf330753cfcfdddec41dad17be225996cc20e3646ec1ad13ad9b390f11f7f7d6797f04a31c158bbdc37740d35ddf48ddd84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8f93c511c34259eb0523abe2aba7ab5f382dc8cf0983d5d615ed9fdffeb1322a2fd8d10981b26dfce09bbfc84111c761a6f3416bd2e3a4536e793f172d9c0f25332a1ca4ccf4d481e417b5c58bd9225a41ab64b67cfe26bdea96b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4655f7f688abee3626942702269c515650b3d5883ce0434fbc40794a1fab60788c3a5ef37c477509f86d8da37be63bf7be80da3152303a47306ffc7734430e63b9f321588f284fddc38cd740e1140fbb41c8059d83049616cc174e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f4e1a7d5c09054d4ffd1219e4bf18634466e07a4ab96c379c633c125633f7e8ff488d125af5a773efa8d8aa04c352aded97fed65a203f29ddc941acd16caad4f30ae83294cbdbcfe727ce44abd9b8e2130c8f3dc321bacd5747fbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba7f71f69570f786fa7c3f3ee074de4721fd516a739b4aede5b4a7b2a826fe9ef2ee7739641f544c228897c3395072c78e8e84198a6219f8bea3368980a91eb74a7046cc483c0e1e24eaeb08a69b770b9f25b7b763a4f1bf318c78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164ca07cbd69e3d8457b7569066fd68bd2551ac02a9126d92709dfe8c0dd22624543a039ff2509d6515bf3abd5e7a2d0810a44b64814cd5aa4adfa775c6b85fc05c6995674b8fdec6aff454e8cb27d22c71ddad69e940b4defe5b69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h75b7472e15e50fde34d57738f56b13a6eb17862fdbb552e3146f8e419e446a1a9c82d730bca0628c08cfcf7d30928761b04f757164a4b3e6602c63888d33fa883e30123c97d9ca3a385a664a35316c8cea96dd8b69434c00c26aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8627246f2e55d35690fd420856937fc7ac5fafbfc2e7cbf2fb89ff1c1f3fd987087bfb2cc833d17ef9d5dae460e38876b5908444cf157c41cf5bc995fb74bc6bcad85d6fbd479909257fe95a94b801b9721c2ca2ede95d328de0cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14672a4b90bcd1c8567dcc0585b7772a42756dd2d8b9b31bcbefbbaf5f34b3b093839aa3bd76d1ec0eef798a196704feb06ccd2e6f84ac4be801f15e50da0d1a7016727281868bb28f1aeec84a9129f4936c8aa699a8fc82d1c07db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3418b025349ba47f80997b7769972d67717b83fd5e20b342fe38f65a47f31df9307b4dc185bcf17ae470f9a68b16cd8a8489d188c8404aac39470b27b3cfed787290f87d36fae2ce92e67ee798195b57dcdc4788d4adb066717f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d9390df67c7cb5c9247bb5ba6ce5f6702b22bd44375a4711781cd37b3e5c2782350667dbe914d83049358054f3841ff0552d8fa03dd7339b59b7eebdf6d61d882145d7401ed8bcbecefe260e6c3e13cfd3a8330f8cb6f0bd23dfa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h46872e6adee6aaf663c75ccca4251be0e798cc5b2e6bf4d739bfdd656283d4f3bfce67079a87bf97a929b552a73ba231b8e50995680985625439edf8fae81bf0e6f14f4aaf765090acd7d6441f8fffdd239b68bf9327f45e4be015;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90bca635beb90471d1b43be3794d5efbc6f7aa645ccb4d95f7f07e6b26d13bf38b8d62419d5e1107a82c75a29b72be57657b4ec0c72f1bcbd14ab15e68e7932861aed79c3156e8649e687247af638039a02c0c7e2a0fa8e337ac90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1108518188db6316afef3d1e5be3b96d0a9136f1d759ab5d0497d0c5e8b13e0dfb05639e3293a516c00421715f0a7aacf6ecd4601f2fc0cbd2f9937baf1f6cdff4a1b77f150e4dd78b4d2efe66dc3b9e246f40ef48277324afd8ec3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b04d90a04c9d02004fb1d84b13c4ec4ed25a956436370ccc12d1d34d33c162e2644194642b646bacd060df1cd77de217f1ddb4438b559936e62dad3f387c3e691aee9261d3d9f01680be3e0484d7beb73f699beb996d4eee60152;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h186f4638d2d082a28563f0a5c4c81577cb2ba213db01d5a76529476cfca1d45fbf3e4c00978532b0f7b2b8b7171051d9c3f0700cb6fe07aa3d66ec56c4f97093c4a066dc114b7c197ae9f82469865084be81bb0ca5781c8ef1deb2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f2ee58e5fc63b00a096b7a6b551e2d944ee6103c08d047ceee14f2b78cf5521100f5e3157584f094faf4d07eb720122cf4fd42fff609e2153bd833bf4dc8037be3980fb9be54d1fb8711877f4895cdce18b506bb1a1bca9f996ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14226d8cea91d8b99ec9d423e4a74999a7000b0786ec5dde642c4890ef12386196c74ade9e485597e43f7be2c36e020679a2fb712a1173bfe42a33294de0c5a7ebbae66482f9ebabd5334ca9fa8318da93bfaf4dd7f5cd5ab1b22c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf169ba365e6733171ad9574752cfa4a30fe5f445ac530256619da9642ed322cbdd98ed88e0465e6b159f93ddf3c80c6e2eb09ea12e2a30e0a8a35ff218d19f2d005c39156c569e4c843032fd6c27e9ce34e49ed028a1e1e772b6ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h762b0ba64bdde9d1002a6472f5672c20202be4456966bd1eacb2685d95547c3a4918dd19acece1efa864535c5024be79a4fab8c313bfb7a271ce9a0c9fc1b26311bbf8cdf548e62f7e3690ef2c1cd4e3eea6f5210abbb1a4595843;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b16497fb98d2c94cbd7865b351828883c141413df4558e173b19f091eb3459200482d35568977628bb95d8d298c8d16fd4a03748d0e2ebeb66ccaa30697f6cac8059a7203f305ce3595b988eae2d9550bf1ac9e3c7fa2130517f53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167ca1119366ed67242ed4ff9a6997fadb6e521b7c32ddac16a5abc6b008e595c421de883723428905a560a155d93f1be0788ab179e6b8d64cde270035200a978a69420dd6d9ef540b68a33bf21176c9936b9ea26c104445d60b29e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4d7a047c3b6f48709f5c97553ee760728b437f4ff7b343cdd9dd8698200f0694f502865d019570b321efbf55d5083ea33a207d98886710c437860aaf98a86364d765b59e3a37f1adf5b48c1a4515a1ae8bdb2d461bdbe53991509;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff2fb98fc871231ea8691bafeca8564d524ff7be4b3298d18d28a1cfa3a87118507a0e6a20dc81843353bae154ac1f1e74808ab2033e42fa13d59671071e472846cd53b4a55dacc8ca4b51183834f22d96fbc037ef3014f2d08efc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a681d42d1d5fdff3054f809da948a4ca1069a5bbdb1c4bd3558d150c695f8c2e2f4b0da2d740db42a6360349a18c6621d6bf8117c19b4ccdc3ba6de077ded2f58a01bd9e023029333ed00c1c9c60f20961cf43d65af2430798ea2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h94d1140f21998643172d1648d1a1e3477b3681d76c34291047930b040aa9c6966a21031262d9cd63f42925056cbbcce45ffb9113470d5c03ee6473e6cb1e098d6a3541311b5a9960dbb678fa0d3332a4ba4ea07c4d1f370af18285;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133b262ddf5651bfb0bfa099b371c083425efd36f1ff361466cdb042db8aad0f2efbad77c2609aa9acd00a109e3cf951b064a1e364627c9fabbbee6aea9983be8cbccfbab4d852cd98b3e2d01738ac41ad4853c27a0fdea6cb1d68f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2bb7f271d4ae1362c18d3825194a4d535c0bb4169c20967b01b91fefd1750af8a28c99daabdbffec5b6ef8dd228d6bf3e4d6e256a92bc655bbb350860b84d9af093ca42ff3c41c05e0d0ad9137aed480a71881a489527f1c03500;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bd9c0c77cd4ff618e88210b5d7bf8c584a227448f59183ed734ae355de47ce5bd40c7c6af72f7cc13c08b9b5d6dd80e6cb5949ace20ebafad9ecbe744ae7d3d42cff44df9113f2aa6d9eb96f942927faded38b41e574e40d1f1dbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h140f49393c66ce61b8c6b19739702dbd3b8d521011ecab1343e76f7fb97c5dbbc2fa606c16101c2b51853e12c84aaa0e5fa31e1c2df06a950e35db2a07131c477920aa174d2086f227457abe23349e6405f303c622c3eee8581b02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c391196231cc8e3374625814a3f763da55af9c60da2086bb99e80058d5d858efe5c3b1a044686e4196a7f9f1e1be3b17517be2e7b96b801d3ccd9034f0db1ebac6d8a5159f15e86e6e224d42516486fd5c031ee789c2840d7f9ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb89704cbcc742aa34880a40c32a1a8eef58ac57f3deca81d1115e5da41e3563beb4f1ab64161778861f4e3af22db30d1746609104666815bb77c58a14b38e6628872d9ed9b5df07b33a6619be934a7b3792e3f09becea443872732;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79e12b9d9657201dd703339718f7e03927d96a2c32f53256ab360cb7e1426ba3086819c8dbb8eaff7174bbc7efeb328f0d22b8d9540ecd9d5050236f7d74684a6576c0c0be14f0bf358ea7bc82fc3b19f1e9b1146a9de0cb2ef583;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db1277eb9f9a83b683fbe634b4abc0cb4e5c8ff4423de8f7dd0834fc2cb5caeff24f3eecc9c4cd1844ff8fc5d268ff18ab508136fce2c72176304c5456cd7bb77aa7b1e8d709571f9f8b1fc30de2a484deeed6f546b73b38366750;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h118e9f923f5b501d799f29ed63d89a7564a69a7fe9cc5ecb4eb5aaacd3484f0632034032d46cfc475fbb63add3d1c14916abaf9980e59bc5bd9a78ce8ded443c98c47328d3642782b023f384e054611c1e32f9046dcf432a2c943dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e61723890b0b30cb8fe5a6aa05145a3f4c7ad7493455ce2134f89d54c7e5b4c3c1a0adc98ca4a5a530a3bb51af91df1a209c5b06503a2d564815242dd4a64a9d49cec02ce83b2ea99549e2c432d769be9b0d6803cbf02d5d5f90c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h642d194fe77b41d0775135f1714e7c1faf5fd04b8b62bcd0e568fbd4089a445d1460c875576d24b41fd52bba6c6663195e8a6bfb902513ca20cf46eb45cd081db8fd1286ce30da6d4d88d2f23db81940c7b10058218ddb9c8f627a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123af7a925703bd43f655e2d0c66b91aab1db12c7dd9a9b11d10d936ce5fc66eebd614d9f293260653418a21aa04834bef0333252ce1c3bb599fa611b0de1fc37b9e5588e3a067e94332e4bf21286777695382878f7993a5b69f8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf19f369464f5754cd37cc9f6eb11921c4c8721f2471a829a7c8d76a702587544ab3029403495bd622aebbf957323dfea0af930f7f3a94270af1147fd2efe6b8235c82d3f5bcb6f0686e251372ae5e2f7e6bde7da93717ca5d21300;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h117fe8527381e7af5f9821f86cff5e3187bae0c15ae2d1aa5d72e27f619f912b5c3dda6c581db5e2ab09bd456709ff21c9b3a939f67bb9aec1069e421c078226c486a335f024493dec2265dd3398a5b7a0e84b08e2ee4e50c60db8e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14af0768b6e5324b0d7ae196d9b2cef5cb84b103613453e8a69a7ec75633a100569ede19e67d8b6cf34263c306c6aa32951de0ac952426821ced54f9273fff69e0131db39a5a0dd890c656c71cf59ee5ce27e288aa3900d8966a884;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf19f610ed00312ddc8acf85b5130cc65cee96a273442019f0eb2c746930e5dc549328dcf034f11dae34e3dfe9691b7df0f80ab8e4d877d316169016d36ea67cb934ff89d2e66c587b126c51cebbbc80b6df24b3f28c397ccc5e43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h117f580097e57a871c1e156dc325795515ee36f1d0c8754aeffcf26b7189be46d15cbb2f2f794e84d740ebd82fd2a9aa708fa5ce9043b3412aade37462a726eec3dd318918791df97ad104572bf7e4ebfd824b06705a149806f9ea7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f8048af57f126b42516c62eee9b99cb81e8dc13ea5a1906064a96ad1cb0041d889070e80b81e227ca7b81f18fbc12cdc0a4e6b86769578dd8bfe16929ac7933a9861a032893b94ea8d23e7a9fa1dfbda70d9d5961c09411a935b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2142c179cd569b4b600134e76c2e79762f2cd437928f16db65d157bf8e452a54a411f4119084feb4afe886f5e1f5ea2f0feff960fd44072263dff9c3ed9a16d06864829c74c9704569d814651721dbaecf1a7aa97dab8164ade27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb52538b0e7d07553d21fc2107bce796649422c1b26b112eb124e702250f8829a710fb9bf27e754e1512704a81e7780cbeeaea4bdd1850f53b6ecb17c1a1ed9bb15764b180dc3842330081a1a16aedfd5b2045bd7aef47f031f800a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c9f060b85c7b65e33aeadf8f705a5b31b0e2daf20d46d6537bd19d465349cc01ae18c087bb13b005eb281c9e49c1ba14936f0da26eb6520f5ecb39d2e2cae0431f808f336a5fbbea725fd1463204e1889ff08b1f09712d8a82304b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h84eb97a3aba35d17b197aa51c39d95ee6c76a646a0e2b2810a7c0e77950b772f3d9937b799d2bf3b9c096e77a23b57cb445ddea09a496925d3c0c8f2d34f98d015208c2fbce266e49f97ece4ab29a9cf7ae036308a463a916a9a90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177b28bb04c7a5ccb8d3eeef87d12b00f4ec6482aaeb10d8ff7b93ecdb24b6f181094e1d61d1295a6b9117825c0b5de9eb9714f441a16c28c5e0ad8b6fcae51283eb73d4da88a4753dc9d7496e8f2ff2cbcd9b247516ac2cc86770a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ff889db60ffe52743c9ccc2a16d4a77451297e82901aad11b36d0acc34e660e27bf042276af88748fa01efa25f192670e50be599ab80606039ea86771470c8ead61dd8a9718526eeac7a90fee7839a27f774737944eb6532046e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a638121991a3a95d06175148733aa29919460114a7791b920a670f66aa51d1427f18523f039d2e25af3eed5c01bab6dd1ffd2931e07738b169eee82e0c7e5f7ee40c39b4ed136efc47d9b17bd73f1195d1409822a5f6ec4eb9d316;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1191dc823daffd6afc2589ace714f3a691c42cc80a67ac839150b185709cd70aac3da57ea293347d2626b1847baa7a872ce8d9315fc218639dedd4a0baee25058ff9d9084fa1732ccca35b985a62c998ec786ce7643dc3914f0714f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3654eef16a18159f5962b50e9832d09839cf341b1ac309893f6e817a969eb1442d6884591310f4071970cfc2621cf636fe2c4efed45cf9949925a4244fb228e7bc3df7bef21cbecd49110df60af529007e9bae63fb4552d8dce7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a63703aa6ee587a5abe2a669121f79d06c6768e814815657e1ce90a5226dd2f86e36ac356362fee8b03faa33a7cc37a01e86b244cd2eef3f65abd7b9f58969173ba44d4dd5c157d9b2d108d505da1a35c9f1ae027d21f3125e863;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e93f08dbf5d5e37d67894772142774d6a0916fc19f802222595c436a4f3f7fbf782f6e06d8d41c4ddda3edceb343e682d4136d8075de0dcabe165dfdea3804c3f3276e07690cf08e2c706bd53330ad77613fbc81fd6773d8d9124;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h401eed00c11cc33806da1c111a6a745d0615d7269a9276c7fe9a2ea282cccc5323d1e89098f62bd55c693bc5df05fd1b207095dacd715c5ab1bd78497d751951cde80e200ee79480a4f3fe28730de06daab621c9eba86feda5d1da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7345c065350851c77a386873722f04995da7976aaefdf20c8a4bb4d8ae7adc668c89f728dceb308198155c41469c376f7594b53b61dba16839d22bdc424a269d7808f5951e1a4b1e7e64c2f8688497a480804dd0d74c451742a52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdfa47bbf300a7a569e4c8f1b0756a42e8890c9b0caa44e166077aa00a24ec8f70083aaad455ab0407e0875e5bee0364248dc7f20679750a48bb8687c83b5d0d1ba98931a2c168158a8e0c137192f835c80b575eaf9551ce55c1a4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfdcbc01f66e475c8f1c300bf9ab4436f4a8865b25dd85079ba8384f603042eb9bde20247ea96bc41ed081d414d2ddec6a2bfc9f3ef4da5912bf861996146faff8c18a20dee31df5eb7d1045c22718f68b804fb114cc439ac41bbe6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b42b6b4dcb4442c12cf98ba3cb889771dfce475f7b6c81bcb4119d84f5503db9eed292c1af778959d9b6a90a4518770ebc855282703b8fafb0e00f96ededb14d4c46054dd749a25832c4b73455a38df0dd60398084ebfa399b8f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b50cbb393a7a38966be689052e0cc1af20e79f5e224333045058a153a59b9f97ebf05b041874d7d75cd19b051a1d44cb9d6abbef7761b1cfa63310bd1d3d12281c6a3c3c6df26f4aad1002c71d8e378f46f37ef7e9d79af6b68283;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c80e3aa6cb906162b5ed974eebf12b80bc00bc5254826c6538103c2313f612e15279ff2ebc246b818a8d535198771a2bb98a239818eb74d81fd27a1bc417f559b280bbdb01366aa9ca2f0437ce17295f1e34abd0d3b59c71d09c79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h661a5afbeebf96fc1e045cc0644217c1ba15946bce7282f5a915a09f6f00fdb47dfa87269bf04efbdb77e97b396b3e836dedc29a9b9c4155f7f61cc5c6bfcb53e0b2ad3d97fc6cfa022c32b10a9cb824a1c66c28d33e2f3b81e131;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb783785e3b00cb6aa86bf4e6e9e305d16cb7b7321e1a2d4bf2355595014be5f7534e5a43b2b615b9a1461c4a8da4cbe643522abecc502cf166e4f1c3f4eae3d2e190dd406b502044f88bbfa0869b9975381afb681f7dcd1102db6d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1974d1b362ad35581b12a6685230a502a65a8281876a534c87c56274273a31a9b69438006f665202d59e5a2fb768d65ba98cc20f937a3a48171069ec9e592a114a9feb5ed8c769fb58f4e8f38362c1b7fbaf448103ae482ee0c2f9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d8f2da211ecda001b4560af2a514ddbc2a93f44a18c1c3d0cc4a56a8c48f52ebcbe50f4bd0378bfbec28571bfaeb0c65cdd4c59b0a2d2db1f3d42b87e69865827cebccce1b191a70481567cb703d7539e4c18a3db33ec4c14c082;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b609afc4a6cb085e6e3163c73ebe396ec6caade4ad0beada3eb016b8c55b8edd814c74cb69e65105f2eecec57599a7d4d256c6c57358fb110a94a35e6d258ea0b7a4d611876ea0834460d7104f0bad314fc02aa4dc86720cc80c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17aff7485c16379c85aa88e23c8e2ec4fd6bb0e64134460890cba53ab97958d4b4b842f95dce3d8b76e3458720903a25a57746561c9b00e3f5ac0003ac4abdd440f7c8adc68e602761dd05241aee72c98193764234ae20274992b51;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1430c61914f5dc1aae05f97d4a77d99309bbf3a629086fe625d96dae0465548d754d81dbb7076583b90d9a2c1629f8bb75601b11fe4955560d57402042f6fb6de1e6124c5c964828a301d256981a4d0c1d4b5fee5c352f63e742dde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa183c766d4071feee19b03a5c579662a0134195ec07bf6e1ad81f28687580ce0ff2e838ecffd25826eb7d1b48386f99c5351adb10a4be04a882cb23d5e416d20a49719cd27b4ac04173dc9495110bf358c2d24419f4d0ef531876;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba22669e02f2b1f7bf92fa58b1753a41ab9dcefe76fb027e6c7f0076af29490a1e61fe93d0ad8c0da5d2061b7c18225a1871d122db42f7ea3a5c889e07388c18b0bd31089856722783479073524915d4e61d7747cc9b7328035053;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1969f6e4e17e64f8ff501f84d08752a7153c323c74950ee1a0287080d9f3cd939c39a6fe663e765247161bdf0e1761c5cb9d359d021ed962828af85bcd72af15438b4cc78fdc603ddcab1cf9d7ce1c32d9f6a4b692d5d29b09fa7b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d458a7735f2753b66ee1132044f2f7c778d47a30f06025ba2a4e431b07eabd64ec887d16de25e4c12dea9a9b8eefae826e89f8f329f8f301d9a6c18f06d1fbf7b867300d3f72c4327799bd5d00dc2059f6840f673ce65b7b9a3ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f96efc49d7bc9e8daf206947afcae3d03759e743a563bfe2ba8c1de463c4705219864123a31402eb8f85205bcbdea4cf6edf2abed220638e00fbdf6e8ae88469c13b2c5c13567fb5bcd9be7821801c9ca3e00e5d7d80ffb4bd9b28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19089bdd4f317b48d2dc2107de2fb1460b71634d52031d68eadf7a3b69cda23b7c2e2461af9e983f4493b4f87451211b25ac8b51ddde7d99b82655d427c3fbb99973ace2c9515f22d59ab566e14561a6f6008dddcaafdd88a59c1fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148a12998f4223a4cdf20e5840a109ed2490d69ed3744b268c20ab479c710e37fd5400385c5820d69e46af13d9fe59c294a67cec11dd21e1f19bd1818a4035fc8a7b16595aa92d9d805ee671fa4f597c21890a4b86ee31686a873f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h497808b6c873ee4433be6125e7e70bb783a1045e9b76600beebc662b8d42dacbd0d95e420343b2d2c97b7a4a37ec2053bd7a8f4198860e35e8f111d800bdccf4797dfded49ebf90097017bdd536342b860ea7c3620e131b0ca3c13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f273aac920be76b16f3acedd49007b855a87845ccff7291d04fd451789eb3f2952c3d6d82dcd9689bba2797dbfbbad7aa532769e3a2b138805b8aeca6938788bf3211a84cd81ad380782f902a866cecdc530164630206c1a70a78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a18012f54161a67908ea6748b190ac32a1d6f3fb64770042e9cb62146e42da6f35170bacd15b8c9721a39bcc030ad26b06fb0d611b5fc6de303e74340945a26387c10f51599f541d5eeb64df8c576d80aa05c80bb7cbdaeafd32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cc4707a141c89ef33769e428c99881234fdb9cfb27008f11da18d7b1ebbf5e145f5bf97c23942f77001da244145930ebba3fc6ca9279e329842e20e63a644021ed78cd97bb60423ff04a8d74c95720669170bd34d425c5ff1df3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25663eb0477944c061218485dd1b90e4b977a86266346cbbb796d680aeeb546e5efed99e45d5dfc35bb304ae68f66831b8c3ec6e8c8d654927ee1e7929efbeedcfc1d4f8664370c1dfb03942f358d167d4cd965cf94f0d68b6a4fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd936466a4a8a97f62956b143cfad08c81b7ee00b535062ed73d256474a3de889132244cbdeef4d432ce86c39f44a806c19190485adea077542c200f90192e0fcbd049b67a44f996745ddb6e182cbd50f94f10c1a12eaa73629ce5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf487f148a9e0226d2b9b105c9fa9930469b36ad160621d788b6ccb6c78fa2348d0672d6732cba772137e3dacea9af5369cf147466a49a3ba87c54b158abdc20d7a3b000d445a84e9f40550a283443283a17c2715d364c6ad6ac3ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1720ac724d9548d7220937d0d0937facd9376bfc14cd9c8e71e94914c6f89e3e5464d4b1b3332939743aff209f62884b4eeb2870b45c06a527c4b88d15805b1776d2ffa2d969117904f279581ce797148aed6313042d0ecf11cf381;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1abbe3ad905f36c30feba0b7a83403298647c13359268950314b2647fab2c9cf5b784561f5b081ff45701a5612ebb44fb2304c66ad5aeab9777f4c8d9f9fce9817329886d90b1b270676496b02c8bf589d555ce233f0cada810d589;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ce55061f3a99b778509199ddd2376ec027382a1f13796a20cb2c11f05b2161bf75eb29d7288a7c55c611e3f50b57b71dc957f32be42747f7d009c89a81ede25635a13edfbc362e4b2ee9b9bd1e8e8b97b4119e57e24626adae307;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f307c120cdb4e9ea76c554aca67c114d8b91b9dae40d9456aec88be7db9a0a8e103bd8bffe91bf3b4061063ae2bed19a9d16a2a507a9872e0e023f727b7570948a03b50b37e30e60dd0361f44029569814caa190a72b4595a3113;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hddacff1060b8c2600a936312d2c0f07e79c4d4eda9cdb0278db0654c31f88bfbb270ed1b0548dc3aed6901c6e554857ee9253e13043943e410186d448dfada088c7ae0e328b79ff8eede0a0c79e9cfef8aab1037baec6b054adc84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a48bf97d9df083e0c582dc25c069055a778ef791eceb47c714c7e89a556303a75fb98cd6bbea22c5f3552917134a52d3bdfbaf32a19f24e754ede24bd22f47b0f2ca82f03b36360380d3ead852a427e5365fd40a5d972a5080e18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b454bd756881c6697d5fbf5cf6b8341119a5fe4bc960e1901ec12510847004ec088ff311ecbe353571d6909f7cb9e93eb0bd982cbe29296b30893583f51e00bba52db228ecf7dceb0b90d383e858acffdc13a53c735fbb575f036;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3400c574ba2f8258f2e1b2bcb0ef4abdf50d68e9732b2905241cf191651c1cfa92619d01e2cc683c60189adaae8692a8d6eb1d795b22c4d84ba622cad3a654d75c197e96e0b8c0b58c83532b0ea349d66b0d2463ff3ba4c74010de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1145ba1b80a6c90aa6820458363c6d34c11b91bdfbf8b3406cb31911f7fe382e0c7d180eea7a9f02b38e59e4405b5edbedbead3ca910f45f645367d7d79e25b879781d5045a9033d48daaf74998e9fd17c72edd4cb3eb0433f1ad55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd659622c5c533330b881035e3d6122b2ef5331954bd59e4314d33108023e1ed31ce0a19c9e138ca8fef4e2acdeec995db318b6ff7a800cce01947693dd220989643432c78606e39baa1394f41ddf458cdfc41386c018738fbdc2fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2e18e78755bb297b438adff71ac6a5df5816a3dafca5d152bb8f0272a689aeae8a9be0e07961c0d0e17331cccffb83ed65705a81474103af398abeedefb4fa17840e296efaf1eacc02be9864f6c03d723ae38c2b5ec7689371b45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8856294a1dc36365d05fc44c9f1804f7d31a3c2819200a93a19aaebe1232972d95601549897a7bebd4124afaf87b85a458b8489b8942c006c297105c926b856663bad433cf5a6d29f29db5c5fba2fa16187a270430add7a7cfa3b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0f3da7cff694bd8f5a8acaeaed500f09d7dde1c0b57e876fddd4e8be4f3b13de79d4dc4321628f21d1593c2fa05e2ee702928fdb74f9fa6b0c504c3274351a409ff978532b705b1ce7da898fe3ee8832e9d724b52eaf373fd3bfc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a45abc82434f0acb75ea029da5123174b0de5277761cf935583a8c2357590654a4eaf4bdc86ca9851396ea0343785090d2f38f39f9c901f884717011e9e9e511c052d4f3d44d9195807352b73beb1df11078b4741b498f469e400;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ccd2e80478477cbb8566f5fcb4e5961f1afc157ad0a0bac4e535fc28039eb304daa16a79baffccbdf848dc7968f794523d2aece62efa9cd482cb5a60386ed6296e386529350f3d6ebdf8aefe4c5494782443ba9816564390165ec1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d554cebaf1fe8da5ae044ced74a7abefc02ef7c7c6405ea287168b08a3f81d379ec7c18a6424a38f9d58e8ac23004e97cfa6e4e4fec0faa22e469436db49fb172ef31575e5f3b5535ad39a051273f26c2063081dfac5e3dc20211;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e85f98e723a31b9e5156ec339962cd4bc8fdcfe7653da2473da8d1ba1c2ad8613d5b7d91ceecce755c773dc561935710101496d253f896f112c645df68467ab51c70612cd72a665156a461981277ec885d5873031e68b0c1feee8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb5b45bb30c876f73bc20fa46a878dfa8e4794e356be0095a2032eaa8891fd48d47f57723a1640d89ed8ed1dd8bdf17c900322909281c7e2c4ba761372b8d81e08bf46696dca96f99e2f80d249b25df49a4468b944aea3a9160834;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb6c5ce576d031e165976e8808cda567cfb6b65a61cc51c2ab764530e5f1a90bde91a141244153a055a77a19991f8456533370c1f08a500a0dc50cec10b29f2297671872afa51dca4e0ef426b4ae562844f0a5c506c29e9a6ca11f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h804783a6f8feaa44aaf6ab0af8d3ab27741ede3019345008f510fd1608cccff0fd081d061933ce5ce3eb19f6a2da38e7433bebec7d3a03e5995606121dac06b2d0695b0b3b655aa4e5499c62634f8de8d9270676a62f01cd1cf095;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h433e267d2d26d463d7739dceb2424fed593626972e5d59965ca9a200119a3352902eb06d9fdb04f1dd7eeea33b1172c3edd4298e25ade0f30a4d6fd5db09f2f197571f11460daf4fca12140a756abd9a7be6ad57a177e296a2c5e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7e22b47e1e344ad0d5e4c3a070f04348a242f180d71647a912edf46c16dadc391d331db970bf28ea5a04d94aee9c34a0749186dbd7cb9504d335ec3ac8322e68f8a2982ee47a500f6bd4bb38bb8a88b3c4ba9be4ce65b5f21f469;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e7967eb3d2756a8d758fe8acb1e35d3db330de0e1449c317b279bfb6c326d1a2ebb5802ab613a14a2d9c51da14fe679f59e379f3acb81616e68eb93bf2605393a330601e4ebae47bdbf179f67b77a6bfec79cf6879e97cbfd3295;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha619eaeae8d7ea259a815557756b2eee8e7edf9cb0189d726936255d689560bae0f7c8c16833e629206e315f0617e0cf98903f925c0db8a4afc0bbae571f1b7f5af9a48ba32eea1e9b8e4c92be94db51af4994ec50b6fbeb315558;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8490ae083f972d3ebf9c5275fa1ed74d203c41c16a015d169dd883ea2951286cbee7d4370c21d2fea7779b2a2099ca1bf877025f0547f48132a93ef49b7a21fc82ddfccbb2518a4633c253ba0ada67e909aa0ce99ae6dfa42280fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2ff45d53cba140cf30090addf2e051003f1a601f9df3437ee04eca27ffe5956038a7bba52107b658e2ebf78eec922f36769befe6e6b22d716b198e7828cf0b6a6975b91d9fe4fbdd99eb476f1c43cf6e011960524fb4362301f9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1612fc86a0972ef72ee492dca8d1cde7b24b5f2675f577dba22c01cc404b9653a2c6a6b0201fa11322c2940828d28d14340a598608fa67fa9ebeb8d360670e0e4b5548b4b5d7a4d8eaca0756480d6f1c50b31223c17f5052a88a5ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d270369c64e66ac6c5089958fd1ace403a80ba34330a1d7090e84869c63cfc98bb7bfffc331a6c94d7d12a280117bd3f2b6ad10176acab9f0f74fd3b2e06b3157d12e5d989115d346df388cd56ce8c6569133de4b461357bc7ef3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h988b6b0e6ace795c8d6866488f0c420f64b013c493231a4433800c500f64333c217eeb0fcf8676610d6231394c69a0a3b86a909d0748c2cf39f7309eab796f4d59f71cf7bc4703434859cb82df0a239a62ed8993373dd53fd7001;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he09490409d4c815c6b934097dc80e2fe33eea98822f69a2bdcd3698ad4fde3e167ea4dfeaf7b41165b1e2c9e8f14751e2fbb20791cb64122287bd83c5e581f105f5a78efcfd6593c1ff771396b124a6a76d9229dddc0b52f42ed0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194e5e74752539b2f4a15ed480d699f407d9c63380e3edae9b1ed20e42edf783642d1a9570e66598693f6d9367fac8b7bddd9b56abab5c4b9610da22954c322f6885402ac4a6b108bf7ebe2fd13d668a6700f9e510e7b2f59076d05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4f89de297c17057df9f7e462ddd3216a4ec47aceafb88e397bbb8da37f791acc2d0b8a58a6fad5895927281bb4bfdf0ea57340cfc8b1ac9e262b0be8fc61db549ce732a40a2d46d021fa0688ea8938349f63eb13423be552ae5b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7941c99739792a009d6bb8f8dcc5f5beedef8f96fcf28cb58ac81c4fdcd8ed0e7bf65ec0087da5643c1cf17928a28d9e7441866727b232a48d2814d63c4ffdcd28b96424cd307ebd7263af543f7f4d1a1e25fef4131333b66eee8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf5f5bde9a0206da5788d3c43da83617105ef1fad73a4aad31c0dda2b3ca60100aa4e785f3c6f73e458a5d6516e9e907178173f7f7527f45b8afb56b71cf175cd873ce0683b0be7eb79626011df39854061a0cae112a5e88fcf251;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13e83d48421e6380b231760ce9c25bed2dfe3b84304ffccdc8f5cbb32a0697e83b15176caf275b5e284d1becdc2409557bff33d815f09faedf725afe963667632ba8e7000df5bb1901d0b2a65dfd93ec6ddca0fe11acfc3874bf33d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h149eaaa8cf08f7658f0997d6ed0fdd63401d7d0ac05adeafe4374b483f4c05f430dfb2f7b3d349a76e6fe66b8a85a0da9dfc9259f494b6875b10688415984dc5d2d0454319b6aa612e3ebb9aaeb5c2d32fd9e770a7c315a4134e6a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9cd7c8a83b49eb5ecba8e61525824a575a253cfa16430cb3b4983453ccae979f8b31c58ef8c47a6eead596ad2b12fb662a6276a8689fc06e8fb0e67e21ac582381484d6760667076231c13b855a950986835e45b2c43878cc8e2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c4a8ded2de3ef6449baa10061efa37d7050f85da85a3135a7ee8553e6b5e36170266917636ff785127df66854fd8a237d7519a8fdc20df48500816ef47b29b1499f1f2c0d9a518e8134f868c8c5e8649a42c23bc988f0d713d782;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd73baa7da515c3d2a3a2dc0f56bda7354f6d5e57d544c67cfbd07eb8d1684d2f7c0dfe59dc6ef99f7c8635efd9266b03f3c88d2141c9d670e3e7d3c6348e73771597a87df994578cb716a4552064aff0d1efa8b59b6455cdd908e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10959847e2cd8c4fddedc6f06138e837e8bb65a30df61002f6798886e6e2a0ea5664bd04886a5625035c15330230ce3623c2c16589f2b547bc8c9d1fa925ed8c2e4039afb0c58a178d6bb611ec6b42c149326b77f0a093c86fde10d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff340133dac8a4720f1f5060d136b51808e5557ea4578ba5b30791f22226ccf1332521cdfc26b364891a1a1256ae75ad3af78a34c8d0e8038407c42eda6367bc04f6256239d9ee902a38aee409fa571bb62c4753f8d3a31f8cc171;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc533aa7eb56d0e820934d4aa0f6019a6ed89b0a4605ab88791b450288f633877be5108bdc24236be325b70a7af615af8a69c5996f8374e0919350ef809d361edd8a2b1678f89beb54366f270b3294fc6a8b37967125e17234fb3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b78cc32d2133a8c09c0e8266ccd8a0b9c6f57c56315a795145656575b97916c3255b70b1a324b0d0df14e2b1e0b195d2630702301ccab1911838be34be6ca4198c219cc157ae8240c9ad6d5de154b2ca4c3711e8187fdc5ba61a1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89eca1644938f901b29dd99c77941f2a75935d96c5cc91374f1ff054c4b592e5ee91b77a1e520b02cf84fb2bca6a8dcee55d4f54d6ab5c1fbf8199df3d7b1665cbaffa72450ab812611d7cdaefa07af7d7440ced3554a45d5f4323;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h28c35762945ce547a093a900fb97b9b11fed220c3676b6ed4f9ce715a5e1a8736caada9e9f4dfde895a5a5b6bc14e69aebb772227677d97d80ed947b09f1531a7e7becd51e3abaef8b476e996c7b9ed7962b4881330beccf7ad717;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h844c4946e18792bd312dc2481096d2364d178decacc3e0e9047373cd9e64be3dd45e49a9cb6f504b304b0a990be5012bbbece6c94073c37fa56c4f07d43202137f1d9ddfaeec5f8ea18b93d212ff1515e6105ff4415382438e14eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1268151dba476b46281479332c6eb7901548453e3a1975ec1e7b3e383e4f90863e94b30a2993822f2e07cbb74e45a5fee3866cfaf7f91aced11ccdab3ce35f4d78f6ab81a5015141bcd409e51e53d0a72bf51f98ca188b2079d9c6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf4f89896fda53379dc60233ac014a9fa5e39a8d1f3df366d52eb62ec9563af714f33d8d2f5aff775ae1ede1a9ff707058526c99212d9f974896e2cfc1869b466edb5f4247ec1cf057310349d0068ab36bc78214d642d7831acebe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133c012dfdbe5340907d3e7b5454beec3158ce943bf42f8714ada78de1408fe95c136c16eff871fba5b0485c7cbd9f2b891a72b18d31fb29c7c192e092d42c0b6d43d6a7acb800b31a39b92adfa08abcd29f9e43263281e086b902b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bde8ac9de57a2a59509ab181ccc8fbd4026ec62b029aae28c52d7475293f3d01d1142fa46170cb9fff2dcd8e6b51effe00db3b5d0f0de49bc35c36f977f3c453d7d55b2e45f7443167babfab152b52551b94a9b7115df069a20f4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d60956b848e764a009ccf9691e404e175add1420a00e156d88b3531ee8eda421374700588132d4529e72b5e687c0d5e05137b58f72e2accababc514f08dfe036b8148c5cf13e31bfeadfb86626669f7fd17fc46543f92b206d6dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda188251e9237accb98020c7b7c1f430b8e005d311f9130fd29e32d4548d85628a54bd1a88f9c1030e7d74c112d9ecc2f31db3f42efb516ef5a5882f464204ce3bd2d90119b44d7c21efb158188e23cd1332756b2cd45b64367d04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1699ebd73430f564164959fc9fbedc836ffaa673a5e883d8e0dbec565b84d02f676f03a49ce320e478e2637eb284ca3e8bf688165f745747f3555fabac0e71ff148c490fc8a55048b83cd8708c18ce4b55cd092c4f157c7aae6cc92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ad6f504b6272f07707c440361376182b34898b5ca3cd579374277e7e301cd0ddec966bf5c18577b701e3bd6e81792fa6e2cfc7052912f0a40b0a3ae0217e7744d3ec418f72b66d24d2744ffa17cad63cffa9e7eee10b5026a8290;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11da6a4f448f948bd809e9e0de4f1fb9266d096e4b1fd15c2285d884898691f3dbc33bc1b380dc94dbf4b7f660792d5c37fb7cb99d441236ad44671cb2bb5ca2d93463a5c33c9227571b2cda23d757ac21d12e3dd662f7b0c4fad7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127106d5907901084aaf79eb9e84cfb1b200624f0d0719510fc0ba4afef39a32a65982e9c2de3086e6323c55bd1fa362611a687f3a8239227f6d36ec362484a734bd9d9ab769e3fa499b04de6cceed5d535293b3ecc01355ff2b877;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19485f6ec9514139fd46bb5297206148e13a71e6fc4945738d6b18094683e55004d2bcf43fc084f00f0f6abc42204f075b380e49b8eedd11e4d005a5febf3a68b3a1d59bb5b8314998d963ce1859dfd99d8b488e08767247a2f2426;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1daac4ba229b8d4d2072532fe93fd28b31c74fa76203832ea15f1280e3d16543f0b4188d8882c86c4f801716e860fbb4c261c60a6bd96dce3c23b21bc2c1cef6ed39846caa367a1962148511f2b03252c7058fdfef6356cfd82bfbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ec5431402d5111e472acad7c6a65413a4c0d7df4c7fcb9d96692ecfcda956058e3daf5439d1fc054ef8a564d6fcb252950c56936a3ee99c5a4dcf3dfa2183995f7305086d6119ef4e43ede71e7c430c00a0c4e5abeb01268968f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9f820b6c1eb08d9854865e0d8cb7399608b4eab0e908315a173a40d4c86d6697586149cc59ffa72eecb3ec026a836fee1e078bd75217e84b56051202cc4c98d6d5281dd06422e854643357b2b51f2d9b1d47d2862c1d838c67a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160a21444c36be956e1a74ea8b2f72d12d696d393af17076f1aa75900b1bbee2537db88342cf6965a0dfec8e80ea09fabd8375c9ae0415df55fd48efaeba3e814a836c5aa45d9995e4e659590eb5d2d181ca9c120e48a55c9dfa5cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he721be55b10b737bec36539245fc60feb0d9a85cec73c9d652ba6d4c13227111e2c84f2c8e80b77e14c3d4f26a8054601c65c4eaca0972c4aa2fd7c146f8610df08ca8f0cf48c245b12ca768d3ca51b966c2df775ca2b3b8943c0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b18ac9ce0aba5a77131de00f3c1a67d3c85a3f16134ba2459592111cdef010652835d2b1c1963b73f6231f908b20e4388e2cc043a84999cd461e30af7ef0304ef06bbb149dfe1d9f2dc5e18897c4b4dce4b1630406794ab59bf83a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38c12a37fd944ec6662aba2dda268cb4dd219e75897baf66781bc50f80b38de285464baa96a78642a446797c77ed427a13f79e95b40119cab34a6e495bd24c38372c391859f899057adb800f029f7a5de241204177b67ee0b7d238;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc9568bf462f21082d17672692210f96869dd59fc74442993fbeaf63aada6cf16dbf505f733caf70184f373113dbc9a014ccf80670deecd265d7f14108e209e54ae975375e96b65e0b2be29e651b2273c030f1185079444b99bd35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f2bc778946581708658bb2068fd76d66ea5688e4a3c65cd38ed8068f88f29004095aee511990fe38ca12f47d4b49d63fec471f311a525c169fae4d8b3040aabecb9025a689a11c661955b653069eb7a492a972019b2d4346c3b87;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0e4f9720839834b33bc922a0fe5e6349a5fdf1cd8e0f67b4ab09a033b021422dd3934e381edef44258fcd90cd65ab8974b4f379c008ff3c8ab52526e1d67d8efc3642851bf62006f6724ea2139aa89971d896334c617b8d85f99d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167947e90055e9f97ca9cfdbf53da5f806b49d1291546feaa9b6656cc2eaecf91a28c609eb9640aaafd2b39a3aa1bc9f7d2c3b92ccef091d3be9943e12e72ac12163e273dec142d74081d44054cc8801c8de71ec2e232d6ccae4088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b829718c5f9d3e765880b3181be2d6ad330242f515a2c3d1bc90ebd0725cf18c5355662a6de3eb2538870f000a3faa01f5867b0cb90508202022078fb0f03d21efe7ccaf0392e8f717001f08940b439d6cef15f3e3e46c70cc4d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13e3eb3e403a219e3a77b05c16a17d9dee5ed0535825e2685321d64d3342fec68b800c4e44d28e031fa0b5249c0ea6fe9bbdec4c46caa4be6324996ee78b075ad82bb61ac3bb4b6d311b22c1fbdd651df6ade5024811a5102c53fef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5095f671efd5e67dbdd851003aae34da2010204ddbd75791c034bc9d17f117975d62c360d26d62fe967b834cb7269c4e21ca6a4cf4865f5fe65b0a0f4bfe8365cea41662d986484b9a79a238216056f7dc1e14fe36b1c07c51f6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192bba46046b7cc3ced38f94d946150dbbd90c5a60ecbd42225b90a6ff57061755bdefe0d9728cef8b694fc326b8d4e6afff3942577a35ae30e0b5940f76c31a50615b06ed8d85de1bb7cef46e74a8f68a19e84524a800d6f43f80f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b7f02fdacfaca5f11808c8348baffaf1b892ae399f42e918ddd6266d76679cdda3cb28892af9ef1b16f645272d0a84bd91c8301fc978958d8390d4de8d460a722f62440f17440da9651c8dedce506d25e07af53e24b467f41b2d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f3836ea26e5fa1e2d4c4fc28935e921093aa66ad670f9f973fe5f6e5542dcd02f07f94a675a9b0e8844888421e41b791aea65dc77a3e7092168b0188db4c5c3b817fed23318002a6720f7dd5e261626433a5ea2e3ccc5d3c4cf3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e957faa8856f88063c220b223f0ccb62b03a2fa9eff84db2ec7eba939d20a803e52087a623a69d164d663c1a118919dc422572b7f5e3fc3641f34e5f0765318bfdb1eecabda3f0bec3e05ece220c40332683ade5e38b778799028;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e9f52425f6548702ad151492af6febd7b78aa10a8bc1c65d7cadbc3e2375614304671152e68bd6d9cc37e151e54da181029d24ce2e0b5b40e1d06587c4669cdd9d1caee286a3bff8745b243b34cdb0e3360d520efc6b954fa8a14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1066b9c03d84dd8da09308acb8332b9dc78983e79cce363f5dbf477f9143fc432d927bc2cbaee19a1f403b039d6edf64a3ba35e019d91a27b5fecc1a9254452cc80a72d7c926d68766b42bc1fd29a5424dce2678e5a04591024e2f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0430731df183270ad95e540fbd57e8ed9a560617e1d618c1c2e2669691892d1cd15d6bce5cf0d2214903cfa020823a9b2091687b3909f85b33b1038a50bb8a379c9ce9dbe61c983c7d08f8b40f436b62e8d9de0fd8fb708875fb5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb7a63b840fed792c1b390f5835ee361c15bb9ffab667d6c2b2c0dd10c3e0b0d48db26d55093fda3f278040cbd60a4e4c9ca89e6e44aa4528d193af0bdac580f996e8946f68c4d1604358312712f69734b8ff0fc20a487f3d98778;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80b2e393db23a8678112b9af2555a47885960bcde044caf8e5433856d307ac480143b2243e52a9f926a933ec307ab34ff74bf11e1f7911b1ed45514246f50e3d6708c0c7308cbc7b9db2c1f5898bfb42b6a7d8bfb2535b57128ea0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee8c6f4528b9297b7da6a4e4e534b49a02b9a474559e20d5cef731c4fc2bc15c8e136b0aad90cbcf3ac2fe073df50d5fa5f0ac81ac2cfe1d02fd809270dc040475d18898a263d14dca1453965233368ebdd425ca29be6555ac7524;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2d190f9f79a56c4c057b35d99929833773e4204bda9cf12a208bf9aecc8a1b11fa86ea8f8b1d6590164526c6a8016c296e8835fbd145661277eddaf624cf3cf5209af2872ed5f98f8d0d17fcb3e43a619590e860e199e7c87d4ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfb09d2a2cedc70051e5eec0773a4dbab34a4f0ae299da63a1f4a8a5f3b8c831379e0a3098eab5aaab4b34a87f7c040eca9e4c8e4ef4878abfb298c4d03681177f6bd2dbb4b048716590810a756053b541122b3822d911ed46747cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d4e884b78e821d1f0ba0f8a548258a05e5b5e6abd7f5df5f56da5a675b9fc79df7316780f2f173a4127d90fdc918ea3f18653ba8f1e09180687efbb62718f094b80002389f9b7fead5b14938032f01b297e5e073fb72e2b6b8518;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hced0962b759ccabebd5e55f62043c670c181a1d2fd355d65266a1507946925dd46e6423ed96c9324c2bd2ec52c509b433a76cf3ac652284653564000a0c113b4c168b54318ba97308f092375a24aca7f3bdc3a4823f06e273e169a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc5f306bed0f9dca72b0452537f88c47220e81f69d54fb48944df2c816b57771109286ed02c09babe5907c337898dc9f56fd1b99fe58a0dc6a0ae674a1266c3faddbcd9e5822356558f697aa9cd0b956f9ad858599c0c966b6879a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha57a0569acd12dfa14c7e28cf28508b4e9e9693e2e684ba43a4183ac3e7e43347013e4f0762565d80f3314dd6e41568f17c44a409812dfff0e5ca65cc688509af1a14909a2a4ad897550f7ac5bc4569010c4ca2b3dd145f6ab7e3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f69f057b8291c8d7b7a669899c4d154e0f42fcd3d740dd3d0fced11056cd9fc5144bf608af65c2c304c2503645ff3037ce8ae496758d3bb26ec52a75e07ffc11f0c88e2ed741f125a53889ed46fc77d398e098697a38718be1569;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5acd6bec82ac58d7016543082d55ac3cd1dc48a23b0ad7c9801b22ad7fd05ca2ca55cac085652dc979310aa1fb861aba50f7a8bb9429928ec08a512750cf3f55c01dc13baab67ce130d678a9bc6ecd0f5d38983b00fbfd5246f35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a64339c72c126fb46469a510eaf29bcab5f9fa411bf4b03fc61d40de9c9014923ff4548ad0aacdb1cbe075a021a8e8cf07213ef34e2c0a9defb8dd5a10408c901d95f07811bd302411308059470c759cca97fd05ec5fb001b729b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16367a127fd8e136a72486b19036ec963492ae73a9e4b89703e3cbf751660e73d561085c248342172d8d531d227d7a3b3254c00be0e317991dd1dd8498d7e4a7a966bb8a044e7a86a66e58594042dd5ccb96145ee4a540c70ab05a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1329a5295d0a0bafd091e5d2d774dd86388ea1e8a9eb90c2dfd0de06d85f6eec0e8150b48b75467cb866d9bc521b68c9afbc98b298dd73edeae921749c927407798e4eeb55c01d02f3cfdefd30fc9d9bf1c2d53f4c2b7296727368;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c4d3013db18e6ecf8c49390cde2104c308b169ce59bb7b856dec6da9e0680d214475f6f91cc557561226b5237b965ad81887e4799dbca2edc6cde66918f691b12279e74fffc7576df7d93c2d70684e0eda031900d32aa54635e0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b81f5af6008f7c4a5a1afa36405c903ef07ffca74bbaaac93a290781c804db213b9573651a9bb48e1b001596f968d5e11a6369bb01b14bb9090ca5375267b188a1ce5ed21f79e3316b31b57a372e98206da0f6e66a21f625e86c4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1652d3e3f50940e6fda20addcea986de826acdfebb575c9c252f3687480e5e0eab811dbe151d049b1e368f852bc625e9064b9251c00aa17d9f777090bb803267c156f178eaa1b51c08a824f164f866cc44ba73a8f3bc853708d5b25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d2444687c2e46b706b1c6da47b7b8d969b2a87b0b82d7d43786173ed37dee63a8bfc74f9ab9af0e7cf81e7f8a94d1483d6732514890ea64e5c8ad7a140be36b7a21013125367bac7512adf24a313aa6d6f333a71c6b9167979292;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9703756d93f5597c613a7676b6a89aa0379ff39707251dd28eed03d8e9235c04a64792238e8caade485af7883446f35c265e31eed65282322fb80aa842d645c6d05cc27b97b06da0a4ca9ad3b6655692f79891e997dab52b958049;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49f04da38c4515773b57422f9b2537b17fd440f70990709b1589639af0edb06ed344bdceee6c0eeb4fd42f135754208aa958271d5673dee19aada5583900732a42d94eadf2cf55b9c4958471471ea313ea7a11488e1c5fc38b4f9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf83b18e03b5e75f4a313cfe86f49744f8b8fd225d24315342556d891b256c9ff0cdfd41d0d9256996ba615552eca843cc6bb6bb251da41da8c023f14d1d36403b34ea6a42ef458362f1b92d36e787bafadb30b72f79cc40c52752c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176663c237ed04e8be59afc759ed5861fe455b9687bb27604c8416588a20b993cc4ee672a170f4b36544e8d75576c6034a59bf174f6bc8521df7903c5c2c752626cb42e3ff2223aa43008fafaf32878dd324fd1cf533b890618d97c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd344914ba1c2cbb7adf9347d96b839f9c0e56fb5aa1211838271af282b5ea8ee2d7e00d6942242b12354c67025e2c356c1078e60daa3436b1fbf5a0caef8ec5d2a2dff585887a96ae98716f44be9afcb2ea07717ac7ecb9b57cda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c196990c415f76aa3371596d66f01986788d654c00bfb399045d14704cb32d2a76b2e6b7392c129ccb631d1360116b43007e397d1e5accf1c9551059c9d90988c36591b1330f58d14577d0f4d3e59b56f5afb3bddfc7983633842;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haaeb9ab78878d676f07aa8950ec5b3db31779371862636d76cf70d8cf768a788fefee165c55f19f216a04ddba65afd1793371ab9845aef009387498df5f51d2b68444d828939e5a5dff0b66d4dcf324a33dedf0ccc68a2cf5e9c5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a2df42ccd8e1c119badf1c9cf661c5e2f03e364045d50762867616754a5a434907c8ef81ddd94386bf2759b72088713cb78fe5fd3e7892f426b759c38f11bd5f1c1a59ac628dc98a225ea905e30ba1a3c69665bc7f24408990a01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13619acfcee53f988474162cfb2d72ef6d5c546709fc6e72dc9d0b6a9526dbdac8e180cfbfdf64ce7ff6fc2651516c0d1a90e522162f9b05ca41d32d16b14cc8939ed8322a6a5d3744b67452ae110f78c649f1322474afb057de2c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc6fd0b0d2170e0216191d8fd5ac98adcf3c34341c8ef92e78d8cc95db0f2226aee40c16a4df355241665dc4ebb5925ed36a5062c805cbc84401ccaedcba9a429554f3436e80fd5adef628c043d470e0b0b542a4d7c2c7ae9c45428;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c98d108a6d7cb227485455a8f6b475ec7d156a6927853cf90d5dc929be2d57477f7661531182d03a000c9f81fb7cf59990c60d767ebc9e155f92f34714a7ca2dfb99052bdd8746d536f38f24c0a47faf85c34fa7ad387431c1e15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7b7536e6cfa80c36a3e1af831e538d2d2644fdeb6497a5528262db313afdf465fe112afaff0243b0b476f28860641c0611344cc124089d89a6de16d4693bcd7f9ce328283affa45c34c60fc86de87c890d1ab7efc4159d4a32a95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9f72582aba962a3f61e8dc1358d49924fb9d3d12d9d7a25ff80662478283a54329b29e05f28b60c794674b3afdd9f9cdc3cb2202ea7aa43930a714bac3838170fce7c541fa7c28f252ffdc379b11097152af8ab82bcd08d7b03a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10db1c28472d5e87525eed4f2306e7ecb86e7c3d04eb3fafc4b43f4e70966a94feeef2bb74058e050f7c7db61ee120b889ba1610bbe8ef44b50597cb3b163b82d0b96f1a25395d7f477d10e5317581c2f084632605b0f9da163253d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h112180313811ef97c3d8bd94e83a4051f74971010653dac2a5d156cb86441a45c0b944f231385091fcb94be92dd5a12c2214dbc3e2d18a44dc35ed4f62c153a6db007e55d513b23b626f10a263f6f1f0f5a0cd01f70267fc0e0916b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15537f9b673ce25445b061ad21d8e603db4c0a6b370b36eefdbd7754ceea612631882d737b02b895eb633225dfacbcb93d394288d6f27427571bb5555a4030f082b8fe6bcbf3a9c86c98ad41d5165c597b4baf9b0114c03cb7e5b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb996537eeedd884ca958773514c0a38e596b79c256c5a978f58c463bb0ad6f59b67a1ad3abfb8b7017d8e1dfcfb3d4924eb43897e376ea2b45cb36f5da63a051f4effc82555a724b4ecc39ec0c9e8f898956c2c6c24d77ff2de53b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fdfb88d0c588c58cf24fb7c240646e0413bf2b7ca6ffbe9ea7779bbac57249a5f832a25168c30cf04c006f707da7dc5e6f9ac86200ca19fb5ddd09fac0b72da1e9e1c3316b98c772931d080f220a654925dabd86d2ffc5e5736129;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2353316739d2f9c1f4503a023385b1e719a646e7f7f22567a7b90e335806466d20a4856acb3aee156dc95bd5f2c54f80c606a2a0b84d0a25910023d5e4bbfe144c814aad9c31fa109abd5bb3b4ec82c5be17d134e160812e83f42;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a88e47d77ef58e60bc3456bcd0659afef638b5b41e8f3f3630a712e44e4f44f50e5ab65e7830634ca582b47488cbc35c89c684e0bad000d7d25c1ee8424925f984a65073740a0927544cf4d0cdeba0a616a8e7415f15c717543cce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c45004c2e20a970609041a4d03603322e129ff5e12f9bc3bd5818e055f04e8f865018316aac5c3463683592ef1332e84388509c095e4e03cffbfd5a8ea86a5b3c1edcf3d5859944d2d6ab20e8113c2f0d13447a6ae04e6bec17dd7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he77f7c0ddfb2e2a66d9e9df8550f2e7aaa482306e07a3b0c7b85ed40acb5f33aabc43234aff9b43c5b1ae74bece397df502f044163d9fe1ff03241c1df754cc3e2f683ad7e0510089eeb3d553e5403993c600cb8859a701e949e3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd675c05eb63e59f4526a35553ed9da3b7e416ebb714ac091736c9754ad71a1c00c5e3c48421b6702b54ce760721da6c79835a5320b44141869778d911c584e7457e73924853924e47cbb65c36e6015f06471d91e8c5e00a277439f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e852164da92dcbaa215764762c4c2e236d092c3f04873e36fe283027ed0cdde3fa97c1374b2acd8661b5749ccc7214007a8e881193a43b4beb46732707cac887d4c2602db311840374b799bb99edff906bdd9a23cd37ce03158c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b62f79af71bdbbf6c3969f2f148b33158a6d2d4314c5f02d9c9e280b232a394e3e658c378a9548a24b2f3dca9ee4256123521643f86f3dbc24176f5063a14e203d22759240ca5befe5c5ec6fadc1fd2fce4f89937d000910e203a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b4a354a620f7c9dec0d779ee671a2c60eb879b532afc83ed1e0041156ebc4c36414bf8a0e9bd67e032d82143f620e337c0aef6ced3f6da4909c2a12ab0a7823cfbd7f266609dd351a20f618e0f2f549c6916944b78dc0b2da5872;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7b1fe0f8660c25755804da54f28756bcf9ff5a13748f175282726b7e2d8fb48b4e32ac6797cd47c0287260f9bc0b744e5cc6aac586d3d983a49b8eb9ef8b65cba811ebbbaeb7f809f67f6e1084e7d496a05f34da339bca0cacc59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9265caf9abf97db764e4a5d2efc6a7213f6d58443c4e9339eb773d6445d61cfbf2678712aeb2b2a704bddb9ececd3f4f8c39f9e7126e8abfc712797448247b39e2975b90d7cecacab50968e25e6d1073c927a32f9609c69fa63316;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb477b804a3fac17506c071a0a6aa8d6cec87f530b82b0b5517f59b3bed2824f8d862f5712d9ff979076b2ccdbc25d6f7639dc57b950f99c11a6c5396a0678f317cae41b774905018054a0f6fd5226346e4366be93be35125461920;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15cba0f635376c9a167b1650109f1323904f02eaa009d85aac891faab2e978d960b72714f056c23a83bb6de483d46251985ed53d741cc7e5f03bfc43b817e2bbc1b6b50ba5b06b9d8e5acd75f103ee5fd1c561f18ef38f41cd41769;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11de2b3854e56de561ef2945139f52c92caf19049d3e80b9456d9d059f637067c5bd0203c8f31cd83ccf0703b20f0230e4e3afcd8a5ba5e318ac6aae949917714076e476b926762b65165b0cdc7abb93891fa0a42d3775510626aea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c94afb2efa95978e0e1de5c2849ab8c5eb25509261977a69cc8dc0f2aa1b5248e7004aaab6e5f804dde8e9f82a506f7973b2debcab766184a310e9cee46711c44cdd959feb5873042e7e6126a51dd2c2dbfe20b03addd4954b3c53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd0e4950f86e4bcb93c2f0600df05d330bf8e4fadf345873c77a0baa75478ac8246931c8301e69c6c502eb1ea05845b1b8a588f4c2920ba834e3cc383b719b5761ea4335ffaa14e31bc74423c5e9f6d167bcf31ceb5f4cd4c14666f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1619c1d577edb3febb4dc4beffd6982dcef695fefbe6a3b7c17703bc407623a1f6ca2dd0ca6b8e770060dbb8c5583dd9fae05d6782bd54b1046cf123311cdfb41aa3386c497167083d8b474d7607ab2e02455d58682f9ca2c494152;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f57e6b1c324ea954b04592fa08b19f6545d43f2701d5ad3872f846761c2642519b7123bc602e87dce106939aac7c88d1a1dbd93f0060d97a3f41545a1d0a0edb54a3a2465efc01faf064278ca849d0e0a13110d72c5b7dfb373168;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3951022e73eccd2db88dff4152200fb2addb5e36b578ae50cc304b5f1e4d15edab3596909577401b92dc54317f6ae0519d00751673c15eddd82036b30487221d76a3ba1b2a04ea676cb30303c63256762d6adce1be5dec1c38137e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114ba01e7ae5aebe4c5b85eaf2da671dc1373134995fd31a3c195225ccc30ee7db910423969be31f23c551ab6982d100e1704e2d08f844cb7beaf5e261bb63b852bbf75fa9c08cb77a83420a8c63a41712c5c7ec10213d379036309;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hecd741baf0573edd74935723dc0df69a1f6ce2eba2915d3503598bf2aaea6a860462966eb13390ba07f68b5772257d4984c1953d70315854ff61c0628ce4476334ed2c3339255577fffbb8b7c23da0fecaab297cd43864cba078b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1234a6dda2a47a9e3152637dd2d135b25901df618b63312934e467ffcb87af900cd0ccd09c95ee95aacf3258ba5b2446942773d234d7f3116fec13a2a599a096f22a283fff9a66af20fef2d7af8318fad57fd7b2ada4e885b0a3601;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1343dc8eff6ae0f11c35a1a23e424296d7f2c931be049bee2b36c218661188432461a62091a86188b116082dafb3ffa41cc62505dbde784f9f2d0a17532ce269c38c9bcd4ac0e704391215e4e75c401cf794025b99af1356ce88d61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h124a03051fed94e003e11981567527b9812818ffe10324bba486f072c5aa2aded52f867226a6048e6c56792411d1a239ca6f64cfea25461336b0a0d8cd3ab203a426e8ae1095a5b3db9f813579f277be992b13c1f02918fec80b9e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc15390d627b291e362646a78ff0d7e5a68b1615dc9e59ca817310957d976d8ce05cb66637e4fe6c4773eceed53f4c9a9bcc9620c0e184d86971b4b7560c3ab974699a20e8491d9b990f86f44d0346ab19565ffe4b00ec5ed3a57f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb61a2dbe0e91bc3d847ea769b4cacddea9a280001827582e6773688c13791e1729b4dd69fc4a9e58e37fe0e8b2bc061e72821476f315c6043d584cf4f11c5fe850fe16ded5000eb05b5491f7d417c0788f9bb5f25ef298c16d7309;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d55a34f8f84a45ed8726876d2844d500dc277144142935faa6ccf03b2c27b24d667e047138c1bb81fddd3c709dcc22c592ae5998d4ddac4997603e2f580f6cf99b253ea7029d3c8d28f7e8871eeac3db112899242ce7319af2d543;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1879decf91021bf32924664b3be72aa691897a3b0fa4e5b44c18df63f79b5c25239dfbf80b342caa4b7c0a650df2069e7e0488223163639f114f8b4a3e98ecba0373de81111bbadffd3da35110581b0d17a13280840b7558ebef432;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa6b1339fda6069d05104d95b92e91cd46914298195becccbdce1651ae15179031940b5d15e42c2639100bcd770b95f02d01bdd5c502c9815a1b58c284be87a691ef7f208d27d989ea59f9170c5b204649ad3b284943e3922e5110;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c02b889f237b40f0d290c8f841ca888db405b6b6220d131c326715702e4271c0f0ae81e6d77fe6f565348711d921e33b4847f34497c21d7033925461ebc3c6d4ed12d906dc00c646f40e77c6eeb12e1190a2b8af6e57aedb03d6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb28bfe03491a6483beb3317bb1d1ac5bb6a43c7d73c076368810f75541674307c853bf89c2c1a04f1c1528ed9db0b63661524178fa0b6df6e5a61fedb9328dd60a600487d1f713c65484d18bfbc8bbe3c2e53d7264d1f4ce70b9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa12ee47c41e8ce2b893dcfb6a5294fde5fbf713f357d55bdcf2cc26cc81edfab51d90781ce917d4f301a9c5c828a2a8c8c63db5e81c89673ab36aeafd42d56f299113c78130cbd525885abf184822d7019c115c67a90982301da6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37e5e470713ea6c2dafea3944fbead694526497d4404d576bada632d18961b9c7ce632eb601d159e15c1fb19ca64f48462c3933efaa37e12eccd7032c8876f2430e4a9d3c090adf6e86aa06413b5209f41baaf18460eea8e3e4cc4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe445abd686fb56004b12a39502649c7bdd7e8d8525de2ceae2daa9804ec868f189cddb22b5d33badd1d2a6e6e52db29276c0e354d2f36b8c2721cdb464fb8cde790d0faa41ac9581d0c1874dcb808179fb8b134af3195ee68964f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11051e815f93e5e41dde8753a949426ecb92d9a38b574a5bb6c683d35427523d8d356900a07e283a4609cbef2f1c822d8597a700073eac0f643e55044f594db4f963166d449e70e18fcc6a4dac339648e36db5a8266955391245558;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h198115d2eac906f6f46d66966171cdd6d43718370c2d703be3d4fc08d30eb69e069ad0b59661125afa0c4e1cf26ead16fa75ad8790d0bf0f8ba0866a6e7e0b73a498a80c59e062d28ca849be43a5a1e1754adea29c5ce0c4641e3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe13a768111387eceef826c1e1efc9955e8073dd5d56ea5e09f844afb4371210a297804a978858b6df4c116d27f898e23a5d622194bdc5e4027b5db920ff10945960f62aa58208fd40131b16a51f549a33d28d79a39c1f4fd6ab80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9b0cf1449c9336694844733a73dfa69708df842a2b8f462d2f5f0bf3126f2a4101823a445e374238afe779c40cf647b47df6448b0bf864924f67b525b285a9225ab1cf5335fc86e57603cc492ccab59a9ba2190cccc73322b50fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h42ac95ffea965da65c06572cb8374131fc8efdae9a99774b31e170b814f7641904086005038d1887b99e77bfcb76629534dee1963d2b801305d18f3ffbef217f2c0e888f86073905c5f8aee06b463164b59d10f0e301b9af0bd024;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b11502bd106ca2c97d3472be646a34366ee0b028e141ef671756bc7f38c94dc8f0da21683cf7517065232f9274e95b264792195cf6539c67c9ee67e5813642a8f2266269174e87ec19448463f0cf8533c066fe4d3740c16624ce69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d715b886acacd96df1be1069541cbc03619d994f22b60d99223443ca011a68202386543dc7e743792a20cb0b17876cd5d36afd8e1c6c2059c13742bd773708cdf370a026cf6ad464ea9c7d485fb6d77109dc9b3d31a6ccc6323dc9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h94bc9ab26c5779eab96ba28ff9ee9bd31dba8053b84a501547d2d55eedc0073bfab6f12a2b4c11f896b176afa9d44a62ffdb62112f5431b800dd25ac46c0b1192572f097a865b049146972a2a5af2c529047b47f5dc13b04eff0d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1965148fae2fd6381fd465c0f4d2b45c20447cbcf9001f73e60a01cb20ecf906ac269801b4808c78d6367980acd57f2dc7419c710e0df23386a9e45799e9c36c2b3b62140d9d7f23631f4f6f962b825767da81a74a9038aab887ba8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d268f05d477d5d0668af6b6ba14056b78f9c894b3d8d738a758135fca1095dd0969ed5663e96e78d6d29aeaceca10b94054b4c6a8ee7af2a9833ed2bbad95b44b6733e0dc4daff2703782bfae654168a0ee5088e004a7efabd950;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h66b06b025f8eb0a881e5a29de7814ec44a05ea3d75bb2ab338662f01672e5b180d6c4c57e3ab02f406f481bdaca5df15576507e95557e78fe26547c59e92412d4cfbe45a79ae09b85d656d070847ff9000e124357a103ace6164b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137a1f043752a3606c7f7d8001ae831ccec9a911343b68d13071e5f7220a6976d6c11735a61aeeda2b61654705e4113b8896070b6d2d8e9f703866d502ff91c65da82b7c3e5cd9ab0eadfd7ab3a9f9ce8e54d0ec0ac709eadd92174;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127f3b800e7e9d169285856fcdb6a2f49278a81cd62ec0df412b7ba838c79e2fe307fbb2816670e79fe163c765485459ad20674433512e962e89a483f32d19c851ea22bf006acd30ef99988d34c20ea5ebb7d70864c5e53dbff5d84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12967bd11a88d486c4b77869b8c4a3610f9e73683289c86cb3118049a0ff5ed384c1a5e9323b5d65f2ec42124d476cb4c93a618bd97225cc4b31ce9b50fb321b08e6d85176d97015a47e6300e1a69f59a5702c5a8e0f5ef7e9758ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4e4030bd5bb007c7720f877a8892587d01e2f5bd0859e6465027be0d87a9bca50821e78a24ccd2454d9221e75db1f99596f4cc7668de2ec66406e11fe61d43320bb56b52b3584772a790ee4cfbda6d8a21a185be302cf5ccc257d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c43076363691d65a4dcc573a028968e102bc0daa33fdcdeb16506c011018bdbf35bd8223fe7c6ab449a6c4f409e0680f05fe1d1a2c1440fa853ae2c98722dfd30a15265001a88acb88701e3ffe1fa55ba19cadfe4ba6e73f85bae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbbbc1844b10a7c777eb39ddb12ba051244aaed25723c2e9f0477b48005267e1e2c30ccdc17d939202be2dd107360c04b57a2e5d633f9ab8bc7438bc0b36f6b9f99429de50b6230bd503c00cbb28f80159dd9fe52a02a05c4c5f489;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18dbb75d4a3526af27f575cf4003cc99df53da5767e91c41e71f1a362a286f296997f7b284b49064774cf2db4c8b1b8ed9e0539fc19fb765f69f13f5987e2937429ae314719b943a9af43385e889466e976160b8bd36e031074affa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8732895d0e46bd3b5948aa6e7b6d78d78c249390b93aa14d26904771a420a5136740b18e1de8cbc06ed93ae38deff6d0fc8f5cdab17cbbee0611379751fa76dbc3173add787240194d9f59f77a19363602302db3a089d3904a600;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c03b79f27567554cc35268e7f945a38132eacaaaa01fe39246a3f543f2f29daf45daed5e5cb0e7d66f820316fec7f715466d349a00b7a934d281efbb1661c5587a13e03b48db09c22c1d596b5988319d78814f0756c7c05e689d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3405d10f22e22d4ded2a3662907b47a035bf98f4db0421781964815cdc231c078693dd76ea42df883930993b22f3c92917f1198e79a2d432918a66ff79a944fe29ca08bd1bbe3606e899c10aa07749ba909464a191d7340bf5da1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha26f0dfd08f03262be1cd2a3473e56b87a09603000fb42d5af0b29ec902179a139fe035402a35b74f02d6b0cd383c3b1d40774b1c2f8038402a4b30322d1d6a76995356538ef7f2add8ae9a280e7a301c0cc4fb5d75814634d7ef9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he3e72238e9261e1ad3f731611fea2bebe42854a85412c563c0cf581a3487238449235137463c100ee399fa2e1eb358559ff72251ce1a60498c1b65ba97f84ecc6162c8ce88f747f99ed8af2555b2c498fcf5f6b1e2a35f7cce07e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa8ec99917d76b232e6339fcdff210436855e6a1e365f2332db19c040016b271c1c56a5227ece469b30684433bf3981235407e341cd0ae329ba0c619ef4131061a20dc74371a3ee5cfcda8ff1f4f0696d33657ae5a21733251bbab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19cd029187f94e2c595e4aab341b207c3d45c86709a5448793c34127128d2923ad64574687046f85f619deb37fd2a74d0c899b848f796930ca2d8ed484c6d4cad722d71ab77986e4f80a025371a8bb9319c6d0b0105429bffe9073e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d913d5bc100316fed3429adbdf3122492e0548c8454040885fdc215fb5d358b17f876840792ea9a60ac39b00f76208a3720a0725e7d33448faeb0e05b9d57e1273f4890d37326ce86e7f35dcbf685fac8b8936bc7084c9c864cf5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a7e3dcdd92a629cc5249d82a2efe77a855ad170f07cc7e53b752ac0f96ebbb71ae576de9eb6ad330653fc09ee765d777b691f1ff7bb60722a99f40f328b2c552a1eeb3e1324219fa01ceeb5308f2d3da8c63edd60421a3264edbb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3833dcd12f78a9f44ad28adcba3d5df54d53c0024d11575296c377d45af2c1b4b7e419ad28a2248b740b4c15548b5c18fabc62cbc8fb0ba049b35ed9e1b47f240eebd6ef6fcf47726d18e9c16d368edb3ac902e68f98c72573eaad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a3446a170824320bbbc3a18effb61e01206c47f3672ae2470d04735e985c149ce39769682abf634d2542b3c5393a1af10990005e93410db305879b657916610ba8a9bb940e812457327da4b40c12593b8d91ad210fd3d42978dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e8956bcf1c3ed7462d6b756e617553291f1b101190c9c8f6fa9729b04045e7d1b624d802fec2b36ce6c10c29b9571d92d92b8807b150030445fc857f94a5c926dfca344f90a7b65df00cdb745dbda8e303a876ce55eceb6744f54;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b79f2641c5bc01f21848040e191a80486613fd19ea56dc006786a8552a8640bc566683553798ade86ffa71c7e68638e1cef3e7e32340c3becaccc8362fcc737fb332fd9dd5257c32bc20b4281c19d45c4c12926d6fa9d50a85b835;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3fb04dbf4ca94e73e0622fe8ae41ac5608f9a34c13059ccf0f8b3c4005285523104f7713cb7daadf2df22fcd8557859bd921353d903b1ec6e048b996be23047ddd4cd9b71f060832f6e7e8599f252ddb518929e9372e5278aa3270;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c1b02c81f0554cba2c4524bef4971de6d9cce9b7402f71764d086c9bda17e2c57542ace10a674a64b90de0bd3d3e2e0e9470624a3c68cdba9b1c3897c9962dbbfb7fe8b64b2dd9c711537b8eaffc8bd8a3157ff7bc8fa09810750;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff610f42f7a3d2ae93a4ab7245eb8647ebbb4b2e10e8e221ea3571c1d6949336d0e9f3225e8044f012b2088b304c2679fa997824a47a67735e8181bb0df01e1fb191af264c7987cb216fa022c62b736608c15f5ffc86806ce818a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f70c285570fa80f33415f4f65564163d825eca848dc899c2574dccc0b035c59e46f530dd61abb6f0856c3eb954115efe59c3a95bb8887a76c06b6b01c10c5c9dac70e111d40f237ab781c50393495002398f2856c3942daddda25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1184d158f70c3ba97e116327e984548580e0a9c42a69a374a7426387f4a4314d18a5b3cfae26cc9ad590b4e2605ba456e85808e7bb259826dbb1dcf55b7b4075b760ee7e0451a42034894c4bbc886559fe5f2d612bdd68e95e7a32a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfb4c9919b284b8bdf2d2ea059f1addfcb6a7612b63a71fab07b935f0fbf45057eaa7f4bd00d4010bec15b7edcf9d72532f90943f85d6b65bc4a08a5325cc382b12e39051d41383e61698f1f6d1ea7f834dfcd18b641b0d284d8eb3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f386fcb628d8ede51c45d906de68826b240b2cc39f751e15fa013b0b2ef387b8f282b0e5eff926e790f7dae1045d918fb3bfaad7b4398a5648f82230e809fbd6e77877794f8e6059565d61e8cd3f31fa5d125fb4628247bfe9d9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2b59beaab1ee5906827a8c2fec3e369e2fa9e7b0ec1e6579a6c1af5a3274007fdde698e16eeb4fc7da21a70e9be18bc310cf53f77ce2ade1a6dfa40182b2530024298b04c4bb451dc73096e07aa4890e6b319953efb8bd160419f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h42d0f8baa31f2809103dace4dd98cfb043dc2372036fa66591c52eefe328024a8f53f7a4ec2cb9a6a518a71857c101a3a588d1ebd8ed55745d2acd9084fb57ab15435116a8de89b7fe6998d539f262e5f7af5a7e11dc18af370b68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1251399e752c1fb51912da9d1538550021fb03c2b4f79c22e394d78c57f0607768b23651fb5a6000627b044f47e2fd85a4c0e0a218975dbd524874bd2afc89fa07ccd7c0df207a235fc3f4f4a2c7fd212cc6d0c67c6d86d59ebdb49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17835baf80fdac69584352b1b7f063a43232db173599481031477fc4f88f2e6477e778af7824a88a16d371b9a006071c6d50c6cb24b6336d3e6538e60c22e36667dcf593f56df348d0d0d25eb1e1ccdbfb30b98fbd38c4ad54e88da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4cd9a42fa9c7b4a0cd74e0a0d2e90fa03b8ab40d60ada2644e77096b3a40b96f328a9b64068cb9cc521876f54064896a5d083db61aa5ec2ce7876eb7cfa97c2e44da64b12b3187bbfa9fb99b6b8f2a95845abcbb5b97ddc6a35774;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3237eefcdb1eb9fa05bd117ae09feb43b25d21309610f64cb2bcad0be1d97dc39aa5f5aca92f34187815ee9c4818f58395ec78fa99c44d2f84b8f64d6f0b06c702e7584d3293663de6532f0451596235d5c755056221f0a0a1fd0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf8913d51464eef4ea4bd7921d36dde075bac16829d5c0db7fb25883fddbce726d36200693b39c98d1d2ff28e663fa71fda9577c3d6999bbad150be60ece7ee183f2ae2e996e6ad09dfd332a6e21881043ff346af3a907d2ae3425;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbddaa16f823cb720a4c95278a3ddfac4bbca8e657fc5d530aed100f02b0447dd9714cb44967f62f539669ad17d4db708e39b1c1a24d7444bcdb1cd8e9f5cd1333d909ca3595c6f999af7f67dfbff580e1aa054a57d46072ed62036;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12cbe4a0cbc7f6b134cd3b6a8935701fd1711ad3cfa4fe6b7cc47e5b6a47c91c92ff4eaee58b5f3be70c0802a2e39e3b08f8f22b360955fcaa3a70d6d3d943ff0ce611204603f37ae2794b30dcd994d1b14afec5f2b6248cdc4fec6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e3c7efeca162d9eba0fdee00e9505e7bbb9ebf33ecd5b0b407bf1e73f0887cf01eb359dd169d91a2ce922e3b921b8ac05e19a19dbb2d1f1c2d0ea4edb5efa50cc29c6f09a58e5a61011270eca64b25bfa60d1d20b909dc07ff2ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12dc78aba7923ab229ebfd6f2e870cb56c523cd20ffdc6eee3ab0371c63bf278d9d5505b23d66440837923efeca391b06fcd25be8dd6e85d0b6dee825d01d627ac12c4f8d5848b9384033ae635a0bc5b26ed3f7b10ab316a0c16717;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a40df0fff74ab8f487df2c287b07576c353744d971d09d96e331703f661908ba76085c0f4ccf8df963e4a87bf8586b0e0e09ddfc726adde122fc6d9f91f1d2b55cd965f14385c7954cbf24e10be91ce5d98c36b4c3230bf0ed25a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb2b8118b6cc912a1bf3cc00e07882db93aa215c39e9a6fa3a2a8d9d95a9d5f674a56173754df0b80a0cf2f399445ec07de749b9d3f53fc2a425dd0ae4f5af4b939dc7e3f5ecd884d13c05564beb003b0513de023ece550c4bfeb29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a5f50c3955236cfd5ab093ac02405eb9bba08328c5669e93b337e6e989d603c7409056428b2e41e8900f249ef8f27f26a09407604dc7c95e8e5e7fb3c32d476c7b604bfdb2edeb3fa53731ff9a7da8fd71a5aca5f57b69c471d58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hadbd1fd4b67222ad176708872bae8a4e98f8dd41a7cb9ddd35fc5fccc50bea0116a2e8be43b39133d0a5b094e2621a002fa62b67b6c57d2f45cbb3c4ab46597680b3cf82d9bc013e60d02b9715d1cb51d097e3a592f7bbeeb24847;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5dce69bde6e10e326f5806411e0e9675f3664606ae68de3e507bd1810cf80e5a8a916e84e8f450b353bf3b99a1f614a147b84cffedef0412d6faf35c7602445e3ee5ad902bbb65af891008653a8ff448587ce686cf2c501bfe8e52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa07b8eb57db647ce7c51cff196290499bb9b8825eb0544b10cc794045cae053c87531373d37f7a4accf02866b1d804c9e502cb1207540627f6d67491603aada73d70c038a481500d81902a3a643eecd579b18c48749e30ab42746;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7260a1701bf47204877f4b8000f6565172885f6d62b359756165050a567a998c20975e158a0cb13f5532f5b5995d4f940d321a583c0921b34a08227a8058d1f937e80f6256fe726c23bb5948689d6bb1f9ccae30c6e914965601;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9996316db2370593363e7ca3bc7ed41de7aa8865748b208ba7931d18ad010d3e90c56c41c6200966e3276f00a1bf406775354a52603dcc912b7d33cc1d4d422f8236955e3b05687f36a89f8bb2b6c47d0271568083d9cffe2c0111;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a97827aa2c65f46fda692bb29d638fba0c3fbc1c3daf9598003686902490af50f462f6256193df6021930dc63ccbab929dc3dac990366f264809e56ff524b1c2ff69eb4abe3ac6f523fa04749b1e1564b77d98e8bcce1cbb3f822;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3882d69726a94eeb99ce41025657d36bef8ab5bf1cb5c3cda4ae5074ff24e90a3721e0fb15bcb05556944d9251475fd16829391e0f1ce20f26ce4c01ab4fcc7816a47ab77f70e57d78c91b2e1194197cc31e717ba30bbf526cbdc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2793cfab28e026b51b8a0fb8c12e2f916c6d58e031e7670fe1e29c2e49fa00bf062b9370155d6df34ea5b317579274b9730077b6c1da4bf92019ac277ede9a2302264df275701a6b92fe8aee9973c6aeb86708e49e8ac20992df9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157ffb43a31f00f895fcd9d148760496238f60677432022c57434cce4368b4511dbab389a1dd138ce0c9b87d6bf792b8fa252171064379a8be051cb42a4047367e8a791803c2ea148795897a06afe5dce5f4cf58eeae17cef899994;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6242827dc61a072838d6f259d0a8c8a9e4d43e59193bb233926da609891a81576eda723df11fb3898fdddd07457d67f96d4abce927e67af660cd0cf44c65abd8ca9c4b5b318f3ab1d77bd384c41cb54b8a85b8359e4ab34e18fd01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c154ecc54649d68fef7e0a6f3544ed45dbe7514dc3fdcccb67eb9b04df9b113d4e4aad052a7ba44c248f86bd5a718791e5b5b6e26469b0a1e7992417253eda22842b4da8cd7d21d3133094364d5a85a1f91a6877064552a25523ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ac422a5650086d7ee40a16a6f9f482eeefb6c9dc3b2fa2c8ceb0a5180ce35c8e2f5c8bebd19113b238e4fb2c94f70548d11105f53217b2f2cd0c3431d8ae11331913750bfd7a7b4dd7156ec9da5e6543f4ed8b2a47ff54c5f0a38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b1e382eea593d9a2cf8bc0d0f1cdc2e4e6a78b554b4b1840582f610f4c56d0a50b7f45c82954d993f8ea3bfd950a9e1236367af7e8bbeaeca1725bfeb8090aaba2feed49f7f9b5321c33b98f9cb12d8e2cd5c70fb54c9ce5201a11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed282f4e5c1f303bae5d800d4d53ddb7e301a453cc3bf87d5e4b2490ef12b6eb03a0972c537cc51ba116dc101183c013d6e7f9afe46b279afa2d91aaa42bb55cb6e0596ed64e06ec8f3e4ec71bf30d2f0df42d4df3b1171e7ccd3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1854ac35fa5425149b18157eba1ab8301f727de1b21bda8f0bc69a04b7bb7547409f10884649e434cbbc42f1425d22f77b1b511a9fe756b8fccbb0e649adb9bae1ba0258abffc9c3ba4efc13cf1aab760e3e15c3a4e867d2722b42b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116f9dcc0bb9058828a3d8752f8f90d386be36dbc159010b14c7fb3e2e80d92e87c14ccd70f26378b7f82be85a22a023c534add839ac12fac36ecc6e8b054af54559b9019535d161537036dc6c38b6753e5659aeba4ab73e0de172;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d06899d36fb38edee9516fd64c7df7ca5bc48e79062fca2b9a2df8cf0d1cfda6f4d9ee5b6a99a6f8e429efae5afc8f987ed58d03217c4bd4856b8e1c893c8759b168376cd5186ef4e51cd2dcf9d8f460d243390d9abc64d391281;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4dad01d367bb51a5961075e2cad3b06aa579f25cb71b529dec93573d7d975cc4e94fa145e8b14b63e6d31e63338e55e363a4ec2bf154819743fb98cd1bf1b686e8cd6696fc026e2ff8103de79e2b7dbda538066d0a166dc73ea1da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fc910332663a8b43b7d6fe022953c25021f4842f8863a094974c7ca7dcd3b10fa023a1e6a8c4c6026189b9ffe1bf49513917671e740523a181d442c84b3ff9298b6b5506d4619f36709b53714930aa54e60ef38f03719878517d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184702c9ae273c172476ebba66f7571d2181e89154025219722af097dadb78c649141aa9e77e4766289281bfeec7f41924cca3ebe3073fc81c6071f4ca6dfd23a15023fb1050a9c95c9bd9486d0330b02701801a68f72a27f47b045;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc37dd9c741548405c487106b02fedb0cb14d76b2c4b8f153642d39093822942c328739e865f46aa767350a6a4b9ad1c633b1ba0adde552a73be523d781e2cbf539c9c6d20d668ef2d8304e67b4b6e047b66fa71aa98868bc738fa8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8974262847d3225d9f570013c42e71ca6585c543bbe439a8754c23eeacf521205fe34f3a677069dae7d4e3c5ae5dbe8703e6a7d9016248f97c0cc2946b873da0b6c65ef0b8aeb4a3e79e18a3b2c7f3d98eab89c00f9c7dfe89a15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9fb404f16d7e74c6fdfe2c0df7262527a435bb826712ae274982f9dbaad41db5c16fdf8e6a88c818667d773f2b21fdbcbf6428095163960752bbab9d472e7e0e5b3c82c4ea453883f0aae3dc2438a29ec9c103f86ecd68c0fc67fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2d0460023d399fc935e5835ab7ec0e86626505525657d1cc46a148bf6f7b98f0daff7f4100e6ad959cb6a5924e49aea5ccfffa4570956fc221b2df2068e625dffec060f97874e0cee26fa5f54abeaa755c2bf43260ff915ad9ca7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb5587d5e1a38f58db0cd457bb20fb38656c68db4e087831875fe8fdff61be730796234c118f3dc4b50b7e15607a2b143783d3908e9b5689ba8c3fc137c1f19336e08a5a413c80a93301dd4693e8defa4090507744e269e96d6bdd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff68f191ac3e7f33e49db1fd92dc77909f44edd88a569b2446d27744a72f5c7b14739e4729c0a72c5e71814e28cb2efa91a3c9d925844a9abce4a06cf3464410f4d905b30797429549df363d5939cb0fc45d6ce9e452eef8d6de78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc1f7cfb0e4a95cde9cae4b8073e8dfca0330af10b655d286a6e5fe73d02d7c41507ea9b9232fd697865a1bcedfe0f3647e88d27a489febb060598eaa830bdab85d4a2262532e9c3137471dc29775372e9d4d70636344d25125f9c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1776a7a80d4e4b72583d3e82a805c7f6bf89840f9be8d670c243e026b3c523a83f31d2272f3566e2c5069ed811eafa10b0b2ed78482e1fe6d803c0a38fd5997a4ed646c5d858537467776315a0c39db31526f2c63c66d66de8250a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fee03817980849df4eb0b820614b367d6d09c548d9102ea7909136f31132c97726b77ed0957b5129c22aa7cd9e5ef444ac126c51a781ce1d1cd2e95a901654efa6a4263320734fc420c9bab4fb24b9b1ea61e9ada9e20fa98a9ce8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h71fc35777cf35405a72b747e6dd9181e75b290c2ca351b2db9a67a8b936004d1ace07fbeb570b29e252bed93df24c49e60d121f5ff066456cfd9fb3bed39a2e8afae04e283850ebbffc165c3ca282f20dd64fc10fbcdf84e2ae40a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f36fb608a342ec80d32fe377c8ab973b852427111d5780418c746b828e7be80de44dc2cf8b47ed645c116d249d82080ddbdc71b82f8ae5641acce1833fefcb37e27a2be90a3dae9edb525ab305c1e78b8aa9ab7338f81027304e2;
        #1
        $finish();
    end
endmodule
