module testbench();
    reg [26:0] src0;
    reg [26:0] src1;
    reg [26:0] src2;
    reg [26:0] src3;
    reg [26:0] src4;
    reg [26:0] src5;
    reg [26:0] src6;
    reg [26:0] src7;
    reg [26:0] src8;
    reg [26:0] src9;
    reg [26:0] src10;
    reg [26:0] src11;
    reg [26:0] src12;
    reg [26:0] src13;
    reg [26:0] src14;
    reg [26:0] src15;
    reg [26:0] src16;
    reg [26:0] src17;
    reg [26:0] src18;
    reg [26:0] src19;
    reg [26:0] src20;
    reg [26:0] src21;
    reg [26:0] src22;
    reg [26:0] src23;
    reg [26:0] src24;
    reg [26:0] src25;
    reg [26:0] src26;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [31:0] srcsum;
    wire [31:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d153a6a4c6ded75843cc0285114db85745b7b647a26e4e59c8ee2b35eb56a7f788a7fd06f24e3050525ecf6cea08361667c2ab9c4395874e592c3e4e68897666f61be4cc470923a1be209f7c72c908bb660e726388e1955ebb1bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11baa743006d3c38cc60653a34a3476b73ae0913ef60423fcfdf7265b32bca562891b8a40de4be83a8776c946101be12c2379fc0f8ba496911a0b42b0779fa81d9abaa72448ea2c09330f22a9f080fa7cae42dd198ff9199b2ab55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193ee063578d781143204a9e7041199796aa4b9c8955374a1c59196ce9265d6e710feb4ca2f01b4ebab27fdca6eb5cdb1c88dd00e288e9fd8c3546843888fca1f275838dbdaf015951d14b5134c5d28a5c71add91d6c51e04470822;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5cabd8e99cf20c5dec6127a694fd8c90dd28096d3669c7d8b57283a41c47fd57a6a72257a16072cb1ac76d6517bc79272e2d48534c1cbd127691e8e61bea87e6161bd72f1c7bdef3d6d3a254c5604aefa2712bb30eca9fe2e3680;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18cd24b5d85187dc7d7879eb23314f0ae6325101bdb4d4497beb8ceb2df0d705268247b62c63ea92be13bb3a1a30e80e3057dd339cd039c66da78b9140dcc0bdbfae7b41d432bbee3771f1d1d2ce4e817e0e677fcca50868bc8a085;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h887815e92fc2fad7528557f3e332be7964c8bd75d638200e7bd50d3e87393b6bdf83c774b9f7ce9108713c199ba49402980361a50c57acf284efc2ace013cb03d604b401b874ac2a375349067932d58dee2b0cfc11d9c72e6caa9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h666ca285395f78e307e641315248d9bbace057c54500acff951f656c1f94f3cc6a2a2cdcb805343837060bfab57c1a42a9344812c519b68ce907194378f81380855a477165d3695c036a6437bb859110938872a45fdb429af806ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b7727aee118d13b6b164ffaee376770fe8f34bc3cebc7aba01a94e996fdd5c3715848a7a50ab63f886b438c74a65606bc9db8e9cfa15207b252d9ab936724dddd7408d4fcf391d572e85ffdd3003315f20e01d5b1f511becdc004;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93c3595f0b8db0d465c9fae060133ba26efd55801921ed7c04d3ce994b4dfc3a5260759d40c799b80d8aaed13569bba7957c572b34cf154f57ebfd1683ae6d23ceda0096086d0e29816c91f953b2229e882394aa3fd6c9d7236dd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24e9bdfd55b0418efe02329ce3f53480cb26d19e73d86541710aaec1d2d90636957a9d41d9fc2812620e3f5ea2085d27781639285274e73858e89ee6f36efeecc275d909dda03afe88dfce91e79e9e2c66882a14727de906606daf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h61cb9753164b50c54ccaf7803247912c6bbe0ca40208c6a9b03b6bb8e1349eec235ae6e59ef66683cd3b6409e0d87eae1775995a2025a7e9dd18cb240fb504873817a7455423732e957248012364ea83d49b8267723e7da77b76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0147d5bff8209f5894d02eeffacffe583560a2a8dc89accf0ae824aeeceb387ca58f72acb587152c6417dad61e163f0ae90bb80f6d1f09cc3cbae60ef32668c2fbae8905e4f8920195c5de81f8eccd9ecd74cd725b0275e91cb67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30974e0a127d33cf550960a20beb1099756cab5df5ba532d15ee2db4a5589841b003070971cfa47c9468e4cfb3fca5797527fa1bc050f31a351b9b8a57d69cc83d6bca11ce50afe4d7a121c8993675922fadf6d53b9687bc308a14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa5f6978ba91e43564152ee16ee352f692a83276de3da43bc80b272448bb8dc6d0555bceb02bc6b0a5cba29a6f32772c6289724cc828c21d89588c80f59382851b7d7b7e2b09f2f3f84a390b934a069b3f93ebe7fff463dfdf7742;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb54285f63c3ed73738dfc71754dc2df0d50ffdaecbebf093f591b97fb53bcc29059f81429c6146cce4a5904f45df4fca907ad3ec3b9268da3ad30a7bc119fb7b25e8a93aadf56b1f8e38c7a7797172089f12563a1ebeb6cce27af3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d011a5fb69def8d6f3133cb5388029640d70f02c8639216bb9290e86284165a56d66ce80d3fa9d7eceacfd9f53eacc1d9a7da247c24aa353e1e31e19a6eee1b05b5687934d8fdad89259f48026b11616fa341813a818675e5db35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15da679bec8a113dfe67240ee63163a017ff545f6fab16922d1f9623737cc029bb163f81209df9c74f06759b28ed12cfe97b60d66d8cee2a5c5a051906bd0033a5d49601ab5651189bef22d710108988c9b2cfd6f4a99f92f9f99f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h71aa00b28b11af1d526b7a27dd1976ef082a14592a1122b3a3a76d30cf628154996e4495ae6ad4d0d7e31eb98333221966ab173237b083f84bfe34f9c74d0aebf6fa2d14b4e8880c1afff4bb5927ff6b9856baf3aad2f3b38cbc28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50183159b65b888d3efe4cac88901e2354ce775929e1881a68d1031e21ee8576c9312eca59af266a36d6a4e840cac1c646dfc5e1fac1d1ff99e7cca542eb7fe77d209c94e60244dd64e4076c266055bf4fafb507225b7fe199885;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1169b78afad50486a45cc78f80ba76e555b9f303c43a6e022b6a57314e85d31c77baa7305fa0a8fee7ae60efb80bdd03be55ad9a54ec9953bf1a6b1ed5e4851b5a7bc4c844e96ffa696ee779d0128dc8bbf03a244848400c10004c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha869d7dd1ca5eae9bed80a54d965fa3240e561fd1d97d2afa58c5996fde7a18f3583160e47a51506d8734f49f4ee2e2830c39069f0e1896e9c44b4500ad8b2cc9c63fcce36d6f74d933f1e964acad305feae5e48340e7f75bc0f18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a060d011526c9e318839339c9cb3149639d6462b7d0540b5bfc035958d5ef51344d7de8f19f67294bdf97629ca8c7a3c6bcc86f8f1237595ec2f9bfe6f282d7b8c353069b29f22963f167126fbf05980d5aa8b4b28038a9563496;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122d5ebe72d352f4c0bfaf9a1c50ce063d241499c4d63040683e6bdcf9bc19f97f82e051dc20b0688181a8713465c0a1682195bb3e1d5bb95580720cfb17ec4184ad32ab47329895a0048a2b278cd74245c2a20b55ce21d27ad0432;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69cfa8b1e8bc0f24787ff992fb6b5786810dbe51f0b8c66a2f36f3e6d657a5e6609805459f0a8189bb68c46ba631ae39f9507c3b5d31c7910031583200c8b3a4c7ba1aa2997bd1fd7f10be400ab28134db9a55eed5b1a54998df55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db88083a0089a8ad8a96e69a7354497cfde014b9dff1f300c2562596500d958ade65ca76f4380eb2484576910a80160046c911d2707ffb299b8d04a4b66a3d55c82861fbf8570140f9b8e59bfac2019ec7d2db9141ad8965bcea93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e6768b2d011be8fe2c826b37bd7051d45599c265062d0baf462cd99b3225d4ab0393d7e75276d5fe554ab0f515235c3c5d2f0be6a9b812a5d006321a70dc313e2a86479ef8f1fac350b3f65b0ea1ca6800326a92838f2860e3d4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf3345a9c4ef975cf4430ec6e0e4783ac7ba5192bf56ac0af4bf1bd765f85d6684fed014505452afcd541b06e3da4c57d65c558dcb04efb854cfad6e01bb3c1a0fb2e979f73995bed87e5dbe4a5ba96f2be4069351a35119f0807eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91e57ca0d981ec49aec79a09be3cb28eeac1e549a4691656a8af7774f1f4cb9a5d33e570509dfea34e700571e84f45ed76387e2eeeaace0702ca9183854f3d647cc8c31ee7e7c4b77f321dfba456c6c7f9790e8590e04796950ea2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7ed2ef69dd0b128bcde1be94d21dce8ead48dd972dd3ed2e8f2449e1c2eb974299d5ca29a174e60ee7a27ccc699b5070f430982031c99778da9daab953eec5694c3f169ab2519b3ca77195299b274723ab5a5571e540a8d8475d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14171ea6da99ab6e5d3cec039e56a7fbecad2bb3be5d448ef38e3580528d6f515d1bac832a7db5ed02adb122d29bdbbb65149d05d34c482ebc0f1219dd3df83daa88d5db9fb1735fdc280189d16d675a1928d60d2657d3d31479915;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc6936fad06e13d77bafe763c6f5d673480ce6bb83aca39d860cc688458310b616393524cab365782eec88259ba23a63558c7f5cccd21bd59da79e43a9923b8f27ec21e111a1dbe475f949274bf0b0353f31533d288c88ffc9f7750;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19be2a9851438ced815c980e1191ce799159e4374a161e03b2989b3c542b1bc04fd6f67e9f580643d726c169bdd0260ebf2fddde704200cc838f0cee225e94caa3b2dd279ae11c3b9feed4b2b433aa1c520d70cd48ded159a8785c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9dd3f44e357f18621c61f0717f2715ba150bdd7671756b0ec00dcd1432316aff08bdbf7ce7859e272a2b462ed0b4416a310227cb9b0b0d3a7add9cb306345cb7f6b1f67b3967a5debc4e4fc64749271a8d49ac1f6d520b4d37139e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d8a36232ae508f40cc395818bee49a880ad786fe8746022b6058d8ceb903b9d861b14c2c74f2bfe05cf9090e1b320b786d5872a1d35bf20941db6994181b74b216def0a7ab694f16eea6dc619956103c419e7ee1417ac6c0c7e22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h21fb5932470e1d4ada2590d22ffae6fde06c335e3b963eff1ee0a9333b7bb4d44d591400aff32561ca3e1d6adeab8e51168aaf8bb61a2631d1defede3d61e6430f6434c9523fa8b068589b487dd3d8ad1b1fcaba10817f563e691f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h820ed38d8205c690a04a0d41e8470ba75fa9a5841b7783985028e7afd1b560d44f0cf390407e9c3dbe56b49468cf2bf60050a749de72336a8116028df630f57ffd6a1cadd4576b061a7d3fd8127c807f47a982c35218bbd3c36ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d011063a2aef846dfc235c396da01ddc5706c0fc4d75173115f95cca4a11921601ad8cacf22d24f601bd9fe84c8d0899c00c902d362fb223aa3e7bea24b97cf96b3f9a464ad7a179f1cc6665b85771d30622773170191bef84488;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1243ca78877c03ec9ed3b7b0eb51b9e56d05fadb7f287da433b9781498c5a54551df478380f6863968992790ef9d5014e987edc5a5b530620928515694509386b1895746a6dd47cf14852d69ad581cb5db6f99d6a62c2f07094c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa634003aa0495b8debcbd8da85807de9db5009581625eaea87a62d83bbd021ccb8698d5858ffc8a6fe4f94532eaba5c5ed397cf6dfa77772e701790c868388b54325066bb7a327dc70346de4a75e1c86552406ec3d601e9b9cde6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h21b738817fa55b399dd560514f842e5b51407990ce2655519eabecfd866f0848485a850bcf2977fcf8da183fc9f3429969d1ceff9e2277d7212c3ad7f069ac90cd81417a96e81ff93d121108c16e2e65855f6c97f5f34c178646dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb69501fac8c1f3b615bcc801261b476909c3de2ba05ae9332c1b44f1e5d6408074278a16be881ba06427e108df5aa80b4b82fc45a66f4ccaff55e0e4979b5be49a575348520eb834c568c7557b0dfbdfdb83a6af669f95a53bd3ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b8b5ef5d9caf0d4b40120951f3c7a4d24614e14883a7eab7159682ec42be9b065e9d1c48186bd011e0c1831f7ca3ac519ca17f19bc1b06e7b7c08787a7f3f02f78b5a3ebee57768d2ddc642ddd39a225200cf4173c38ac055391cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1412c0e3537dc82c6651bb355815c611596065793d83af9776bb9f7fdb52b9a3a6a312813f581ffb534423ea5fdf91af612e208d09b5323c194df01516c5432febbc4b8b3ce7266a78970685e554a89b559cdb7445bce5872b0f3e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51cd5b1af0c48f7c6830c3959d5ec7ff148cc8a62d9e525ae3a4bfad0dc731699e77ada03c60bffb96525de986e4054123080861360f3e817da31234beea833947de7d543114112e9a2faf9dc03936a9cca9f14a6058487d55714e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad60f0e2404f95786321259840aa85482ac8f6424d7fd6e3a7e78f3633acf1eea774b1e8d2e80d90b24fd11dd4601ce4c7d44ad098a0d2e9b2b94f33200d0059689595b023f78d99fbeada39f4be2581035cfa44ee8ec5e8fed3fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h449f145ff52d05abef0b628140271acfafe51ba6007daf461f81646e6db084beaddd6b0107d4fae7932768730313da65d5fc7b2d0b3744ed6fc48382f12fcd0484b2e14b9c45971b0e249c06697a9f4bedb8da8f98127aad0ec9dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e040cbe070b8661840c327865a80b9d8869fee259c844dd3c550ed6df6a9635190a3542058bb06e60df0c45ff6e4768ab18d904eef86e0c8107188bca9beb4dea83cc92ee22e50123a09c86098ec1cd69ca57a03bea5695fe7464;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hccd58d4fe1e4c9e84db21cf740368fee6461c3e1d2b4ff9f6fa166d08fa5899c57100aef6a993e8a76cdcc0c1d23b5aef6878c0ae0562f43dfd4e20e1561da231189dc2d73e4114046bb30120efe8d0391a1ac11c2dd1f601b4ed6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24afab53cf021fa998a3ed5f690d8458dcbe22dfa30dabd31ba1babf66cbb12ce9181e902c7eefa3517228fb541c954df07a7c0e8f566839c2e478b3cfba938fed4b84a96bb840b0d2c4c4f2770ded4de484ca281a245909595dc4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1912deec6f1c0d8aef9c1bae2ee5ebe48f1b38260cb1529b75fe3728efe9dd7e9d58b33e3438e54021dae124de3aea3dbdb98570d2173bdbaa0081d5a4075c762b113bc097057a3b170b27725a416ba7623d331749be0ca2b9c7e6d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef4a82e0c0967c3623346e1eae084c2734de6fcdb7007436dc011ae58ff2cb2ad34318add1cd641e460495ae3079d1b79f1309f1506dce69da9df8339017ac314118db6aae762b97b7a0021b18a9a81023485d54b785ee507b4089;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h868074e554154f7005b997dbafc04841ec887fe5ac355ecfe11d6e2718bccf3de4f7b3f5f35e6998134498fea1383ddd0383eaac02a5c8477914c9e4a2df889ed8470774abc6d6ad0478aa5b35f540ae5b3be8d6ca9280cc3efa27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a73699acd3d5bd754930bb6c1cc24631feaf74ed5139c311c6fad4c443b8aa56632f54b91123eea2f3a95fcb81f7ed4fa0dd58b40a47fc4c2bb26ef51855fa3928aadb7da31e330a31e14e8e28a4f034b995c85987046ea89e54c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc79e7a48974a6de98063b1a95d6570d7ca65bf86df79584220b4ee18f4fcc8e3fed8bc7c0bcd23b93c8e804c93690b958475f3fd90984a4f9bca522cb081f6a8d6efe0aa5a7136f4505047002a8718dfb01ca4d280ffc960e74aa6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ee84b90d8cdeb59e25e8325c6b13cdbe7fdc9ef542c35b64332b5e738b3c194e230e529536aafcd3a3db398a93025815f472e5cdb0fe53769c96ee775ff5b89929fc14bd2525e71c7632f7d7051022f9199136ec86f9f49762452;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf639d41ed06c1df7f76a342d2fdbaca110b7c0a6e355fca20c6e5d33571baa69bece7ff7681a8da1b1db5a10c5d9d1a1e1566786d08fd976a4ab143af02bbb6b179e2ec6e401989b49cefea57a00d57e401fa4acafe14508aa694;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111fd7f10ce4aa1d664893625aeef32774bab93fc256e3bb2dba19c9ab3dd904242640e6dc38fb7a4cd462452889a5765d3737e77f73468a4ddbb8c0d9987ed47da6f5122d06bf895e7ca7f88f46425d13016ca8ad66425e459c579;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed5195e5d25985ce20acdc81d41f2e3bc7b56b4130f5b51c017d4a2341c5ba8c2454d5d73ebcfbaca761e1f13fa442e065b078bde47970307ed0a2311a9c0e3d53ea849052a6f5c326c225a8d895e521dc39583faace2eb83e919a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a51621319db1872da69174a9f342dec1267b9103c49669b125888f7d92fd40df59a0c99b07b8efde666d05ccbc421fac446aba8b5cda104ce7e974413f0fa1762dc45fa74d4e44079192f0934c86c7939a0bd0bb45677e3d6f4a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h730538d8df9bcd8377efc5a9791b8b6d37f9bc7b1a7525e743910cb028d320f7168783ea19d9555851f3a4e5863b0b917dc1e4492d65592b9433272f9716690a02bd428f89e83a90a31a346e1603539f2b5c4089b5f0b82e259738;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a26be11e07dc690dcc151fa8b359a14bde0b4a902648ec7de4c55fbbb24517fddebbcb760689aa047bdd8af15b3bbfa13337f5af4ba789565a25f4e892ab78137e38d19d46787e502e59eb2dc1aa3a7e75fa6106a1f4869ed4e274;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b86bb927f37b6684751e7ad6dacbb72787e18971a38c7431f3b06325f0091e6a0c2fb6914ebd5a2efadfde59e6bcc8bad4c06ffbeaf227d03e12e247cc3ba9073dec0bbf939f2a0a3d1f5b06836ce782189a086149175de897521;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1245ea376a1ad5cf1c95a86cac53444aad791fe407a205e4d539e73fca8494d7161f184f88f11924f29eb50e9b7cd37085a52958266bdc4e964b9bd422b087cfb29efb57fcaac9d12f049a90b2bce40cdb7030afb70d17994361671;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca8029ceb488b228514cebee4667e7b8a1ed56def554e73cc8d8039ad1dcccebfc6831de97472e2b5f11e57bdaf424cfe41085665d3c64a8f1afffd18fefaec893849a628263aacac9931709ee164bbb2e4ae263c0fe15042a36ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h268ef7e7db9d062b27b99e463831a313255196d77a844ee12b7df8db8c8055a28adeb8995bee5bab12e9be6f6ccd0a77fb4e6cb4bcc8468e255dd74501f688519f96659948ab7d39f8d691d0b880411723ea328ee7af38ed59810c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haddd81b0869113c20e28e6283975e6f1479ba16b604358c262417dce3476e2971ce21c72dafc3382a6c7e5205e4ad86b7f06a3397ba6715368a7b9287ab3fe791eea4637e3fd3b9c6302b0b75c1f4f1a47ad2b2470410a480ac27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133ede9a918817aeef24bc2e8e80b9b18a500557c8af5092efc92dde7aa2ec7e81cc27fab8a271949c8d582e3acb046eb421124437e7512c213500cd98b4243ecc59646280ce0735d5d02c971f1f00202e991c4553b50bb7201841d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5fa869095ae19db0d76cb64ede154b4a01af3f2371eb42ea9029f6ae4ed239b7be4cb22986e2ab6fb43944d5c3c964f7f07e7de8fc76bf22928ade1473da5a9e1e42b866b1d6ecb75871ed3c3a0bff3146edee162a14ccb7c077f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ead8797c13bf349f94f96e8ecca418b067c5ed8e458ad966510e328cc44edbb2c051aa10eff547682c1f7df074ac871e0307c63002b37c6b2e42271c8da19af7624543e5af1a3929ddcbcd883ef6aea94f0d9b66a9c84c4b851591;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h82e258ba562d4f7a43e34be096ae08e799a55e131314ffc5bfd1ab0405dd432a1863d77970d910f78bac3fb948a84b3fefd22e47964a3fc00b5a02cfb55331674bf9912c660c311896c98bdd08a3befdf95cf146050d2fc7342a14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c27cca546116bf1a6feac0b63b362985c75c3a117dce48b2804e4a7d42eaaf33660e7bc2012a943c387939f6240a8ceb78bfbdbddbc2c53df3877b281334db9ceefc12f5404e6442d1081545d3f286a51ab1ad41c56634c9de4ba0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b876f3bcf431f00d6f6848fb504ff5171242e84f3a75c882febc6f6111a466b50c71fc25328168c08add971f8d5bc5473cc52532121ed77be1bba7b8a70a1ae8f7dc27ecc50c1d3f40a3ac54832b3b4203aaaf9693c7aeb3d55411;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c70b49d0f4d552cd81c8518ff5bf7f36eefde3bae2a619f608c595529727fa171edc515e8c7e53db1d956f97c39ca4efd03ac5f34d484117aa79e5bdcf2708ecc7d32fcc64d819966892c95cce88584462095b090c595257bc728;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a92bd7280a8ee1222a023f6a31c76a2e8a45d017262fdd9eb1d4baf5900969e40db87a677b693d7cf1792f739bac28dfe653b6508629dbf905170efaf9aa10f4ab1cfc14b21b364ffa9f85c4f6a1c66f66fdc4fb0d825dd12c09a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5cbe5d53565707e38936d68cb78031243612dfeca81c42839908c9d6c41748e406739fd67768e4866643b4a4bc1642cefc30415959273d0f640a1dd89b710f0ecb857483e458f39e9d87bb7c321e7d013cc8dd3bfe149a6b423278;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6e357b202675c48a5910dd59738cc33ffefcf0594a45dde76e52f0dc52bcc340227365368adc7a9f2d09a108f8714bfe6f7abc8ff5e4b62b912547125b557b7fbf08335f46cbd026f1f40485cf1ce727ce97aabe7cf5bd4a649ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e4e23edf36631bdd10f27c8d2f7e7a3ec6a75faedaa8cc6b871f86833645fc299ff5fd439b0c50ac06ce45c44811179d2b1808e75418fbb88e2421f1a4c664c17d3be36992f298be4e3f915a9588716252f67e3e46d45122018a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a31672eb7b74ce994d4fb350fa0b62e7aca331d5d49cce3f968ac1e29943e04cb11d608727c51cf32b50b0222423a2e75ba1f669aae8be5a5b42f5a93c31328b4a5d37070bce2908b1011c6d3693714f135496b2cb4eb071165d4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4c3544ce900c466f1e93cd359c549323245ea9f3e2c7428d88f0d08f2a75d7aad17324f2034d2495bd7afccbca5bbd131d1ced5a80b1929015ca1e3fe09d665fd753a368e6334200066eefe6e58f712b2aac614218cd8e5f608f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a9d2e9c0cc1506d4330681df831e12b908e821b83ecb7b6eb77067896bcbd0ddeab19e2f67f8f371445a624cf44a1f784ad34bd7fc4250835a14018c5a7b52102ffe9d6c3dcd4865542234ca05f351bd8b4e96842245edec696c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5557aa4aa5a72eea8618df19202979b8df3106d1cffc0b8f74abd300b081d1f367078114319e149cb894346f8a666e39fab9b91e38ebf5fbe1465aa23c614645e3176ed140b895b775fd741081572f85e93cfc13672a8c82f8f52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f861a94711e094acd54fd0a3573131130eba871b93df32eca83359b8b8441774753ba86689b78086b637f2142c88f4f424fb469c2cbe5dc67b98b984e92a16010882843b7bc3c47db089144cd9da5b376facfefc4f2ba5350f54ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169d722690f8945ae67ef99cac210f9a5a0f29457b1ecf55a737a8da29158a7cf50a71ba44d030fe15de27c6b89eefa7aac015c2513990d714c94d986f0efb5f72d8b9e006da92227aefdc60e3dcfb68a1e46bfb6922d83142ab3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h830682434dc44b01be39f6e436ea5958a14bf85b27a63c69a1e249c0301a50662e33b55557a29321c8894165a9e13ba1fe07ece264173be4c5a994c740e6418b6cf637cf244eebe5855c24c042f3ce53842ac25c2b65a9af427a9d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2eeeb6067a57d7fb5567167224344f34a037d03b3818c74aa072b03e83212e951d98ac4a3ff08f390df48f2a9072f62ced5bda25b5612003559784cf6027892d01776a7a6c6055d387a3158a4ac0d6650f880f16c3f9cf95c05768;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h52267aafabb45c24a3753e7bb6b416f34b910dec0a289ea439a073ca96e45c94a11190c80a1c9fdbf606e321d995841a3146948bde9ab7273ecb57ea42628f7d9111f9c704f592127dbba47daf0beacf92d4df0faf2be34511a1ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa3fb7f70d4f001010e6ee82c430f0cf18d2daa7c36294b9773ded39a41e28da4ddb186e70549133576f48b0125116c5af780d68c7004823edb0676bb2c6f8bed72e6042301e33b6b4acc2fa2c85e80deaafccf5951f672b9dacf7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd42d6bea69e917a18c29e03b2fd18a1fc8014c654835f30c82bd0d5b38d66ee47b39bd060082b5f897966229d38a624103636d58e760a5b3fa6224f8653e730ac27c5cdc3fb606d11588741525a24ef39bb42fea7f7bb41e9abc3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7dadbd12e966e28cc6f98f94914c9ff03d1668578acb134069ec67bcd0630fb7930e3ccb6b28ce318c1d8c724c98115819307f5f97a9cd46ccf68a61527b97071c8b5846048c096c85a352d22153f5926b340e3ee426f11cd0f5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2605f141f8483e557445495756c6eb38c23e705fbfa8f10f99b03dd915655160211f6f258f26ce24718897a97b6dd88eea90285f7fd1b90f5e3417d5849737bdccad240e8ca334a158299a757694b5e99dd8b47f048d6c4e070bea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h341ee60c362b6ec3113c402f98ff1499532ea4b3c305aff3b0902c7b37023b7f0d801b042c553d4162146809c732c2975efdeb629ab2eaf3f72d8fbe017c26c8fb5f3b18e5e77aafea5bfe24579c4be271595edf76c2c2d1a7ee0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h159bc81201838f07e54d22ac3fb195c5b8e17c3e420185e694db8a7a4a1a283d94cbb9fd5c911e1a5742c568d2a20286039ddb709bde2b6ae532c5def49166ff0e74e32f7d8a43da9ea8b421832878234849b432c71ec56c9709ffd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9056152c1b4e419b415ae42c4c8acf24630edf4e540fedf43983b114597c79a9faefba2b5fb7f3541f1c2688614638a8a2d1ab6a781ce846e06bc0fad54d8c65993138556dd76d6abd62eed0a77676fa84850f60f335d09fcfd69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha93b53b9a91c1ec88217deac71dbde0deae7dc62d4006dc1b4d419d2fc9ffcc6b83ca108b768b19cb0ff8e7c9b38f29c3d17c70857fddf129554b1856647b8b4e1db4ab5b73ecb8ed939da1402c69a4bf8d2d3eecfcacd3e1a3616;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h151eb82f50bd70d0b913e9722c897b365226188dd4d886358672424b4beba801458ebc87c1832aeafb258ef14c1b4c490ce4d1a3e2449f6419ba8ae86c424973e7afe71b500e977289b3852b0a135e5d9bf3462e2893eba3ebe0fd6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8e27c9514a888a8181df2298d6e9742d50eb3fffd82b613fe32f483c3b9616e43d60f78b1f48f88bcfe4fc0e3415dfc971fd1e2ef2c8870d0d18e6e2fb2df2325e910770e8e371561bf15a14bca69b72f3c4da7f57dfc0c36e5b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e36e701e7987ba45713aa425dbac29757677f97b0879db0d6c414d144aa1bd3e002b749b6b3a26fcae944a3daa1e002827a086ee2b81bb1feffa6866c1f4b3806765ab3a5be5dcdbdcefd4128f8aea8bd454405f04be284e944a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haaf2c687c97779aaea760044b1d0649c630d4f790ea71cbd45a084d839da3893b8d0708f8b7efb6ada964f0024d677d878c832f022bbfd2f241b4012b4a1c0be40ae598bd3401b3bd28f98e52602380c1adcb7d994dd3525fdde79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf1c9e511fb60aaad5662aaedd915f418b7700960ef57ac21e80bc34d97e2954aaff56fa33cef2d9179ca3c881f304de0771c9061d362fd75af0c9cec50f1381b117f52a255bfcb75ecd5811f1b585dfd14736f61ab4b5c622685a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h703b3cecefe215ff6937776f99af4ebdd6c4d88f7ca7d02d1dd45f519e2dfa71577a4d226e7f4049d3eafb273a553ec019dbd50d4aca28b58a5e8c958585f4c71cc9bf60819ffcaf7f42ea607be6883db8bc62798a6e83f595f0ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha3c9ad32bc8befd6331ec4cfd0d8e0b65459ed7ed27d57fb7f76258f4022ba355acd625e8ba6b2024430479722f7ab49a8b548b64104b85161048bd52453c43f2465bf36a92a7d1546683031d10243381782215cec074cc5e1f56d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85f4f4c35a6c5da2fc3b8770e5f1867b713123337c81994ef06854d16a751a825368d53ec121f9b2a991e4c1fd9e492557a026199efd6d338ddaf2bbf35b129cb09bf16c16521dbac928b0f62284e36173a91827fae6d125adeb7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3f7ab5974e743cce5c4df628b1a2f43b3d367d28710c35688a5ac20d05c2ca15ebbec2118d74af75f6cc48d23fad2e7964c0a696bcc745742144c2f827f0b60b6c443af3c29264827cd53ebb9403c77266126074e5d464c62287b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he2ec07a9fbc4be36c5b2538f3aefc133e8464cf2bea59c9edcf2b2f77ca5e3f9a80c7690909ef375a3beed6d2f4694bda7b4e53939e30bf8d52a45bc15a506e2a5bbd9ef392aebd36ff9246e9a9032cf995e40edd947a54a2fb99b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed6e7ee6e0e291aa5be01ad4f2e27a7efc27da0cb1ff1928e15022c07d61c63c5386a35a0ea48f9e725f4dce7f5bd2dbbc8385415793cbad23ead327fe4f225c97b8c5f8a3b3385098b8c4bd6f42ab3e5d6c6d90e543a931ef20a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc5883995da4d43e94b3b9f3f59a38b1f4c4a80e6212b794115f1df9476f7ae0fa3970a28df6b18a10ea59bb9bad11ca9ef08af81d1d13d3866ea9d12d07aa0d567c652b61d4266f221b29acf010ed874281fdab520858ae9ed914;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1397fd4a7cc7869ba3338d80ef3940b9c7104a76b972c470d93f1af5dcdb66ed73630625f6fa58749a41375c5444d8740c63a44efcad35bdc8ab43e2b716cb0676706985ffc26b63212d4fc9e9eb8eb63f930d8d1c290138c90c9e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha15d3f450e385235dc66d31bcdb99684bb25f4b4c5ac5f3e3c41f5da2196cc5d581d72ca2049fb184cbe7c1b1e22a034f65eb6859fdb5199f64d8ceec6c6f28ff384f79bffcc267b4a89e9776087a5bb759f2894657cf8bc2235d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1546d48b8df5d7d2966dd5eabe177dbe1eac0c81cb7ec6523f1260b2180e300c43824c14b0ffc09ba7b4c9b15c14df0eaa70f77a0d9c7bf49b62d36e5b7a72f5073f1125bc8804411174ad0b454b2ecf238c55b9c5e61e44f70636;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he47fa8473495142d1d70807f8f497d13092aafab33e758c5dccae9b7454ac9f59f5cb157a5da231f04336a7a781c33a70704a0d2bb0ab09752a0a88526d536e8808abec32a1f84eb3f5ebe4730a7ee7dd156f012376c3b116c1767;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1858dbaf8ce2a6eba2c7561d3428040134771e483e6f14fcc02c4259bffec60d52fc2c8ce9187ba7e863b14ca245de18bdd9a150842785ca6144b89a260ac6ce9455d7bd363f1c1ae3b52d2ba79904e13a4ef807f69541a5fb1e56e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152207916f7a69b9f51a3b7708555390e31209b8fb543be358016d25b101bae303af1d24268c3110ed4e1ba635b3f05a8c5f36c1f9faca2426f4ce05e1ed51987fca62506ed0a0628a5b12911ad5302659e9ff0d40f2ed6e541fc8e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e0160194887b9bc49eebbfd9819711e21505cdc23d06b976df8fbd9e788c7caf74e54e40f650161eccc5fb1031e590d93ed29c9835f05173194dec13400618630d729c89b56555d3bf28b71869b5af6b0b4983722724dee084852;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4bd4a4a6424088e5a915be696802eb4eeb0418a6fd59ad46449cc83d776de577c42342389b6d85271e4ab6ad0a2b7403936588a16c1f4ffbb6099f48f1912ec622c83a65e237b2aef93cab2f6b6b7bc137a40de7d8ac898cbab241;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98f343571ac66fc8bbeb2de2849beca6486e1bee24c710588a7ad94bfbe358c66335426caec75feada653007e168e8e0c5d8dcf7bf6cb81594a38a35a0cbf0cfb6e7ddeb70415cd2dc09b8708ed56dd0d1b55e8fb0fc37ad72478f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda942536eb9669e1405c8bcfe8cfbedeeb7a60d5c795deddb653a9c967bca3db8d2b1c2a5575fdc8c59b9998fce662428dc173ecbf3d2fdd13fad24063b1ceaf383fe614aeeece229f7eadfc5d7337be1f5aa68ac3ae2c16a4b417;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a88783f87ccf40351dd852ae2a0019891d80225fe7832a79d59690cd5e3ad7079eb2e1204d8946518731d96621e56efb2b2e532bf57780f98d4225039672ec419f778adffe6d2b1e21e68666a7f1371a1d569eb96049e6bfda5d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182024d74e6587f20e0ebb4d70440a838d85d0a5ef99af42c7fd6f07e6da3317fa7258f978568e710f2c8e0631e0985b8d0b27669f83542725174831528be971868c62ca70358d0de37e0a6f71bbcaad70305335637bd008b2a744c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc7f9b665421d71a04a8c3cf753f070f4e006e047bd4a68cef71adb881774ddccd49cedf0e10912315da62ca481c1017b3c45cfbffa0ca2a904c6c1a8e41463dda4e598cf946037c1a40ebe4b013a4448b43b6e18f3556dc0de4f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a289f88ff8bf0a7c8ae6afd0d48c3301144aa054d00c6257af32c81fe77eb01fac5f15bb82de2004826d991360d488a0681c03f16ca26d2bdc107fd5a5d232de8e7ec422c2e7f7edb084a213a6e09ff5eb3363bf379b9eea628b8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b21fbf1d22b6cb87c70be6a81db0e5ce41a8fcd1773969533668f1272c38e9a23cb69dd3783ae49c54e18fa82e951b9a390f787dbeeb8452d6ce4dc8f9a643b34c7999cc26e642f958afae61145a30c0231b8ed4ed8c7819f64be7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80d57c30b56104f2368bf620016a7cb7f25f8a3393ddf1969a92f5d96e62e61718e0e751ecae1d430c630af4fa5cd525b5728be4f3efebeb42d0249d6b9e6e119fa712416016216cd4277095295b9313ecaa7e89c9f34f930197b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27e8c70acec457a21e293914608dc5d49feb14af28810bcdf3bf73ce229eb3757a7d0e09faf831a1bccbac4e10a3f707e8948ba7567694c6dec151934e1f5ef94dd5137817e24eaf21d609072ac63cb8a65897c68d29db31a62b50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd5cb1d38d4ea3fdc9f778e6dd92ddd720f626d956d9be0f9520628fe0d3e873c2e63482f75968fc00bc77a95c8e9a6565a314b97491c264a1cfb5cbff3fd43952b9637d52e59d25d7730f99f5a43c26e17a4991fb53dd7265498c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5d6e1a02cc9b8c4c45dd347ac5a8c98dcd9010c9266ab5117ae67acafda0515c315e1114871c807c2ad2a3576488233f4f621d42ce2701c3c3d3eff88d431d2cc14a8e2159a4c97d61eb5e9b221b527f183818c86033ec2b36a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13cf882063dafb0a786ea3f920b4786b39ae250187dbdf0c4ef7e62fb651f89b7a4c31f5043b05ff08984cc3ed0b40ed1394b081aa4ab971102b18318ab120c006cde690ab48b38de0f85474683f6f04b95bc617a4bff012f1904e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfbd26209ff19724d39da0dbe1cb253fdc69bc24f85f6a3c650df5866c4efae23f719128753a73f11f534ffa7ec609b780c5b5ed49c7e78e844e6e30ded13be5d07839d9df83fb406d6348396f025414724b4b0c590e984eade8efc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1814e1e3db6ed2c24a0f32f693ffd1f7ef9621837a71f5db4f7cef71912506da33082e4facff01dd8a54f10d7763bdcfaa03c95b65a60541fdfa707225fe68ac2022251cecb412d133bb0383453da55ff37d59ff31509970ac28981;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d65ca790173994e2e78ca27a13d7ae963ac052e078d0e84149551640893b3806a88bee221e36a4b2c47634e3692d13f98334bfa40a8b34dde9d9c9c57b2711ed334e7d8d67f426be59d5b840ae59748f79a9cbf09bd1b94cd825ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd8bc92571dcaa8c9e18ebc1c3846ed83bf879b47b31f69a3f91d6601af5d16af93759b73ad3fd515889c2e2ad389dd8177548ebe214c03e55a7380bf0425f5732c423002f68b5191b548494561a5d37b6533109b420b5b797c7511;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9b21953e4b766d858ea2a9d2270fa0fef1fcb1fb64f971a4cc853b9bd3628a526628c75421f9c4a17b836608bbe2b9c5a2704c6989e00f7c373b9b364928fd0dd46c5bff7424ef5e08c5ce045c81705b99b54a6fd1b9eb2e24c1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13321ae65464ba7555707b30d45129f1c6d90dda97236e9c5450ebb738dff791b5e0306529118e0f306934ff0201af425ac49ad71035670dcc03707517d8edcbebdc70fc226d93fd7927c22cb574dd39faa8a1d1fa80b24fbc59866;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18cac76e894fe91e08e514ce81762ff861ae896f0cc46fc55f997543b2fb8bd674880f62e3c73c8f6b2b2d0b1fb92f99fa264bfb4d278c18a2b0c7a4493b5b3f48738f0d73884b470f2dcd44eb0e5c555ceb5de41d47b50b95e106f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1986b98e8a9fdfaade9df6aaa13c81cdf8e0edb7137f098b5dff254b84d82fa9fd56ebd23d7f3ac7fc4abf79794192fffdf98fc68c97400e5b215696313a33beb916d93f642be75e2e6c6ced7b7123ec37c2c3783b6865b35151ffd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcbde06c946518467b135b3659fca2800ca598ddac518da14119d2fb57a75dd9e08065c6b5e696b0b04def5f11d5c606bfb8501790d256af566e2e365f626131876539085f611513491e570311cfb6baedc36b57ebcb1a2541cfd00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a009f98d9a34639a9a73c41fdacbc44a9aaf48b5502c952967af48775884670c9669d15b17d91efba53e3b960d529e00f6a54c4d1f487bf0a0da7fb9d9794d13b6c992ae54b43f01b5c3441d74ac5e4fbdfb01d64021bb21a6764f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3a83fafafa7fceb9a22df76c1f56369d37a0cdeb81f1549f3f2d3a2e426d19efc1a2bdeaeb9f14845c77318e88942a637643a5702e6c8aebca8f30e458db2ff160e1c0f07c8c43d545640ea62974d48fe511c6310cf3d4be28c74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf937b9c38234e817604923e3f5d6b7493234e59d2281b894a08d9d74e2b02748048f602f117b96c220333fc9d98d58d43db86d052a2dc2bc1b1cca9de47936286769e47f0ad085b072a515a10bf048ac7640b70a59decb7cef01a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8fa8aab03163df7dd9385e24dceb926503659de125ab375ccf5970a968c2a6eaef50719b8cadeda8f50ec67b89ca15bdd0c86225c5c40eb71d657ad23c4e7566d17aea394fb2f5274e77ef040d608bb708fb314782b3b61d9c3f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1260da83dfb8c59501e75c39f15c8b03b2d851e51cca8767a8e5658c6adaa778569441b8c2e1c834c8189c358f8f95296336b27b614b03cb8a4b42bd2170e4a10253106d43446721b283aa72fdb16f15bc3c3d0aa575199f1a0280b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d640b5f34bab02478156b01c33a7566f7fc9d0f785308ed9108717c9642852ad7808e4e2e9f533ed079faa4b4bdb1e9d1a0b9162795abe205cc6235fc2b63dc0a982702219caa976dd4e3666b854028319be0832fddddd3c7600f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188aa6119b4d4083a615f8850d45add335480cc61782c8af5f3e9408865af1c10071780d671613a3c876896f11dedabec858133a37ca0a18739ad99112b5990a054a0b8ea7409fe3521aa465b4834a66625be1e6d2ff5fde9b74f3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ae3888193214da5820c5bda4d07d3881de636bc9b02fa26e543e89f049083b04f792a85d42307b7e2279a37dd010b18f9d291cdad1ea5b6f36f887a77697d3caf219053a1e47971a87dd4ea7eafb1e75f0440cb3fff01d08a69a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1edaeb1fbc33b76616e174ecb99ba2a1d464deb5b9445f64153b23310124d0977baad87982f12830b0a08c6f1387f28c00f1b85c07efc8bedb3016c8b3f2828436034bdc0cd0855dc32a2a5f1ad83264fb42fe8fa09e288460e8f88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb204ca55f010dd91c6d3e90706873a927b3332967025bcd460ee3658dc49ce63a6dbc557535c794a4681bbce747c5fddad6940635578d79b4c0978091c6ff7da07bd6aa049db388f97e9f02aa454e189eb6b0687016b8e80185949;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3db5fd3ce385dc3740db5302f48a0c0abf87720154c470dde43280d713c2502847fb6ce800ccb7a48728a51aa3a0c46a3c9c0ed1491691ac1b9ae316b5198ab85f2befaadc4f997688c8da681f110af646b55cea7e72f0fa3c64ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h938017a6c54c9e87e74a53e5f5a784c8c4cf0b2eddc6a4db6ddb7ced161a6d12c1bbe8e5e8ea83d2c8b69c02b7805932b4f685ecba06ff1e9a904ce0bf17b38efa8f728a787607f750c64d02cf10e60470afc44a6438b21f467a7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1662f627ed5ee45ab59f88969c82efd114b8f9f4ba5e3c78636341ee9c9e4a7d18843fd4cfaf6226da762de97cb905f37669ac774cdcf9ded0ceddcb3daa36bcc936de9569104e245d4c0448cf5ef972fcc85787b81d934a37dc0fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ceb87c5862f41b85f1425f62be1e3abd61d85e4e957f00a3ec5a997a5a789025fc60802515e78629489ea6fb359e60e4c8582dc96560222c874ef31ada22248ee335a47f4c8bf9f7741d4d494900791175a101aa819d788353f820;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1afa678a5bcc7b35cc05edeee6b8e42611554c81f94e8c3fdeae37fc5fa67a22c4a7767c63244dbf95f8b253c27e5e352873643e0a7de2ab28d1d9bdb05ce7363c48666853712ded425d53b2ce52fad91a8d29a9f27a16a47de0a2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he34b4f78acde9f1b1e3a6b49f69b5ef82daa472418b6b647c559bf71f1c2b813c1034bbc109ce676d4488bd8c8ae9ab64522c28dd0e575c504bc6c579d39b15e508a12060f0cea2958687fb6f01d5cabe1302ffe692963ac40a041;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef4a9ab7c22807189a0b08c4b59b283f08571271f548d014b29d48f41174f8127ae6bc12a1dcd42daf95e8a4890a7f57586c70e596b5186a9424645c5e7a46e3f8e672431cfdb64546a88160150c9b2fdee96b4a025c34fa83ca15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b1feb1725e117e537e4bf95269373de51e6e3f4d710a7d5e5640ec3395720cdd630450b77d84c72dad26831810e0e36b0b3ad0b4b3756f959ee885b2d6b7ecdb4b99049ba4687068e0a3af72aa6abd8b3798fca13daa9fd7f42bc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14deb373dd75ff0de6a01e844a275d8019c414516cfa73be54237e8b84412efa04952aa8538be35528e479a114b74b0fafd6acdfd4a20672dd7c93f51d76a54e466b7bfe32219601c164b1381401f9a9481908b317baced2f974217;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec97614e9e0df6e665b26c38475c6511341f372b50a2be359ebdf87517651386d382200c99c111737df48b15988570842f55d63912985c0bafb7ed322a4441e45dbdbf925c5a35f57a2cbd23de332b37543c49f491f3f3116c65b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f85ab7166370fa127fb76ef21394b89e909b02780ff390fcca9cfbdbff7a06629df18b85b7e42509204ea9386a0e8c45d1941fa12c4ef3110d628643a907af4c7d282f06b6526ebc048dd165e442b436a8741f1139ff77ea2f3733;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h135ee96bc0bb62f4d029f7b8c8127d379f73a605a26e9d61873abf755d8d4698d610bf1661d397ea9c72dff1b9788d06dc2c00a817684f798eb4dc73a175493cb2a8c3d9e26c64fb5717822199bb5cbe4d60227e560d5046cd5657e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cccfa2bd69b9f3fe08ccc70d51846f39448774b3a5700c3c07c96dc869b95f99b48b2048d8db341d0ab5fe22427f9e5f4f913fc2636e8f91506db7f3e2fe16c2ec4749d000f677bb59972452afe02176d691497cc307133e7e3ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h138a2e90d019cf1c3bf0382a1c3c74558692fd5b3eb438e6774bdbf188635023ffb502c8ed40bb91103e05f609acffee5840fac08a8620c4090aa40b9b09fd05ee419f72edc2bbbd24a07e866eeb7b60cd5e30334cc247afb87c9e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c13d89f56d7a0b5f0a1a13f381d9b18386ea908e74c8f8cf5510452fe757aafa9d4eea9e93ac5ea500c5e499f950b38fb5009980c09e1f831b927fed4e457d629a47928bfff9507d18be264882c18c30e628ed4d427020280d82e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5456fbf5ac34c07d035c4a269ad8fd2b218269466a2091a9a1801e938ea6b798e536a8c923fd28a3bc5b14ba9790323ac07c4fcd16e586d736f638357055bdcda8ac847ab5a672680cb1d43a5ec6b4da7160e335256564e42e253;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc901fec55a88d17518a9892fb1d2d36ed5dcb39461df170c02d00aa7ed38d73d0f97797f9cb62485537f32afe8ec9ea52cef3395d8caf5e0be31e28f79264ccb286a6a21fb6d902fd0cd31a6b9c58dca3958b9a039a3440ee6760;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be7292e78d1df1c9e5ab7906a78ef43337d781d45ba58a5a11870b515b620fb60d474be8d7a332346a97bd289563ff66896ce548b3d290db2dc76aa6d1eca62f96568693cbea19a7061536fccfa83fbabc2a284ad9248def4ae7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19bfe9ce32baff8fcafafa6d87ce9b9b06433d31198eef55a915549f19921de0b6977666aba8f6bf2d68f8cc48f158f1723f7ade53d4af17bfa5229f62c01be74028087de78f77c72daf9447a4a1a861908d15439798cb6be44abe0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1064f09f45ce90a8c91b441dd72789730ca1c9ebd6d50f7982fcf97651e43ba6d981ef7810c696012aecc717b06f26df89eabac7f421fd16f1c1a283fc6dac05dffb05b1e147ebea263a7ee918f5b764dcc3e48555bf0068111799a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h163c86a0c055ce9693a946d419377ce203468d61f489fcf258c9dfbce8a3c4a78cb6ea1c64343e1df887c22ed16684945779b4efcc016fb53caefbbda870a507b86e72f8ccbeae84e573223e0951b2e11125e622ff9ab0d662c5c74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79b3b4e3c655817028d661b00c2248288b12981df705d2ef5aaeeab397a9386db6f3456f443b74f60b290c8ae854578656be66691ba06c053343d84c80fe20fcfc8d4b08fbb86f85ef63f09fef3ff16d8b34b11a28da59621f1f24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a4a659e731c6dd30141770980fdf975c3024f73306c2a1dec9b5ea7069e817aa7b6f9746005fe1f8181c9bb4ad901db1881046784acb7ec599dcc3deb5bb8d7a5b80b8808a9c3b7e9272d6355a6fc56bbc92946c33e2fa82d0853;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f072fe3e9fcb859a3c84bd6c64526377eafd2a31bd533c027a687be9143acc7d98e88e775fe6d5b110a6a91ac284b22d81d1b2c40b191ad7d11ffe217a2263648b780368c9aa2d2398f7f4a05f6213e596c86c8c7c7dcbdc7f3f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b61edf8f9c9cd34ce7fd296da526c82403c5ae60d2b87956a07661dad2261b21d77cf651839aae4512edebc585b74cf127064f193d8ca4ae257f168fa388c99879786c16bc201305901d2caa0203dbff43aa5463e92e55852a9979;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0e5b42e50dbd07313fc4249c4e371c118f5d76f6bf40d383233572c4682c00dd712bae5de5fd2f41c6500a14a685845a142051339e8207d453cf1456678536ad038866819395baec7600e0b94ac05d08cfe2b5a50e97a3abad8a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18733dc9d745863d0861271a0674de32e5c3cacf71ca76504e5c210286c7a230ff74701e98289cec2bb3b07e3c2ae4afc7ce4f980a7ebf4c08c1c27fdd5e7d3d959f2059cce23437f780afbdd15f81dcb7c8934306d2990f723cedd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ff15bc00c7269c07180f194420321db76261835b91db60072b09d7cafacb0332168d98d9894c21b4acfa6420e42c594eeded1492e9ff4afd37d86d3447b45ba7d8f310f63826a0a03018fe3ca84a7ef5339bfd814fbfd5e8c6245;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a6c5366c0297c4221fc6a9fa81bfbf0290940b348e79cf79a35b16f41c8629121e8c7b7d14e512ab9ad522d578b70985002ff778440b67ac4866f37e878b248486101583665abc3ad3f991b9f831a1262a952ab69766cf0c14765;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec9ecbc2711890894c202bf903acab43064643bd2732d63f141b90bd55ab5463434d60f3ec2b9a2933dfd6e3aa38d32354d40cb2186b45f58b4635fa86b4fd433294e000c8774dfec1fce3374573eb65eb8bf013d15d1a929b9b63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90b5fdca61bf687e244990620f3a00a4e6351669a1abf3b56c6037c46388bff901dff3eda89234a1a5f35a6609844c334724f7c2f72f89b53ff18f5ee5aae74c2dd023ee43e5555fe08929f3f403ac2cc84c43d036d41b26a185a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h84c0ae563f0c6a13249f80eca7dd7c874d70949d1b0900e5f9fa3a14d1a025ed48a7f512767ac0e8fd808d3d2c55647f3194642741f6a183db281982376fca5b9c6ddb4d53a4026b150f3dc4fedf2ad1f452293e25653b49a93a5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a462b9bcfb7bd832c2e177420ca8cf9adcaeb7bfda875242f12ffc1f37d7f825c055d1b65a682b346a87ac7d4d0803f5ce6f26f196034df2e29d0b90c4c24b8c6ce9c9fcea555ad769a6c988bd636c5f05a22a68a5fc133381b5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2bc399cef7211aecccee957d9f1b9c62499918c58fa6aba532c70574705d0405704ebb882b32a248b0b01cee84c5c4057b6ede6d7b4e2a688146870bf50cc789e2d038f4aaf5eeefd9c41f9f92f4653d38e899eff83d2d8522a2de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h118e933f2a1f9366926f5848321eab7f4240bfce1db119b7a0155c38543b807ad47cf2ab57e08b58eb1ae8ba70b8c545a70676fe4dfb575b801bea9737371de4821f06717b2fd20bd2863ce2702d3183320ad322f907527cbff42e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc299bc5de7c9aa4ceb6188b19de4d2b347f135a01b5d0b12e13a6fc5c351d50c9d3ef3946ba924ac5d60388e61dd9e0687dd62ffe790691c27208a77f96a9a26d182d3725421c5d4c507cfc9c0b77b57fffbc90ae171566b3482b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa3c6e84a548e7a07abd0c0550ec6422b97f2611c7939a5232eb73c81108a33fbc43d7fd0dffa445d35a40d1c309733847e9820d40cf1d5ad509a1e57cd9e37fcdc8a2e2c58840962b55b23e1b7b7415eb8584fdb4c805b21dc961;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9fe2083e552780fba338f36a434b430abea5b25f2d0a6422705fe9fb50a3ef82abcda423715ee9dcbd2d5572a18ffc15da733caf059eb53ba581e027222d75fc93fbea0ae52a3b928632769a955a3206b3760422e685678a553257;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c43140aa85e2a0274dd3e336ad0af2e50b17db7a85525799f772695429c0dd8c9e31aff6c7d59efe587474ea6732ae830d48564cbf1f845cc5edc85654e810c11e8749f2b4e3eb20a84062e937596cf35a00b6f80b4a96636a113;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db9ffb1abdedb541b2b57260fb2955e708c2e13b811094a2b5f347ac6430c295b89e274dc5fd49a4bd61930f8be9df4ef74a367c27efa7d0671dbc54dacdb48985b18cccfe42547cefcd11df32045f572bfc683ca4b14d89f515ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4a7477d38b7fae30d27d0b66320b53abdccde748e15b187b918a24cf59c69ced5fa1b9c22ca2a8b20e5473dd34e22bf8a0b63da59adf8ad7094a4294eeee93fe62d53154ef3793e477911b3235394bedbc9411c3cdf8d6e4c5a5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf0c3982e3eb61c0046ef32efee035096f369f68f9b2d7e9c77721c07a3d2034ab3239c883c0e91bba976873c1c8e9b61a4ffc8de87aa1c47cb628db50497c36d72f4ccd722c384b187445640e0f51b2a19bbc9b719ead5e6b45a57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h139361cef01f3f0ea901329cbd138dc69c149ea8c78cca10c968891310d363c42095c35ea373cf9c6e98123215aebd4b7c9c33c8d47fffdbf06689061ea68e0e5a0a3f684e2b8985f80d971e7dda86c00e4ab5340190d48ac2ddc1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c423c4d075ad71385986b6b65e1dcfcdfe83940e4735eab1edb7d4abcec25efd86a9d6b2114540ac840feb973254dfbad527fef4803b03b7a2f7d9d4265ad4c6ada843b7a776f95f86292f0ecc4a37776fb71cf140745988765bcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa3f123bbd6c0e052b8c3e7f73608c29109ee84a40229d7027917b8b2c0d8e5d35886069e27ef52f048d89c64c48401fd837ae7aa0dd3b19a545c0264dae3a1ed9ac3067148ec1acbaac54fa63d8fede9ca08c52526d43ae50ffe0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h894814ec98f4422364a39bdb4a3b58e67506cc8dc9dc69fd400c97d130591fc1a28caf2d4f21ed1b652d451afe88130b2b867627deda1867edc5cc4af19abd31bb7220cdef5c5763bac6ee55a7625acb601c2a33a763a3497225d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h132c4a75fbb1ef6f9d402a3c2910bde033365c66e26bb5230428f16227c577260eee862db1c2484792b08c8d25349fa178ecdaf43c96c39cce8bd61122a22dd644a1ce93b9a69edd48ecf54803138b3316139775fbdb6c35a75194c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e6fced63832f8b4f3104a59d208d18dcd0d09a9ba58efc057781dc4f9a1095a792bfc822d3b4cad61f8138b661fa9c4912d14cc46228c01e9ce5994940cdfe01e0ef2ca7022b2659d20027a8cc728273e34199a6953ce4086b15c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab0beec683a785ee30e4315a8aa5322cf4b61dc702c126404c39738a2df853a72655ce9378e66a83f04caf37a0f513f1b946de877c9b11d2d00cb8406864ed19b9ad76b9f4db96441e80ebfe3c0cab65ce5729875125e87a06d2d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7ed2ba8f7a271c900de16a94b6ce81e386830f48b96ebc00fb61ae077e0bef9512663236fdf25c4c58284ae04256075852b184c7738c25232e529d53578d4e5d3ccfcd6a929b8aa04c6b613bc6f50cccc0c59198ccf5b3f6677b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h159783930ecff5c93a4c0a0e989f85f95f6e8853d5dcf26b35a6071abed4e302c148d481ae1b53f60e9e59a3adeef42c8814e7476201daf1bfa0761bfb42e5b815729dcbae8c631b47e666273b03ef3915e3a936c70f4cb7f9b635a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eec49f566865b21115bd17f5fac8b9a54f04f1b0542714961401a3701f4f341c3ff0c36551827ddfc138c6155db89948753b790e0586e2bea2f22a56926d3f6ac3e14b75d2c476a19746c65bc63a238dc70bdaa59cbf637efac875;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95171a25c172d25790e64fc7faa8e601e0e8fe2bda9bce2da5769a1811ddf1f744f38d455ee6764d9ff407a98cde796b9b55030927583f08dfb0be07c809d4ea5690b3e3478603311fcf667d1962389f56672d75018b9c12e475c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b6039590bc6d8b8ed07b3eefab382926ea8071943868f2bfb90b11aaede69f3e3514e7ddba064c29482b78c460eb6d87b3e115c62a2f97b439ea24ce8c5508fd57ee4b5163ec9a963c4f8f11bd23b43f5143b967ca1f673bc68f05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h430b366f8a867f61e0f261ea4ea47aadd5df4add61f31c1cfcb4639d6ccf1b88f9de935fdebad16ab068b35eb81efa6926c038a8fa92ef8d112a7ed9af23ce7635b60935704055abe696c1e8fe10c9bb996bc65ea1e728bc34692b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h132b405c3fb924b66972bdd8f9a7a80494a4a7c4837f13c4a297d1df97a9e276e3c414cd2f21ea61884ecfdd50481df0df5971384b5dd5051ae4b6ff4f4acda53383720edbeb889c66759a2c0dd9559a1657c40b3695dc349e6d7b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h140fbb8ad1e0df7b21ba5d5c871b647eb2932a12e3e7dd688375b01fc09dbbae3c9442467fb3831c678a5673ba31fb4e62da8b3685eea81fefffa14649bd9619d2da07cd714783b6e1e167730684f262727fce5c177a6f209828768;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h448e95bd2b018c40cee213e62815e81adb25029348adfe7bda6610d081a72541d2ba95b96c076fa944fdf650047300d58a400f5430a29ccb4a23085937997277cf60b903ad064fcf4a5a14b0909ded4311f36f50e084537b1ee299;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8aac7cdd0f07bdc325b12f3e836ec0f3d459e98014fb8cba09c6e3284d561101b51e69ebd8c9221cadf3c5938e5d7d90c2c0d371e73bc8fbddbe212cd911472c76999749a2d2c61f164dda3a9d8e858a42377e02ea9ba20d24a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c01a87ae01ac6f5b37f2993463bb224f6c13f7f288bff5023da347fcb3250115adbbabe71b6b21c59b1114d762f65570e0cc831fd41aa2ce69575924b0c988b972f83559005ef967942f9106fd96953f6554adaa95141727e8de6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1679aff30f296340ffa9e9d0b6c777b9de8faed5169eeb53783294a39efc4d53852c1a8cc7bd2bc52efad57220ff0bb4a7646e659c83be05de8d3d738bc7a90ce1d81432cbc1d6272ca62e76dc3ff7456361cc32e0d8f3e90ec5ddb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9593a0b1ebf27e77f9311ba8c82a8150207280acbf7d0ee9d683fb313361cc3f588ab7049646cf86acb1c9396fa23675a8ecdbbb7daa69159ed40c6548b35fbf18a1f66cda844ff7f7bf39f3853349fa29094db83cecc64c11887;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h132dc4728397420a3d2bb6c1572838f93dfcaf2ac8fc03786c2671556f301c8f01e08962d38d12d8c881203924ec7fea5991e7a925a3cb84b69e2815bc075e222b4106f01b90ff8cbcd90b93f0a767bf59c19e4edd42c04eb444a20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he00c65ccfc4e09cd7d74c18a2d28de258d3e450c266176c7a32f9c3ee72c6a976d649174c421fb3d6f68a6bef2db0ecf3ccc3f6f752972a3bccf9be24860c12979058ff04b5dc703f1005747af9a37a8d27fdc32d71181e90f4e64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h21aaa172b6006638bff12acec1c0193e0eca75a1c3c4fec4071a684372518344a3b79927850da46c176c56b5063053079c3e980663e17ca7676419c8cea4e7faa414f4a5214bce1ab708ffb42b31faacb90719e2010fc1b32a5ed0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a3e6ad231466522ef128f299ea3a76512b78764685bc5f1473c3aab4e22924f3b45ba09b5478bca8b16cc27453ec4c541a26bfec8d7bc7a63c062ff84724d1140aeb7da58b83be7f3803fa6f5a5b6e30ba7f4935508ddb95e8cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4cf4341701a9b947c1ad57158376da0cc1e481552a380c2265b784d8c4d1e4cd0c6d2e39c3ca2798a41f5548e0ae07ff9b7422f6a8a180417a7f9c18b76a9fc982928f0d80f2c476f7ee44af8e20df576fc6abe5bdc89b51afd98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1327c833586ee200454c9505fa3c257b3fe66c482e55e111b441dddd0edea52628d4bbb7014e73c497e6f6726d7c1f4f2778f174ea59e01f4ac1a85c20c41a4bc5e39c97e65314cf3c988ca5666ea7ab27cb05c2877e80560ca39b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h117bc86ee62b64c96a773222b511e2dfb6c54b28b0a8666c29c920da66a039ecbb25cdd97c49b4ca443872437b154f3ab9c5993610bde551f4015fab0c6155171e517dce81cb8b9fc08af56f2844f4fe919d3d062861258121797d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173c70ec9c90e5b4dcb77dbe4bbba16250e57646850fb2494ab9d6f080d5d302cdf2ee55936f9f489cfa0aefb60262195ff3f73a3d12596041ab0b4afe9335d8fd2809a4e1b7e93ab4dafb8df80a81fe077c0d257c6051b734fd622;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195980aa50e3b054db88a2d7fa39a022654783d2f50f1f52c8cb28f3d58e29263acc79ade925b8c9288d53aff22ab57c3601be3c21b7d1f4b6428ea376c1b12d80362e1a9fbe6da6f381ab6553b394d67f11c94ea086f366f7a7f06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he3228abe8e3baf99c6d4c209088224cdc9b60a4131c094399f252060d97e5c82290b0295aecba903c1a2b1295af5fe08f8ad6e16bc61adb4474a947e1dae9304f160b7bca54ef8eabf365b7547d81c00ae0ecb4d6ebfbf639e5db9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ec2ff155088919f6baab774c091156d13cc19c79f32d70942e282bb4be7a9163a60ddb262b045dcfcdebf60a03508d798ea938c0b80c488756f0a6e283530be2b5bb7a705f4da7abac21ad7ee7bf91c62dd161ceb8bb99e9552d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1999bb5622f3d296fffcd7958536451187aa52e58a220f01e2fcf4219c702764bb0c133a82514f39b5bc27f2b834bf3e84a806afdd2d1968e212925b57bed2667e92fe5c8507b2fae360ac7c781e8f43f31ee1893218879a8183a3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hccf184aa4ca320d19735e655d6e35e3c85af81b289f0aec6b4a87ba3d27a4d7d29b4548ae333cef9a913bc64c4127a72ace09f8aa9b0b3257b37682c8f2e9e0a63f2a3a760fb3b3c19a7c50d97c3c443cfc9959b302f0e3feadaf7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7bc8fa6675c7cea73e77b0822f68b1c4204a986e65f0b41f31583d573c08e67542bd37cfb93dfc8b26525efd2cb3c314d455a817ea9024a1daeaf5ac286b75d6c98e93b4886cec025231ee81fa8eeb3c6eff73bd23b197066ec555;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fc1fc1af1a61306bd9664da985761ccf6dcc81a6b04574fd6231f82ad88d6ef22e9d78cd6645c240fdd38f31a2c89319363444a4288187526f03fbc92b1a1d26c92f7535e49569e9e5a453bc40da7d9d42b02fa87fa0c5d35144b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbdc4299ffa751bfa52cb2f57d469c985b99c578ddf6516b9824cdcd6ff641d4d829278c67b3b0031a9a4c4a5d8cd2f4a28a80327824f619f326c49ee98a03d17016b55ab16f4bd439dd0ed39f0375dc657bcf1001d3201739c7732;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d6c48346e6921c6e7ca9d616ddb9ced7a206be19f27452ce2c790b7161de7195efef08602fc44deed6a16d3068cc20dfbeb66032a979ff0f5e146b323984ee3421c9e2feb0847595bac57ecf80ff4e0c3e0d317995aea166b6744;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa57a6a5dc8f7a1ff678f7a2c73a6668b4a087c6e8f60e7bfbbedd400ebaf62080843cf006c826b823dc10fad62983964ab21e7923f36c3f7716b19ee2b656e238cf7f7c1b65902b36cba30a6da73cc0c887e98a9a40889a70084f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11138859d68f3aaf28c30e73497da84bf8eb05991addc3b7fdbc5f8a7680f0b65ea0a601dc379061583c3a804c3fcf31d7dd6641e435c14b055f2082240a2211b9ce93cf00f0d1db15dbc133b2c90caa1a07beb92ef90a478f8f6dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef2ceaa106b9acc6f81d67c8d7b3d3bd63a7fa589640cc46e75247ffbc01b27fc18b1c179ee8d619d89d8efd65efd8070a2625addbd52559300a7058d5750c3f6151b17ad23c8f59c6f3b14afa601d562020aad8b67189d4c56646;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha581e4f78a219b5448aff1c8fa9db8dc7bc96772ecfd02ef835c84455cfe7002519cefd6159e76b2241991577d8745a20cf6c19d40cb4e3f01270b12ec07a4d7ab2e417886c09a335b0606c57393bc4bf850adf239dcf409447aa6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0c488012b0e4e0943a1147ed6341333b1ee08d62a07b4a781a8173902efc428030c3d1a362d7792ed9cb4eacbc38428ece81e9541ec9502d15595f0a621e841f9be00d25a0a7b9628d8e3eb870b91c44cac3f7d59893e11a3aac9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd05bcbb616e24398c3bd968734ebb5277afc436bb6b56a781af58878ea227dfb07e9cca649e29c03eb6717b25ea535b2670bb03e1de03aa8626914e78c75cc299011c5583db4d1e142c242f195dcef1b88c6e9b6bac4a45c8f9e80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1508d53cba111a9ea6f122ec3d2c395d63aed10c4aa92b242086df7f2840513c2129d501a28a54114666a014196ca299cff428323e884714a6edfd591234a797d52d89d82a5c9e077c9b1b93763a08c2d5c0cf4eb3f30b10b4f2511;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e345232805ce4fcbd7e4f3f8d68a4a08b49bb9eb7ecdc76305cd2e96cc9c1fc432a0969ed9b88e995bd131819d26735309fe037e497b6e709b9940216cd1783a9fb1298a529ba55f61d949a332e7f20b6277ebdb7b2eee0cbf58c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15de030d01b01f8a5aad03de66f852b3881683dcf63a21de9ee2136c59abd0530aec0c1a9545834873e54e6d4fb5e46f8a1fcf0873788ce08b828f9e787c5921fa5f279ec58a049e8e86ee283777b56b21ac358882af82b35a75245;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182590cb98fa64ace6b90835432695f6630377d0f2a49f06635abad1f52bec46e5e3a3de94a570ba0c6e36cb52f937b6ec5ce39a5b80a2aad4b4d1bb1f1a0d978ec918f9ae1f2fb1884bdd23a2b4be21d81f98e269ea5d52a443541;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9738fe02db82ca3b2ff16aef875e3c79b920961fae1cca9791f21c4d09254a3a2031631d7eb628349322dbed51e2013c6ff7a0ce6621f1757d84aa7479e7b263c0f0e7136c5cf75a690a418472d4121655f0f7be5c2a7f4d33ff18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87e88d28b2fd60bcaaf727f8787aad3f544e6193fa719143b9776289328a5a76cc2ae4185615b15614e211a2a3be61aaceba34ae1e01769aebd469044deb88baafbc53893ab53387b957b87d0e7438af194dcb9659b7f89546511a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7cfa6ae6b99dea482580ac646485db64179f367df8e991f0f234c2f199dd5d409836fe7a61fea0d351375e34bf62a5885d06fe0bca097adec2f935aca05ec0882b22ad7ca767cbef36b5ecf50b44fd295b51711b4b9586d3b59e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158ee15ee3ba84d5ca73dd0ada0735e09003edf43c85b875426373157c10afe2ed301a0973c6372bc78bc74f98fc52238e944b43ff3c9ec949d048b62e36ab2d12b69816673d2a05cd31473a20baf9b84049b99e5933db4026c6d0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb6fc96d240e480db00524aaef965c0e913467a65cf490bd1782a72d2f0cff6fc6fcb6ddac5ce4f436ab4ad56f84fd980e66ef0cc591b1e97922d38b411c8e504f38b8bb3368ff55d72e6e681d7e458aa2aa07ee53d641acfc4908;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a4e7c741f1adf74dedd1125e5fcc4ac404428c375c029e37623a8e99d69d68a239c760761ac09fb8139938f7a8cbc3839c5a09f53428bea22fb5b2628291f4664bbb2ab60dc7189b074ed93ae1f4dc15729d5c9d2cbe2c92e8305;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13211efcabd998588c5e83e1dc76777bb7db87ce927f34c8d09bc44238cd3ce7d9f331df4333e87d6b6c6f7e02daccbfaea0162ce65b116532415459394fdc4683289c658b1ffdbc166930722c849a0c63564595cbf6f75d0e60de3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h952923957b061d31cb5cf46c10ec4939f6c8e6c585913e54b8e8d4043b0b2da00266010b637c602ec7c80be7ed5fc208613bdecace80d35ccfbf016506aee952b1eab2d5ddc5c356a712ebf1cfcf833554fdd36a17146d2e1fe41d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fa6c344d8126b6eee2f4df0e3b87cc5b63f959230cafe82a3038975ed4899e95a59ad8cbcb00cce9e74fb996899ecf65cb9fa401e08848f1c12395367586106c5c155c6d2d4a033ee7967ca3869388bb7e388fd3b574c2c9754b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1761fbbce68723a7e43976006ba1c71a96b284991a71fbd02b27ba65a5a6be8867635541aa3db4456142af7783be631176a05790dcd049aa9ce6fcb4c1a4fc6e24f6d2bc8e9aaaace50b9cf671f5de37506018eb3a7bd4c31ae557f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9f7460f94a5afb45119d5fecdb86d06bbe87d4b2168b7171e77860e899a28b90e9cf895263eedd6e0325538b347752891f25db278bac615be164eb8b183228766fb9361edc3367505f89150ef2a1cb5d373cee2537da9e23f4167;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ac1b2b629322f60a30838430f7cbeadc49f9eae340b340cb70f94d302d8646d3969c9e2bda5d0f99c5dbf2622380893cd121137cadb99ebee2bdeb8310033a3f5aeaa35d333f18d5555993e5f25a47853c9c3b819d846a40dd9ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1419bb72b292333d7c5996c3f232bd9794e1cd6e7fa8d0048522ce7eadfad64aeaf653305e277c2ae47f09916fe9d849f97f18c339b3d453c6cd05ac826e0f7213594ae2565e5d0ee5ee0d9bb85f87b0966d871a42718216ebba91b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb90a7170f4ab3cdf333fed5df87ec580cd4cda3dd52cc928826b6e0931834a83d8a74edc231ee34a3e8ce407ca6816e33b8fc382cdc2459d4368c5e38c9a4f8871a9a8d7b8b63b0e19d2989113f1b8e6e9c596acbf8cd6d2a8f56c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be1ecbc870a950a90fad26a03576dcbaeafcf71ce12b46ab34d6dc2b02939d136b2f0f6a0d3ff33487d2071d872438dd9927219165ac177d9e5f42f54463dd808decd06f99d0ac5de49d362df35468095159e1f2358f718f34e0a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca367c80af0e67b73ffc9270ca8057103b071bd1cf27879157abf6962102e0819604c723aa3f43ddbbba8d0352d0608c1a6f5048bc2c42bc2353b55dc732c42a9f97e3be9984509cdf0c8fd5591a1a87508f2731573750be6a87ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a95d7d28f40d27d904027bed67151d47e8fce01ee8fe604d08394714ee62d424fe3bdc1c0885e1683ba46fd36c8212edc307d6b58a651b98cb826e28112ea4fa0a6f6570668e6f4eeaaaf0989664fec5685d144af9a111baa4aa1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ae71ce221a93e353f88a1c1f09aad24d7949ad94c3aae6fd8640be742ecd771dad4c6d3c660b14f35ff9c8723d5f070aa9a0660c9cbcdca44cc6b81c4842eca558faec2b7ae70331b505d3da00073248b06e86adc90eb35ccd816a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8e649239b6921426974497ea1b2f076c31597d88c7b5baf0eb22ef614e3660e1570f291d8cec94a54a82d6bdb1248a1ba4c6de20904b5c762e048ed01892537d1dd4231d0bb29a5f6c7f79117012609f3ceed9a9950e49d4f6867;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1303255df3ff235c8cb4e41eeccdc1e10b60694b900f05787e1cd8f206f92ea35f7e9b880daa16fe78a84c80aeb427caa5d9b7779aa117e98d23cd844438f6c61723e54e5c85ad2a32d7fb87117f93388d26f3bc5bf7d8f4e1af46e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he54f3de89d0edc5e0446bb42e4e40605f887fdd0408617c0f67291bfda7b8ce015856451386d04ad6fd3bbee3d4f4ff5bb405a909525066a49081d9468947876e8ba2017a46a473c54df9c58b2bb65ca054ee79e872042b05063af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12110c78e17f2ef1e5437fae68c349b9c81565b2c68abbb21c60ba4227e926757ff269d08eec3bebe4b64c8691c744417c87bd630399401d6ddd1b3365f734c99dc39c9e9fff71188a7e2809fd2d1a84d74c2c4b9b3760434a49b97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1027aa3edc8ee505a4e3f82ce00750d22af935fdea695ef30f6b80fb21f9f01fa1b049b17b6cd0f62343abfa913fdba0ca3fc993fb65f0835bfb9bc2ba42b5af51f8db6554f0b9676a5d0911aede9aa6d4d9b1a5f7efada5101fcf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc9974623341a457d2e46a7deae7c6a77f161744b93cfa24784cb92de81b6312a45673dc71044f4153527996dad9fff78fa8a1e5b9783acf703205075a050a55267e067aed6d4da6a9c7aec68311e798c686e5542c5ab1f6ab9b594;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182ada65b7f619d510c45c1164dd8143d5d8a1dcfcc632c48832f3c920ba1aed653b56a8629d8231068254ad408acc74e90985db8b9dad37b6c41430b0d813763ce4990257fc4f9a00091a7205a8fdcfefb43da704242b11fd3673a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h74403d0747320e32ff60a6a3534f35a58b1e64319129fd70ed820a2d3c5d3de902243b78a4a04e8a0453c78a797d8f2d15eed0e604659b0fb402d019eacdcf61314e83054ddfd5fa99fb009269291679fbda821119a4118a9cc6e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f6b37884d7979cd15ae90896078f97d3db122e83688f77d9a6383b82834151b9234bc6ac9dbd1c6609be3efb172b1aad7845991921f0ea9f8139a04824c74c344378a51b736f626c9391ff0e102cf182552a165cfbbb5fdcf2aea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2f77970c52ce1c6850865cfa0973840a29a5f7c44695274ede335be86072a7cd32dd7e3c0214bb8893e556a16736d95d08c44767b8573239c29f29de146cb2b35d04e8ed1fbf755c75fa03d2354990b55e80c0ce969171d4fabe7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bff3b3ed40be26622da0ff0445bbf100f3110d5d1204c84c57db986ee470ec7b0a6e00e79a5601b37dab730d60bee58b9b9d7fc174933f5fe29094b3524ef0c54b983c101a0312b4a105f1a8f40e5745063a34830ca54e7a91090a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f4e567b15d3ed412188b94e1aef9975784ce1b0ee7b19fad70015012de3c8e32fe6650f99777920b73161da77b95e68e1e1dd27858ebf8b8308b8edf49696476ac48105d98e3b646cdfb1b9af553543ed89d2c4da4d6d28df3349;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121e20f10b9d8747520107995420cce5517c42ab7613a760c71cf0156abbb83f5265d39ae818ae8d4dbd6b90e6c2ec1e6677efa11c41fe609fbd3166e5b3d806695e0b58818527c0fc5ac5a149e7719f6a9f09f833d3754df1088b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb77ff70f270faba66ca66d9adb9b69f92aac40a8b5922947d390fe2aa90f763b81a5b80feb79b53395948ae8f66792d48397b31b65eb95f489d222b2aeb0477d103db1301a548b8943efb35e87f25bc444318640592ffd3305b92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27adaf6ffd68329e76445f9bd2e1801ba88b1ef89e55c8e532b15d034e2588572615977be4b4948da7e1d68e977702c53b1094e63cd5ad43ca00194c46cfcd27436562a06c91532bbbe21b2c2e8ce0a69bfadfd264f261147a7add;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f0f22c9442eb26e3d7df8a750cf7b229a2ffde3be3387b27736ea9927ece461ba7c6f989c08d680529e78569390125dc610ef91259923bf9b25607b04dc5a6993ebfe7ae7e1632b1e109175b8fada92aaea8ba578771cbe90b6416;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192255fee388f69717fde4ef92f4f1cddca99e3ef927adb947763f232391d7014f971efc2b076b0f0bd3d0f1d41ec23a9680ebd060f6dc87108d53b6d6acdc26500b7c9006ae7d20d00a5f96bdb25b5f73a6bc830031b0e2e72ccde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd110415a0ad9fda0318301a161ef8cc2157e7d1f60f223bd806b313469005408b04897bb045357d675b0cf3145e3cd068abb948c014655717c57a4cae5577e937edc54104c68cac56a6cd5fce928ea5ed1b4aa1c57ec590460d264;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfaaf207c5001fcadfd1d1942f6bbf9eb40fe670a79eb3c28b1d9bc8c98f1b6bb4e22654e887edf67ea135f488e2eaad1267a7e0f601fbb8b0a9b0f4e319eda2d8db18996d60cb94e98a0feb0a86a287882b7c53b3eae14adae02b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114ccc78f5c1ce5977e6989ebfebb297ebf51c7a715ad0522ee1e45e777a8dfcd948e76642394e95e2736e5ad047411f88cc482693497892ffaf2f66e0b21f99daa864fd95a691e73648f5c17daed5853725d659f33b6510b016b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157896c291163bf4a2b2a251217bb04d0e085bd6d8be9050630acd116346ad795a1b1b979317877aa9b597508907be9571503986bba42adb4b178c8772c27c3f24f6efac11f014c0cae2ef16d8a23541e5d8d62dd8e6b37ffc7c521;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9da994e156110de04c19eafd1af6cbe7b5662b423749fca01b311dcccbd1f35f5e725d9932ac95d9c19556b48ff9d0e4c10ca06274aab1e9f46cff71464421ed70e7711a21abea9edafca69b874ebd106500ff3162c315ad6af36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10303d44a094851130780966ea017c726468f21b1b8101d39206731cfcf11ab48296a209f40bbd7f18158a678935afd54f0a178faf389df7de20124007ef3c655b03d1ff1095f417a8e4a578c7bffce97ffeb4d11587fa1d66e1322;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1740d7aad80ea035580a14f0b1c22bf55ae27e819e9d00b23d8361de40e724563b12661e17d27c7b911530f25039d61135cfdeaa887eec114f88da3fc5fad41d7d05c4693bdda399065efab0b0abd51d4a3cd138fad4f8e8991b083;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2d63e9a76eeaf0f08e4819dd51cda7106e8dfe8ceaafbf631d05be5c26fa0935e5d79c8458db290f4c0a6e07a791196a0653faea6cbe6c3495c8d0aeb5de4c753b5715509feb45de1e558f10cd37beb86e8f8817ed26d71c5fe8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7e6104921f58f43f052ce4ca40510e7f5a6b21fd0a181dab36d734c0cebc855c205e566a028e6689a385150ee78e26fd3e40bf0b1b469f497bc144f26f8656517c5d09e8175fa3fa508858ce9dac9e3ec6dc83509866edb04d72e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdb0e4b1cd802e1b512c31a97d56c8817bcae238fd1a9299061a980c91a73459a63e596d2a3470556e7deb99619e285f9be37abdf2add600dd2369a756bc6ea76ccc11ccad879d674d2f551662f1e8aa36cd57d16f4f1994b6fd5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67f42b6b04872b1db11a3ae04441de3b82aa89b49bb62b18a52fd5c884ed6f36291fb6455498e99756f67253da8592546dd66533b28c032e0919683ada9d34bf0662141e553b31448b1c43597fd73d6d159da6daa2929fe22ce7fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee18f01722e2985ad6c6ec10609eb4e8a5345a4f14cd3f3565785ff24f4a661cd65dc8d8b4db6d0d869ff4e2f5ff4d216e9a845aa3a18c9646efe0ede91ea0b1a4962f73c3a0b36ed40b22d1acb77435782581c1c658a01375e325;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5a58c01d4241c07c9ab57361320c129fc27bf03c0fcaf5672094ddb09999f7ab9d633604f2a6822c8979f3772a26367ea21d05fe7a838b68c8688d3b84109bd2b0494b5e66f4de1e197acb21afa05b6689280723492e924c777e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19349acecf19005625105b3da1f8d509e7ffc63ac20566b9a652329cda22542e02554214c558502055c5b556f86e2d28e2beb2a95ee0bf588e6d7e04f98cf068bc90cf03105101359b2e741df1a20e91061fb6c21c44a987ddd4f65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b6e9f0a5ac92d65a5c5a4d4d6a1200677491e49d0645452a7367c451b0ad2d06866f440fea0415a64e0fa2c107a631200221b249a37f5304f3efa85c6eeb006b3dcd968a3f99966062d9379ed73127dfdf83c584df60c2033f93a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58755afbdad35eb89a6d2806ff9764474d7d1b5377d1803b41a148b0a24fa9d20842b485ceac4c9aca9a5fb6651ba6fb11b9a16030a88ce1ebaafabb88c4acb67f286b6482bc7c382a98a7371d55d7fbe7fc34ae81c6126ed9afd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c134bdb8b28263f7e22a474252c3d29d34f79fef44d51591492bd98ff55acfd9105d2339c5bdf7b374af32e025bda1db88e9b847eb7300e33eb000b1bbaf322fb26a2943421a89a0eb06f2b346a59141065319e63f0ad72077bd74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1371434b78c1898e9481eba1b144376e1cffd18e76ebc8c418b973faec1c42746c586ae9bdfc44634d0d8a1d654c4110ecd52e0e1b6ada852466000a68dbf5bb3daa1b5a40d1868cf877898b25525ed83b288af7e10f851471f3740;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6665ca7130b8e968d85e93b8187e0692d88457fc8cd9902fd7c79c2b09755d55df37f884b73e9b263bdb3ff5e7cdbc5798df29c1ae170cae7ca508b2c42e701282e0b073f4549d6be24cb8a18ae38ff24762a43c096ee77873f5eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1021f11872dcdc8a30cdc01ea78f8285fda0b15e2da24e33a5eab28da01f4cb62db9dbed56c3e8566638603cdcb9e8fa642ed6f0ff16e6749868caa5efc67a6cb7b1b72ebd1295b0d1df86144558a3f77f7a59a67c4efc165715d24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14976265da8945b34f878365e5a9b5d0ae68736056952f658963d2cf7ab26a3ad79cf7ac06a1c9365ddba81560c1543634d36a23cbd554a101a39f46661595fc52035a2c40d8f44d710e9ba06dcbf7443a4f1c23c9c760d09d74c09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3073f9e267f54d094492f55dc01edf416924ff528cbbda9e3ffda1236abcff944b0e7468b62279a7a51882cd3ade79516eccb55dcc1ecd14ca682dbb62d216389d1140eb1897cf38240e232105230e4b30c393c53a6bdf887266f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f4d25d9f88921032a26dd90bfe855f59f2a4b33664a0eda9e69d207e6d4c34f0b4f9d495402093bec34edc0188a71f76f586f2c4edd6c6eb76629add9154e49dd257f5e875824c885605c31ad6732cc1f2062b1de6229902cff180;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4c8cab8df24b58733e1c7c24c2a1b4e019a43f51bc00f2ccb8371c2c1d976708b0323561efbc22a3fd72fe4b4eec0a1d74e52ae23e5efbd64e1df85845603307df1cedd5619fba6766d0556baa8617c277e5ea6bdbae5a8478965;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d65c871515025d37979b82b3bcba0e4e9f88a58c408dce817c5c7b7cabbde34f7ea3959b48ed318f8fefafd47dc2b7735d7ae56da59e84f4fa2e64945a3ff185f38639a2cb0040ceea1f9db310830dc486f2ebc3713bda1055f5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1898e970a20cabdf5dbc8f32c438c9a4851d05d71019bf1bba4dc617d2df041ca09b094722826cd3ee44414672b0e506c7e9cf0b5e3548eeded0f6cf2cec3e4c36185813fb26021802751bf392607cd926fb8c851cfa29d9b77e862;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16dbbdfeaa756cb9be813ba3340eedbf3906af26215ead73ec1860927df58de326c61b8b9cd2ccc3f2f487418b8941dd60c2fb5bed17d12616dd50ff977f2a3ddd7040caef99e8c624b56fec2b6fa0c083f06835f54331a0c9dd53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16cd09c8f6769c685ad2554da9262c7708ddc2050a44d056ef65876a5db83ef2c60c50f2c09b5abf253a41d58d4f0b8236f8b5e727c634f695e4fb7b6fc0868564e582c6e52457c0ed7b6da904129a1c5dcafcd564006ec7c566d1c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d58262678fb3dd711dc7d1b46904f24174c73f1b8b8cfb7dc6bb00b9b79a4eac2084e4e73977b751d9cdb673006c5fc914cb9f049f7a7b3fd3173c5b61c81ef86154dfeaf36fb478791d02bf8ce8a8021de40ddb0e244f48ad9a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e17b75f836ba8050aaa63435d09b71d3a7393e47a2a00d5fed138e95e123a1ae13497cd6edae7e8e50d1912795b20a40efc0cce1b48b01d1477a8afa5589b2416aa862e4f80f87649e7583be81bfe85115c731859d57cdd367845;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1255f453ce278c7dc04f6d2dd696352c2327d076653766607a3e5e1a0a4f1346720887c8896e03939d51dd3b6bfaccaab443b6c1f44cf1ad2e7f8f0ee92436cc2d16988e7c2b36e12529a82ccd365561aa73ff57abbd481a728ff59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be346b713143eb985142ac7077fd9a290a29dff8affd8f9ffbb7c84a56a75d6770f0f8bd8d92721d8b3cfe8b24244f35daa59b71faaf4f651dc2b55943656ae82371adb23bdf74c93c65f190038027fb8dc704cf4df0293802d10f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ed30777eee5daf09b228894da641bc22d96429c6d5d8f43d41b0df5fdb6fd5e9266e0cb8948a5004fa3c08e3d4749543c99880d2a6e29c1d3987a2813cfee714ec6bd891276de0b27cfee2b4dd18b341154e1dfa915f0db58439c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4dad8c79d7e08d612561202ab9c9f69761e55e0df9b5dd7ebdd743289b93706d2d3ccbf8178f11d486f5bbbe37fceb79a1570d1fa5c557f4ba195430b30108beb8dc08bdd95c84505532808151e0ebdc5a140a21d2a672395199c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6f32299c0d35c8d5880a93597195f35170c75739adb7f8029179fa19bb057a462d13faad9f5f9690b1c5bda638c583fa1d29ea8287c20ccd1086e5a75eb1d471d6d18c12f4c35f36ff307154b8a2a765be49ccfa2adff5aaff1dfb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc21f1f87dac584638dd1e96805624f33afe009cf97167f74c9e321df4ea1b941a80c123bd2cc743ae436f5320bd38e3f17cd2fe23ce8248dbb1889aa5150ba8566a9c4dc6afe48d274ec400f9350984869da99f15a7250fd7ef311;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107fa49f03556509946e581acf02a6b49e8ade57c7a4b5c70acb30a2ffc26c79071c586563e86cf4f0e045832f3666eb94fc43f92cd07643c1aebaa4f8c7f331a32391a47c08419e986f777a98e2dcda6db3769560aaac38f3f416a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4ed14b89706bb36ef35205996acb1c238268cf994150281475147320d413eaa69a507ef21caac082a55b8248d3154bf6c4cfc1917aa6873a1f12c531e5b6708823b3158c2397255e1ed1ad4268a7689cf7c89eaf13791daf0af48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1127fa7faa89bf6bd8c76aff649d9604ca6e1ed680ab5a91239eac75f64e8dcf783a128e244c827f3afcb601b6f2c91e21b644ed0c51024ea9fe62029de00f6f41c80a4f0be8cc00c330d7fca36dd95eb79acb0559f6f486c4c00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa603f58cfd92db866cf0ecbe5e947c2cea0262f8843d33296394349de237be2ccfa004df0829d92a360067376b15c112a026bede90eafc60dcabe40bab2e5c94d72f9ff0b002285201e62c7dd076c54fbb43303e1967facd2bb91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c01b28fd4f8de8a579450187893813338b5578d9b99f61dad4dd568d1203790672ea6b39327944383da80b750d11208a8ee40bc3c8933bec5427112519ad89411a869f3788feeb275b06949db9bc6b18c3b7a91a10ceaee8ab226;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38fcc62a272a2f8156aa5c8ca826b440b949d99071c331c44c421b4657e969d38b714bdc978e57e86928bfb934e2d142eb91d6b34bcbba7c80b8bd749ab7777d42c4adc33e7643c45e32db2e855769e4ef0e49123416b3c0e1f7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7517dd063b503fca55a1c2b1f101971942ce2a4e4a62341d331cc26080d15cdb150566b5c1e0c4c81f7eeb108fd803bda9b7fe6d8b8757fe2c90c9d56b1d38c4ceb0dbae39854e3d737347778770ea5db3cefa97b217018b54e13a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h55db8a24d2a1b4b2d38b928a200da319d1bf7deaaa096420e256bad40522c5d02a7c2546d5e9a9b4d3ce41ea4b5b4feb2e5122864cc29ae607a070ba7786a5672f4a4fe8eef26a657e7dbb3720ec9d6312a55ce57646c5b5b0673b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7424286874a0db7d23fee09947ca6262a1da5cce47277d342416d6dee232ddb7a2fce370d0e928877231c1ebfe9fc863e5286f9cc58fb9d64856921a635cf43096a3e4018c18cfd64c25ef98d20f27e9d6eaf2234a490e49a2e1b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ce8eaffd3b49fe17265d7b7d88de290158ddf3f6bf0f5b5938b5dc1f849afc958a9923ee9357c02ed0404d51364124dea1fb27bd5ece4b5c20e82e2eb0d0e39e031173f26347bd34e2533869143d51ea58ca13ca646559daad30d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9bc5848100c244bc0f60f3275de8cc1287715773eef7bfbd1126e64c77379ef8b29c668208ce3313decec1652a48f33f4cf972f59ec4c921c1acb7c5a69ff91fd4a7bfcd6d927c53403d2faa252f8e5452728d79d8549bb8e24e74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182f914eb39a6a2d2d7cf1b6bb789859a7fa53f9a9afabeeb53e266126f2737b6475cd542fb619dd521c9e51bc8bba0801713a8507aa53cc266956af9abbeb9b9340fdf33bf752f82c5e1737346b19de06aad19b79229a3378b05b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da42db9056394018889641f7850f630efded0af5ee84133eee63a253c9ef22909ed362eb3434b687ebbd20e262e62f552ed9c4f63f97151c2a7d64fbe6cae3fe4ca751add85eb17beb8ee628dbba650a2b47a3fe7adb3b244070b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41bf691b78a867c7d4c4c73af8ddab4a41c1bf854558e9f53388c9875657ddc456df8a81461691b88bf1d107e149d26515b403ce4135611f53c64e912ee4f49c0800b14b550ea78143ecc9355970b4bc728354cada3194c8d966a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h132ff8458c33e499be4da2133573f1197b1852c2008724c2f80f2837d95140b2085dcdbe30ca3e1f321b06960efb13ff08f5046f6f0fbd0595047fd4606a0a22cbefd344906ec5a5cd2cd763073138f84ccc4eea27b8328feb3934;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6861ea3432662d78e3a68934a158cfe2cb0bcdd6026e6120271972719569cd58ded6dad21238ab8a95aa873239b5e62e4fa5b8b200410cb5b47c3dafee33ea8d57a98db9a88547d8fbac19517f5f7c5ecca0fee85d6396a45a6496;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff6ec35e4a4c20bcf85fc76a5479f0e67c4dae2c78d1870226de4b641c3326ff89caa0cf3cb6ad69ecd48e2950f50f72546fa4b81e29e82f485e73635b30b16d5f16d4c87923271839fc7d698ab354caca3e2bc78d21b752f08dc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1809b23cabf1b3eb1e9a9ae278fc932e7a220c04ebe04b3f04926ee54bdd8a6ef146cc08e97737c1fdbb2abde275794d6e89928646cef3342a526ec042b877cd7a49520f0de592b7cd86aff4936072d0d0a408e51bcc204d24efbc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9b64eb44b9e0fac02ac50fd9815fb195fac1e8a7e4db031ab3ef2368cb1aaec73a89e1f4245ebb9f35867531327e7fbbd211ccb27ac9a66011e3fb9a9c3d20e2a3d5ba1f66f1ee8b5ebd1480cdc0c1711be36c77f442cedb70eac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c940d7db6a30d870d45a5881a9d17c1b8def2e70ffceaa11664483465d8cc5e046c474373c60c08193a2fba90a4392770082f7f6d686a73fe92e83bb6ccdac4a43b2abf8c8dcbf9b52cb3a0f3bbb04900528c91fdcb4b920dc1fd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167b45eaccfe8e81ec3e557ccf4b3ad57d0ece1186d7236834b90b9c4cab29d0a72621a934370484d739a2bc16f846c42f6ae8f1a35d6f718c78c01f21725f0c53f2297d0b5d993a7d3e913cc9ce485faca3c59f21e9a1ccb5e3430;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bbdfb45eab3ae0a7125efdd5d10a5199d867426b21cad10381bcac465b5b43ab8e2bd47673f1cce74daf56a81037a16c0f7a5593555b2da40523574f22ccbaf4172079986f2f7abf09671e5004322e9b0b1b5542951f111c4d516d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6ae1dee7679bb467fccfbe09fa3b833b8bb0d69b42d5cd3ed163b16f1dfdca3609ada95079f1f9a35aaf5ae85cbb4650a8aca15a9b8d74c4d79a4a99be004f1d972a621946bcec851b8b68d8012d52f0eee9597bca3fb6d0eb8d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143f827326697825abd064bc8a64544c59d793cdf75212481dd7b8ad7d82ba37a924463bc6fb4e5b2f292b8f4d2d842ebfbe9af2add7c5c4608d08c67329b31b7283fbeede3b4c785b4e4e68b3d59a16e17fa708ea9cef2c42ef911;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18ab809c4e1ed89600766fe08f58550807576c3c1e29fc80f72adcd37b5a576722e528cd516e9aea65fdb665f64b2ba0cbbbba9baca96d29e77843173139a209b2683c4134ca4c973439025c2b45c1bf3ab007912c4a11c29a1afcc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1693c33b4da79bd72d725493881b0943037da46fb4d24e2cad98ecd18652f5dc479676cfdc18532f8686d236638bc50e92bb5a2a96277865c1602323f8b7d30a61f699c14c788a7f2d20f8028b0ff5efc6096c581b754d9412c8392;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a42b1239c40d0f1c0cd12a7dcabda9450ba10f174e2f728df86880e332eda25c7ec11688e8ad269de21d20dca32e5aee1eece01967d419d4179dd5e1b9ce8a8097b841ea52ae72d800a51f9331541e6c1f99895594b4696d8ffd49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c1394d76d0db08c321b96f37d1fe95a460e3c46cb9b117d2f924ea4d7d55b72853f7b4694f521c97acf5bcfd9e11991d4e7ab8c012cf9b07be2a879eb81cbe32977f38b572a6c5b29884bd8fe20f0d4a938b80443436053b669de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1242ef9e6b04dc1142a8b8407a96d9b713786d51e089168a531fb0d14b04d9b5ea55c8477b8eb8099c93dbe7312fac08109db5aec4fdddd7f625a9fa244a1bda85967e84b260bf5cc75817a99847b343edb533065832948742f3c3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha476e95c624412c789b5ab1d45aacc93ff7f2b09aaa9ba986d4805a4789c4546a64df328fcaa0eef0d045cd617161b7c821bfaceb399c94bfec439e6bb6db12e7b311286cd21ddf2078b18e6c5a8a801071cd69787754c6a69666d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1931a655745549b4b3baee2f5f1a5f0de79c55f6a92177312131e469c3fab3e681941e2f8b7baef9e5d776003fdbcc26d0daffb9f5d65f3b20bc257621f56a9e04644c4e9177bc706aa0ab9cffdc472bb7239f426181efe34356bef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb0b313c11ae6d919d1ecb746e35c7482dda13a7e00810f0267c40fff71e4cc5faa732fec2461820ffea18c515421490a8717d023b060a4082893291e932f3c4b2ea7a9b8e704655dcc0f5a3ce8e69b2353c4a32a241e8b0a47de09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95dbd652681e182d84600a6928ad81f61d61186218f3ff367e05650bfda88339a75ef283a1b532711c9cf1b898a21853e32c3dc30b72208ce6fc4abf361c76041d12be35a269ea447ae5f6e8543f5b7d4c9b8835ddebf052e9b26a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1955c484196e2275958106f52d6abd099e17b24bfe164afcd698fe711b1a0ed3a9b2beb322ec189386a55f4701c99805e408c3f058a22dc300b9ec9fbb95ff7fdc28f64b960b25eaa583088ab00e345ce8f0931c2e4c9af78a29cf7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d92a3df7fa1255ad04702c96d48219cd1efce34c6b003008763818372e0a66da7611dbeb9a801727429348c588576345d38b3a53de2bcafc43a26582f8af3b8fe0ebd6762b5c92f5f67b3e27f570b702ebf01628f3fd57e04dc3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had68bd314d607c2a7ddcfd1a5161e2b0ac16ae73b91d2f296100026bad33a0b169aa52c6f15be5dbed433c8380404a1ec9810f54d9dd34a44813a259bfbeb143b572702d7f6d74ab341c56ca2ffe2e42ca4e40c968452fb81ccf9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7496be3fa9e54654eb0c20bc60a6608a3d6568dec129d053522b72332a00591eae68f46d4635a7788f8923412b5519c0147cc8d5d60691eac2e5f32160a9cd4f4e638818b13c0f7383fe9beb63dd3a46559685373b4125a184ae6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c8213b4211264762402076f5d30d652abbe67ee19a7c3cc2fb2dc072d5b5a139076e229f131e5279959ee42936480e259e03ba702b0310c69250c45e4aca285dd8eddc8b1071c0df3c478196c20980995d7b8bbef2c19dfd9a01f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h888d37474a72dae83cad2f502dbf8ed28466f3c7da36e58eacf26f10a7b1f83e42ce79fe5785ee345e51691c7793a591ef1dd609c8f315259feabe0b57a0474e795869265b69f831ec0d35577c8e648cd9f2baa0d3a256c9cd7b88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b56336e8818476c229e484b5290212dc4dab17fc50dce7eae6380b08059596509a350c29548a4558370aba02e915e6e9a2920c4adff71f1a4101d3903dcb5c143d3a59cd5e5d32d5318830bd0ea9ddd6105b5db042234a6cf6a6c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb83ec4da5bea6f9983f85f3808257d2652d7cf0f778926b34fb071cf5fc84e7867623ad9ad66f5e0f41c595400406bf84cf539db78041bb577cfb02aed3ddbdc9794ab607d1003a3b9a4ce1fed54f6ddb0f595cf7fadede516f0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a75becb8b0de9467bd80aacf726d1f88fb66ba705473d69471981fdbb8b3a20ac000e51fc91ccda1c64b8597458a3e7d9a4844e853fc3923d371d12cb38b1a796eec9d10198c27fe6dc6d8edceb322c7e868aba3def3a862e1f255;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf07debd61ecbde4e3fe3e58b548766857bb0593b223b42899314d748b1d59fde182a3e4f34cd6a6e0b6cd75319169c24717d769521e6ab985b3ca6c9b51ec491ac8e90f2fbc01e7c7449befc19da077ebf0f6c50b65a7e87cbccd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2c43b7b679aec0c70de0f29c821ee89d48a0c668e649f587684bd5403dc55b18e9b97395f475683c30d4c3c5529fed7fe6e6554764e7a253711374373a94af5f775c0d300a535d9402d0aa1afc20525d95e84089d65e2a980325f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1653902cae543e1388a29ad7e9c7aee0f856554d6adc9116b74a9c01380bfd9ccd56a863422a58369d666d3c14b12caab67ed92eebff4d2ec74e0c3f970600a137a4c6eb1693705de59ade9885b9fad0ff7568bd5d94a4963d1dd80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c7ed965e992421bdea8e7401dd61d903f185badd7feb75d38c570889ba4a82064477f8e65f340a2e4a3495e3e9b8fccc83430adda89d402e708740528ec763a26e9be32837241c010cfb4a973a56234b337b3f9fa29c80e96e57b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef0dbe132c1978e5d0485a3783fcd81ba274e2a38c6107bd01dbb4835da5cdb51831c3de0649964c8dceddce5f711067ae0b6fc7a9161c35f42561ee64a60289a92b5b5cf40590a46ae0a0850a0ee97f9c42f69769182a7b0a7178;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d2036ba40837a7ae7b5f6cdd29746c797ec92a57aaba21fb83f18f39f2ea8bd18472178c4a044a892f36935c018144d9811bf48c5394a9c204d9be2b68b2e153a54188d58084a67b2ad9e81cafbfa95f1827ec35c3a7b1da57e55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12025888d2c2e10de4fbd4d4f49cc3f1d5e32ece8a717fbe0673a271ed8b8c99f980c73e6ea8221132c327829ba8605741c76962005011782fa43847bb60414483f1bb15be08db44e64760718b58050d380db71eb12da240342430f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c6feb9c5052d5f68e5826649c07567569133f9272d8ee6734e9a5612aaad673a2ec6a9dc1e3f6332902700a1c5bfc2ab30dba36dd2a7e5b2aa7b703b44d313afbab73cc08a262a8186cdc9ae2077ecb90b340eca2f940d011e18f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h74711bb01f19d5157ae323df0f890a091a100f5efb7e2b9e0618f04607a144f755837baabe520478b347161a408d7a14fa1103feef9621b0c97ecdd224edfe535a0337f1052d5132d87cce268fff2aaf7cfa2d078eb2441c405b39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2d3c221b125dc58d7841736d8eb6f1a4b752c9cfe5abd7a2ddcb83c368d51db68d70339480f9abe5aab8083e238425d8958b06387922109e083bafce7fbacc89f8e7fece22fe9d06501c6ee3dbbb22abbd5c14413e96aa5c2ca52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53ff95b2d1fdca8a3bbca64f3019a20e06f1c68e111d29058588829bde19cea1a3d3da57b7dad3f652092ed1e212415ec00bcbcb8146128c98fe5ef7e8f83bd6c32f4e3d654f47930bbb665516d55b8fecd15468380b64d40b47da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176aaa0aad9b1272332c52761593f5637ea9d86e5ef02bb3e021ca02fc9f039ac43f3c821a77930b6e15eee1ef9cd2654765d350bcd4ec326cfbe6909a1b2c9ff1e6f99432a2c04c9c7d8d33423dd27167ed0a7fd2323cceab64af9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17679c21cb7ca0b599252b7802ab16b96e27b93b9c9cbafcba7a69ad32a97de911494a206d38a2a7fbcbadaff0493324773e9653964ff7a58ac0a6a5160ba0891f270cc2fb94bc28c7795a0bd77c88e0672e0df30eb2bd1f2e4f225;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c38390c575cb6c371706180fbc821ba33ceb85e37b4a45c5426b74f8474801631dc2dada895c89cec3eafc17fbc18d088fa3fc064fec66fef9fb216793926bcf6fe0a371b804aa771c375a89ff69e743c7f1bf3776cf6d077da00c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11647848c1f64af0a460400b0f711b35539dadba000d852c16c07d12a8c26a3c2781300d65510517acda80123bf967c69178feb5a9f98367308e96b595247200417a6d87b430eb43b1262df7c19ce804a0c66ef9da4f54c91cc9dab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c11623ee20932e78bccfbcf602c47a321858f5be44020e1d89ab634b083b9a77c0e233452a0f90e2b3530717e18ba71ea108afb60190d7ecc7aa0e9bd2819cdbd9fcd3811c8dbd5ac65bcc5adfeffa999a06e9424373bb8cc8aa0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd74274b3e465991a51343c44be0a9e0614ed5812132df90fe59f6b0620e890932bdcf113d1167cecc28d083ebf837cb9224116352fb17fcb44e309f9d096438c51948e165cc15b5d67ff410ff0ae5360e37cc3b6e0cf1866c4fd45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd46fa3e7137e631028a662c3a261e74826a3af56b92e03065d152f680ce7913b105fb2ba53aee5868562891e3a424d369757931725fa4035518d966916b19a7f9025c07e56c18ecae14df2ca260943eb9f2c3079f577560fe77b20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h132a19fa44e0732bbafd62f6ff98a8448ff0a4ecf3cb78326f951e7d9a84315928cf17cc67c2a5820a861ea1117b268b1185620a00f66b394389bc3ea5022b01f8851a2b58a823fead1f031816eacc386dceb08dc427d38635e3e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7824fe5b78f944408cd319d8812b3d281280e590b9c9a832e7469d40d9a57140be86a1dd0ce7bdfcd1ead8d7e18e5e45d769379453180755283545b068631a6d411dadd10b2cad0f562de3e3146b782ef30043e31772f25a4029;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa5a93df10cb549b7c0f758fa81693c77ef1293d5d919ae485c60b8ab1dedf4935ced30e1190e34bf68a58e9b458d53415868055ece81b02955d52f7d63d1bca5d97e9c6e3e137c952aab6e4355d5160e7cb19d66638ed0d08f156;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e286a343c38c0b81c2f19fa0731ca4228a81c0a16226187fa60600dad11d36059d99b54b17f3895e1c95ed63ff856ef47d1ed75ad2fd718f389c3cd27c8cf299df7f0c474cddc61c41dfff44a91d8fb65ed50e14cb43a3ba10398e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b497f0bd311397b0a58a3f30892d8f19ddbf4a6692cd03fa6fd833f752a4d4085f0e3bb28e35a965d882f6ffeaf56512391c85e580814cf2876338785c432f91586b37a8b38377b978b3408f067a168a7601cd445d2dc01a71893;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1784f3057d9f7c587768ffe788c33fab43dd686f8e51f0fe6b30c196a3d446c719546d55aaddb628863adacfe8f37b69ebd069d7e44e9886ad78d73b42d671e3d435c9a7f1b0f99c7619eae1bc0903cb588dd91575a0a2ac1cbb120;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h487c52f195aaa595c6a64fd7c854e2dd615425cf68c4583f7940cdc82eb2146c4a26192d2b18f9a9ca51a844f81852f1632a0ec0619fc3694bad1cbba2d372aba2b15208933f413e3502ec105a0ec8b1b45d5565310605e1d46ebc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d8bd19710a772f515c6c9c8954ea7a459261d1d01a0f2b59342432d12b9567add8fe85f07e3550b45e8f6e01295fae0e963a83d2995c84ef4984824ce6fa13cfc9989c713fe788a7fa596a6831ae9959f310d41dc65caaa27cacc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf27d1b13c28eca94307c00fc7806c793140b7eb824bb224f93311324518aaeede83af82f9e90f474c0719f1f858d820ebbb9eda026584f097b7c94b4a919cc9cf9d6c5a9b8a3f55c64423e37581e4909572d8f3ef3454ab16e79c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192bfc3f413439b59b8aac5815fb10749d9cd13263b2553280a953d94be179fd7d8c72797a1810dabdf317d29494616edc9db9fdfca8a7354892e4196e0a9089c4dcd4d94001800007c778e80f7b455eb384e8bfe35a89f46abcc41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1978a9160e57d30000324b6924107686c0329c73210857a08f5883dc2e0149438ddb8cafa623a931e2338a1982b8fd7701e5ca23797d07ea5b3ac5849d750cbedf13a82a7216052c5d088c0ebcd8cac104283f852fe246d8b13fe0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c049a427e736e8744acff58f3eae9322e2644639b5582d1ba07b0bd8893e3cb6f40f3ab15370f281d411aeb07849c02d4f86efe7258f5a95ee29ae7c6568725642cb6e4bce7bf54c59602a80823d00749634494777b6df9d79631;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c69370495799cddf56d77bb78d1fbfeeeae609c0cf7bd569ffe77b3ee55d742bb7a98e9bb514b83eece63e593a4aad8303f1e5976306fe51fba3264f9261b09f4121c5c364b8082f373a2cfc333596dd7c687accf2a56c85419459;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2328152f18bbff0f1efb5d2c96c580d9ab7d8f7212e9a7384cbdf409a1acecc88827a5371657c0adb343645f504691983f31ef40e325e600a59c178afce7d4b76f1fb11ededb3b2ba3bc8200fad0518898bb58c262b880a7ba5f80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43538cfb7b625f4f85f56daf6164c581f2089b1303ea6ac4fd30280c64ce448ab8839e6e981bf40505d9127c79d8ae1aca4e2cdd1ec85f8a3df96c1ae8d64ee80bee1e478373f8feea51f3a8da64248af38a8aad021a0ffeea08e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce4a26990d96f98fe91245b66a6040059661305d14b16eefec85214e31fa62084dbd35dff245fa35f03811324e4229e3daa022230c05a18947369db60223df4287f289125f97b5f415178b020d62ec7470409d1010ffb983c4a61d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9f542f7c88ac1b7b5a394a2a02103399065d76ec84a471ad7067bec12d1d75f28c2cd1c8adabab32c536a378bfcd538e7a36f5638765ab25749ad7e786e8c1eb49c6948b25f0541c7cc767fc26b69830e4f74d6c4b1c5e6af5eb3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe69f50401dcac808557fe693648e297bb9b1565a89b98cf6c119899830ed06794737b768f47831cee098b43019817e808ac0c7b2d889115b24b6f5320e0ca2ad226b27cc4b2dbb0d7ba62475d6e445863d44e3469a8f9539d735b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e0071e4f9bebfcba1e7ca5c4b4d537067bf1666bc8b04624cc93f87e2f1ec6e37944cb414c7ea4e068f83ef10596f8261d4ed25baaf37e2379ed832b64736d265c0aa42c02f32d9026f8480328135edc8410ac31b7eea1f450243;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34a467fdc97959f6b44fd2a8b317c3e517f2415ed13dc2f26811d39895749eafecf68e849523130961a9071cc6ac49361040f35562f8cd8c36b65d7987967112840cdd26ebd15e404e11812675ab409dcfe478ed621d473b599411;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af8a25db654ba0525625705bdc00f7ab90cf8e1e7f9929a6cdd920bd15e791fbe54ebe25b17b1c03a4b678e3bc513b07e87421798e115ab404aeafa76309b4a523761fc4ec014a666c5ee521aca368e2109184a8f22c986e5c783b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e5e9cefa31e5d6d12b0a287a881df232798f5c69972c632a0d1cc72735918c66742a93879cb96b51ffa22e5048d024a410c74bfb9555ec202848211c0c7f1c58ed9c9af15b27d9b69fbf87d3bb5bd0304b4e8eef8c7dc40e50b4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h464809bba66ac01f1f4da029673e100d7d7141e5b538828b91d17ae0dff399bb78ab01ec015e219c794c808e0b7fc6de0c4f88591901f60eee4fcd9a09c66a866775e0b0fc015a3c2adf1ddbd56835807c196675c6b56d26875311;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2fad7199614636125cb4627735a63ae8ea71812f8b733f2dc4e2338672492bf96f01d971d516df57115172531238746dca322cd85f617f03d2573de4d92f314c68d043796569135d382b3cfa8d8d809e0dedb6b210042ccc53fdeb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b468e1514e8cb1e3fb5cdfbe80e881c76f810cbe5cbcf7d0b46f0cbef079abfd0c54c8654e6b24ca9293c33559a54cfa144f81a55c7f1d68a00a4864827ad4e7c5353a54ccc6a224e14481221bfcc4ea30e6ef2dad628be0f5f9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b68fb4c0d20b606f4de2b73ec7a1bce3e42cd4c6efface2a53d8f9f1578e718a2a0c7b715d9cfcd813751284bd35dc5927a28ce52d552a5d1f9f4e774c35fd43d2579e045c981b2d6fe7a042967fd94bcc6164d3443458db0309e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdcaf8f76a74529334ec15d75180867d6b6d0214f655acb2646980103ea09a4232a1438b1425f8c1f38cc4ad496fb9f40711d19f0321b0fd977c08466fe978b5a7761df313baddbca49766f399a3bb1e8f3f0bf59325e9d61e52eb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19565b0d294094a146cf24779a00c6ed1b1310f30b833e86b53c0a2499d2e1a25af7b832ad4a5e4d04f2af075144bd562a4ce62cffad70b20fa063e71fb825f83439cc90dded8f50690487a0bc7747010f17dbcf7ca786977cb2422;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d5b33fd3681ea20cbe8457618f46ee34b1b6773350e360e4e46e7468f89dfbaa857b64ae71e97710107e905f47242f2cbafeaaf8f8313383e4627549debfd1c1e7c38d2fccb3c1c5a3026571a2437ba57ad816035d25c323c98705;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13363b2628e098894faf41de823caa0216cfbe39779b1a7428637b84c8ef1a2b6be90b300a16d00c5d29b70a91bfdb2980c9d3b21706e783d9574a332e42110467a0dbff9d7d57419d2a781782398aac958795f670cf45f8e4f298c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h360f80d1d39201d6346371101710983f637680af8ed622010ba74e59cc7c724a0fc68bfb6f0d4f6da5d5b8895fd742e0abc48209ad81228f5faf54c91ef975d38a25df127cfa4cd383f0d138af2238ea220fbff42f3b74b864b4c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca61b07b445c47c9e5a07355aa12f66e34fdeb10a8959f2621c02e7acf43b57be6ee9a5f0010c040319bfbc7fc7f653753530ebbe29f32d63e902e12315c491022d4d3e0e6b01de53650d3a52216d26419645e89c6e10ad4121a74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bce7c0fc625b5c4dca4404e56d651780d20810aca90564e6dfc440b6ef03002509cbe2d494bc46ba6b839fd6b4f1f229d4dceb58cc6ec37acc43c37012c93583897a3d6cd58090625ff573b833b633e0ad0b012e711fa57b22b4b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5476feaf2370e73099555d2359b0d758844340a957768041656cdf570612e5413c7dedeb69fa884f7ef198edc8d60397b4ea1db024900f6c025d3b0f48b30f7104725ce4d2cdf500cbb0bd1fe38625ded50a754c52c66a86ae64a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b42747929e1a876e8666e4f4b49e366d180610680234520c1900ef3be0b2f3b0894501b2158398eb7ff133fa36da7c5c6ed3250e27bede595c6ec5edbe209392b650e6c4448fae5d915956883df1b7b237a59864d2c0b2fbb23e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f62799d2767124b5d9d04f9a7f66754232de340771054d2904def61a04ee8cbaff99a1377622ec2916941edefedbb126594affb75c8a606450c0eab6eb59b4284ddf343315e4b5059f876d4b2035fb6d89e61b5fbd4c6c78f3c94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6a6284e47caaac097842cbffebf45ef1710be4b485f3463d99f2f756103d71b125eec6aa8e410d040034fcb7fc47bc4915bee25225dca1c36e8384e96672369d240a7b57a67b9fc3701252cf0dde51875a3d515aba85b2fd4fca0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab70839fa55d8f4b882a5c92df3e4dcb2776479ba4b3d7e6270dc5d457ce89b43797770a6e1a3f4b401bea98fd636f50867d34efca01ea6652b05440374c7967633c80dc93a7577a3372a3e7844e6df6c7e75202aaa29086912693;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d2a78ccb95cdb972dd13d31d614c3cf40c5e4b8f695497ac7d111e10cafe80114227d3de5cfad20f885c074e165b4ce755b69cf949d21dbe14011df23f10c170a365c13a754e702f2ee22eac8f624d41a89901254372a8fddfcd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d96f0ef7aff00ee3a771bc6eb4bc5b9c6a0e89adcf9b7f38ef8bb3b4870ceb1fe728a6f429509af7522089ac33df2b9e702174a2c24c57c1cc8b48590668d2ce479ba1de614be3addd442030224abd30bbe9dd0578eecdca1cec3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he3fbea5c40102b4321b812927952702b7e5bb02b03d05c8c8a0dd618eb886638e67c2510e1add5154ef6346feba2da93fe7df61dcf6a68dcdce61fa351bc7b94acdb322c6006f521aea71e52ee046a274f42b26eff015377c695c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1577dbe3975a81c39139130f338daf14f3c98878a1a9f0d223f8a3655d1d71a1c347c5510c135558165d736b847a783139faa54d5f6e4100ebc40d45b4b1a2cc2506b014624b2ad25835eb5360ee8d5c50adff585443bfab37b0dea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a07ed130fa3d6e9fa430fff0c073712831394edef0533b1e88ed6f86d4c1f6b88530241b60a8761dc8a8dd39ef95cc5de8105c39d63688406599395dc63d8dd86860b60014c137fc0ffc3b10b5e101f3bb04fc85c800e2b88d448;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90b4371a6951d4f8d1f127ebb56354c56cda677386b484c2f8341da34659ab85b9adeefe718b6b79da816509d7b0b453153e2da4533add797bae6bae71fd1877336b7f99fcbf722104986da13a3f6c18456db6409c921d4d28bbf0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17123b50e939778f4324ada9840f0424f7e4a7ef2d4ea668916452ce6576c81895ca5cc0382a2fed6a97e01d17848da590f467790dc66225051aea6ce22c44557b65eec770fd3ba562eee5ca33cb313bcfe70062ae9bdcc30741cc1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d5d39998781b95cfcc0d579c9d9ca03e4c24deb99ac9cbacd763b6420fdda62f86b7116b0cdb3dc0f9a0b012e84a2d1dd3e848bf1335f56167331822a97d2da8cec6f2e6e71eb6e0d1173b89ca1c846f5a449d2bac25e8e5228b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7dda02baa9e9da6c8c3c72dd219bba09113b9ceb838f550bf0f78e617da4f2a561a1f90949209383af6d5cb8242061360c8006192633ce290d270d6f1038b5a95c98be7983cfe3a4c2452c1daecf2c275650d24d35d0c12b41299;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8ea150ea90893cce4d9e29ad8d0d423542293b046ba63c71749c0590b42f68e2750b379ef6a5381bd1ccf51a975efd72135b29968dccb125bb580e706c4a1dae9347aea613947af51529e3189a075d111fea6adc3a9d3ed20ded2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d5d33febca9be8e341d0e795a27ef743d01bb3066b629629148a636ac1ad69136ebd9f44af77d9a3a5fa4749d8452f5551a653714d10e29f4004ec46d82ebca590437361e4e10bf355be6ca4ca89267d98a1985d2d38ebc100bc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130a555f976566d1ffe25c4921e035c894676682c2e9cf529aab3df7470201f640289cf9990ca170c1c28c169ae09760cdd0e03a8e275e00e14d57edcacf3a6352d470ab6bcb7c3d074e84cb314e48ee4140afbca69004a10cea54;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0bca210ed5407bf8adbd37379e78af2f36f28171b46237ba2af4ae43f2c9ff89c26898bac90ba7c770d81e95319a7de3532b98225da361e7a20fa52fcc6862814a7fc3419f888371892c568dde3b65c8269f8e8109485cf100f4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3fb89a46329545e86667fbfd9026643d1046456fd8a618db6acd24f50d8ccffad3feb3af56251b49bff09e49f163b5fa3db28d9a45a72ed244897d6398e34c04b75c3e7d1c2a8cfe4ff2d792c8ae4772680b28841f6315072df5ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd3a6f2cbc996b55b748cf711d36d82878149d256f8d44d68fa0c870e356edd5157ba9ff1fdd86268c9b18cbbf94a6711ca400fc5e1cb6bfdf37981bb367aaa746821eb23fe5fe207493f7578da10e4bb7e81fc8a6cd8f7e245453;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98f9052822c89e68f9e2055ac0251a2f7b9ce066002874e6373abcfea0af5c2c0b62ffeda57de45d9cc366398fbceb3b50cf1972cdd50892b6cc20776db8f05dd1cd61f2c626f9f5c21f8775861a60ee0a52b1903e7d4406991c35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h763e7226fb34645a7285fc57349416b5cc3b8490d91823b3d27012aab11e942aed42475a0d4a0815e033db0cf413e3d2bee628fdc109044669415e06597d9a95472fea5bb470b8a0a86e920d27c98f68b87cada6cc5e871addd374;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d47f0b41eaa1d76d77227e8b9feab74330d9ddafc1d961fecabd5d1931fdc5841ab4bcbe31b5edefa235e9a8372dcf85c884d42a17fd2a4172a88fc393c6c891e6e9d91202ec6368618570df327824de88e598037c610544d06ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef653adc79fe9a750629987377e226537e89ffe08ce1ecb6e26a094a82a0c633c0cd627fc8db50cda9282abace27ebc829086fa5ba5544fd447428960638277c591b0370881c6d41316da76fd4b3996dbee632e143d2a1ecb1c689;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173f6a8d794fd87503fb289d898ee8cbf86d9c99b118fccd781a67b4c43adcc4fc6a6ac892f2dbfb5905110eda13d9ecb56fea15d8aa5167e0b281983846c93cee7ddde96a36d336a583ecb75a914f4182d8221bfd5ba1d1f4a6e47;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f824aea58f006dd9683c2906da5f4ab2cdfe65d4c5cf5cfedf2b5fefc08a60497ae1ae1cc693b380da3fd9b80a04d4d9832a03ffd4233318d21e45b1c2d509247f434489ed8d24fba6fe8346f2128bb21214b582e24e89cac6bec5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd21a24646fee82b93c143c8c8e97c34b52ddd34e637b04cbfbf2d3312fd4a83462feea677d2ea5cca8afe7c3322895d965becb82d03a8c942f99c0055dca8b0136ee30039d1d5c4f5a3a0a182bbe9f2da3a3ede112831dd1c51957;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13db401bd2103a7bd22d6d9d3f7f8af951c154eb963dcf28f43d3bffbe59ac7ff4d2b3fcc36742ce16201a1710615f9bf60604604bdcb80cf0746699d96ad9dc68e86f731f2a1ecd39ab65c658d845118fc48be858f1f34b5615663;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefb20a4082193bcbbcfc7370639626061e4ef124f163a021fcf66d75a9902584e3a7812b168d28378dba280a778a77ab5608a840d938ea73ee0b709138dfa0377e8c9f542740be0c0d3d35256c6afb12c57273835ae6f93ee37b89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147d79a12e13a15a4ef06150072deba4acd4a4cd12eb27e8ed9f2f991d41f85a2fc81e6bdbe3a0c39de75595d242e47c69a9255565bd8eb6feaef78fcb6b47c8d20f4d7d1f72c06bb5347a68f03bb7fbc5a2a2a504ec20d5c963a9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha0c238d3991eca7138ad1c6d2c1877cfa31f2da389286b255bb85a24d1c8073e95cffcd0ebbdd837dbc0e919f9ab9c05a84e08733f218e3ba7eb7299be8c3fdca271db6996920863d34ffb323a915e546a569c9ada05d7840f9835;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ad1eba8308062f0589e18dd70097bc3e10d1736164a274f954d3b64c8741eee5cd28419e3c91374ca3475cabc775ec658cf5f3744eae233ef08140a8ab50e8362ea0b2b8d8d32cab328313517b046d1972d33f4c34f1e78b24294;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ef93ff1cc601839e647fcf44a66b25b47286b43757faaaae9ead6221048f711ee8ca9095e590171ec3361dc8dccf384607c2361f43edca878a3c5edd45ec5ebffb16722482469bcb49716f73ea37f4124095f7395413df0f64a28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h870ab9a4ea4739149c55a5b02bc5df7e1d06ba9f93faf1a993f83349aa52b807dbb148519398d22689ab8797de7f8558f81ed36823d96b91e75d8906c834a4d00202c7e67b80372d83760b5420787db1bcf622bd3effc6f060f21e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h788b9b76c129f43b676d8fd79201447b810c5deae22bd9a301170bf940b093e6f8a63e1f939ae5baf70b61b0a5446daab4030070156b4f4ca9a3cb67494b94f3a4d85ada6b65889175d654297710cbe323afe5893b893019106a8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea470c61157e46d5aeaa216349f380bf2f3d6b3091155f16737427dedb2224dede01e4d799bdfd034d8f902d30373b1c68b08fa2f12c9ec19487d1afd1209f415cf18d0b5e74b6cb789c158a536dadbaf5f004a9f69c0d7dd40301;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefcf7e580c563bd2adb9b72847c9d87ea5ea50642f42d9bfb96eedf374292897db50241d41eeb0341dfacf01cdd7143b49013f6696e9d3c3dd67eb5ebbcda0ed657e58b4e38628259b4dd2a34be1069518aa723ea2ac5c3a038ca7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ac2c379df099196feb6b7fc025ebcceb02079bba81bba73c1677c2f0556445b34925c9475ad04d9020f75cc6751693081a56eec4c0411aea814bceabd466da5f8ffd0ef868b48091c7e9035919ca0739876cf15194e2aa6c407029;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13186373b89eada22459071788309d42b48dbb465c76fd3e71c4d89e56ffd1bf035a5093ad3a56a0b0c398a7f8ed30bc9bfb634d6e7f5530382e08a7350342b85c520be22db602265a2b64dd8050f6d905a79670d50230fd09efa1c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8dd33cd1f000b2a7b61662d2b83e125f90dbfe138abdef7de1501e9500601437c0a84acd275816fcbb2cc0369475a0ae646ca45490404bf3dd2ed2ad9929d04a35dc47250e10fb5ad9d7456d567ca42ef4dbe4285a561a83a8413d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11715e27453b7c95434ce64500f975be5125402fe855f55e34220f4fb03f08c2e106393c974f8ee2bf269030c9d5b58775208923036392ebeac9eb1eed7a09fee91e579006d231ac935dce6e15b5ce91eada39411e9ccf6fa1637ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd4519a14f6c977bd320dd4e54bdd53e766b7421ad5f9c0504735f7aa5bf6532ac469174740efbe47a3ab9983c573f3bb48865f6407ea0e191471bb79f3486633d98e960c9c57bb0619cb71743680bac44ee5d5d2db2de151e4330b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb522abe7b93aa528400943f61ce848e18e58143193142225832f6c1bf1ecdaeb502abb94d0657587624083a388629669d9aea1c8d3c2fcfc675cabf1387e6b9b589e9de74207fd858c2a30767b808e21bb34054661988308a60981;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a8f3fd99d8c18bde025ff8d87380f044e0f1965648be817b5ab73a10f532b938e1dc0e59ca02d8809ccb56e15a163f9513dfbc7686fdd7ba511819a8d9637067be1f34b3f5ef8d7c5847c8cbfb8063458b7a35c6a374b832bedb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1249cfece08492017ad39e9d30e5dffe6de605995f13f42daa507b5044e53aed1d46c6ec698fe86e7689cc3929aa84e13c1a74bbc996809ecf3f519683b17a3608dc014c59b7036fa1e45e4ab32ce6596bb1041196e5b07c6f3ae7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f861ae1fda6dab243aaaf40d1a8f2b2aca30df290bb96518f576e5c5be5cf46f011dd52b1b68ea48fbaebc767defd3dce29f7d1ff9fc5fcc82e15ce880689dddb8f72faab8dd67b6cb591da2b647bf093d16c51ff796115610982;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d9095cb579c703ba18232cd187c57fdc91abd3d4d9d65cd1c97c584446eeef7d00bea6a290618f2276fcfcda793b30f6faf98985164217f64dd9b044f62c916697de46fbdacd5e91435ba45ddba53ecba57ae16c9c1b1ba8f429c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1afc840bdbea5a26dfd8db25470c7f15a5e252dc4775ec54ed8654b2e82c1decdb1278fdc04a76bae82e8d5910502e1224198e2bb177cd22b587ca67ee86f480c49de08d17d9193f9e83f87bedc4aac6d5eb600f46f719b67c41d03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed2cba96f2e039c04b69d1f3f8d704c56db1de8b3e8c0e9eb2c288d85ed1b49f488ea147764b03af425d6db3c1a1b6b4476572714d3243e16054e3c030e5f7762f24c3fb9f73f121271e100e24e819d8eb26f4c668cb18f16d37fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1077b079207fb164bfb28647fe39380c27cc167ad2dabf8c42e9246145fefdb19df0aa3e46e7d0a0c90c06f157d0c5eb318c80f64ae665567159d44c8645f2f53267e842e73d35518b6abb3e030468f5c9e310aa97f928cad2bff05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a997bd30a4f23b6d2462fce7da6f8629097b19e54b043fb8155d885a2632f5bba2cef30f06500afd496b9bef4188565dc84f4a7b72b698978e08ca4d202540140bfc68cfcc7f9a2cdea33419478de85ba9efc27d5ef8b94f77477c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h640edd91d49495a49ea4c6198713fd534683d6e0e57fa68ee16ea10bba66935772bff512be761bbc04c0ee769e51fe1673b20fe73920443987ebe62079ba0ef3f45132e7df632a0b7d6b9203d4d0f583e8f5056e7755934dd9aaf8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5d8fc80f43a4aea7c88dbf1728a05150610af5dc7bdebdd7819d216f66bac45d63c9efa72027a5da850428c327d38ca49f6ea6b28e8521969e6d3ef3dad726e295adf23a5a069628e3b661341d2a5349497315c8e9a18a6fd4013;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a85d2295a345a10748ff1532fa5b85e323e3da8cd4efa70f9fc381e66e2d4490cf59a543f09dad82c6ea739f3acdf92c5d89dc51d32baa4e13beee0ed75e001262acb39e0f1ed091a8c169302b939c50c9322ae4707a44248527a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h719c41e49166eec7ce61a272aa5c184f87cc0871a1120a5b0907b12d1e2502b0f06513ac64be560cb86c5211124612332296262a2011df874fd20c0531716f77d7eaa14fb302d56a87b8c5aec24f8ec9ba8c15a424ce02253e3d80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb53e922f7a88dd5639e79309e1d2de8012f9d7f55d0659a9deb16af4054428e70e127f87df6dea694d80d336fb4a9e20b3e3cdd708184076faf904ebca7cce26bd5a9422c7875d42a75b7ddd52cda76eb3971f0792cf4cdc09f439;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h553d6f111c6217cef03df67517ed990e0fc7ac8d0df636f8abe73ba5ec182945aca8713e8ea41abed61305f53fd85c34a1e9d66ea0df55d60c74acf1e53675151989bf5b8ef197259ec5b939356a3f30ef54d76ec66e81aedbf76b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18eb25c98253e9e9f30fc0a99f3cf4735f6b88f7b33b04255c0112767a2e776be76d17411e0d89eb445c706dc263a38a38c465afe8d555977567eeb6d5d5d04b6661ecf2c4884435bcd8e7597945825710f3be9668f638b6855e1f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158a6bd31b3ea1934db3e7cad80d631bdd7e3b649fea96e703ad92cbb09ce1f59095d5953a8101f3f30f7df5164280ab878383630e07c97fb6f550ee19d4f907a6151aa450ca64133c61130ff8f3109bc5dbe75b1a39fe2f1118591;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7faff11ecff6f1c6148b0e947708025194f69d00fa13f1fc39e0c5f618222a6c68ab2d2514fa947e830c02858cfc4b3e0242ad6c00cb99ec35d50d9a6da56e9fcfc27cc6153a8cc71f036f46cf8e68cade8be27fac265437b941f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10aef38612cef642abd9ca8f158e55bb0d97ef1c0b27f2bd2a3871f35f3d2154d50be64b9bff38950b9a6736cd876e515c410e1599752381d4bdf97d3ef02b95fab9c98da2b094b2d519405de47d6e3187992f35f553e52bce16fbc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd869bfd4409a90dc1c9c3de77f078d481b3c0efda7c16a0241c27eccf8a76ce09574e15ce01e660c9cd691e10fc4a5d9e8ac8f0627b642637166968613749c410d1f2668932869fb9d17235d63defe6c162db81d555e9cdec192b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1425b17b450071a7a3d6642f4d99ff391ce875eedafa23e0519e08ef4bfaba4c2574cbc2830fe93f7c047a2b4210ed759979a2a25f66c5e7b262a8d273715899a9253322001ae615a9976139fd69e5d3ac49682c78d52b85215aee5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a7079e12f46d0b2423b421aaaa313bc321d2753ce6844c73d5ffdb54d398756deafc597d9b9c79f79239b1f3ecae017d30a7df1966b5209f314d4e9d8775a5f0e65957304a1501f26d82da27e873b4dd6e16ee6da755c1c85e0685;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8411095c97fe4d184463d126f5b8c44bec823900fcc9a7b65190014e52eb8dc9e3124f49410d86e7918aaa89ae25e4dfe1f223699fdcfe7f64f22a25a22f94943436590716b140eda4862259c23954ecd74bac9d6fc6d46cc46a99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda6e7483346fd6d7be35fcfe2bd274bec5cf1b867a6dae7acc6fa38abcb17b477ca5a6306aadc168918f0d8ab663d84ca57dcca0369211e05132e0b99483db81b5749f21066dcd95d1f1406d4b36a7ee036c4fa31f159b20052434;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha80061dc709a5a55ef74b2bc2565fb0ab0bcea01a660890c3cbde69acc83300124732f4be565ab97c537a0f6e3863be2e0ee1ddf713a9f54c6879b9b2832d7e8e952b535ec6db270026d6622e884a4b87802195799cfedfe233290;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1396c3516b4873a7c691063a2e1be94815034bb1b44b7c5eacdf314b713eb01cadfc326f72bbe86430e90239d157133adf06a772f7e43c6902333935f86b985a26b3ee9c613bdce7da22644517f485fe0e1d0a91b64d8518bbc5509;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a461cbc1bfde361467cc9dcf64d56a94ad1e0e196e9d75d75c4a9eac7572433cb2d42461e3165f64f6a210fa84868fd8864794f453b1e4f82c81c3c84215405c4a11b7adbaea03fbf96319bb3b7422c917d57015f8fb5ab4bbcbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha3f3fe2a3a260aa332d55920da965e2955cdd9f3e7f5c048a558bbb68fd89dc6dc7c8b801e7ff0e118d4ce364c9e8bc631b0dbfe9be82b9c84ceb5feeb2e61ed468f39b34b21c66ddb819aa9d403e0f0d7ba6378d88679ffa4b35f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a650c6a89adf280698fb1379afa428b768de55bc7ccf0dbe518447f0736bb85a92313f4a516683de173ed897f948b2d4e9d855bb933f6e2e537fab0a039e97833b23ebc37d79218b9f4ee85bdcf2e2a620bd3f06ac1ab81a848c57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172ca2082d31f1a4d5a3ddf906b69e9874fd0b1bc7be4c31387cafae5a062090499b80c6d736cd16f9b70ce1150f3f308f2001b18a3204c11cacbf59c3ab067d33b15e168bff28093b296004d92d0609703819d2d6433a627a645de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h52a81e768804c05b378e0ec3c6511d06e0e5c41d43bc287106955acf6f9dbd5de3f9d316062366556d74305b5966178108b0439783600491c33174aacebf6e95450218be6c8238827cdfaded106fc2b10b35bf678ecbefb2f59824;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf529faed9fe08c9a828b1a1cb24fd064fed3377ea451d9d286da8ea787449ac515a9182f807b990a1210360717d7dde8bcdf7b634748043b739f5fb9ca9951e00338196bb231c3b509f27972d9e8cfa22c05c13d0a162ca8189568;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f3680893a40098087122a8951dbd4fc954ff3a7ebd0d460fac9d29a555af3c09400ff1aeb69f5f3a16f1ab15e219bf0231c491eb39e7de582172f51e008fe5db613d3d16865d92bb2340c30b5af417f1b12752899c06f55f87ee4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113785d0bb3b0ecec2bf5dadd8cbfa3f5c01670053ba1f7a9f412f62ea8d7fd63e7e412a8b2deda2465f982acd67939aecdfbacc2adde455910fb86aae5444d879d921668a8c7d23ad3b6240b301625cc996112f8217911d594154d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f15e57067112f6b2ad13a2f0a72430833e61154a768ca17ac79b888cf295b678243513bd07102e2fce730d78db76f646ecdb8d1ee5a61a167128fad35508822900e7e48b23e7fb016699519c371c319c9814fb1753bac4b74d884e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c8b06a3ea9715b22ade9d06d6807eb02d3938860213c076f25e1223dda0825ddf1bb712d9cd0e5772d7c4f703e2e541ab7b1a969cad4e9dadec795eefd94153d6cefa79e71071394eaab2a6c91e1ffcb942a5bfc52cae3ef5872c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6777616ab0308771b5b513028aae9396dc951a5e6fb22b6b0fe9e80998acf6e8f3ac14901bd4853259018631e53b7d7c87cda82603b8ea061e20cbf338205653b96e5c6b7921361ec29d5a9d24d4ced75a7c2d8c5f42cd7cba82c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a86b0f5c69a25338ec4a2bbb06c3022775bf7c7f82b62aa6a16d61b5ee4d7a29e49f0aba6d4097248959ee834323b0902df5787e469950caea2db104096a78651f22364c627053b0aceec60af501cbce9520dba4bcdeb41c074ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h102ed7b7f32d17fef7eea88a8e145c3c07bfbdb0882d89e675ced3ad8d79917d8c4678743ab3c55e46991b712e1e8620f52d30a4c5dbea12b32bf6768af9eb18414cb5841abb5188b747a575cdc3fa88980596e5b0fabc6e4aab19d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125799604d25a1c769d7ba5793ac50724302971749214bc2847e2e24bf1039cd7cd2822bd478adb355e665bcf92ec27420985a114730f8002d9e73d5c9c32558a7dad42dc0b994f171d89b93c3371384fa0d9d584c6077639ccac1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c1bf2647b1a8e31642c1d399d838021760cd426c1b43cd7bca47a45ca044b0b8d9489bd8004b788e73cb8e3152fbb5a6f205ea59ccc316944537831c8ec7bc7eb8af6bd7453903e58189ecd980f4471cd1c45a117ea662f310a77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7e985b096b8c7292846da7ad399ced271039fa205a3421590cc8a9e4553ce4194cac2533a55dc7e284236bad0a3c07427f165d32851316c256030d19730e89ca24803b693831bb41c660ccac59ca92be59e26898bdb36853b9642;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a1ae600fcd9165a32182f39b5ac0c76295fce51fee13a59d33132a97236e90a02439a89272ebeec2e65841079b4f43ce7ebdd875d1dd2270503e2a471bf655bb9a4b61c790cd5b4278c96281f01026afe50a3f56a22a2064b9725;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6d82ece720cca07f8eb3c4abf0634bb01d7ef46cfe25c8cdf30ac4fff4978b08596b8243a8d05876d6af8544a9d9fe7d443eb205d9e7cd27290041ecdbdf3ef6d3b67abb7f99b14fc1eb2a763ec811832cc1bd4fec08e471cb40d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h77dca6584c4303d49157bd5cb7ee20556ac66d43832e15381f34536997eafc93c8e1051a151ce3009fa6bb8c9d890ad0fec831e55a5d88f1f6928fd53c964ada0eeded8711918726a43a4e4ca2c6a91be179b7bd2bb161329545d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h372235303a185cff3e13289571873dc5645b4878acbf78631e23dc96a7e4af657585f3657c57853519d37fbba5ff037b405e46e46d8095faae61427dfe7025abd714953ada4e2f2e1dce11426d42dd75f459975bab77fab62e50bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h175aab25ec3e44360d5c409e28f8e634aa39f5771d38435bb16f22ca62fe4659bb2120281793ff08b74e3076508d04e9f46ae0d4354a2f8f5f5ed206b9dbe68a29b2cb4f1077f5979e95eb0462338038b7870685d66faab0b9d699e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0daf215cbb94a06acfcc37ae8ff04dd1fd4132e58797137a298ff53947c4ef683f1d4c02487f0f5ebe5f8b649d86bc3a585fd937f71a683f077d82c4cc5ba525c7315c1612672699378cf226731499af70299898bcc7b4a3d10d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haeb62904ee375ca579e10cbfa5490907d6de5a10c65f5c0fba94c6a6568098f0538eea3dc85a3ef31d38ebeca9fa888cbac035284fbbb1b99bca84ac0c4d66f9769310517e6a2f9e19787c78b3092dd8cb90d4710d747f6a7354bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b7830d5502f1c4ddeea181f5de33a9b8508f328f7289b5195579b58c86c0a95d6056b765cc8b634c87f7494b4e97adbd501609ee842f17b9924598c7dafaa353d58b9194d14b5eb7278124953a4a8c9401ac77d7e336f51d5c007;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6410f1aace0e2ce7807e80969c56967584061547be9941cf6c01981035296c77a3b93d69dcfdbe63c1d2bd2994abfd2e28bce145eb5e917447bda997ac77672c19db1fdc3ee13df45a545ed15e87cbf7908f1a278822f3b96f41c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19cb404b2409ce378c58c0c93a026a032e20966645fa9bff99fe5e2e0dd14a1c39e753282418600cb6c4f64c9c049274c622c4df43b859545dd6b208712845d11824bc53d367dc5bf9044de806c60de706246dd5dac4c9bb73472a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c9f0fdf95baf45006b0506eb8fdea4eeb19fd542d7772e1ef9c9e18baabac90678be8d20bb631c9f007384065b27f6875bff12bf7e1fb676cac4c81941b48bf38a33b20f94e956c407cf75368cc9a5a649c61d98a5ac77c954559;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h92577aa7dbbb44605c7b875e10a4bf48f910994d7acdb006a26bed62c3245c353c4032046ea741480179cf3aa88c3b2ec69f7990de17830a41b68e2e5f761decdf37e35c00287034f19823c1885251f1d0611da0ede079ae32d945;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h888ae059927701aa0fbe51410148b435d30a4bc2b1462c415b4561c6c47baab7cc4c8bb5d275304fff53b89b3e68ec7b481a2f8ca2d268e42faa0966cc21f0f3ac1ce545d5f8c6ef5dbd84b8d80723f279b4fec3cb4552ba222276;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h790f37aa17fff8d6dfff8ee2c5ea679a77db03a96b097cad19510e744c9b590db9693af68139700e41676473543784c21476d017bba594461bdf741f9962a28403db5ef2785d3ce68b3126ead8054135a234caee007cd5b58437bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4e2e06b6754faa8fb305a255534347ab6ef912a98cf6491af0872ab8b5eb87e17965fcb39da5440f5a83dcfbf2213130f6bd4765a64996bc10b6998ef861a6c0e8ac846efe1abcd751e3b96d30e2645019d9736ab36a1969a2f48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7366508c4256c051fc16e269c23a143f576cff6fec51780ae89e03ea85aef2cb162275a14e6867c3452be00b4ff8cfef464d715cdaab91aea21a83492e6df71980f2daa35ea0f9af86aa919ced0d4db6c60e0c15c651fec0d9c7a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h73c6aeb9a16319abeb9088320067bb982c59fdef6f52ed366b57c59bed26cc3d02d460daf2c12090e3b6450c63142281c0ea017200d2abbc92b53d88053addc0a56b4dcb1eed8cac555cebd9ed73b411688e4231a48ca99e5f0cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd56bf665866e18bfea73849bb14c6cffb6648222e3e2f1faef7a6f79e367ff649f1b1da35340c8b6ec7d0d407e0a189706eab4448660f239161ab5dfd649a3f39b0b5f702ed8aacc4fe5f07929370bc3f196ffdfb312e41be4df3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f0114f75fff622b51ea358d34ae3aec11cdedb527b1cf72eddbd0102104e38f6873cd9e69c06949c4a350735e1fe176df126f72402904870069973213a31089598f82660074785baf707e85d724a1f413b082ccfcc9dd90a1a50e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16bf539008e29e9cc37a7b793c2b1a397ae72f8dbc782c03bdcbc9d33dd333faaf2210efd5854892a7519aecc8cda3f18d3db6a36168c86d1b57b7c5e8c7395314aa26b6aaa46205be7829fa13c1ce58157f682c56b25775063acc4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7766c74166146a2060a6b687ae33526c3f6d4b45fbf36c123ec014f635f0489263e50de263f939afab7fbd30e9acdb43d44f793ad5cabf3cd00787836775417fb070364efc1c1de192ad2b408e88ceab7af8e97626aad7a13d4b3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b51ce7151ac59ec8c81180a909eea18e813e3d2d5d09e8270e7ab995351407dd0ebf5999bf098e7f274eafbf863e2aaf390ac1f97c1b8a515df164e0d88a304210c627882a7b2300c31d6c02bc769bcc88385d7f48a5a0f10dc04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70e5c8a58f7433c3c766dad8a0c84cccaff4e162389146b705ee7d76fcb2a635832e8bc57610edf2b1384cd13579b33a8eda2ed0e4cc6158f082f3aed97e6f34749d5b1229ddba3c7237d51f3a298b8853837dec874477f7df3f75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12706ce9ba78ae9adbbf8e062899f80fcda94207d1efdcbb72f292c98f84b3e1d21e7b4bf17f3194db74cd5b96c062192c76b67b3e2c001a0e2adde41de0687dc69e2410a6d207b254f7c79871d5e8e1df277aff1f5fa05ababc86a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe66d91e9ce012ad553824968a8703df661517bd329e4e8d2660bf07a2954c55b9b3f02d77382b1064ed4eec4ddf3e4229beb9cc30f4dd434e2626eb3a821f32a8f14339817509bd57d69be6f6731f62c8f7863fd17b5d860fad46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hace629da0589974a403c840c94cf6cb572ffb6834c8a829512fe852b51c305d3be6ae43633d3132aa0b8b5bb4d2f66daa95b497a22561aea22ab6749e49ab6e9ea9a360db34e38ea423d31a97461553b46856afbf494d2c74b0514;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2efa8d29021043244fc7cf3b64ed62284375277c03b8e1b5744e264a7daebdb41291a0c6714b4fc3ce07a5a8f195f1acf3f1a9e49ee4546ff7c5335f26469da8245f98de71eef12d8acc846fe4d9dfc56b8f2c1cec5b74b19c3b0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b69bbf3db7fe9e9f9d8a510cf2de2eb919239316ce8fac210f88ffa7d8049063e304b4040e5d7bb6af8689fb67a164367ffacc237ace4b9ec9a2001c93984b60db66b31539beb744eade945a1bcffe34b522e21dd2017f5980cc7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe9285dae6bbfc519bfbaa33fa454199b2a504d43a209ce731bbdfb6fdc612c579989cff8818dc8514ce76ebf5d5705c3589472ebfcf8809ce3f2e05ee5be67ed68e9187495b773ed35790d7cc7fb0e3303eb50d838c2efeb31fda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13040b9f191e8317cf95a94f94493faea48a4b67cc5465aa95bd2287f071ef5232d11e36b1fd955e396397098e64b96db323d2cf9a933a28cfc02296029c1b109e20c3fe209c514e25956ec0b37b054ae575ad240a58fbd85c4d1ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c7ab03bf2bce234417c9b767f0088c11f79915610aee66dbe1bdf319640e7f34564c3e2b28ab31f78dec179fcbd4f1c61c3be749e587c6e3a1eb3a6ce73920ff97602b5d80093df37b8314a4c7026d538b07ada2779a99bf71746d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h109a6999119b512745bcae4b3d16aaf0f827f20ba25a54dd37b9bb418995e98a0e0a9eab9d3f4d06beca8fa84a4f87d31b82ef372f2472177698f54110fe08ce85a4bcdae18ea9920e017aab8034351d3b8c69488f96a851826de1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ddff77baa60367281dd0783c36d55229d7705cd045c040556fc777cf12383d440f362bb7ce44dc8b751528d68f7e16cc2549595dbeefefd06e957e370e370d403eb20b8e91be7177f14b106cf2e641f4b96483a50a398c99a3597;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cce3ca9f1485af718b0ad76fe0f37797cc6deb9cedc45e68a3d634cdb13712b3f8d01be44d79218d0d6a853ebbb913a6f17396276f4ecfc1bf684923969c7265248766f9ab98c31eab488101ccfcf6a82ba6a5b985ff5458af750;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hedf0636ae20d7121e9f045b20979ce0c944bc0dd9af417a5f8defd17536b38f84cea2579f6be566233e2513978f8ddd7f451532d9f52cf14fc0f3556075d581311311eaac641a8e7e3610b7d2564a037cc10362459a469c598155;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfb19a6ff3c1fd897b5ea1b31d0bcc6528e59e7b752e4cc4ea09530d40e9e68654a9ef859f3b5f9f2a25b76a9cf18907d31f02bc0d1b65fcd7365db86f8f6821281062a1186e60210e2665531bc81941dd98f29c93881e370c69f7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h151d64c6f8a5027817c2776cf5edd9677cde1599be4de968239617a9165609b9ca36b737fd3771cade8d94d09d89396ee1fc1bcfcdda63bbd6b26b1c42c4cc96ea1ab1f3e7d7a73e26796bbb0e3325551055640e7b235aa642ab21e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h178bf37c1acdae0a8ef8d164b765feee025c173f2ed23d9dcbc42f89af11251f8146f2c8f0823c8509370bb499adc6ba49ee3fcc3d3e3168685915c524cb85972fc36301619b557827057d9346f77693785c1626cb0c0347e93feee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd08381c3dd6b8540d7b437d33dc35563dab55a1a4893578008e40640c357c418dbd21a1de7022c328aa4dc17d9d585a7377cc5bb4bfae12ef63e438077c9f41a44490567ee02bf2ca735bd0ec6149b0dc44488ad5cf2b2bf2c27d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116c0a48f3929e718945b0b307f146d4c321df8c9c444163402e454b83dd24d75ab7f8f9207a39b0744941e8e079ec14ddcdec8d4c0948b1d159e4943f9ab7e96c880c4ec3bc42f3c30a3ddf503c35e7dc3a8f1876f27b6bc54b886;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h77e147991f3d7db57878169daf03d03e0fe615e3cf95c63b0b089b95d8977266dc139fd471495193f6fd799bcd1068607e2a298b681d4f93aac181f16857c51847b2b8d282b061a5ea5e56f92c9639a3a6847e146ac499d1ba3bd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184a11cdbf111b4570c09605a65ad3193c6f1184836cc39187bdedc9615fc0301938e73150a869ed5049423707c7ff3ba10f1f55b32ffdbd761ea1adedfff13423c997fcdcc65c59417d16a482fa0c9fb8000f5f02826c62b0458e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha070f3bc956ccbbf7cf14f81254c0398bb42a3ed26f45199868742a05ae160bb9bb61040b349bbcae8c292fc2bab1cd0585c79de38ed6f5ceb4c085de2f7ff34a881afb727cd251327fbb4b1e0af91864592bcc94603e803e99722;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hafad49621c35b1f6aae14cd8306491bbdea83043fed96481d7e5dd953a3e4b589ee6d9e873c8fa8b12d9bb64d843db8024bb7beaee3514bd3b36f40427a3be1f1f373deb38365af15987b457df7513cf6e7ab98137e2820909dbd6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4faf7d4d0be7c56b2c85ed9ac893d0ce7bcd77b997a45798320ecd8dd1938a170e844cd8c1d25db8d94dbe5ccb7a480f1b2a4a2c04c7b1ac992d28fe95eecc3665e6d00be2d80e324009f22c79c392b78bde9f84f3b76f08c4930c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164aa091f75d8997e2fbd94328a7a701b182ae368fec4c615d58a7e4fffb5ffd24f6e1932f78fd10fcaa4d0930050b4318e5f921d0ab1d134fc3a8384006db8b343e2d819d0dc1fe4e769977ed7325a537b54b8e5619bad488a320a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e240a151f7ee51342c5b9662ed59ae3f5e34520a8326d4031d4ee6047a62e1b408b229f2440d0d093d3d2c87f04eaff7b16b7ce0a588d91464d6e9156ad66d153d49b43d8f4ea72548723fe7e812dc0c220a24c486adec5f8d223b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20d24cc28ae7c7df91a4fecf182ba7438913f95dbf7108b68d478895392b0ba19e3de94570f882f0aa89b0a226fd7bd8096c8cc3fe2498e731947d5ba788d7477155730372def82051fd7df058b1712b7309d1a96c6b5791deca44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4059b4964fc719a18f1bb552f46caae8cfa5003957ffc68f455a190531c240e3dd624aa847bb4198c1b346a38e23e8a6a4a485d7c43d5906772ffca1982faca5162e9ca434ffc328238c19c082104c552ddcb18b7a210d9590db77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1988b32b49577cfca6b70c660aa88e066d896013e751262319668209526464e98054452901d4e51d99b9c8dd7e261f12e087393c7a4102a1efa707f4804d35a1b26a143c01a81f434e05fa37fe5c0dbf1362b4281d43fc94b1ca89e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd0adb8ab5a0cc6dd2a8af179320b1cb7209cbc1e283217241efe2f484f980544d36251aedb6a9e11553f6e0e52b0b4d9922a6a504c749c246a7dc082133dd2ec7239588003046334097a582850dcc579acdcf7c0a9014268ba940;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7e1e894c62c88ad962ebb274c8125c4a971f75e14c7a2b6968041d2e3cdf3a5f01df62feeb5774d237ec858fba12552597007b93e8f57a07f0f059e7737da27c501c36208806fa9836012783c04aeb0068227d056c6ff4a98ba9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164ea0882467493ed5749c0f69558a6b7ea4da384dc154abce7bbaf58cab602991d0a2efe27089816bcdf3f738b2d284de367074c92ff330ca9e1d835e9e45a6596e5a5624da7cc7bbb64db92e32f99f5384921cdc743e11b132eb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h60d69960dbceede7988f98c27619dc69dade49e042204cdf81d4f5774266e9e982f9c99169583c08168ecedebd2012e5f8798091412dfa9fd5f18e2729a6424d2ca9c3293f9d684cf2b78fd8f39f6b97159ab4860d70c29077e7af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177bf7464a4331d2172a2972e95d4c69e39dac9349224cb9781b2c2bcd8e178dce4b77159d93dc330f4f57d502498f1c080d4b5f7f70a20c9c42f8fbe319992a684e1c5280f477dab6681084465de162c001f0674dc6363cc020fec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc4605918d1f6f79177252a8d72e9cd40c3f768b37ef22654d1747c26ae8782efd542ea82bea2cf8978b4052e0dd11732e95a312e465bc839c2cfc278d33da03ddcc19e0ed897dcd00669b009b55a4503e4fadc520f0e253515e59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a883e363b6837c8b8fbacf34dbea4e834106deef974f3970c721beeaaf170d8146da74637aab72adb9fee6895c51b78c6c62d4d09ae4eaae90fd6ab3fed83c6e087642502139cd6a1a9f5c2dbceedccf8894a900d8d38f38b7fe8f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0cf7a2bde42095d87d694640204785f0ed55dcacce7f483c50bb234c0b5f16d30ea6220023265a179e7cc73b3d79c8a4c17478e7188bc74ef5f188be8c965d3c168be706d27bc27ab21242ec32433b79b2f5bab6a57e30a585400;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd08cdc24afb2b53f0e6fadd827c0626e5a257139d9a6406f938715cb0477c040f5385b5cef1cc5711f93dea64bddd7fdbd04166c1bbd8849e945571946b79017604e836761169f41cca29dc3083cb179f8cfea164073378c719620;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1490d40144bdcce211b569c85443af17f218ccb5f2ae2a40d94cc3e319489775b35bc1e37ee990a5ce545e8289284099493bc4e69d2475fa04e6d5e14ec06d3d628e04627302e5bd929ef4856448e996fa32156afe57298252d3252;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d90660b41e1eddb734c03b99747823101870c9fe11c5e3c10d749e0828e48087c8e89b0444ce167abed58acb8ae279a149e5b3590f8c0d16c73ec2e9635fa3de9ea82657c6e43f1ebf1588864c10896cc38a69d925e9919ec88856;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127ea59752a3337a3e4ca1a9f70b749336ccb9211888b3643b23bc5ebc67ba5ca4eaff8b79bfd40a164096260c3520bb52890377544bbac28fe30b2564aca7312f1819526c16200a8eaa0cd93a33ab8efa67e1f2736443cc3f62fc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da3b4afed81cd64de3628fc6d3e7df059767cd658fb24bc4dd3804802ce13f6062e11c2afdf665b64fa3adbb3170604c1bfa753aad378506be433e996d75a23a1a03a86e91bcaf97fd554e85ab10b915599e40cff18968af3c35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e711754778220e85f9999debe93210dc16f30e7193f7f52271d692923adf5773bd3c45dfe30adac92250673994d4e7a387a8e3bbc9fc0eba2d7abd49050b9b5867f823b088ee1855276f26bbd4d96fca5555ee57e2826b4c049e95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e5250aeeefc0f8313ceac30e59b67188b5cedc4903d8eeb8295c53a48e2ab941f76eb03df304ddff8fc42a12021a2c7ca508ecd0a44fa17a3b615ad2977df1d284ec421fba3c6d8b5cdeb3552e5bda322ca31d5336089d73d729;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1df744ba1164b9c99c18609f2bd2dbbd9ce2a5b0630b55600f46486b4ebf2faf12a10edd68cce33c7afb42037f3d0199220e9cbae54595348264a0b30d941a82e8ffd1dc664dab3c514df646675c7e9463b6d1559f01d46f2b1218f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f89cccdfab7d13dd872c35f75c0c28c1127733ba68b79c6ca8acccbd4164fe6db0f7a2d48da9ea65728867c935b99624f8a4b56827ebe8124a5b19bef93e69d70b659c464025f6e760d811d28a647ef4756a2f0a464d5d5c226cec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd607320377617abc47da8773b1daaf3a5c3392681b40dcc2f94cf61dc2f71628a55975c897ea1dec243e0704fbb5d5fe718b4bb3afd3def156b1235d5ae57b00930aa1621c61f652fa6ce1d2e1bf3c420548708ded3e2efc7da69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f27660809d7aa83e93b3217f0e6f63ffd4e1ba965e6a6951b07217aaef99727a99ab3584fbc0604dd0f48592196643955cd80d97aa801b014eee3c23890182b2fbe060010d4348eebdd74d4e2ba548f2141c195ef01da5682c6e31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a067babbbee621a8159feb68b9a892710b0b40c1633c77f059efc54647ed49a85a2a12f905c404b265690c8c4a0882e74ad55c3275088c97acd7f57ecfeb93cdc744271b440f9bc435edc6d04eb9b7fc729c31c80518d84db39af3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h191461b23257ee1aa7d3ea6bfa2b8507fe1f0b26c731d08d7214cae65368243bf415a7b9f493eb98bb97483871fbe248443bb9184056536fe06f407142f89c3e9ca2fb2ccfd19c8ff8012eff65cfa699ec4fcaa8dc9cfda332219f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a1ab58cdbe26984cad7f741f712560b0aacea4873bf707ee683d5ceecd83fd4f106e0f5f78766add79f39284dcaa3c5fbd4b570bb81b496957770a6d61a3cfdabc41d5f45b5b7fa9f1429389a942718c26eeafcdc2df519dcdb38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b1e3b2adfbebc54c72a4efb5f24a62f1845f4b2ae37d2b8d21f47e237e32f39ece5d676d7d68083cf781fda98e603a736c99fe3697c85d7f42d148db2f8323e1c7993159682b3bdb50051f3ada7d68168ed06f98d10c1a2e4e8c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1608e5856535bfee10072d8db74c5213d5b12b166fe8e692f012e21c54319430e76bf892c79973eb43a0121f68cd820c48fe23237f1179b5186cfc6ceac67097c72d9314286f2fbed835d2c44f896eb41e6e30c4b7ec218f5aafaae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f508599c943b8018ea74b34e0808105a075ba461a8f9abd7d31b12a38ffc4f2a2eb4bb909ac179c6b70ccd983e541d1454577ee1cbd0d29809eea6be2d8445501cb868bd41b7e15ecd47ad7239126eee2f4dc11346d986d41135da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4d45d469a0f34adfbfe8c027a30dd97055a21ddd6041739e8757be9d5fe7d089f02da96489accebf1789473a915007e27d1fc49b76c8cad10da1d7a68fb7340646192d4594e4cb11a648a4c5bffac4ba4e018843f8e815a73d79f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83ff7009fe88fe6e42d53bfb2566d8286e01e7ca9c867d9fe8537e5872edcc04957b6c9d1102b61b9dbe173f79e102869524c85b06771cfd5f0a60949ab336dbbf2a63c4ceb4d4f08e3ad9a870902d1e886ec9deb791a2841d9fa7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha91f115622a40db57aabf34011cee2d9e31b93d7562c9d9332a425b9ef331fc3421cf3a8eb436b18d181d9a45d2ef762a289fcf1335517a1df8875cba27d3c716d4f83bc5271fb6ba14382afeef23125a679894df07bb5b40e297c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4cdc4c7a0fcfba3d7b1f4148a68c80fdff1d5c9f6bc1155396340cc34a839a06f0444c95b5171b7a439c42acf60fd5cd155f0df4bf2dffdfbb6f15f6c282dde935bf3fdafe882bf4b4b6165be6f40ad5c902c04afd89dda4c32f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d6a2a1337e2b9deaccb7e0d4d917605bd7b9f63c3658fde2632ac944de3b4260c6392fdbb7ae167e6e3456906dbeae62255fa0ca53471decdbc39be0b91ee00698588f740117dd563badeb160e806955203c56fc21e963214ac0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14932cc726bba91095714d8dde697f4240bfc44309b937d5993ecfd164d63bb04c1a0771b8aca5199a7f4004cdc1b29da1670137d6d4b35d6b43fd1b667def9b5170cf4541516666d1c916a58da2ea0cc5bae1de9366e16145d3699;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd776d7bbac51ca1a47013724763d818521208b2139b2a9864f182f7be9dbb1de33382c9449befe0542a7e452edd73d61d19a7978ef1cd8846126cda40790a5a7b0f43e859784422985df3f3dfb9dfec73bd0875d7106a375761f0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1831f6fbc57ccd4042933db84c07f877e5ef59c82c5d6e81b947af6da4b06ad362d21c426d26c3ba4ccea620744f99c103b5dd3b3d7e26e5a62fdf394a360a5d53a30a8365c3972b596420432fbcb86b636edc12394815f8e07a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7521871617ee20f8f74b7e01879e015216e797a1ac4c60319402944f44cb0bb35cd74d00f04c8543722447a133c1fd330c6231a8088b45f781698eafbbfe6c62f9621ac8db589520abb51369caa7a50107c76645b5471c11259a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce63461771fd7dc601fee5ef036156e57f24858a35125aef72d911e8c29259a25d8ef833ad27768e3a3e4fe0207739c8eb3f043e4ec47c3e18708d797918b39e48dd55ae9065a912af0439cd2258b0829e3c20ceb759d4bb410a4c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h939d57d71b97f55c8a094aa226af8e6613b6ad3940889537caf32d97c6e5fc1567394d2514014fa50005fec7730e25f4403f9630c7d07c13d159e73d0564b245b3d4cba653f9053ac3f8a6fd203900394b93d1bdd448d7b7aa0e22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a441c336d98c30569a875084d6093214b3f411eeb5ecab52ab58c97999c7a44a4e93a71eb9316fb9ff3f3b4e4a18981dfd77e65afb481a07e6899c18425d7c9fd1c75d0f4364ecd2771259820938d28f0fea8e0afdeea211588fd4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16bd7a1f4f914eb6e17ecbbaaf83047937f955288959ce3d0ce9e5807b4a154b9a12fb6d6ba477793a06af56307c0950d693484303c3916b1cf5d09ac67506249c2e90fa9a6c23f835bb21ecf31a60b3b2845ddb33607322ca3379e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd0a6fb0290824da92909666a4e2cdb93119d579dd145af8a24ee780498d1ee5c4c87e3fd89c03f4b85a6bfac631c409292c7d13e1629c0f723053c1beec2e40178bcd0a74c486505320343a06d3e6a3d43e67278fb209a1c96d00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5de838a839654dd802d238162c5cb69810562c8c4cdb3bf5e9fad2583c01fa8e4a7f382ad4140d8b7650ce3cabdb3cea9ec89f7881fc1c40f5f2408491c5372c60d591b86c5e849fbf443a63845461e349f69ef09d90d5d41ed696;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d01c176beae01a4fdc5382eccfdda0ef7bd721f464930522fa165e2fd30f659c48c0839469c173ffc726f0ba2ccd49ad47b7a2bd85c9e920db431a7118a904b053ae0a41cab578e69e986e6065cefeeeae727434303124d9b3ee7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1abd2f1a7694d8f944f032604f481ce6839a7822cff433558395762b300c1feac9beec5a42e8b5519107337c8b76dc35a86a6a7590f52ecb7b8b22b534a9b64ae47cdfd84ca3e68bd3d87f3020b6713c3ba524b2ff6bc09ed826fdf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf590ad92debb6bb623d9a77031348f5567bdbabc327467553d4dac2dfbfc4453c5cf45f389fefb1476f0686d8bb15ed32f33f900b74b31b096e1d3ebb1ef7df6666a90b1af42c653d981a5eefe1e560ef71c861edfd3d79b8b6d9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d8a781c452303d0d3cd4f80d6ff601b770da2ce64195c80bd28cfe360f19c389631ba5fda11fc39540aeaed947e67d9a4e07ac071ac467c4f750e064e412e6ffa868f4a2d25b4d6a0dc13e1284ea3cd00132cbd26b8fe570d9748c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h74a46e76f64cddc2ad893977743e62dfc9f7203504a4793254f705f1b0f0243d97ee06aae884ac08e8ae98eada758b47a1f820eff9ac0eade5b4dbd35b2446f8674ac634b1bac2a1eee14d2631d40dbaf07d3036d40d7844cb8799;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19097b1c051db3ae573a201d67253f9e6c84a58e0c9296a30f7e4b797c51f807cab16981806fe640de220f47888a5a526db9fdc5ef9cae63684def87abc2fe17b0bde65ae0a708b5e8266770ca825f2d7faa414d0054cf360c27a78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85b353cd6905559d2fc2028d779ef3deebb71151e2f70fec2309bdbe4a5acace17fc6601373fdbafede6adc7ed5a4818f15519252027f6807872c01ca13600d83974ec0fc377ec47629fe9c377a5f0a96ea8ddc2387cd3c92a4073;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1a3023c114ba743fdcaf029c33a0077333c9aba83af25626548a2abb45cbeecf738ddccc794d4f0cdcca35defb6ab827e561b6632c8669c0c3aa9ac409026aede10e35d892cc60010b8289a5748ccf01737cde160812f42dd388;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62e7d54fd7ac2d971ab285d49643990a09b3d3034e74b47d6a96f2fda822e654f92777d44b7f5a47c0e2d5128377a17adc23b8055aeefe2e6dc80159fb0b9d2afa631d0f18c40681ca77e8ebe43341c9c718c7c41957472da701e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d8c8a69df99b175905d48468b11905322f7bd53d685acb79eddfa0ec18de312cb20d49f7f9acf67160deeb33b972139861a034459c20d0164ad365ec58e1ca1fa09c65efce892da45f0c241db3a463f76bab9f9a3d228d828e4ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160638b1f2be69dfb4dc6f3b95fb37e538630107d62ae2d259410df453a27529d72e9f3aa838b563c92a524227de0a8a19147411ee355ef1f9a34af6a4fee43a95da193da56d61efb3982179058b55f5cf06668a158d88f01b46edc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e171380b3c66bc933d7e3f75f5de2fe22542b1f9cdd2a11a0bd7a56ef984910822e96dc9f9189d4063ef972f1a42bf4e6eba03db69a38482fdcacf712249ebac9953f69c05373917dbdd1cd2c2ed515ddcaac45cf834638afe883;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb0bdc980bbdf7d7063265fa9ee81a3c851c7370babf47b113d880a1964f2e096d8e4f4323b05657a39d8a5d4c8b09fcae88c133dcba8beeadd79d5a573046d77db507dde18ea647c01f554ba6b0ddb6b36a5d58496aa04efe9d9ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h981fa1bf4a785c51aac4cc5a526c07a401f6a8183cb045fddb705c9cb0746a60f27fefcce0bd1ded66103e2441a6a1e3ed60546e415e893075de3ff7578ec97c13caf3bd143210266ab61375266664401007fc08c1fddfb985eabc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1992db8fbeb898eab498e1c87d2e326b9fd6cd01e75c2f67b80a72c3f28b76b9897de33900b5abda5fc530bd14a7ce47e25ca684ffa7bd5d573640f0a0811917c8abcfbad6ff70ab7b04aa8c09588b20e4e11c85c8782e07a1d4e0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157cdee63238cdbc822701a432fe93cc0a042db4f02225d5d4a3d69e834d165c2344762d517e0e026792a043eda4304b720127a6ca0560a032665c1b17df8c0927cdc237d8720f6fb0c4c827e3049545e6aa854ac5411af0ebd1236;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68a4537e988819b818e11a3624b74cf85c1ede60085209f6096434da9d173885187efb2f7ad27fc08ea13667c9155aee1f8c7052cb4b6f7dad787e50dbeb746456dabd7051efce035ab75502a5bfc0911d4433af0a8a56c319f2d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4836c886ed55eff12e6ddaa72e04ebf95c82eea58ab083efc87d3e68a177330d4a63e2e307bd424f5823315c89568c16e5e50cd197199cfad62efd769ae87f602c5fe61d024f6f73714e2d4a50e5d26aeb4c56c38bffedcefc08d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1972ce2759a7b6c0d9edb2c8b059d404af22b2e367fa82c4b18c09afec46ded9f108f8d9ecbea5a617bb717a452a36826f033036c0b419a67e729eeab359c7c689765630bf2d89e92f02480e23bc1a60f1bcbe6a113fb557e20d48b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18461489a49747766a9613d0f17d6fbb3bf047a6b92edb3057fd9e98ced75362895115e8de5ff5e464c14f2f497cdd23a8a9b02ac9e069fe15ba9eb0c89deb64517eccf1222edf8c99306e339176e02ef9993b96a60fd89d9ef0b39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67661e556b41ee5f7a7d9c70f10c826be8e0f0d44e0010185ef016ea2f4d384bd92eecbf4b3d6040f501da57115ca3713fcc36ebe36bb9e55dae6219b29ffdff7158397bdef85837618d51dd103e81a644ffd90842aabe3e84ea29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7170952c1a5ccffee3b5eb655c7967f1e8d919f67abcdff2e9fde0f7dbe546e8bd59ed09f1bec6aafc54db5ffc800b33db9b4d10b6373efaa011884dc0fe1f9355f5c4fa6ea85938400007ff09532559fd71ae841069f99dc745e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f617de3b99dd07847e7459a63cf738a50229ded7c1871833d2e720b8a5e9062d69ea850dc00a8fa8daf68d4b1f2360b3d6f355bd2276679f7a9a41ef98a599d8c5e4effc530f2707ba463191a6232c1b3b39abe6c1cee0d124d0d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f79370c464ab4ef53f6c50f411799f8450b08003cd09ef29e39e4580b933ec518e2f4b4f05776a5a3fa996fbeba9e29e56438764cd19118d10eb90d6b1daf32d14c0affa78c61d31f5aa50697e3c800a3c9bf772421850248faff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdca0aaeae3c6dd4b59e6c353e80bd60286843eac5872b5d438904b793dfa6a71787bb8265a3b458709b0f1cf7110f9c6ee75f1357b66e85c0944aaa9a9496ea900b81bc083a2978f723c8833a6b8691aabfef6e152fc168f93a8f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d1015608a71af03ce0385e312a050a21f3f10b9a480a75e3235d6ef0310a9d5772c227bbb800fe762422b992bd88fdfd9cac644a87dad5afbd19e973094deb8a253a6832ac0ab761d4d8721459958bcaf23bc1dd3cabc0c24bb969;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha29e7cc497b1d5a2c63a63afeae460bfa502c894017d604a91feaafca67cbb43650ebffe13c3122df408a686ae95be504993ecc74793304df14e75044d66cc985f918ba55693aefddd9053524cee6ca3baf4cdeb71ed839099b865;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1173e1b5c5c20c5a489f1d92eac8f6bc94f5300d159655f61b2bfbfd026291653900464f22f6cdc7381127cb2d9eeae102c2b854dde77641e259c1e6c5cd4951a0f323bb94d178bce0aa2a6f9c3716446ec8b928581a9ae42578fba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a32dc5b73af8496443d6a67e4d7d7b2dd2c02f4ae92ca50ea4a886febd945a303d736045fbe4075868d1b2c20282bd5d2287ce17f37577c800e163f06da57f3b43e4bf6234d166aebb5d72a319014c7c27942c8f331eb3e96e086;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6ddb1c66f85dd605031d8868d5153adf34fe5fc0a91542815bb007960ca649d9a4e8800ae6ab3f677df00a834274e2b0aa797f466aa896ede0002cfa3f340e39e0b09388e8e6f85122fe43fab09149680408d2f794c4ea5b25568;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b071d2ed0886f0f0e3e662715f67c60331dc4e5aed4f3c1a85fd32893f464f781b2371b3784fd4a212f061cd642cafd6e40ce365f2ef4490d1be8907b41a841168e2080cb42d8fe27350dcb29e8bdef41e2d6ec1d628ab78c3eaf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e3d9c96c24d9a0a0b1928bc69f763e84e311467604e98086bf85e99eeab983ab3499325ca72e8164bb6a3cc04f60104fb1f9552b1aa0e466ed4bb86a0739322db566377acafa38b0b8f034df9acf5f71a6b9a62cbeec66065569b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h44febc95d6734b488e80de209d05cf178f1fd7de886e00c0879823f72a3b4f47b860dde46f425a862c8e248630f890745a91282e4ebd0f3d10c8f0b2aa0c05a2172e341cbf907a71afee040bc4ace9faf45a688013e183978720b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha45a7b64fcff558dc819fe9d4759efee1124ffbd756350e2dac31bcab8ea404bd5111043f7e23f69308fd5a6abcd90c5abb8663ef72faffdc75447b10ec889909c61ecae188086d43d4b88db57b99930966c12a32e54f79dfeee14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc1bbca37fd15a5d6429c1a79b065a8c8b7bf0d9efe74a43ee023c66e1deb342424b8b1e0969175986b104e20fea35b9a53675420bc8d9069a88f253b1b6fbe67f7226e675e80d3ad235324055c76f8df46fbdd000c1f554be63e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1b267290a19064194ae29ff176d5744070d56f5dca7850bf122c638a85f43a32b3132ebd9a6101b8aa44c479d8c3c95de7f219d26f3df4c66bbe3703f9767417b364758fa6778411cee0535576844dc98112980c3149fd7d8b9b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f478ba76f31dfdd94cbae17258b1a25ec2cf5e2e5b6450a8c9f9b43f3ca93cdd99076ccf54d25426e22c89e4e625c9f34b7b12fafe9f1f171e810d25bbd96c8558ccc5f19dff812e665cae46e31ad20286041cfa4afe6344798062;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4f4f102baa88c28d52f07758447f2b7f53ee4a0fdf1aab9b4c141ce5d15e98953e9457e495a38154386fc99cc4358c8c7ab5acb1afa5d3687445efb3e100f29fa3c85bfe2148bbd451d3686579b0c2cff3db4923a6bd2f91f2052;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h760104db6a1734078f137b000c83e48b7f7c72d6c484b75bcce95fd0a1415f21a26ce1e912d132488687037b16235f964ace01969c10f8ea0a65eb4279640f45c1b3d369e78e12caa8e4ffa071b9ca5be55656815fd22ef3895a28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1901eea29ab55073e8909ac87f871c9fd11fc7356133f32eadf52fd9cb99a9be43789f72a89062fddc5730499b64f3a04bd5ffbc95f543614efd758ad336643036917ebc6af82665665931c1e32edcc588b890249ccf78cc149f3d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc67961b3c74f68056ebd4dd6d687155fd5004c8026af9d14f21ef2a052e41e92fcf0f63e90135318cd902c7948286e32653fcd62c28850ceed42423a617aff9f7741a4b25024a33e3e93253841f81ac8c33bab348b371b4091b66;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce7c9d5f3480da67b5a42dbc2ba55ac8e52f67e1a0192cd5ed859dee42e1861a5f1ab4f85e09cd99818b01e4480c99b14628342b99bdd5603ac4ac0c8d5f7b2cad9e7e3fd0bf495746320ec0318cdb1311edbf82036473ff1248ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7864fbe7e62f0c31b963c23f428242b30de83c8ca90878364bac2fe65e4dcc1fba34eb83165c80c0d562eb90d2e3d12c411cbccd3ceee9b71854e3f18a9b20b79654da06fee1b2b96e47ef0cada8e3e0d63ed5346d6c60746c2930;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde378fce989b7a13204cf817fdbb185b65fdf326a107e03cad81ab9b2425750d2991c3f6b4cee96364d778a6e2e0ea64c2922d19a6dc849f08acdc4ace0c67443ae34b7818d5373aeefbb9df910e75a4b32b0c3b0594c0f0dd633;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e354e2d729db6d020e4a8493e6f26f7eba177def1bf147abbe136a3d28f401738fd24623333a9ef5cbd4a43ee44efa94fbc52df41bb71408268e8de0cab85888d836a29ae8aa5d8cb9ca2157d28d6d0c936aaa785e1ee99582b837;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185fa19b21bb00e6b2cb2cccc836f42ec41db1dd6558206f431ea9cbc2ffb37ae4ef62dd376c33ecf53e82fb4f2e677edf9f6fe1fdd1c89f9718a7c1a6d9c441fb0b2fb859d671049bb921cbb2c5c15e009ee819b50bad5541d92db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h819666ac9be89eaa609e0bf66adf8bd3ae1cfa0cc987b345e7441c25ae964daa5ca930a4e5aa161f55248ab2b67f128225e1ae5d06472becbf054d77dbfe1aa1425856846176c6fc0b4109dc0c79db098984cf70a4d11abcc35b72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hacde423543f426473f00063f5ebe9b19d6f7cdc7ed0d9cbde0382db52e23648978f7afe2defa8b58b1d1138ec87a3985fa34af2b1591eb358e12469538f26f66ffdb9c6814189dbde8cf762ecb244cf568d6311db5a8c0ef7e08aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193b8542e864a670771c7fc942e72a71aba98b5a46bfcea0f6e47e74361d9a7ff9bd2c7067d36a36a92b9f1d92534dc1ff1e1ea5b0f13368d4e2a1a58d834279abc68488258688c07b6208572b865ba11ea467159009a6f513fdf4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba78af3eee341e3353957403c4909d20ef89fa447a6c66d05a48e0f8a0f1d5038a2cbb5332a4ed834a212eb49bbe2d8179c1453b842735630a2d9c4156d6d64ba020325dd1fb0d99e2a7d9e1f8fed6837059608bf1c7d0f0c0d4fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a25e26ecc8ce77eda9f15445c463936d5e4081148dc2c11bd7c525cc408f0544a39b1fe87935baa45f142dc1e84c10e143bd58ce5ea1a721db55c51e3c318ccb0d1ab910e08aa629490a31f8a06d392e061d8a6b5c22b549d2430;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f36e7e138d438bc8d45c1fa256a475731f9edc8a2d5bff3523fb5db38d9bb0f7f62f958f6305ad035b3c22eaf2f654295fb17832eef3ed2c5875a6e4fdf9474d68213e1df809693fbd1690c2d465c6aa0b430d5b8e4559af50ef9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197924d7d1d9b941982ad2715f3727509edba00a8bd969594b367c1bcc55e02d90dcc5e479ef82638366c786c0fa82bc41af25333a7ee0e6653a16168bc13a845ef3b9e623d8bacc40303f9c2187d9d89ed526fd57c4e535600dadc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1801e1ed5cdf2c21007a8d9afb35619c9ef151a11384d1f1efe85b34caf2f7b625eb87c1c84343f93f4c8e7a02d1480dd8ea552b16d9450c1af3b433aaa52421a6f6a1047ef6755e3354e50a176cf3484e5940e95d2da124e66b71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a079a8dd4dc07e45aa99f4218b4f783c80c1ed33c2a7e98af954f7b76df8e379e5816eac6de813f135b98c07339f46789ef1f7fc14bcea05a3e94332b782751cccfafdaf66ef0a6def820852439d1544337394fa55ff62fde9f789;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff6c06511cc26fa465d1d57fc5f10a1d98d1fad0688e8a7375701636d6d25dec80956ebce9035a8f17161cb2db969874dae69a6e95e7213002d3d102b79c7514bd5534554db2188978eb9d4b4f3346ff483533d6091af656c762ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13daae539779fb3ccb733d1febf20abcaa3fb2d4bab9b73f7a2f2c13e9774770f8ea8cb89348140846c3b84ef7cee2e2dbd9bffacb760f926df392b74e9b6162bf94950d4f5e1414d3e3e40479af670e7de311a9b0fe91e6e5b6893;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef612f27671825376de21aa905fc8989a3d66c770641c94a987847b43697c960c68cf7be9383215b4bd16eea4a82c92a99f0b0b7575a8b40145ab3a456247dbc66dd532b31a369f0a2891383935da8fbff46bcb039f347a6143ae5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h982406683b7931040c68491386f02d9e5082d43934034aece7ab4b3e49d1ad55b5de3ee8e30ae774ed43a2cd72bc406e64647adbfdfab2da532c045f4d1397691f5930c2002534d7d925f3781df863f8dc866b7e1c5058dfef0c06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1b9d8ed7a002928b5e8d04a0bee408f61932533fb31069bc0329f86c2196542213514dfad4063fc63ba14e41dfaf887ebca13a8955182f2020638e082505a83ee638816cc50158166d1ee46f690ea3a12d68c1bc6102580007518;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16cdc950d8519f6bea6241c45235325e815f80b39c632ea63f5136f6da0473b0af1badbb13e22b138dae8e8d29590d67499e35b91276b030ea5573851cc300ad198dcfde7346017f593fa1a745ae5058d17f508ef7539704e048089;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d12b07ea6e4a61226a8d5df718cb2cc095fc58fd8367b9125f54146ed889a33ecba79fcbd1597e2db5963452463d716f360e8b6971065ceb58b115aa0de9df13e3d3292aa4f6cb385bf2ee8458462004d6c757dcd8831f9b19c7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1096daa7e228bf11231d1461c7fd0482b7ad97ee7b66f07fc9b4ee46f121fca21527bfa26da6391e711bc0501149b0ecc9a5faf57ad168834bb331cdc19f5ac647077a160cde888fdeb3fe95bf00eeb39b36a70d5274e0a43fa3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0ffd23df9b3c3e4f9f1746aae2f74c85d1fd911502143ca489278a4fdbee9c0e9a581b27e30e9f8b1ab67826d44758568ae34d3d4f74cc5c4da66eac132b13b214d3fa1e6031a67b2b9b58c4b3df28b488f65d103beaf93900a5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd91c001cdc7778557d14263fa4b357e09ad94ee9abf6922993b13add3c7f8ba0e180aef6a7f1ed83e5632a588df753f75627017d2dd288ec85c04f006f3ee9ce76aa0a4683dd1a9156b9a5b2356d2e62deacd3173a4ed64ab908a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h66684b2bc03e58272176da03f755aa18957802df68fa3dc25f024f57cd350944e068d175dcc36966ebe9f8fad48639291bd36f519a77ada2961964cc3b232966eccff537c791ea3d45e9d7044ff223f5d9e6eba34186dbd7898b95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h997147a309c211ed48bab383ac3c3b20014d944b641b27ad424599b9abd7bf85e8892d3c70e6120daa180320555a9cf0cc6302388cb996132d565e9e2b809f2c55b12f43d2ed32a3071184483bedd6e973392657dbed365781d9d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b4c9def22b41bf4011e018e1617288c64546eddb5bc824e0f8d3e0ae4333443430743651199d3e484054dbf26c8a5daa9ad3093953c8513f3de2bd6eaf16414636cfe8613b7e685286d5a1df9c91f985871c33be51dfd026d0908;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a54fd7cf8d687d394e1c1946d44956f0d8f6b84ec4aa188a90c4ae28acf681d27a1fc3a38e59b74f694db2ac880aaff86c200b36e0386843d8accb9b6402600237921584cfd36f7bbe5f37a46d6bcd701d453cda83cccc43022fdb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed0e1993d9d6a19eaf7d7b03ac975d6998f000fa4bec085e1fb88509435262b7749023064b4d95493d75a899490f46c5f56853d3480199b7f28cbec306318ba8b88a430b2dfe629df29b4b3109e0addbffb34247c563fdb027c24d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2339fc566e363a064c00bd7b09eaaa5a2557330762d0d4c48e38378497f10e70d089bb0b652ec772357be4d805f212c0c317a778f7fbe01b057caa6481d62d5db35333c39a71191fbc581dd0eac627ef932a4c2c9e9983312b546;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec183cd14d76f04a9b6fdd522ee6e8ce4e04099d05909244a1fc6065409697edf8d4685a7fdc3f7e600e18c774eb79aa86667a6bda95be3f2004cb3e4b9d433e6ade64f23593667ee8dcb172a504de7868698f37da9ae6bd49fde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5fb886385a724bd80a628fa25a17664047c38910e6a616ac9955686ce5f8b331770a7817516df720d28db22ffb245f7539443517a47c71d7ccef7285650c2840e65ea80e7a6fc36c96af9b40e07876593ce2e65d5d426a5214841;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf67460e0f0a51d18a254313e6dcb1c00c6fa72e92b5071b37541d439a6d77fa958626196bcfd2219eced369ba1febb953d386e4dbec520b1ae34bc8424725ca552da053715fb315caef719593210ff44582afd9e543f719e05da1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17432c8cf66d3e6b9cc38021742be14859ad01343ee30782530e3461f8b3cd18a08be8de7b314952c02f31d274f6ad41f2d011596b0d8db1652844f3138d43f46c90d70f91d58e8c9baa2a5f86056a7e2a619817fdfa4d158f63577;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190329c6b4af089e5e8eba939ebb50507a5b8a5e0149ab0f492c2801193e576d9c9696f3f30b5a04fd7f62a548ce4bafc0192d40db848c60f836741392784597a1f79c21d98d7c72fbd08b9f2722946aa6dcd215076587341d196ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126e4a3991be3e2a567db4ca0729321ee1b3a427c316aa206c7fe34a93cca1740f7437a1fcc8c7f5661d89652e47b601962552713361db28724040a833330fae1da93cb2499683a237e5776f107ad69b6f6dec86e16be7ce75d17be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d1b81a09db20e8f42d0f9b696e590a7e3c2318fd7c132e126e3a14745bdcb5e7c478d403ba0b268b7b3bc12528b1ce0be1bd3109e92f5901ff1f764cfab1091151640d7d4f989a200aaa9ff705aa93d632024fa2415c73e3761512;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h588ae239da5b206bfdc9a3a35a79e06eb8528d67dffc4d76224e9a4ea45a8e16076462100133f2e67d1ec7f3007d35dce723d696cfbc4fccef712059d5921c59e8c814d3de8cdbf4da075ca5f0d6af1eb7c3122439a6bec2b02d03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h381ba020ffcb1dfe3d9d6415f63b60b36ae317b3aa3003fda35e8a224e27d73e39703c167599f875528f5ea29195fdd2acb4871cc67a80608a9141a96f54efbc3fc45d5e5f15a7ccfad8aa829ce471825de4f97596eb1332dc6f73;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15deed4f84e2285b736aee2e8930e0b89be5c1f9e1ec8aa10a19bc61d0416a6d99709e25cbf71941f03a1b10e10293901b49ccce361c3d440e5fee95e98c956b80b3848bf8617892c0b681ef65896c88b5a81ac811108bcd8e98305;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67347b0d6a920f0c872d06e416b519d14b28a644a7cf8ee11a7b667d25e50b3f01793d912011db3636fd0815186c50836ace0366b82367c626bc42e49f1e111525bb3b2e937fae9c8fa6e815dbd3d73ed5a2294b3a01d6d247cf37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h162e9f0c7c9a70a3b4959bd1af0f9fe7a5cfa81d02365483e9e169b0a0137fbfe882547e8f093ad45b91d0f55589487820b1e4840d60098be308c3ce91bd05744cebda2f9a05694f5b8ee64f67cd0ef74d854d54cd7cbb164be72c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9f5ae6270cb08c09d6b5aff64c5bf2ca7430f1a0f511a3ecff107e6c1efd1f45025c220740694c7923d8a5b95ef831d7818d7e0316a9931a902db772e4a1120ba158d86989dfc069316906e347f2751aa72fb3a6cd5be50ba8686;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f2633e57c9f950d34341b509512eb33343efa2356b0ff14861d240dbc7f43bfcbe25108affc9092fe051f328addeaaab82651e7d87e71863dfd9453c931963520288ca658b9ac197dee7b0df4e334e09c81f576826e619e092838;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e9fcb233b0713fa2b8dfd05c1b1273da78151bd17ba2b02f7fe4eec4298db66f1c89832dd3aae06039687806c20b983dee49057610503761f6791044f3a329537e36f39c486c0da8d78e8890d68536c6a0f0293bdbdf06a118b01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14da0f95f2334be967191577ec124d8b4e66beaaa348ac3267ec9417b3a7ad2e83aa3509062052f10030ef388b576c5677ad4688d7cdae498dfe4f0c863d1601d5de2160c47405fbb47bb9e8ad678b026c44abb8df36066dca827b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54e802a62bb13239b60e6eb0c268acdea0b02fbeb2b5821462968330678192ef069700a54856fe343254a459f72d545c5198971694e161e10146fd8fbead261823e8ea12e3f71e8bed9a90f6c5bc7437e06bb7ff64eefc42433e9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf1a799cc61a2257955aa55a2284173dcdf311b3053ddbd0b32142d2ed257016a9589209e3eb794602c09ec02ebbcf5e44c7d60b732f0f6ae0cbc7ae0de287605328b6f7fc680de3d525e28b57cf177bf7b2080589503dd2f3ff16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hac6e3fbe54dd152e78936ebe93c6ab0e4a11f8f4fc99ac9205382e3b3c1c20f3f2e72a949677895547c4fb5a71704150ec7df709a3d4651979a0f6a76ab833c257262f04951b373285b6928ef9c6ac55a1b5c532dd9bece4ef8ad0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he699dfde423030c05a62d40624ad011b5b487ae9c57c6fb47209b711cbcced8feec44e750c2331e25d97c4d440e59d69756d9f19411e9dc68846fdede3d90baa80b6b69909300dacb85eb04fef532cf325e2e01f99e6e6ba36f83;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ad24a59e93ad546044e3ab4beeb68470c683da3ad207769ae051740cb22543dfc1b26bf973360eda360f257f6fa56ec8d3b6cf41661b65ad231feb9b1971fd839b81f7b31ef27244c45bad50c6738c811a97c84ff22767211d59f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1658655da212317863194681709787b91262cf99d057955230f4ea7f0210d81a75677d7fde0a237744130f529ba80e3c2f42823cd884316732fc1e9b8cfd00585579ac05f6364dd917f5149ba1a872a709437360d7f121e61cdf615;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1e5bd4703512b8e73ea3bbb536deb07bb77d240d215eacb1a29029695131ad28561bc5598ee0495205def31929f6f018df9c808b58ef05f27202c861855d0d8a6b2421a5420ee5b2fd2969fd608ae9267ae0367f416b351f5706;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19189465ed773197cc2162dba052b8afd844437aceac914e54ea14261b7078192891396cdef274d36fcdf4f9dce5c1e80360c36e4798dd8916dfc60a37a4f0e0caa13c946e44a768608293441c62bcab5e42df842eb83686b74efbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff9ef5bfbc31a249287549e23023e4f199a3ef3b61db7bd26835a44aa932f00959b42083b841fb27395ddfeb9585847225cbe8e395133b7cfe0f55a2a01472e504eaf9fadfb336e8ec444d2f55a6b72b318280d3cd4a56b8b8bfb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d3d6cad04c70f1137fbf07e72bb649f4226922ba1e966321085157c238dd9fd4adfff8a31962a1863ef87a82382eb7eefd82d28aa93cc193a6f2654a32e0510f1ec33eefc0a68e91e1e9e179e469d43d7d973338d95fc1b3f0df1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffdf788c197dedaae4c449d10837b75bf3c0b54317117d28509b26b88a4e9147bd6b07dd3af0d398cf1b090fd6b4e3e543f42d4fcf13b11354bd84211ac55cdc558bbae42b4a41f2904b72512fc28a3344d34c3107adba9e1409a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd876f0a7875418f1b3bd1fc4a2a759e3f21f73af741ca58767f886274f6ee468eb315d7734aeeecd009ff8aefe04b9c320fd46a67031adef1d5722041c7f0bd501fa74bde1f702ca86aabe21fc9627f6608a52bcadc9eb759dbc1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194fefc3491296a7dc3e7a8d10e5bcbd427a1d0642c3aa52545d019ab05a12a8fcbb5df54865d7cf896caab7775b4d3dcc26017e471ffde99f0614408e7e8ddcb2763011cfa5ef88b77e9a983fd50b24897e03e23c753fdbe58195a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h92a2c6e5184db2fad52bde73042886f3b944dd6b18729aa406e7d519f5c190a5f792ef3edc6f427be0a4d44d43627e0553bfbfa6e8bff9b5e118c181d777f10701403ba04be3afb2398e6b76ce92549ac2ec6de7ca8a642e73c600;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d886f7cc546a2f85e282322115444500bbe3cb8ba43cac4e20436e5aeed1a1a1cf51097bbd6e982d33888fff8f814f6ded0a122b44d6fa7b94fd46e18f1e634430768c1bed3dd2aba7451d7266e2bcee3438bbd996e420830317c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1033b2338b9140534f64d17d254c9e18a452bb8ddb33f3d1ce024b88c24dc99aaf5e365e042c30aaab8fb163953bf69ea6bbfeb03c0d038b16c65c56c1ed57785d8e334f32de45d90d484c9239ce964ec2746f5b41eb17d5df6a998;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19386de0ca07459b67aacf2689a3f83566763093e3ce7e0abaf8841605259d2fa4f9d6865d7b35a8ecf38f7e62cb0a9d52286413e3c3efc90aa2af9605913f1334d3bc84c6f3763f9360dbfa83dc4aa36d2000ec6832d090fdfdcba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190a59698e31204289a86c5ac2f4d3bdc427b05c5a7a417f74ce58644937860384d4202982eac674407ccf299c47cd2d0ab9bdc04a34ffd9f71c5a84f08182fc357542bf3f6f583fa4b3cd2dff710d5f54aed118fcc45c21941aef5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h198886a26bee09b39b59b87f1ee1c054ccc87b55ad962dd19e510851bf7fdf2feeb3b1270da969712869c0b67bafd02aba4a4c84b5ca9416ab656462b944cdf9c9e6da9a0f0396488c5ab2cb14368507584f15388847cdc565105e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c283346b9a264544aecff6e13039406e1beb62058ba214c08736c9f1dfb880ccfd463f17a09396b5392a501fa606fca00ee9023f3226ed100e4a45a37ca5457fab45eadf5d744e13ac0afffb37177e9de881337cc733064778d0ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b2a373454b1b3efedee6af396e504a84ec534566a105b82c416e69529d35981339322fa5f3bcd9eff20c0f8fa7daa7bff712ccfe102514c3d4ab84acf273a0a1d114fb562adba83752b558490a02dddb0ea911ab5115fddf7428e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe07dc493fe8d820f8a692e9093641743285b2b27627c7f3e3b5148ca344b7914e8cd44316db418750fab7a93ae2e70eeb49fc0333d2dfc5e10464a8a0e30a7730d6dabc20c251d435f0c03c55e2e47539d2dd09f31e0e83a20614;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc7e963092788854e5fe5800587c39120a848550f9829fb164cf031bd7e77f0d9e2e9f865eb2783f77c9796685bf4044d33d9f19561870ae0227386907536ad63ea41415f1c25ce14cbd4dcddb85f0014869ad17f7e9f9cda333c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h698f450c86d2e10bd52e710d9383ca649ddb30be1332fcc08883d5b9f4ec8747bf0b5cb8be06c603d2d4270d1e41989cf3edfa5246dc59ea3c08c0a5a15959b17c4ee8932774a32b0126d1d3cd86edfbe8d863a0d1408594babc0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda0a84e2689daee35a313a1dddea3ca7b6bedc615e8598a35520d89a5815a8172093771d097f31266f5fbf1cbdfd329f192fbccc06124fde44e7dfd5fad35bcf28018fbe2c12b17bf015b58dce1c4b5de2a60c24670132a16c9a68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc17261ea62ae7643db7d438acd7a3bcc70fc0f291d763878bfedb76a7a0df4c2ebeb2df2ff123f804422a7e363c30aff7ccee013a0f8c4fce4f38236b84bfa09d93546496992e171af7ac54597f3f24b46aae793b8faf6ea4e6658;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc5371a50891c8bc73cfad725d7de7d7253285badee0ec06440f5b9c8e48daa1c538578442d5c439860f3320fb8689fcff1dfa02bb68b85930f2f1053f451db322fc88a3123527a16ef921eefd08c9b6f25767d0abc8eb14ea217;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h341a3db618194c39500b2cb448fbb098d1181953ec48135838fa30e63ef1835c2f8d7093bf5b55804db7787b1125df958cd7f6bc1f67649d9d694706986b7d364715784eeea5bcfaffbb86fecd798ee9eef92af03cc0898d4bd2c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35a6592242edb0272eb3614a580222ec2a86ed19b6b97002eab37a64e03d71e427c28be3f9ee1a90cd13ca18da9391a5895f942cb975a848e5368879e251b9452594bec0220d42bf4c62be38bb346cada8f93e3bdb69fac996ef8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1702cae507f8804d701cd61f2b890188397173106357550ef2d47cd42400f0a78dfb3e9b2ce629b25c88a4928e81c9e4e0f5d8893397f878b720a877f5e3754f7c32aa77c7042d6c2709b853a3e6dfc45de1490d8856f6b36b48996;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc8302239167addbb1ea73e4b2ba9fc772751242447deb3fc781bc82aaa7db73d815fc90dc9138cced0f9eb94464307518e830374f2a37a74afa3a96bc70941a4f3c091273c63bd84996e21c329a8370588ef788c6e7ec13f7496d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h504e11ddfabdbb8c4f6c84bc6a2c4265740190ae9e76f9ac72249533534ab8df572cda202fde02b1f8916fb192909007ed160825748214922d50a66b70d2dcce9a8be39300e6a6c4fd2f8a41333824cac26f1949058f83ff3c6151;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7f55da07e461d7d66734a96319e610850babbbe731384a19214a9f07c8d35d6354783913f975f7b73e1f909fc36cea8dbb46e226df753687f97f76daf4a41ce7c6ff52a8706bc0a76329d68df6b88523ce99993046d474d982882;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e31ef812c973af2e929af3ee7b716e4cabd2b2b7b7f1a23317d4f46b8f70226c9ffb6c202bead64c6f38064009cf0cff70e304f63003e4729d416927ba859ddccf27746c69dcba914fd559f28fad82b6bd4e0e3dabcb13eae1cf6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190ee00e468aa6672ad051ddf459e6250c75267386d9381e269601f66bf6c786ce9d299e25d703670856e8e4e0a1588c13bf53b4b45ae7db1d67ed6afcd3351a72c99d497475f0954e95870ef8f8488b11f063fb0b4d84dfc00637d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ef67f90785bcda2389aaa9f76fcf66aa94b0f289f3a07dffe736248bf1c11abae527e956074848e2f49931b8b81c377ecd614fbbb3f37375a132d3ae04784f7632b86de164e674a69ce729dab25a38fe8d692f291db9347615650;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h59042ebb5770b75d605a48ee1c50ed6e1bcd68f7ae647a5c577dff650586c878d7dbeda5fb1b2530e7fa3e0e9a6a5ac95e44b67c47cec175f7f7dba9abc8e3b46e9f3205f5b8ec4652bafb8c114b2669c1249cd2c3ea77ac83ae20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ff6ef45a4a3ba1734a3d757609c96f3a1e504445a6f4c0597d95de0cdd8d48fccc46e8675cdb82fe12773b7380f21c0bbcd4784f3bdb0906f0f2b9311c4a7c389de1dd3169bef9c54d863c233bd577728b168bc16d25f7301969c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1675231fd9b67258b15cbd08bec48244b4c7e7221c608876a1543f12b8c071800ec04bae6fa1129efa575e206fbe79c42d81aba8fc55f6bdd257a46391e19c31d984a3263f45c13425f6cf2195a9209304d9e97cef624d791916292;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e91c72e0c1843e201bcf6faca39b7b2c818e361a135f4948dbe5db4fc04f23b71b9cdade46350efd2f3dec576fdd9b497475d35deb2528626df119a4bfeeac1429cf848fa2eccae04ad0e785b64ff17663208257eadd228c86e2f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7100b74c0b82c2262b63b849a000fc52a24531df90b5efc519219f25442240d0f1e3e89b344a3b872a7e71e38a2ff7898ba5ebb6a504358bf6f650d21438b9e2ac2d6a716af0e4f71d49a5ee4288b3fafcd9d046686309ca5ca39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d904f86489e8931869edecbdb069d8b003d0727b28f86ed0b6893f1644ef57c93f053a14b125cbf81206b91fbc0528f724d541b2f2cc0a405a241552967f5ad94d5e5c1a92418a8cd5b23c348c3e7df0d79e2118d147cbbfb5354;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c53e8910c0c026b0ece1531f53ce019b2160c734d145428d61bc400b33e98cb4ee0dee7c5003484b9081913c5b4e79ee487baafbd9ebf2e42f0780b7f110cffc5d22cda0183ec475fc39617b3da7a2c0ff56baaa2d9d6f9b5b7fcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72c169a80297a351d3c9cfd81ae81fe6f56f07a6edf0ae846042d2f5c1488ab64759ee399f369ea8030ec5afe629b97767351f20d06bb90a5846c89028c69bf67b0547b0f285e009fab7c640b9e4b44ec04d4d1c110ac77e610892;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h199e75a80b4fa029ef67910e2fee5466e66d5bbba26794d333b0541e23cbdc410b258433fafbe5c44566199e2d088b1885e808fa3a7720747d1e4b33cc84908a93502472d3afd0be58cf46e93c7c7973e79d6859d9440c19c3ea98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0acdabbf159581f62b54937be8b39e498ef17b6beabcb7a902239601245f8b7d260b31dc8fcac94cf77600be704b79a586f48c70de15373c9dea4139d4ef1d9c00d3483a708277b08538a81d94a681db569e280d89cc1e67973a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea231393a542fe0e67d621aa880487d11d0216ade3b9c63aa42b3f2cbc10ce94cf0900de8bd623099ed510b49fd95eab1b252776ffe754a0b822a7a1a12c213e78d9a73552a2fb69aad0a483e77631f680e8a61ed87e690eb37b36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5970d4c903e4807fd28e5e9d709a9c9dff246f562650be1fb339cc04db119abb9aa8c8f6541eb513c5cce3a404099fddc91bd8e969120cd6d9a8fb0a0176aa53444c7182d253a7435a9db0229cb03fcf0806a8e6e129d922a165a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bdbe2f33b05901b78003ee8a30087b4cca87893d05ff18e22efc8a32e4907659a765096bcab6af4b68b92ac6b5ae6a0257781a41cfa0b0b343311353fbe46bb0ddbb5285ef2c88d31c5331fa8e0746d57f65449fc7de0d1172614f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1479abfbe8981e0a3cacbe3ed5cafd594a9f5eea36611952271b13b81b17cda205f4208de201235a1c96b75a9fc1fd80fda212df2ddc0a9e68028e915443d220f7b989ac0e48d378f2c97d99538304241a53044a2e623a2b9a78767;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d337e781c93279b2e33d0329168760c9e7d9b86ada4cb095112d7e8757386f3db68697b8e46e8ac18aad31fd5e156301a0a97fc95ad2b71ceaff3ad26a65b120cd05b17b8b2e158b647db98037298c1a083ee4620a2dcc16551b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h162027ce4bbc0b184b666a5de29d4fc0ab78d54bec06d9c6780e65e8b18cf4d7c9e50698f7af30b34f9ee55bda5e72c744048dac40b839a50fa240676d65c26a7cbcccbad91e8a4b12323dd7e041bf47519d398387a1ae114ab03ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130a282ed6f537d58a8140f186298b5d731c1691d754d5bc2c9406acddd6c550250c2e686481ebffc077a274180f41beef38034d88b4082fbbd5dde0c6f5dab4a970817d15af3f59e86b7f327ab4b38b026e056191c8ee585ba0b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h138e6c1ef67730c80bde60db27013b0dd719e52a2b414c53aaa5f25d266d5e7705e37276ecf777cbaef0e1155d837fe13e6f53e44ac8698380af29f436a13f546d3e4c43a8efc624a1c01741ca7026de8bd88ea888619abdafcad64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8be0ede88c569bd8b8c54e3bd73c43510aed341c2e24ce88b9a00cfd1b74a627abaa1f4e912e103fac6a5ec71cc9b935e32d86c6aae1b882fa8edbb140595a7333a3e47ba768563c95e60c6751c7fbd227307c36c02adcecdac8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9a9f8cfffb80d714a6f146de1b784b5e32646228905367e954d2c5f41873743af788172267c504cb136a5f551596bbc5624aee4818122cee6a8a78d282101bef4b6ad85e584fceb7def2b4c3332c5606a8308fe233cf9d8768f10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78aabc9e7fe2ad63f67be70e3714fcfe1ba2c10df3c60e87bf8b4766b8d627ddc330f1bdf2941216d18656f9a13920a38c0cbddec2dd0f188a7f8c7885690179f5a60b81431f82f1a455dbd054cfa52418af355a0e7641eb332b31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3da83b3e5ba37a850195ad937148cf81f83ccf48eb0bba0fbb4e435a6856bcffb66d33b769e6abe99335faddbfceb3455c75dc9322bf553a8afad9be76f873e12c80c1b20b5b147c91b3940071e47d90bb98f894819affdfd5e152;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf2c404a7274147c87f9cb8ed95457f78ede51b776433f39ecafe1ba9b8b11b5d783b4e7b64f8f1f73ff78abe71ea710a6529184f3d4fa986d219973601aee2dfd553f339e5a8b9cb5dca50f54bdd4368c6269956630095dbb8e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14dec51c5beefaabf669b6756cebcff66f9fceb89539fa755cd836d0cf831311bb21cfcf7e30922ccc3f6b908d308025128b208dc8ed9eab1b2b53f635e8de1433c93b6b2467df8cf6fcb7d50879b75d3e6ca7798903ec4e8717f48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd6e38e7f553bb14d9381636607f3121101f6fa778ce7d9971f59f379bb4a45d3844a4f872ff3bb1cb653ac12d44acd3eacd639904b32b603ffb973867fc840f7b969f5c7ef72b89d6438cd07d7021c3d97b3713e6d7e105b8eef75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8edd67198644c251a6baa0512499757e4e91cec0dd83c15d79a13304a155d27bece9c926ce82b84b462f4aa7051d910c14afdbf5ca6898c79db2e317421d6c1da6da54d2bc9b4a529dab63511dcc90ccd55b3f6c8df8a87e916176;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b8324b2acd7c184b7b1c2111843003955e638e533c005e4458c4c60b2be4af9002e5bb585dc5cc544a0119708693f39fc051520ff9ed91bf612d0cffddb4ecec6c4ff8f6673b93069c0d4305a4bd487f88c862d3781abb6ef968d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34319af4ee800b320d8eaa41a5fdc4c384c9ff2c8e229d146fd4506bc8234a0105407a84c568aef710ed733ab323d0fd558b3567c63ebcaec163f7665cb9b78b17af76b10fa0b8938cb7725ed36ed9cf5c83fdaca5fa73bd9eb245;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d07533fd806fea3d44f1b1dd674ae086f9e089684dd29469feaa87333409ea36e532982ada0599757c0dcae8a766765108609ed4edb80d3cbd3b9be48c7c1fb0a64cad83b287bb026e6437cab0c601a25667bef6546b164bd9129;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c13afe597c263c75970adb857649c9bd710604b5b3df0d743a123cc95451bfc304af51c16246044fb9b7d62a9c46c9dd354757af134a50d6b22d6d6e44b9f986e46b56c2dba990c3282ff5a8eea4a9f7882dbb01dbdb74a9e8e80e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h65a37572222e358c8734cfa7001868d17a3d1230103013678dc8cd50de003f6f141c9aa2ed9ca692d62a2b706a7328e0252ee0b26a4d056249d3266f945c111674d3e765854f7c7a9f855285b1242cd3c3c85b92156e6db2d669d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf48dd0d87cf15e8f1a6394cefbec0fb75182a9042f7a59f93e09250af03035560fd4a0d62ec8759270c17c739dec5e40a99faa88f5e48023b388ea2c61938ebc0c5ac2a4fbc8023d922fce711aca51b6303b254a3c56ea5bc8c20d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11bb41a332e10b5200dd861281ce1c6a78cbf7d2717c7e2ce6c00c1503e7aa4bb93daed3f6a1528dca7ffab8721eed8202c360a8185d61256415ee6ba668cf436ae643ae725e2e78cb9daaf14f583dd1c5841f5674ee9df32eb9c3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h956386fde5346d74ca834c8cab59768e87c98d2a32f2bd49c05f074b60d8b9bc0144fa91739a3809a03ca7219935f9ba29666493c5be8ea39067e6c8a7bafcd7e2d3aed99ec6ebebc662e29810218c894202d89209ced028b5be47;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2fad9c380a1a544b490080aa5e194762435744ee33a907784fa1b89075c51d19436b7f3be0012b9b39425ee94bb1b77ea7991fd414da1e205e841f95308e6c44b2445d4b977ab3c5c48a315f94a97c54f24a62164146fbe8a5757;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8567e0cb19ae01d14482c2078d8af98e956782704c8258b1834ba7c34de371314e43c1c0f61f7fe1fdc9f2f0eef569b7d3508d9b44c03da0d9b054095d922ccd552ef1c7cd6ba21d98db402a1e5d559e9c44462e77322626f7f56f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b31ccf8298c0200d3faf3d6710480ae9f3368d0685b629828bb64f38cc8b7aaab249fbc048487b7b978bbadc34d11e0c1d6f518e7ab6c16819d0d8e190b3c03a90484706dbdfb95152ae954dea7c6c84d65b2fa2843ecdfafb75f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h561cf5a325ec93ad10aa6645e1d0c7a52a08c7925d7cdfe3ef54e1f0f751efec3190970295cce49f3e62bacfae11b5f282b1010642a24091906c2552a300e8da9126ecceccb32147db86d4121b13eb53feee22d7d10571e7e20197;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a128125233dcdf4ba2e6383de93b60ea3fda017a6963fc6013811798e78f1ef52affedce28a4a056b0c1efe9699d93f859591ef26075c7e55d35b03eee50118d05ea54e077415d55623bd6ab0c23899037687a8a0695542c1c82b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf185cbea0eaaa33f1b3c802c391ac04629a2a9ecda21ab1e56b89e0110cc786f7f6a94855a88ea0a76874c45ecf0893656520de7b20fcc3c1861b382dfce647d3592b5ae8f6de80d09826688d676ca6bf9b6bd592b4351824c183;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1957f42755ae9d0cb54ca168c2da46edeb7fc6d49ae260aa885ce1f70460cfa99fdc24ad0c18fca51aa4b3922c98b1bb9922020b9e704b54c1252bf76260f0708b911dbc1f992050c9b69cb4759277824bcd98cda212bc544748adc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7db8b7b27528281b48d81eda210183689b1a368326c139d5e22ac4b5beaf8cd8ead39701238d4fd84c65568fe52b9b9c6923fdab2f681a01f3ecbbf4e295cfe754a0a0471c55bea0e2080fb052e3cffd008b31621a6e169fd2de3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a21a721a40b24b4916bbeba0170ee659e2fa38ba2cbf2f7d0c453b912b0783a03ca71c6bd8621fa566bbfdb71e811e5024f66bc07cca843a94df1fbb51b04417f277bdec70f1b0803109ed0d3e581c692a865db38f5bec146faa6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce1a635226daecc04545e96f62b253a901ff8d6812e2c43d14934949d82982d6e17d86c7b9e4b89148c0280ae1bb6425ddcb92993de84461d236a58e0f41238d170f263cad331459d059de4c4e40bbd107ee81d34feac9df0826a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a46c288232aef5b34f76dda5cb64f4332c7b974f7af875ff5fabb340151b99f9f3da24567024bb26f5921c3835e09e01913a0a7bf0dcd8aca664c82d65a929656dddce5295fd7052ff802c59042928ee4bf8415f73da26800e319;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97ae6b96aa4d9db50c713cd31f066060d7ad6d96419b29c651bfc383a012c1a3e06a59a9f0f98b04be107b7fb1d82dcf7978f6a176b503c960fc1319a076574ad94bb3de7419f656cfb266a6773a20d6f281410cc7cf67a9021a37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ffc8f3da7a31f3bd4fdd43d300275a2aeb5dcf1d69688fe4ae7f69e7e408e07876735ab60d8d5c23b67992b1ada1863379ecaca3492371fb5587121b511b7000b0d2a06b7f727dac321a1e59a7cb190bf6f8422957648567ca1f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hffb7af4cc2ade51574e12bc72f33e782370445ffb7f5fb7f4869c150f7fd7bcbb42de44930d71a0ad543a7cd95813765fe9f2627dc4c73e2948edd75f5a007e709baa0307d6f705206ab3eb386967cac6d71d11140d9e2fe94866d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19971d47f0498272f631f2a78963c4110cad01d5ac65181915c002a9a5d7e2682ab9274576766e3d75ff2b9a0bfa4c5326dd07032069dc3e580d42705b8cc7e4b63bb3c217de5e39385cc96fbfce7279d950a606789a0aa4fe21d2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf73f59b53c32c08d71d84e6639cf7ded7001b5591b37d1de71d802c0f81a4c12004ecaa9387e70805c9e29483eb8aab1dde6d6612d8e8c648d0618cefd5dd20fc624ea3d33687b7648b346711f5ae6384a060b6d9c20d2a7f9b45b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0ec10533690f3d18875b1abc1d2fb0e42a9d95ff724a8c1dda88ac286b1bacd07875b923021aba6d3fdbfa7b31dee0824c1a199c48ff8f32460bfd257d74dd8c745b9dc1c693d30294aec7a09f5fd98a1305055a7d559d08d5964;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc78b37752f942c41ac4e6831f0da754011902a38f9038fae4a8f0f3f46390801a67ca5ee5f4ec19d7f3443f2928378905dfedeff55bd41d84959d366fd8da63d42452d5b0bb620ebfd663a8f1046f691337f82aedc7d2887f7d23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h61b59c89170a65229d4afaac2b87ca7e1422479950a75498207ac3ca6f9683fdcaf3d56c07d9cd093d7c082bab07dc672931361366518b34a923571608a54682921d5f78265a06764c6fb295b6830a681e238032fba55621ae70cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcf69c42604fb6ca57a62b23d2439a01bc073acdabf63adf41feecc3cbfd312d5ed090b7f06366a75fd03ab89c365972661ff85878afd81cd12edcd041307e72313b31feeace7edc367a6278a540d44de3ce3f44603ff66b927f3ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7f45a865e914f389af3f9f5b21b7cb7f2bb6d7cd6fe9660bcc17c25aa9b26f5cc53653864b82b26b5005be36b29259e3352d13a5e0b15f0f9604f91582c9328b35f93ca5fa7ff5c4be4f4ce8202d561a4b2d10fa07b1a70269307;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd736ea3bc98c9b2d37f79eadce449ab630e847674a08a0f8ba4a8fee16366de4060dd9e3a86f601a8083bea6c70b7d16fd3ff231f9c80f1adc7d8a5f5acfd5dfd44eb5445db9b193cf906150f6b85183acde125934edf3f39b27c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9fa295ffc8f08655a750852273acd0a135d83c17ef8f0571a81f4ca51f7c6e49a7e75f5ba9d46919a9ea8e38d28894012b024e520204c02b5739e7e86896186a24183de41d26a0423c702590de83e0e9aea143b1dcfaeff06e727;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7ec5ccf2f8be798c6a051f051728c44100856011a533556d39d346ec5e695ba21b597a182eaf19c46859c02b73e481e75b2c54d9d44b0ec4ec98bd5ba07d8a7a7cb8ff9c5eaacda6241fb3ca2e2164c32de05b3aac42e5121dd36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a055c82554f1dee1689f5cbceabaee6ae173b3cfe12e6087d04e015a4e8b3b5b42dbf17fa9c0934ce09837f3ca39e2b71b9384dfb78781ae26fc6b4fb18b01037e4fbeafde77b4cbc9b82f311b69b9d75a1b012a8c17b393114ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd186475183f1f0ce51dbf5391f971b49b4ee2851daa2e17beaeeff32a8e9a61c0f89ca57e3f99a08cb3ab8acde1bc44bd8b46430b608ef1740824ea58be90dad189ac9d3153edf9f63c14a431fb43679c9cf4b63f8a088b71f4a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20c8425978ecbd82be46aa669af070bef5a7a7bfc92da941e23c63cc141e09d59058e2bbb8e7f1383df56238045956d9fd5f14051e119e1351d6b81c90c56f04795211696eff6d22550a9dbe4c6628aad42b0134d55c180d5bc29e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17685c1ae92273ad58579dc877da9f3a9857faf83d31c4dfa78b415722871967f649c86e9fb93c8f1c81c1c4ff2b51d618e2e3706cadefc3bddd03d1dc8476170bf4ca8b72062736ac1aa4468072875a68aed28ba45fbe8b9ec5fd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6fcf7bd3f5e3d5c561d70f6cdbd5cac49ea65d0ac51b7388edf872e3c84f111104b848337c662ce60446591898731f6e292f144bbfdb8f59931f1058c499d0ca2b64ebbbf0635a033b9a7ce02f9e1f629c7d7da33563e72fef7274;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b360c99b16f5392453eb9d26402603becf885690460752f2911df81ef529c41dbb655d757d587640869a691aeede6696e4a01451d234c4995b8182a20255afe5c6a9f0d2954b7a24797304a6d61cc3719de45ea940eaec1809f5ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19710dca8af1018521b6694f96910d00614216cdaf3134ca208eee715b3d1babdea3876f94061da10715a7f57b3cf935f0cb7c08b3b85dd3f02182c3dc2ac94f7b19fed8a4a1ade92c5ab7d54b82bfeff28098f8878b002473198a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10145806f8fd5ee15df3dc02326d9125ef872e17fdf08c87c54126cf552790fd85cefe1d5b51736bfd670b50817384a726ee900f866feae77f2a9be5c76866607a7c686c843ad79d87c471caaaf10602dc6f842e824f2fa9a751be8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8187ff462d7b3b27891ce2368c0ff2ffecca285df2967014ebcb8538845fcad93b39604d35eebcbf40fcc63ee5d45ceea5b55e5ba6b73981ad7f21f1703903489ff1d9502e0979d077da187392fd206293f61ce6b4bdf6ef601419;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12cd49f48e9ab46c91dc14c19d049d3e1c09913841194302b410dcd1481d32de44e49615f445b53b45a5af70e4b4b46e269788bda3d55cce539f696feed9b1a15dae8d52f895b5db902e39754ca72aa1fda2bae2f30bcb651fb7a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca432e58ba251faef925aef27c781c49351ce92508be9722c4dae3435aefcd1c5832334385cb714f02823ca992d62e1d6cf1df8daaf5737e18d9bb32d713c586ff3f48f7304b9c2eeb736ebcbfef1b2bb75f2a4643d627587a089a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h841e371e536ca5a94d22bc5fd506ef36c994dbbfbd8185c54db8cafe7d7a88653f1547f8f97082ea283ccd69f4bddad95024affad0126f6230dce4c6075c53deb4270cd512800ea0ea3b91e9fa812f2bd30d5d34151e8f4dd0e336;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e1eb275fc7d6313d56454b0a204e2d86f9010ee466f98c1c0de827b79614a1bb156a2b1db6e2f22b43e54712ddd699c32bc9017a4df410ec679a3d31203018d2d2039d2887f9a50421d0b0ff41c6aabedd468c91c57571437bb48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha31e1c89fc5a225d0d095d4265c3d460e28ea6b7c85d50bcfab38bac49480cc07ca203eddb787c54c167b5d7f718d1f95f23d3f7fa7712b4ce6d0db04e8a753052b551d66277337d5ddbd97f0bdc7a3888e35f4f7771f112fdef7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c605c628c33b3b3930128c77423a6fe0c814d1027335ca98245595e7e880b14ed4464284df8492835399f2940aba1e1f840b8556d7662d6f520b020f393b711367b64193c8edfb87e5f57a3b1991d96d1532233d49c4964ec41a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aba13271d1ed35750d39a059247c978350d32c95c06648119d0992d67301db045c9b0645c343652e3601e2ec44a712ed23c6a452d01382bcd448f3dbc472652fc1e49d0dfec8ec9efacbcea629a57e39e5aed6e6067b9c7a28dc33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195850de4a5ec94a5fb91cddded78b086abf0c766291859c8ee2d969372213bcf86136bf804295fa58b5e347a47506b0058156942a4ee10279df6c3e305145dc7f78f535e47011d96af2affc352a20433777a8a7fa6022fb1c607e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d5dfea02e921517ff7730b25dab93c48724ce84068221437daa31a1541860c20b934b61245a583eb0fe5c0d725170a564dd86efef901ac6be9c9c70f2f9c9a53ae4b9c42f62f9722cb597fa91268d9484cef3306ee0cbe8edc35d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fcfe3069843cecfc1454b80a6aefc3807312395c9edf4eb246e5cb8b888b2e363c049af8780fe86f02ba92f5edafcbb1f13f5a26e28a2825a375aba1ebc881ca3fa9a004a2b9d5ec2e070404e0d1908dd531bbb8fb1e3a33e7c59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1579c7e429d45367807501b092438416441c2ebcb1b6346a5492c2813b0ae48b6ba4a952d843a8d707c213f912807d3284472601743bcb90ddfe51417f1e783b597b5feb7e1b29bc829c6f2af20e85e16ae00aa8a622f58d5cdad0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99fcb1b108ce5c54b68387b75bce96f30ef5e50cea533ca109b7f0567521a6df7db743d4471520adeb2d720b58681c38ac70a7584078696bb126132e67c151074e7822d5e16807b1d7f5b406fb898d79ee373c3a181c5e253c1e81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h88456811e5cf95f657d5db46ddc28a362e3b77f828588c3159650f9ae7d11957ba358a467385df2781a82bb4dfcbe8f19ab089dca687e3d5b84e48d675a46ec0a2c7a8cb35bfc63bca1b2c5631cce565aaff688c78c7743933c33c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he12aa67ed1a0c8a9baf741a24474f048149cba38e0c94be52ac70d0a7a5e2686861e64062e5b743a74240027bae2aed2c671441f3037ac506d4075697c961c0009f5163fa58d03622a1e25d589bf5ca6543c0a3663c6cbd1d0522f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfbad9f02c92997a302437a320422866d5c20ddf23a554cf6447700a2ff2c0efc6ccd866b066636953c63ad4a118b78c9999fef707fa81222674a45419d2142cf9f69a289235aa41fa38c370bedbe53737ad6530584e8141657df0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29e65eed84de2395522cb694633f03dd6f21d03de1602405a8a2250febec4d85d51dbeb139f6a2713b8c61af7385d8cba9fbd00325a2130025db3baa12ae297fa46547ef4185267d9af6e7a62adc4ef64af2d95e9fba23e3541b04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142736ac7f616d88f695af3a7bcdbd4f630ceb7f5eb0adac9848072962cecb4c0c4c5e100730bfc34dba64fc63efbe443eaed36f02ac997f20e5c09b20b102daaeb76eb19ce4cf8a19c71c4641c9c64b1d5a5efa084abcae04d2d9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c64c786470b893ee6ce5e9983094d2fa7943862221183b3fcebc2b7c610cb3c2c68780e5e1df114c81b6bb09547c4262b2962c6b432088e649b0e6c6a6f133940baf8574f64538507e366e50e7970cf6606a73c9ff7fd27d0594b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef08d828746e67d622c0e541d4f6bf84a1d1dc4552297456ae17d6a98774d1da9de91a7f02e362fb5591bb001fc6c303b6fabcf8477982c01428bef5e090d61907f9a19611d5b0a25922fc92d73eba98bd84cdbeaa33f5cbb79536;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha54c7f6fa4a0e9edb21bd7d9e943b7124310b4231427b5061004005130aa6b3a05fbdd09a1798e8d2248923d402b6ce261bdcc2a1c9cb1be5a7bf3b2553b1596187f94f3f2ed543b2794e2a3cf9abc09b684d20af1b4e7c2f2558;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cae836133cc19f5e7c8393be46a242f77a4032c32e078ce4e54a8521be28e9ccaa079fca0082a41b9263a313330b270712ef13d7b50c33d40c4fbecaf4d6e8152a900d703219f3dde5fd569ae9abc50e11866158b60af31fc7ef5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37df5d4fa5c7fb87c137168e213c4f3707a73ab8af8c0bc63e0945a615e022e01d7e240a7ee4cbd4d2f3ae4742d75ca6e60421021469e13cce6ce0faa7d21174cc345e6903423694fe522cc61f18a97df063cf08ee57e2812ae82b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b1930b95ca74b531f5f52442823616e3f756154d00ce7504fb962a59ddde1227d1a192253602bff4bcd16867aa36c040491312babb2506a76c15ecdca39dbe06467d9bc84bd1c417f97d3002ef28892eefa159fbc7543790add0ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc6084079f0ec1c0b749315630db35073fa260643552ebeabb9e7a95f24b10eaf5fe16c3123d63fa13241549c4cc9987c7d7778acae8e22d388e3fff8da39ec9a40ea7c78c88feb289fa0e029a5f2edc5895b32be0c3a4fab4a2b8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee1aa7623cc5bd11d387387375539bc66e5a943b8baf421e707701527460022d5cc0f33db5230bfc6dbeb399f652305368760c9a3b16e64b5b655f0564f1ee78109092021b0090241257923442a426af6e61d69c210bb9551b39a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha7f3946ee96dd2f2012079cb3c91c9e7e178299796b6152fbdde1bd085f560db4992812e9af18b22a81ec2b93dc09b1aaa65f8df1087e02de4a187e08345d0f9138f137447487cbf7b74e66e7865ba652f59acabc9f2b1c1244916;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76571c80b11a0af468fbc51ea3b546da4fffad39abd743695188a602e0c871314a2f768b3699b1def796b355fe32674600d71a5c337bd3f16ec07093241b7034e7c7d842abcf800df88f094c8c7daf27a9efde8420fd96f387304b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97611c863a6b1ae7b528ec857f7051e32862610a06b7338cd4aa33c0b18007fdfdcec480069aa1913a7fee4f129c5663343cd093bd61abf6897f6636339d2d0831a715405feccd9f5dfd9e0de447b07e2b60d4c6607278b387a90b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1027cd799b7457760697877809be58543671d2ef407f00e3421668e15894ee47a6790bfd3b8858229da3f4c7fdb217198fd459958de5ac30012adac984a254ed48d2f4c85eecf5c66e5cce56bca1672f6b744576607ae047b29b104;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4ac7e9bbf30ad0465ab5235103bcc509f351bbfeb83070fa1928ae59047e9395498ebcc24ddc1cb20863bc94c44d4c685a3a5965aa81a35fbdf25ac86310b2ddc83dab1c59109d5f71be9611886e9011ac8d1cb15e5fa44f71088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h134ba70e4953340da37755e5fdeea18df7cd7ae821dda131fb915678f5a8e0bf33f43f17ee65e0a60ac297f9e1616aef2302f2f2f210ec3245184bd8060e44854f74395944176f15e9e5fb7a13f03c7f6fc406b6884f40771e71bc9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192ccb54dc6d8ecd32a50b61240b7abcea6c1e59689be6d842ff7cef4dae564052a371a575f045f7ede4a1e97233da3830627ce397ac4356935e380804b550b7720944209a144db2f779da82e3307cf427d80f4b7d8e0720622e55b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b33cd5f37c9635da1c470844e2d58af443267d43190f57e36315b4f3548b6320184789f1dada050f8576c2ef051a3f3e9dd705593826d7edcdca0a6dc079e935a4ca8c3f1555e699ba0a98c5b62fd2c8848a4bc970544119eaa5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb267e4e0d91b47c660f69a2ace268bf4948aa067a04c31fa8613c52f88561970a067d7aae582f607acf75dcda4fa1c80d11190a32c8a8ec4ba54aa55bd5402c1e633bab4fc4cd8aec1466997d6cd006c34492082841627b9eacad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a42af92add0cb45ebae87779487300e84017880d12fa6696a12a17cd27e6ca13aa577b0cccd522d059f7b2ca49f76f592494c19e51110ca8bea9c17bc360bd5e528fd1aff89a29ac81de911632c632dc6bd56eddd0a311f1231a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69be5fe1a79022edbb3552965c3159e4794da3809445edde1b0e53321bb4302524a855582b64b1e829c17eb3dfb38bdb8e3c43b017a0a9e36b590299943342f86b09fe18b987f40fa5bfcdd50a21ac26da356effa1b850301a9b43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1a10083b3bc54445add36221a3bb84fb3737be3f831f2806f04f06069af1b0dede74ff4810815d1dba5906d989c437ebeb786a403f3371506ebfc0c67b38ed466e1d828f1ec70952e08af98595a260bc7e2ddfa4f6e0f11934048;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha87e1f88efab836f2e00a17d7fd461b018ff18255cf2a0882ec34f8329d7cf075e1add3cc6cc717e3c72fb3f72c5edbe81480f52a84059421d536d1ee75a82d680311df66ebf5ee194d2f8566edf745ac9edd69dbc0bbcd5c63f57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha67112907e9657800091f0193d2c371603aaaefd994ac50a6b69381375968fb5318542456d57e86ef2de1b2889cd1e8c36d63e7b6604ef08ab860847aa50d2161f7a229569acf522ce86d32e8a6277655ce532d2d95e5a5b7eb301;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd26202fb29652a6115250753c80d1ccc55b6ae9c63f7666f8b632a956adddecd8a0bbbc2ad1b2eaea2d7f384b109b027785977a59c34e687e1a190bc4b03f149d211515725a3d5237e105c4b45acdb4604f857946e7703dd57a4eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10de1a77c959762f01ef2b5827a31d8781b9ba5a3b33d9a275f106b7e1ec8933294384dab6bde08cefdd1315bf2461e619ec01078cd6e25fded8adc8310b4c45c957343c9b099b9d4deb924a3e1d412615de015c7d183121a2f01b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137d3072c5c4dc71496155ac21fee55fd475610dd388f4abca991cf1718b0a68ef56eff2c8bad0cfeba1a2b5f9c85357d4ba9fb59f0014fe979404b5386ce94431f6442386bf6e1c18e7eeed631aa82c6c0792921ae06a616a20fe5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2532f414500ccdcb7cdd7953f53575301b77750c14dc4190417b120628c460eef839ab0c9b202221682daa5ecdb74434e4cd91bd2a9180d40ab7bb7ee6ae73ac579c0f45439657c825f2bf2f73e03db3d109abe3dade1cce0ef30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h55423ffe87f692651e671d16b89dab94ee9a6fd864175a49f4af8c693164ac074cac16d7808ac3b7b7d15e573037d7a56540d912676795f13f0a94a636436ea155215f4c8cf41108f55f846ecdc6862c5814e47b2ec7fb90dcee92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3035fec2ab6a895c2ca6606c66cb23d149a3e18b9f450e6cd952aebf90177bde08e1e80cf359e40eebe7f9af8b56c2fb214a9aaa5b1fe64fdfb44925da5fd5ca445db1a90d20b66a34d2d790da0cfa5f5523f2c5701a244265c716;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64e22968ad165b6ef25cbee1cea93213ecf1666bf61edf6eb243e4e1a3d90a27177f8f9a41c982c7a11a5138cf07c03b7ec84618ef7158c17073e1b9c81ec04a0d83ed3ecf643e6604376924f939b382588aebbad8555687a4f78a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff78236cff14de8b7c11b44c71b248a66128dbd73cf8d37ca52939cc0b0ff134e055e4fa1b8226f366aadcfecb3c561f417d96fa6e7f746529cafca919d6c8f983bb3712c044d3f4d63796883bedb294f761301dc00fc594488103;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ddc30d1ebd7e7716f3f5ec4a34a38e706bdf2560192a9a61573252976851660b1448446c96335e2c285a5966da20cc9842630cff4c4e0752eb0ae25b1eb842221e7c0cd685390de8c0427443c11e35cd7b7e8bc034e5b0d8aff242;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c2344a5b8e43550140b2e97f4c02264e51b9428448f631aa199aa3dfab02bb68ad467a70fa88a49518fcf473daad699c8b37c3699c9566bae288dd7111af7483c00921fd6cb9db2505513d4ebfed3d64fe402b7648a7e44f3162b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ab047e84c85e23e1e758de831aa9db7f428a8821e812d88d25a2777de87701556c57c4b2a77a47c07863796fa8bfdc70e614b028ea137fa5e4d80033d0404408d6cf2775bb6e9d4efc13668254c14fdf5a4c0ebc1e8946b5b7995;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d7ffc285a6b3f283c99805a315110e4542327e46214f86d8bb850727242c8e0cd9ba43436eff51ac5fe9a5026def89b366c23a478a9ef4e6de2c5a1b52e566179be4a7ba3b614bbe2eade97ef3dedf3d761d956ea63d44f4a077a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h117c2b4713b958607da8ec110657dd1db1f5f1d2deb6b80be84734b4ee50d52377d32872070802c39da58d48cfb3bc151bcbd9dc5ed78c2a238389adc77186f839cb04fdc8b38aca8c9d4f144b946cce1514852a3c1d1ea82b084cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f2427c2bcc59ed59867614a6125c7ba73a9a992319a11427724d6040c213d4b802fd198a1c5c458a3f5afc790903e6d3a5b21dae23c1f20b857ebd62b3a15ce71a4cf07c5ff4ccdd4080e1d7d88c36562b96cb62d43ad65c18bd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f981b8ea22166bec24b32a4af7a28b703851e1226b9c28512a56bb087750d5c36ed713661da281ce874d3f954df7e722b9d985ce921caa9dbc793f4ba83033878fa935e8e2fc0f95a19b53ec978425cfa271060084928c4d43c68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a22097b15f7033615b6d382a6c314ca884ac859f4de04db38131305a5510855337ea5a48050f216e345f513e770c9df71d00b3e2a3d77bdc19f4c9b659ca4a76c8a5ff0059aedee5bfdcc0e8a3c42c67e127f0d404b835abe5e8ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff1eb0008098f0fed7111a1006d83d93cc7eb315ed5511309b0684d1b99cc0684da88f1201fefc31115490fa418dfd5e3b1f0098a12bf1d38244b4b7be1941fec6a730613f64705c16c5575a9f01867d94c3e235bffebc9241fdf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1792a2d02e1c9da1a878e1277740e39216516194b5dea3bfefe477e3ab6c8e01cead67f124d2447d7ab81e884bb1ab8ed67f7abbdfa058fa89c439cdeb7ac54139870fe47d0ce3c152172a057fab198d711f0ffa61990c7e32779bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa5e45ada6bf317e60b1527a35883eeaae593add86239ebf946fdbe6e614dacff039cc77d05e42e2756740bbf8a8a61e456ac4b1b32cbf71ce1287420c6574533c76a227b3ae21e0709817d2c76774e3d6fc1bebb184fc8df7632c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha77b4b55455f76b298f8825edf5dcac68e8797feac169924a3965b4a05e98ba3cf98006cba599a4b42dc8152184cb746c2f0a5762d2974e21c0c503a4d7434dd401a428c8c7d2d249241b222a83e477830113719ec48b14f1ccc7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4bfa07276239f791168034da4602bb85f1af741fb499f8c235145bf7cc9607833c341e2cf542b9ac6f8adba48c9398a8f2e330e29720478cb1baec8bef36ef3296b7174ca49311af80f655fe8c09a1edd26ba35174f6aa586a93d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c73268ed57529f89a8c5f0e703e2b4aecfa5aa82e428cb710845eab489df14d8dcadc26f89fb61f2b38d8f84442dffe9dcadec53716a0de59eca5c659c61d536a631f7348f92a797fbd3c97315440df543560b593caaca4c977c2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca34b14e768dcea628a36b5dbe992c0062660b7af39f46c6db340e1b67eb458a06551c7a656214acf51c8c8f39ae62307fde079e4d5d2bc03bb91624e18b0d3c5f45b5c84420aebb4b9a06c80da3d9f734a087df47f5aeed757aae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a13a09b4475c9962fe9850becf72dd4069de98816bde84853f1b996f81303dd9246a8b95d16ab2b957e6f506188b7e5b682955a3021c55d4c1640151e66e30a8105730457fe8c05b5693e519f47e189b0f2993f4fe997acb14f2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8228fe5644050056a6cd357e0f0c4bc5e02117a54502d61e9eb531412ec3d27e4abcadac030dbfc91717010c18b8c4dea475ae0d94366de4236d37c69bae87547e5ce370f3955f9861257e972cc7835c20af4d1c9744884a5c6907;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4e93e9754a2c4fd17f9c0a48fe0be6af239732da96fdb8e380b10d6c8081edda5fe4d5c93d0103145368bbd827b7792587874ccc9729a5c4886e8b57038843337cd9e1313f812f7b38253492b1addc8d1aa472550a15c103e2060;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129fcc825707b7ca5bf3ca28d7f00de4e7964d57660cd97f52eaf26d88ad4cb740b5c3d73bbbfdf22f7cb126fb8ab9a527a9b8c561fb0e470df876bf6754029ca00fa182294582958661a7335a297820ca87dd7ea4be53b59deed40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d8e42ebe5eb01c919722c1c21e08c62f5fd0be50daba8e2c0f3da6443d0aac089df85e6125548e7580400e8653a6057fdca0def66a120e5f95282c14f7e8012593c89fd85a08621fc33663e40842f28690d9ec48ddfa21e90ef80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd4b8bec8d05ba4d88d5cb39480e7585e9eb188303f58310649ae41743e5674f69f16c849a61545e7d49cdbcea9f2697c6bd8f600c108a278102facc91f6d5f7b82c7f290b384648ff7dc85c1d3dfcb3c6a403f2074f575a0d466;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1df927018ff27da573b203d7904ec892caff2d65a64c708053a8640c1c8c525cc9e1cc962580a1f473bebcd7700609f3aad9dbccef050700b25210f7d4356b6b11baf3b887a548ac19ddb90775371dd77af0326766e32fa9798c284;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36d6499479ddf92666070ae39d6a9fb3c2da3b87fbbe54e7ea8476468610214cb3d31c3da3019b396b3a9475257b8aca903ded08727191b6924590390235194f2887ad21923a2d84b64d59c979d0e23a5a780f8bad5eeb9a069acd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf019f15f67e46554e9662390d3bdfa5be21788036c9cada5993f5a479a3061f05aed47c01153788928f9cd18cfd4b5f809696ef4e74be075384220446711e302cd31735673dbe9d598653e91ceb7e2460c418dc2303e9153822698;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b27a61176b8f96d43a7d6e34dba21e472c57bf62fc6d9eedfd52b6970b3b1690872071c874e2e77f9c2e702b47ba3eaddb948232352256b65c79f75ad403f8626cbb5cdb4757aee652ebd9038125074f216b3c55f5066d44a029c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80d0f752f775d43aafba6db809c59c10075746b455e55563bef40f7069f56cabc35b81b0ad2ff1b502fd91a52fb2545b1ab8afebd69ab5509558235cd3c83f84b8b4313d2b370de9c09b74b26b16157410acf8be63517a65252cda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h304cc791b82c05a161a197fa905f5b8ce47ae68736e62ab450f5740280934c4a66a89f8738b450f0d003bc8ee915f98e05bc5dd88a3d8514cb3439d5273ab200b527c9f0cc7b137efdc7af734db953f720f0050e0733cfd7b9cdc7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3102b5ac6e62bcc12106ab5ce0226b608f21a4798a14d05662e94550841ce5e56fa545e2156b6d8f8075e2467fca47f08d399e65a999bc0112ea6b9a7347a606b01d9dc95f88daa2867aee3acaeb9484d7994d93e2ad971c5af1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7739ba8cfeb897438e9a431035d5eb9d0ba2a2be953b5556fb38a9e078201308f456f411d47f7a9e1ecbdde26c6f0005a3bf6f1b41bf5752bb4bfb8dc5fdab5a9f97bd8a15de9cad0468df5222ef613d9707a3bca08dd3afdd7af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc07c74f294c30d5ebd106db29b39b0aac1ac8a6f018e296d47e8ec93f22f409b2ff98f77dbedb3eaa4cce51ebc6ada4c637cbc35fa74e88580c1d7b01d427713f0d9aeb6063fa52709f7aa1ff8a152868f67bfe3f2cb9653fc3f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb080bb54fe76784e46e9fdb030ec8c969049f96f524f455bd0a12839ba218f92994d342430593ae79e7fed8eb44f72a2082c3aa395bbcea39261a89ebc8d760fd69c8e013b285ba81f85f98746b8d36797c71ae220d666c83ab44f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ca25c7e4fcac6151019f45552a87cc663806d80ebb0bde0b5f1edf21c08be4d332516d5d87b0c7f01440e9396adcabe82a9c34ecf78124f49f548048655a0c5dc494b105e0d2bca70f205e7dd237a1790a863536e47ca37ecfc79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142413c5617be2e01658dcd5c4e02932521c22e9767f54dbccf08a73c96826fc767675b6492284ff2f181ebb5601efa7a9494a2f7875aaf020422ccfe0523a723c9da85e980b435fab51f1ef3fcd339b764ef4bc1c4874ad9980b93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a440ef6212639c8add71f9e0058327bf066865e9149feca38a65146cc563d170b9bc2b08c96c20dd126072e0df0b1ebf4ddb1d032e7af33a701705985312c7c06c2baf64d76801cb8b6a8856a6e3f6f2e45244ec22cfa52c4dfd1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb2af21f54839c3de5f82594f4ebc0c1c53f6d6f9c0bd230c02707b8f5a6d74392a5066b3b0cff20b33be543d389b633fdea904297ef0f654018d992f40288776f6df4564496afcb0fd202cab10c28dda4bdac26922db74c92b86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148446eecb8895bc7b8e0aee91c3158fba9eb40b6bb696de97115f9e4f794991a2182b9864cb5e54861c06d48332c525316fac1ebe588e8b292e22698f6c605b4b5a14851529c0f993c2b950428402642353c850e327560f4ff5649;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1393b4aee4f3cc1c1555993e6076318d3bfe9cac813c8ee1030d099f92a065dbc8562abe427113a9fc529a68d87763a4f65fdf5cccd2de5d7a59cbe3c4dd70c883a85e70ddf652dc4034ffb7e146e138e7b1ffa6f029968ec26e970;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e318f25a79397070571f2d073e39bb7aaeb57ab520b68675cf934d7dfcc0a6ac3606026b697bdbcd779d83fd01bf9811ac4c70872c416c2be97ad3069a134e6d5b49327d9dab7327a6842afe745f0ad5916215ec06be836e752e17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c66ec19a6658ca18342be9a5ce08e17a1c85ec9063fdd59988efa1495005ea6bfe53a5f203d2dd4626e0cd5e0ea82f4ba155b13a3b3cf45f5ee2e4caa9762022ce259e5774155ed5e0163b135c91978b366c2da96eafdb6d7b1271;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d3eb08924f8912dd63dd9ceae4d0bb52fd38e4412d8e959f3c441b49b18fe3c6d1c2c02c1d7c960edf604dcaa454a5e5e2344353e109658c6a7bffa1540a3ea4842a3d19d370436ae2e2dcc9d8799f6829460702910c5bdd7d3f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2a5271f1d6f5f6907af0ceac46453610b15b325cb98870a83aa5c85db42a7862df843685e190a2bffe5032fbdb00d43736b082c22b3e391f2974cff6495fb776d67a8945ea7d169f4e925af9d9850d84640efa124295084ef43e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc0891ed0c5036d9f32aa7f64afdde1d30f5822825ec52f76b02a56755231ec57781c5ce476bf13c0d12a3382f146a643f59d5b8ffa8f835bf4b33d567c8dd7cd0f5373b960cab346fed9c92892c3eb1bf882ec2b7b38458415d360;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0d5c3685f215ea825656805ffcca8934eb659997fc0e8c7963bdc5fd37ad49b3ee7566b18401aad7733bf59500a018bfdf99d6f3910d651178f99883f7c5f109d56013e9b2fed87c59fbf23fd91aecfa2005e2b267d91bc9df2d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1221bfcb113497b6e1636c63e2d26b22e841be94e8bdf6cddbddab215c94918e30b4697954be30618404864f62b86ba1df7bf5a72ec47cde00e395bcfe157a353673d9dc68675c054deaf8cd8d3246da65e4b4f20c1dd4273323155;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136c2257c2a849fb11a2aa59dae0b2a55a36ed489577553debd504ecf719d5a092275f87d025be300354b2e95b3778b8b2f28cee6432b44350c92fa3aa2c47fc1fd5de4dd687087fbf83dd0bcbd3e49f6f0e810c689ee5cd7f260d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haceb0234eaa58332b8892b8fcb26859f2367017f55b3ebad480bc6ff371aa94d54dbb1409002e9e86bf95723fc621a0bb9260de4271a9d7c4b2f83f135f7bdd713996511f1f2fc167315d5f36ab1aced30e2dcdf6611f6b3f1cc9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4e973c9a1d03925dad7e82da0bbaf1c301ebe4cda047cc08524a2534a5da82341ceed480ad31e89fdf5d25c556a8bb3bb0a0fe41eb765c073b0324eff2f532c2a0d082ab5a36c94f79a833a542052295a48941b75d24076eaae15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hffa13d36c2ce5648196f6cc616439b740fb2aa67a8b59e26a24bd233fca5c8cc9c09f72da62c0770f5dfa580e31c3155f0986dec8409c3f2a911e1f05daeeb6782a3bd27d21e2e8023bc125aae0945982d1e019e3622f76a4bc3a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9de1017efe1e3e631bac1d0fe52bb3c72a1936c5c335a2c3e0c316248e1838ace9ffa7d3ccd539cd6df389a5fe21f811457334cfd543c11142ad729bb61d9accb6fdf73be7e47948d299ecd1092b22113f2b9b40da656ecc51bea7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10c7cd96e645459d96959f6d78662a0cbf05fa33824cb862dfdacff7ca5d1a9ffc716d5ec7d2daff248f6d742388519c686802d01eb1983c832b410b4d855592675c75004264d9af254b38b1f635d1e3e14deabbce124cb2fe73cb0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ec71666b71e69dada5511c8f0fe69cc1a69eaafc2a537ed3311164a25c1c87ab83e004b5cd93ef2487a65d8ca7a53ba29702ff1adf0bd8c6c9b902ca57d4cac954fee74fa2eae39aca5722e0a17bf24535f2655f588d43eb16c42;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h433d08ac32b894b8cbfa6d8ca65db15ab2c862295fdcfacab4da16cb34d0703cb8a2c83bd180642b415b6d05a4734bf760dc0bb459a0c21f0db079f843de7503c0a733737f46e16e65834430ee41b8141f1e2f5835a2848792310b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfda4c088f02b2197252fa89b23a3bd3ac7a25d7f535b757d3eab14cac225c04882d9f6a63260d2db7561fc5e1a42f4640b9f07172bdad4b57e1ae2ed54c4a032e448af1e51a2dde4e32cf6f904380131f29b93cb45db543741a611;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130b36bc16eefdbdca9d482c3b3451a97f6eee3a2fba7c9b42d72061896fe199a3815fa18e3d4f37d1e0e91a60ec48d093073d26b0f3e2c6355752960aeb0449a5395c8cb927b04b1ed15bd71fa25ac62ad086ece50bd86e17d255f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179c8b9aeeec25ba8c57caa31bd977df36d9273debc3e5c8fa70485a4568624ec86d70c7d618e0e9ce6eb1ca31e845e6e3e1b666aeb8773d45b0a1ed2cb50f65b436e480223497d7be979e5155ae95bfcd74bb887ce9e2e68b37bd4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17bc7dda6f1886cdb916dbca9b400fd4debd0e00dbc5b6d279b21e8e656f4856e4c9ac215fe0e151c790fbfa516860e4de6e1d7a9860f4c9a7fafef452863d7ef9452390ce09925267e5b1a747d3b3a4a052b1a8c967bf71d60c5c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2c9aacbaa44db322e13950b1d59ef007ffab3e045af8899df8e5b63e5c68c42fd68535bc533b2ac71e904b4289080bab01ed46b1e054bc5ec7f388648018b08530616479adbb15c2983885b77831f3ad3b456309e6f5313464523;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af635a932271e6abe0ad28db389b4b7bf2dcc9545f4f1169bf571371b1a969458edf386977dd77e34bbc18818917b6ab5eab8da67a0a24f6ed10ba6153c0e18d72903c80c09cf994d22e6cb2c6bc60af6887f7de862ab27d7e3f55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c65e408708ee27773766d2969ef4b3ba97094ba53528aeb0ccf00010e9878fae9ea214dc89af4a25912ad41a3508a720ee28d066220c27e958d4acd21d09502811b5d3db0f499ea62be3d1f8cac3d17904cbdc181cfbf2cda9c956;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1185e1fdf6d0bcd3b7dfb2da780e90a5253df69e976204b0aa20557f616d6307941f6e4e08e1d1d656393f276012e736a6c36940cd0c63d09bc1adc882fda9c7b2328aa104b0ebe5937a783c69fd13fb38667046ed9cb1d2bcfac36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb87d87cf5cc7b67292a9d74e5f43401d1e20499086a1bb17ca542bb2b18494ca24965bd22edcfd33f5b72e1a5242a1ded4bcedbc342bbe30cd3cc87746da28b370bb562091c6da0a3f3cb4db675cb6c4f615c1112c1aa8f8cee3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e07b94de99e33a9ded1c541330fafa8b5ca9880cfca6a3fe199590b3106eebc336399132dc55d8b8ae0d2a4890cfdf340aa716c59f18ec7b821be68fce7a686664b1625f6c1e44c525cda7ae9d092f72baf40be352b33e4774f60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19040eb13e8c51b8b4f088a8d7b6b224c0e6b7221486bda75dfe8ef9424d8f0c6645203b116c1b3035540710eb56c92ebd70d65b21aa93e7167faf884b28ad30d2c940f26a5c95690d2d9fe6581c85f4bc21463cdbdf71b3189cd14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2cbba38072f18906e69d03abeafbd8df6b2bf56f29c50cc87dcb8b23ad172717c369e15283324c5652b8cb4eda32c69cb5d581feb4422ed36ded6920ca81336ed119c6339667cdb35de878939ce288e6338835620fd6b48acda93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a52bb489ab0930b05260f3402f3880d0b9870ef7c9be913c097ca857e54548f9a48d43cc47abd228601ad36c96e8812990fb36d90fec3ff04475b4e20e780c124f7fea641c70c888a4a87c1d000921e26eb887d2e46ac11730507;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc50dc04d9a8b52ffbad485fd1e7f438bcf1ee7a72b8afee43cc90006a435eefb28188e2160839b262a9108f4522378313200f0e6c720e08d5d375d6d0ce9d6939801a7ea8540a2c0d18950880f3f0dacff95da4eb1e218f5a5810e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h28921b5e23cfb6ad87e2c6cad6ac29e7c49e2830e47c526828b7728f8dab9549eaf926385a1e5ee64459a757d99198fde7f4e0147d9abdcedeed3595024cce89cae32b5393da1f6a8a1f1f5e552f95d4c8b9d9de89326752641a44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14807d72eb8e46d0f93a4eccb6f469502b9a34fe401b4203d4deaef7150df8a930e36841943be7283cfc9ed61efcdfc18ce99759fc12a934baf0e9ff2f8df45f23b9971f573105b1ec354f801a82405bd649858964e4dbd252e7ead;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b4328934c592e0d243a9b346818c3394d8211e77373990b2bafafa1d7cd1b51014693dfae9f7216a2b1c7b7533bbb833f76ca45b8f9783e47b852d0f3710dd9778256557ce4a43f3051db4eb1be52b8a9057a9d7e78d8e7ccf497;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11730f7b5df1464ec201d948500f16ab2536994756a24de8b1c12e7f2b1e57cab3093dfc308bcdd29af14f49800b3613293170a48731e0d775a9f2520d598b3e4c30f6bf66239f137e481bc91a2fb163d9e9fbc051c77ae3c692cfb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4df46fdd6ff1f3f1a37eb39ce0cae4bf0a4b97c09bce95b2e9da98c7e69ed0bbe56019f1893d1e05f1e92d6275805a9f780758f18748aa35c4b65868b34c74497292b6ce0ac2d03601bab6e6eb4c68d44ad1847d23c90fb5cd67e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e0e25fc858419fb84f645bc8d9d87a0d4c6a1e01672c3a9c74ee412051110f0a3138ba2e25a0261ec56b16ed12d4ed6bf7f8d39a8505851ba6df8bbd83f3001b4913cd0b532f4faa3b99c74662abb75c8287b282a905196587662;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33a0234b55dcc0832216f9d2cc7f72511c01141eb90e2ed67da9cc03c743028a15f14f403f44061dad386d4474e001cc73c4a7a8345d245b812c0f30c2fad49a9c0816e4857113a3a8e26636fca84451c199784313f80c23f94f3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d07b4e972e1e2b7f11882006b39b89fdb561cb6889d5faa0907fb4b3bc91d16a823019e13b69735421a0325bb0b99706a49be76c56e0e6fd984848f6f06a0b0f248fa9d86e05bfdb11f1617974d969ca5138ba499c67e788ff8bfa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2804af0affe78ab45ae37109ea89df35732d9a9e35826c506b6eaf50b42f0b3c822e147bd0a8ce915c9e0e14337489b66625b54800576c453b262e60a7b5526532f3d891fbd662e643ba590d5e7208d93ccffcffafef44b6c99af8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ea259fa5c20b086cbd191a1ab47f851a2f1f2d09453cb85e917b13493c19fbece0cf463adf9410159e03a227fed3e9242ab30f2d99934faa4a16f907bb0ea183eb60f9088506cb9fe1e2a5cfcae43ac544c9dd67fc09f7700a901;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5e7e26b4f7550605de7c7ef1839d7f74d8590af2b23451d7c5cac0054c411f2cda36ed646dc1983b6fa85cb4dc7c38223456be20204515ffe70eb66c287d66c46bbb137300cbafafdbb5a1699892fc0c1bf0365b7c5ccd57f4b8f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e1057909c5ce08c450bf118d7f65000480b801acb4af158222c69697e6d2066addb42f8a3948691df03e7d4ca519d64441245ef6c62b3a2046723050f024b254f4f882dcab31ac63b37e0b99a71c66e1efef2ec1991bcb48d0b33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123453ee23b2fb7e1ce1aa790a7ff794f0a577c1cc9c1f68a3870a4c24936c814960cde1820b201695d88f9e3b837afbaf373fe76d7b6bd123c9973ca3af218170e416412d690cd278b24a5723911b96336e0fd159c28069cdfe7b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h56c3af9612db2b47fe6686a1c8338a244c2a717ec80f5f6c1c762dac32a3ae79a47b1ae9893d16b1bad36dda19eb86bced03f4c47794229117197b4dbbbae5387139b0870bef0652b0ec7d4da3664dafec9e30f05aaf26fd5b2ad0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b6c59481c58009c7141388ec4077045f5ed68e87f94e11848f68323ae48f89c3835fdd8f4827a16daf73f280f4be300503f6564ec3c1f40ef15154cf251bf365da2481b45ffbf19810b77abaa867265af145182edf50ca4645051;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20b821c1fd32dbaeed8aa78f93043597a60b8375c1b48dfaac456b6951d07273420b38f42b9bee4462f57e2ce733b65ba27cfbaab12cc4a2641ef906ed83f77f04c44787599734ef3b9ff905c60c957dbf1493884eb0611b8d8b49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1474a105a1bb0025a1b00a85f2955e9b4bafa1bc4c067ae382343c4cc8ebdf4eaf4c0401e5a8f00c7f7198967917fcfbadfda71d92adf02e681a7cac431cb2c65bb4acd350be99fc6c22659db031e18b617aa5f248d5be27703b008;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f1d668a6c7d0668b4c557a140dd7168bd1d063190b6586849f90baef90ccf656e8059d09781b62ff3e9f1d9a64893d7d6090cba6655f4800580ad1e5260a24f891ac15e856d2b4e318fb793b8437d965dad165cb91c6c8ea04d21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7cc4c615b4bf1b60e9f3a8b473f89789fc3a4fb0dbe1669a27ff737941d5ce38bac3706fbf794e70d9458875cd275e004ff350ef912cfb1a38112d98f71bda2abf27f92bec53cc2096b1dcc8f2bb08d44e5cac41c4f4d3684801c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h198a77acdd4592f890033c0a201871445012c3b1d70713aa883f374dbf984760a81fe3bf1b5da6cf63c48bd1a8870159d6c18861e1ed29610e28cfa02eb1184c672edc1c3e55726555df7dd3d3b9e962a1d53a205f978c2ca40f428;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ac85fc3208cd4507bc07abd863cd951432291afb1d7ab8960000816ec47295dac01dfc19a87b4fca09948f0f6b822d2cd8ec9c81680a4cf6a600aefaddb2509a00ad21155c1b98456e240e5b60db185dd19722a3fae3b85fb2f6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h82b025da3216ef5aa2d457cee8d9b275d5ffc65ac347b9a6d11ae2df85867809433151cc8aea66e4b70fb009b967dd5a972aef4bcac1ecab6a351e45f637c9ee435bed26b6f2f0b7f464b42fc30a44631dcec3e473818211a47c3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd986db92c7820658b225c92423c733baf0acb5a796aafd140a743aa4366834d177ee5b127f1d06d34cd75d23888603fe73c79d64a7b1dd801a5e1f91bdf74f1f1c0da47973367f04fcd02042ef183c64a33d92f91efea282bb6460;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5c4ced871bbc28b4f16d57a1b1b7df6ba8d3ccf8204ae71837d7008310edd03a791856600456e3c132a91b637ead33436694e4d4972bec747365c7a7829e0685609abb52b34205eeecf0f2d5d26028f44a59234deb362c1b4a76a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4821b870511d5a9c24a5477243006dea14e325e24774c5bc4ec1a3b26c93e1f04dfd69d4fc7843279cc6425f956287f823aa2c1f15e5b8497cf62f59ba3288d9997f7dc8eeaeabd08a5719890c708dd047ebed05e9a21295c0e48b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6e8a39ed7c73c044ef50c4fd67487d89e4539f83235d786318eb8a1a466533ad32c9611f06449df7a0c395ac873e077a6860bb29055c1c0fd1d0406dd40dc56a3f1c96d4c782c68f09fcfc0fb694542b326670b954158cbf2f676a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h622c76d6f217f1a409b24ded9e87aad64dfb04041b3e61b1d63bc6bc7c75d422ef314753dd2a444792c73e3d68c99d32148de39c3d39d09eccdb7e1d4e2f934a81af5abc8f0889b3ddc5649d89cbf5a0bc24a44989c0133379ea13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5f377ce9b8ecf933c3e5e80adb59d787a657f26a357283caf32894ae1800f93d5e0deb6d79d050c3fb81f41c74befc08023bca74d373cccc419735fe06817b46f24d3b80588447e7723753b0d22794e9bbfd4eeb91fa0af05f96b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35b3bf2acb3be0783fb412b94cbf1d1e92f07f3ee9e0d78a1acbc2bdf87678d5f37f60f45b96a7de3d3b09cd1ce2b7f5fb98ba7ee8f3226f172c9e23f121c8386656c42a2c85b1ead2a9741e41d0104c605201c6fe04a018255d87;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16abc159a25915e8875b404884ea72e987f3da148e336563135f0bda0b6c8ebd6269b63181c4ad81c129313f612473046b632ca3988de8ea5d6d883ca24bc8c16cf38eb7c32a8df14718fa4d4f476d44025439ab08390043fe8852e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ef5e027008bc6129533db265e7e577e8a1cd81a78c5b92932dcc5e6973d5fd2b1bb37766c945c840f190b22b97db2d1f012fc75c9e3a060916ddffda6ccbaf5405f7e075121b2ad9ae290cc3e7222eadc145920f95ae6eb03867a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'habe6e8bd345b4c4182df98a5c4b7da50c791191b4acb60c91ba99a7dd29997dadc531561f46380e14063d5b6418ab496fdb499881f4aef30288db8a6bf053437935cd7af002e8ec38e0a0e9dba77d850508e4f429307de8bfbb98a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170d98be6633529ab76fe608dd7000082e0c18ba22d875f78307c51f214317ec29994fb609496ae01f098c768780112e94acc0b113d1c679dbade4387581fe45766edab33e6c185439b51d9887b50d007d1f9cd1079c1533ffdf9d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd0be791d22a36a9b6c9ce27d4956332b5caecf92b475bc1ea93593182996b19dda9ee690f3571f772096af0affa080fa821b91b2227d705151e297f07254f2530863b70120debb65f3a36f11016a9ad527b173bb28372c918e1cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143f9693bc836eda268564764186165648e7440924477e51ff56096f1a651aaf5b46ed123bb6d2b6dc4c67ee653a570a76df98d4e06765e00e52a63300195c8c470d859c37c5cb74600d719b3e2514d73951040e8a6bef8f84d7b0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157181f8254a84c5cbdeef1e4fbdffe8b1720a59f2966b23c4933597a5d9429c9c001b97d32530cad2a518e287b2c56aaf38ba59ffd2179bea76b01b41879bd1cdea175c85b40517957f3e16232ae4b2fb7b2b2c42ec9747190071d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f4d16434dea4beb60b1d55fcf42c75661bf83f22a4627cdfd1eefd2a2fe7ec84b4d48683891343e3f210587dca18708a020a57ebf04fa85f818f46b105bf4c5f7f3966f22972226475324138399b08f649c4dca75f37a3be8e19d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ac84680c341dad5c18c05dcdef777f19f1891c9403af7d01f5307f2f900ad653e22ea4fc7f060bdea18be7ffcf3ca01fef8242aec4c22d4759f10970c5bdb13b29177692bfecf6ddffec41bd47fb1dddba8e605a6f3eb094a5f5ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e973cf69d72752f7e595632e9d483309e7d65279159768cccf2faad2f68b3c4d5656582b9e422f98cb5baa63889efeef8f05e37092c6450f602f4e54823233148d583117c2818f50abf181b214a78d39c733a5bf1a88cfca681305;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ed2d554e5793be0dc75a7e27ee005f507ed176e20f23458ab9b6cb46241051217946418a016b268fae0bb9ac64daaabf7512415fc11026438f620a1a9155b4b0de51d9dd3c202fe8df994e1d3816e35b98bb567477a7d42001130;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6da95838e7e000ecb7e15cec63161e3a56f294192c54416b90c49a287faa346a1e872fd8aa5389cdabc4e349d33073f0d6795f3478ec4987d3d916ed2a9a2cd07d8b6150a870e278f231e634991a2c8ca2c748c6501c21d4401d8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e122352e683b611000417bf9d47eadf237563c61868dd2b34f23f84e516a2bbb32aa1cfef368ad103c1de521c63b5eec4a109358ee3ebea3eabb435b1b89d0f9dfa1ff7488dc2173ee2ce07948a43e8314ff00360fd3e7ad8e2fc0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d6f391ee248190b7a3b17675272ccb1f4f317e5b3d132dda0d507119fc6e8eab63a59879dd6bf80ef10740d8673013d1d3cb609ba951627e1f6478b99cd2c4ba90b58dd61b327346482df93c00b2a60f4083d5210dc11c5bb4570;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c46d29f12efd047d542b97b6bd2ff2416fad7e5a27d46dbc98c59bea98783c6c96b204dc94f6e5836b03aba31ce97b6cde1e7b7210f598f38337429bbb6689796b123135e46ab092f81c9a28106e3c080c35231ab7cf9b2331f235;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8fcb89e2ed12c27810447030637dc3f72d82690bb812713f9bb6d2010e066f464154c028896095b117d627c906da749db348bd52c7ad3cff488084e7cec8247dd3f375eba6be5c8acea289b190e03d7a92a072ccd68b52c606ac93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171e8c0c8328b5aa6145c54b6fa5e18363129535ec6c6f9c6670c0ffd4f45f7c4577d0707ab1461fb11448d9c1ff2bbc8f1b68e7bf4c8c9758c98da7939128cc2f2e1757d49de1360e2e46859c667cc7bd15bbb448d6cdb8eaec54c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc7b10bde88f45c6d8300610387c50067a259d01114b35d38fce53662ee61aa9c7e881430800c85bad18763cfd3b59f4393bc6bd860da88d0197f9d2b49aa47fe406be9c59b57e2ea90e36a716586e8590d8ec0934bbab41c51625;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he85444b4973e09ff1cfaf1d144bc35b51ac601db4eabdf1def8f69824b15b3dc875677b5f49a797034cb7f9d9fc495e491263f1b0e4ea50be2c117afd5b445ea57405f29d3254ec54de04b0db96d953a8d4b844d5e479b28276234;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f495fd4249e92350a318d614c0aba03c06741cf942588891d5bb2f7955bcda693d6dc39a8423712e25941d0b3b5fbe4ef636aa06d62b9e0a531c2c9428ded5dc70ee3d1c5a5481f6f3e42f3a9b977e4a8511669123e2e9f6561fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7a9b68c714f678ebd079d35590c9bd9f27e66b537be11321efb34c46f5c0535f5e93d0feefcf2726b644679ebf8950baf8850baa20a27c4efb0ce522519cc85561ff7cf832e16ba322b3ab139264657c733b4e291a2c29f6e36de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104f1abe2f7d764d680facf85ede73a82596ccd3ff8d32cb8950c577dc23e1be06aa234982adef1859b2b96c513a08f246fbefbffc2c86148d824773fcd96fb569968ab96e8e13c7506520a9617c7184908bf73d07ea6a4742649ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd4bc4fc15ab04172931eab2dc44e7c91f63c8cbfd1a18182be428e8796912e78d477ec00634c651206016277f4220cb40c9a0db78ceccf9f585c371f4201b3369ff18a068ed97f65b34367a5dea2e7f63619e463c97e2ecfe5d3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e8edb00935da0c2107577cfb75c17746a6e0ebad3361cfe046c85137723aad2b469ce4783be37c59eb7134892576d5584cea72962dab83e410ae401b400a21980f9c2a870e1792a1be17951ac9939e5f3dcc261f60f0920cd53b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bcfcf4dc63dc50da2457ee34c0eeef2fe3f167ff14571e21974b7e50f0a67b73bdefd7170f9d4efd700472533cc161b3ae338d5260cf8b1bb1f7bad2a62d446bfe76e8e2d095aec01f5e3ce575637497e41d6b50cdc053903aae85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171591a30f890367e053cf86fc7881ba7b66ed5c87fd20093c7b62ca1afb2fc99ced3d3c1ca976055119826fe094983fd1e3598d33d3ed0dc27c7a3beee6da18188665818dcd669883bc54f58855e47e8a158f5388e520245415fa0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c140747e176d7f0fb2b2f3ba386cabe8b2a0085d4bac349abc0dd73ad07d93a39afbe2b9e584fab7743e73ee403dbd7b348e33a4f4395f6a6b5e3c2c246d0b94d470f41bc8f64d4ad6f3e9c5061ec594ef01c4cca1992610143d53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbcc10d16edea7eebeb1c2557888dbc1ccb3a1847eb19bbb5d700363428c8b01f61a5f5f0c5e30cbb23f0fee9095d95c7f0480132dc1f706d52ab23d5237cab1a2f5b59eb48a52b767b616e4d77f35bca651261152a723111b477bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12784fce511fb351ba12c5e8f8ca986a592ab27b73489b16be288703e7d402b6d448fe5f2dce0130ce03f83cc52ae879fdbe4e0dbf275a0ceacf475db9afd451cb928b4711bbca7371ed2f8b0c3a9769f004f0d615b59e1d34ad2bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19af677ae4226ec25a98f79797eb0b798b35a2626c672a4f3496019f7f4ed54417ccb3b1f20e4bf24b61eeadba2e82a886eb505c2eea4d774420e640e43967ea5cbba10541f2dca491305cad8fb863d9a6dc181e435a2794d5be231;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146dd71e8756cf5c9f139eb61d8903151b9593e5d13dafce6a0773a037a4f63ca1985de606fdc3cba1cd23d53ade06f1c4e761d7571e77a4137ce66568d1b018fc31b68e75cb968962c7b5531496f1bd9a4a554a75c45c0e3e4acfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be9a8cf2dd226d66d39fd32ea7708ec6f7b5b1e57b79a6e35ef1a1271e103c89cc3eb8f0395805b718a695cff95675236c0cdd52e872e70698aa6e264aee75dcd506806ef512dbe6b26ce5e1d5cc18d7ec95189ade9685048f5378;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6cf5c43e6410f41d0fe31754b388a88533fa682c6fa4f6403f8846e98ffe28968183bcdacbba0bf3f8c98894ad5c24e39835956a321c084d3c6b1e8b26ec37f78bbf321719d81e0afb32c5fc0524d3e1ba2f5bacaa81bf16e792ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147a486160d0283efda0f029eb57c8c75f13abf37d0fbba44af8392137789981f592f040a88a003a99a48d9631ac11631361bd6c4d8e023c59c1722ba36e03a14153a8a65d69df622aa17bd17bbfc0bc850a317681eba08b3100929;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54682e142ad2c36e45aad29dc53480587058f2f7f56c8e7a38f814f50e0fa1353139a1660c696618ae58363c87044c39c95c8d144ae9f485cdac804b3fcf8e53349fdd29a8dab4c760219e1a3fccb273515e0890f8c8e373386889;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ca6e0e40bbc9d6eb7421ed58b0210afd3b897efead5e808713dacf4a30cd03c08f6827e1f4ed456b9afa5b42edb0140455f7a59dc11a01cbebd62fe51785111a93552870e7e05edf0e6438ab183cd9b1f14024e9dcdbfb98ff273;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89b27de61ad3b7633aa144559d8857f52cb6aa2f734c7af806bd157401c8deb45db48de1cf09d3bac6fad8b6eaa98e3a036e4d3b1574e8ded1b6bf19be4a83157ceae47974f8ab61c0db2f86db68337fbf411fd8945cd7d4b45ab4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c68c7f39e1483030540d7137ae660b9954fe28b115d5f3c94db2a14a8400987fe33357c2d6b3347c9ad0cd3d92672e67433bd359bbe6ec4a47f55c21743c2e3fa11c10ebc4f9e5929d5798f5e8a94f7c3d36fcd6a503ed866eb48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h100536ef3c26e5f373ce0be84791817a04375f8f234202563427a3ea9798bd0c3d8a963426158d76481b765458df336e9a5f47b1a622ed8da424e2232fa3871ba4153b812d3a20ef6e4dee134fec9b73db6f00b80738841a8aaff2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb5e24570ab9b825c454afa805742ac8ff5f62a085a3b6532fc3ed4f71d931a8cdb733aa7b8bdfa67e74ef9404467b95952884347f67aa24c22a11c024adeb702acdb74c5aaa7f53dc9a9fe01d53e74335f3295ad193e884fa5d48b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a2e7f4c6bd473dca629754395947d532ed23827ef0063b7e7e9d9d9594d1445d61653a99d14ff2235b164f915f94ff994f7491ccf90e88444a8e84aba72a9120c1fa40032571faceb95150d00882d93780ee172f73b2f53053f41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14cc1ab04d14eca1a95013f7d4b37051c555e305e93360125641822c07b4dbf4db3b60138acd2c9e074067ea46bafb9574ebf047347dcdbd042007e70cddc5f97a43ff45a932bef85fdf14b0d6f42d5a8e89fce5d54eaae4ec843cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192630d9cb3ed4c05cc455651f83aabf4331a4bbe116da68d49385d583aae007d6deb3ae633ef7440aff601ab796c450f670a076247953e9d8ccc05c7d79847a8a1fdfc6aeddfc1fafb6e209f24b493dacf10f92efa06eb0796a529;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb8f065027c09ce3d50e9b3846d282975a0fdb788d857fff5d85be8db4aa13c7ed7bf177c2eb570fbcbc135f234dd30579a30ebe14576bd0e88323618f2350740299c0bdb41f4bbf1d55599c68ae34d1985deb7aaff432b18feca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1efc35f33e862fadf58874d05c09f38889694811777a2543801c369645e0f821ccb29d5b5a1b420ec34799c7009564f74c61b393e6266a67e2dc875a1cd2db5f4417506142c009ef2fe5e3b006e7390eab0d9513866ca600c81b9b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169bd76f2cd1748fcac43a29691c8e6b410f9b0579e4f86bddb86f58ad95f03543fdb46247a4f59e4669614cd867c6f66bd8c5b26678278f54a6df551e80eea389dd434a4449972822bed4746ea5c974bf298df9482680185961338;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h458d7c95a14c1b446ac336f01b689943535f6cc1a7c0501f95c3d704ae0412c2cc8ffe50b0acaf04a3c2108f6409ce90736da58b03855849326e98c4edebe6e3f66bf43af4c5f4911913285778b2ea68b7ac8af813a1f0b78fe7e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187bf88005d5b9d8b60b37c20daa3629ad3771730405fd8b813d9cb9208dfffd6e32a46094dc2bac0fe6a6d201ece9d87cbdb89f292566115f425f9f4465b1f59aa5e2309b8ab89a0a73c73a39a0941124a3ecc7afa24ac07b5aa1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc5b90ab2667fbffec5700239794d79ab39087494fdb5976c7cdf4ed66f86502cb3e005f0a771aaf25aef1eb309aa7be3e392ed51052b8531b0562c4eff0951729690ccf1984c9e22dfdba24ee0ac545fc97b1bfe4a6b5a7b26ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3970c05408100e67a1f8a6550beb713deb0574ecb250c26bf28bf121e193c63d626bf025d9f321c910f0736e9440ca4ac608fc187f3a095d18b52ed3a5ef9237927443d5250fe7988db312edffcf42f8ee35697569f0c638d2ff43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1badf367430c200f0ad1b99c9e3c086ae3142b074c56eaa550a6ef4d6a24bc6bcd98cf9ccf9b359ea103ea2f00c17cde632ace456bd0e877d9abcda61f1dadb7aaf25c8e38efc8a47f5b19dd0c0f854099a8352b41a92264a4a0603;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7d1d63152a0a551cca1c85b56395f78597bcbf263bd8c9fb8ea505b894e293fb3ca00b6dbbdc054551836445aa055178d6683627989d7fc56fc2d537ee0073b76fd1ef4f9f063cf939ea4b3d806305409a629e2f3406a1acd36e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14493b63fcdf22d90ab2dac205c547c1fd40607f0540adffe23288c7f8879cc4456fcb9a0c421788538c3baa6098120c44fa9c6298e77fe084abb26b2c5c5d06d725e141cc383fcbb1b24b694a830d28adfec5ddde13d7723bd794d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36e19117d407b9cb32aa6f34e5d0ec29db31d49f352f933810ef3d0f39f47dc67d0efcab706bd1f5b6359e62aa6dfbcf96f7ac18d08ace8c0b445fc943d58a3215e0f5160aa5110176dc70a7c62f0273ee25d8fb1d758492778771;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fe388eb7c4ee8a71e308ba4a3fcb2675b396d94e7ed64798fb2c0f201cde3a09799c20a28d2ce424b6f4be822ad3ead76de644a0870614192f1bda92e62be0c0409d097d3ddd8f6ae49160890ea0ff73442360d18cdde9aa671a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e51c9ce484a01f6864fbf5971193a56654093be47125033dce080febbf4b7c2e6319b03f0e481fa1b614f597e8b7dd42876052a032742014762355b4703e13d40d3b2ff1676c04582fc5eb888682d058575d93380ad1ed519ae1e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc6546bdea1473a1dee8d35c9f0a18315b5e42ff6426aa54dc04cd467f5a4b4f855daae38e0d7eea4769cf5e31e95d68fde7054cc8d234512d54140efc6d9501b417a6a14f1676c23410fb873b75a71ece13d7ded13b539696fe150;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h52f323a7880183fcd22bedc62d7fd1f5e90bd885c3fc092974b4cec6ad1943c95cd03528eb9314d21b8e1f0ab7cc4f357f67989898cd5557f1a1998e2774a1c793153944fc75875c79d9c327339b1b3c44b94aa058c2ae74d990fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1779cc2219bfcde4f13117bbe5223e462b26601760f407934671c8c6e7437e9c094e06cb9d954d85305fd68f56e776e5e71df1451882602dae814ffc8cf0743f85020b6f33c28e9b4f38556ad229cfa9a4102b5209d225a86460369;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e58dc65f560a9e6d04cd36ebdfb2a5a53f6a21f4ded05951e27b9fbaf0cb3a5f002ae14001aed86d5b265d92e1a1cd8eb12a4971ea61fe202667fae24be41df1937cafcfb447861bae80375cf59726f1a1acdb36a0dad625eff2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb7a6f4d8cde6e63292596eeaccfd2e1780df55c49afc992c2bbb20a99ceaf7f4763e45a08ef5cc022a3b359e02971fc4cc8d97debc16827915246b1c0046901a15b67d34cd217832ba2a243770e0d489fc9ea1633a2437dc371b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f79adca8b33e45c7515fdf40f8402312c17fb3ddb993f2a9b7da02ddf3792081fe8ed803d2107e179843259215f7d3bf13434654abca9808a6b9839882d2524fdaa301253d25b5860f096347e45b6894c52ea5d03ac233b9089d56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf989d5ca322c3b28f5e07b788206efd59b8401535738a2d9a340c59f6fc76a6eff8f65c90abc2f0e16bda18a53f39c8edd0906e0444b1d9b6090e5cec1ecf47ba2ef029fb340c47d14516c737fede7559ce1057e9556c26e195a71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5c596411f5ab58a1d7cb6b4376ae11267b478c9fa02fa367fa08a117bd1cd715b84c86ab3902f2e939fddd9f4f180ee8e25fe21f4bca0f28fcea278f3ec67e04b51521aa53ec36cf2641083dcb3403ae391bbb93d9a0066f1b602;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38f9e525507d4235fde7395f2c6e6ce7b569ffeee03bc96fa4e1387547e0c551376709db1f604efbc8e5857708ad9b3fa45930146907b7d18bb86f2b0a9a8bc4f3c17558509fb56a95de44673d5f44c67f4fa253b40fb9b26a4e32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d87e1a6cf9022518a50ae1e7c29d22e8fdd5b8b19b657e6083db1e78d05e2dd7ae01560a26393d6e7414886203f3d70da480dd1a92ca08157d67269e72fede98f7c84b3c2b15bde5a9a523390fc81723c03f67ecda1ff5508c0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15fcd637398066634312e69b88d97fc2d3f24d0ee5d6993d66fd683a66969ca5486f6c000667a9d511cd45b6d9c5bde5d2ece063176fc1440bbd593bf4a55ff70186fece662ca249d95ab6fa916f425274d732149743e995b3f10a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f43d3aa6030cde19ad6877c0386112d7a2e1dd8e60f3495fbdc5bf067411572951bf1017fd8f83b3c7156a2b1830dbf080a3d70fc9e46f2fe57d1c092ddb9c0cd83c4bd69f202facf3fec47f9e9f83db9a54d6781267076fbeb1c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9c065743ff244e02fde6100ab01fadbcd17fc72b75e359222bb71a7d6afdbee40067b8fc86355b53b4fa5d71565077eee9c674c22adbbfd3ae6e38d8c407294ad1b5a6000aa2c88ed0a16ad8741479804d5d581a77855c05de81f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h101319fa69b04cbc531723333ce07f9f766ae312068d89f89e15fcb044c31cc21e49f4564e874129d0561afd472ecb9b9a4c21a67a12fe5dc10b9f5a981f7b2467c2f4360776de28bb4805c4cd58315198a099893ee931e3e2a7b88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d78b9899032aa183b7a5cb7824c873092c43a376a8e364da5ff47e378741f3c12b4ac03ec2bd42bbaa343494ac533e8888a6420d795524d72d8e7c566eae5a9f1e1faf5105ce642ef2c3fbf4b21ba272995a39c1b31537166ce9b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d218304a0b36521b61f586c1c546926afa5c4b3fed1230b76c010bac56e5da044be6fcc6350a20697d13ff72ec1a0f05c9abb3a2ad4dd41c55f9a61d4559fcce7343e4eb4f301131436b22705a75868fa4d836803683f9d601bd74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7ea22cd08ab01eb65e25e1c649e077fba90895215416df17d490194b063248c2091f84f4d880a2a20a87de76d2b9f9bf63f26200f304460f0de635713733a446e7c6f80fc7be547082de90af8974321b994d8d4b4a7299d9b4a6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd03e9098ce1751d63a61b7206c1fcae56dc668e8c2619c30677c24877329e3b504059bca3a716092c176152ff2f8ac19391d83414fd02bd8750f2f879211b0039b33ae200e4dc573df8ab86a7dd22acb927f73738ec1479a74616;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190489644681712c9a18ead306afd4f0146327fa67c34560984a6a87522b1db5f2e6da825c3339024847ed22b27e97b9de5d6c67510f323a95e2a66d6fdc76b1ca5a2f82dda4543b2112df14e54cafe47c45323c933bd84cc43b1c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e713fb050ac1e819a099800650a9fc9d3956cbcbd6effee9547964f7e4bd0d3edc4935f0073c1a1a9135593ce77b498ef3240e82069746a2980ea97b0b332dec6f82e72d624ce2285f0ba6985ed6c35cdcbaccf6cf985665df219;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h953eabfc51f09da218021c5d8ca6a1e2f1272ca5061562f03b4f5fd061214dcf2712faabd1d69d36a9b1f1c07246a076a0290be44e3bbd02a64de1e1ffc6586597d6ab6e9346d1a43e0fc212a1dccdc87ccc2b516c5b2ffc12858;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f880917b399623b437916acb8613b46788fc4d7177b9bf81019f87bbd7c47cb2311240bdb375835bfa483428a6aeceb1b944f7f9daca1b682e0901e9ad051a799dc701d26b729590107bd718e8d38e15f4576278acbe9d8e591dbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c842a3b440d7f748f395e5cebaba83c98cf9a5cdff50ac404dbed37e5a0007568b32e89952eb0049f9cfbed43997fd0146f51e4f4a5f1c61524af4583baa158fc6149ce7e41deb16f04b36a8bbdcd80c06289e0ef60a96bd3e031;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c8822af9a7294cb2f88f587f609a666ceb2354820cf986a1fc1a82cb26de5190e72399e14375c1c82ffccc3f12eae7a05d6deaa9993ce29636aaac927c9685e042501804cda080b98400a63321da33c125cb8fa9475eb04a44d54;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1ae4ba13f1c026e0d42665dd04f3289acd61e7e89a1dbc79630ef4280c6f286dbd694656ca939b80aaf1835da3891fd8bd9bd89eaf7bf66e07e7f20b86dbf7b5ceea8076ef9b31dadf766bb4069e5fca70b6493d034cd642997b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ac6b92f6eae0dd82787dd2d34040472ea8aed163836a2e2f8c16790f824ce2408eb90584d90441cd808725babca89ed3b4874688438a1d7ea85fdd8d342655f9132fd31b364d49ddfa520db6d6281f6b093c3dbaea06f59555ecc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30853e1687906647b32104a0890ffc9febb274637f1a2c00a9d3ec3a396268b33e58124f7872dd3fc4103fb4d203d5ae8437a1d04942100e4155058a1b24bff8bf24b3118cccc0be7452f42fc0e48bf72a07b956b66893ce1b7ec5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f656852df10a1eaf1197074965d1bc1739f1e580c0fbe4767709042e0de6da02c91d13f0fcbffc2bb0650d1c33efb0ff28e4b82a3fb0db8cdfae50bf8354cd6eb5ae205758b01f7b0ab732ecdeeaec2d3307c624c88bc72a4cf5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11095f54d08977fb08c75b7f38148959eb21d4b43d21b633faaa7737d8b0314c61f125eebba497afd2a162980f70a321bb6fbdd9a4f204d0ce1148f0088604a57fae00e38afc258dcb55634234f7f1980c9540883252caf1cdc12ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6d4b1cc192b2d5937c3b4728ddbc498108056c7639b7641d67a11e26b93eb8b1590cb79685faae7c6e6fd56190f788a95bcd23d2cadfc215229e927c6d6d344e4c0bb145fd0f29e93e1f8784dd7846fa1fa817fdfe37ce25a452a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he24aba20e08be96cc43ab3c78cc66a78531ddb10ff711f291a0b9e7fc296a8c5a1718e6fd6eda0d9fa320f8ccadb65c3da7fb5c87416585cebad41bd2c9d2cb17b20a73c57724cfefe7ee3b8f0e584729845faa51c60d000369397;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1537f1e4ec4676f8e3e3512d2ab94ac9664654d208351a381714ea17d70268c5f00713150963ac7c44e3490b6628e35b33d046e35632c1503e4ef65b04b815d5e75fc8097b5b23fad109fb0278e9bc4a1d1a4156f932f3ed376e5cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb85383551ef401b410bf46ff00d89c47b69815615276d969c311061ddf04150404133b41ef291f65f40b238a8909b317dfc8a89ac7dc11a095819cfbe5b8730bbdea247bd1e7214c2b7402031908c98c42176dba074e65b5e94d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h178a611fbec823ec6491f4de0589971f1dc81abbbc0b48c9cc23d1b3e03d542a8a92f4d57309c9e80cd55baf1c1b723305292c955a3986dcf4f1f4ce4458834081dcbb395d7a52a784a17b56c951b349dd6d00e4510617937bee2c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h178b7614a6a2196f277f2c4e8e61df3257e59f00bf2cbfae1316c908f9c953f6fcadd55213d6f7d63ce69a2ce1650afff3fd4411648efc4fab5f190fb3500af15d78c6990d77cca47843708327ee9dfb0c9e0f35c2dc6e4023ec1cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd98a13a137129b03a3c3aca7709e5a1d396059e04d3364a63fb9366e3e2d10d058367b09a24a5585646023d1015ad4af3c3dc5506c0363c8eaf7048424107e4c348fe790f4a9cf551e6837429cebb10c34c006fdfa4d8fb5f25d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c63ac451e1ebb9ebbd8613f73fb5cedcbde7693dffe3c8ff9b7fe753a58f84a4e919ec19207271b4046941054beaae306ec733a4a4fac0370a2757c7736294afdbcbcbcda01a70579afbc09de91d4c19568308e351e8bfc470d02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had93ab610156cd1d3926f9e6ec3841054ffd3ec22a8a1f089d3fc397b41f1f4bc70f80dfcb0b4381758bb4ba64eb7a4bd2e7e1e5a44507657b5efa5b8f2bff137217e249ab089877bdfe188b0e4dd77520dc6e1c4c954097547dcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1512902c6d3d7aef22e6d37c562594a6309c015974e105ff798f5e823d8067c08a4f29e4382a19800b127b0b93550d74e43b6a7490b0c8fd3ddca87590652ee8d5deae9063459b2fcebeba1ac90be50af53408f01dc170cdcbb89fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1edd2b8e2a1cd64188bd36b3ceb0de10de15524823c2cf0f9e1795501481415779374996297f765400e260901287f3436ff484fed8bd1c6ca8b846f78129bfde4f05eea734bf93e1cde5422c4f97e9034c384abab73000920d8e282;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192267015e503c5a9675c9b9854fd4fa8924151bfaebbd084e3729e5832942b4fc23f05eccf852b5bfa6c020f7dc5e5b2204b9a463f7750b1df476d7cc7e68df41029bc928209d78cb1d20b18920a0f6e92d81c32f9469f5b5a72eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1439a40561ef969ff1a7800095b886fce87d3b055502ac55889716e8dc81796d17dae81ede8846eea9ac1203b25217be780d217d36b4504dd20663cef6a767d1c1c0d4a22c2c950caac2c4814956fcf42cd30bc0c868a1a43dd5d4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h57c286ac390a0fac713c432ac19e92bb2267dee7a0e1c46a8c5908bd87d9472d11b34a3f58a463e2803a31ec7b613a2a2648fc49af40ff1d2fdfa767bcfb3dc3f6dce26671b2786ab455d22ff33845f7f547cc2593d2d83b5503fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hedfa4dd179974d5d2cc1fd0ecb24eb81e4bb759b43d3c778343c6c14ee691df3fdb62fadd6cb3006b31b8ad355a93bf0504bbd4c3a072cb19fbe28ffbc5299c4dce1f2cf6f5c5b07a9a1834df585bedc41b1d0f9b840dcdb7851d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2b3c92580dfc5df9048722c48b9121d6c7792a462add6d01ff64ff435884bae9cde2a099380cfd8c66357945995d3824b23deadcbd1f2b76315a38e5bcefc237dd601cf1c7a082bfb120703457a89a282c16dec2e801d84965b452;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fe0635441baa50e0ded4a4ee6cc09fb8ddd30ce22c8c4c27302243865ec6b934f8fd9e30ef492e22d9db7d0ca9645d6964ce5a08fac79068c3f7d3517c1f096408a93bfa44f32f3b481599ea6415b70346d173437710372b6fb88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137f54568545aba0ae4c8345bbdf511434485d142cc756e31af8a3e43f13c51e6911bbffb93cb4ea8844438717e39130e28263ce5edc353bc5605e2d01fa585eea0b3916f2556802b44703d7d9e1ff8a36088894ab6f3ac79dcd9ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1531640420269932a560140cf0801c43c11adeb0e48fda9d92a82e07c70d5db4c470e751ccc31c2a9dbe699a6d2c31ad1e75d818d8f7c9b3b298344ed9a2825c808efd4ef484f642aef8a802a060877ee7ceaec59ba27cfe4de2951;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b29f60bf3120d1fc761b6c7b5c77c82653c76e359b6d71406e7de719d6e749f2e3d39d9c00d05ca6b62f706626a183038125973106ba420fbd3fdb061faa6993262770a6799d7db1350408bbb3a5d8c7ff4f6662d41f4203b8a8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf028bfef45c21165a7ecd6d77441475e327cbe0d38f1c9162736a6342e0fffb00e66845b39c6516a8ef5972f60d893d6f2775a72d0d1ddbfca243a4299e6dd01ff4987a0a13d5a67140d331cba64ad9c02d488acea44cbcf6176c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8b87db48018e8a62b71c64c49e76dfb4678c3e496f1e3a103bccbedead312ac2cc16f7342b7af87c109abfe39f74b1c84ce4880d882e25eb14db03c2b93d6fec0c935fa1d76ff8e1e38eae8649e8813a07fc80ae1064042393f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e45e6d3bca9934247c56323f58488623c50c8d3a9fbda6f0ce3c219c677baed9a4d9e5e86ca617521e0f00a515b60211a0ec55af2bd47902117292fb5c354b8040660c10ba95ffdfedad9c312e22ef5597402f91656812d4150c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4413b02fa73c3165e7f429e8499531dfbb4bb32a33c9e4446eae9e9d81f79628ffd1d177e060398ab32157301ddf62800f6d7e856e846a2cf8476d9c3d47ea46d3a2993a1b278153d96011e1e5a7bdab4cf081f3567255ee55795;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1655a5e60f8951892785c53942f3059573d357200ab7dbe6c5bf0ac2aa56f6a2ee8f89a6ac0f161d4b5c05f738782311892f96a5dbad7ae531549c15cae483cbb4ec73aac7d0be35f1b5e661dc546e116f183fd13952f1819e7cfa3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c98112a59d31468dcfc355bea6ab3999e7d79eb1df26f124c1a0afaa17b6a66588634969ecbcf2044710e81abe3202d013c763f47f02cbc99b90c35b106235c1e42925a191480da4f3c38885c81c909149a6f3026aafab6db156a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb5f0a3fc9777f2a5e024b9683885bae242237ad62350cbf5c4aa60bd8d7d56435d245cfb13db7392e66e83ad24827d72ebcb4cd8cbb7e7769d9dc98676b3fa7e5217742d10375287b0a4189509f565eec6777b933521aea7536c3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he60d588f041b3aa36bef488ae5efac4682e5c9c575163c418194db5697457834c5c7095ea24bbb2fc7b309707733e61f920f52392463519adaf9c48fa65cd1d2efc53f16e3364c60de949f8c4a8bad6be24cf225432b8fe361f982;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114b04d7742ed3d4a869850dd8750a248aaed5f09497dcd4e2aaa07d7ba95fe678ad323db7676472ea76398782a89c8670db39a51fc1aa9bb02c98628189ac43b2ee28ad1e37777c9639b614229f7d0b8af25e321fa8d3a62bb6fb3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1915fd85a28044452f888d63f586540ecbd0b8f8f6e078f85b155ec853a4d7b2b391dd66bffb66f8a6235dcbb96688afd955cdba8daa2f414567b791363aa0fedf6c25488478d71474e461b292568ec18152ffe769374724e7e9df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15792a4660c9af84a4688c04c10e6db03c6412582b8d361370e663d74b0e86f54fc9b637136050b09c44ce5543772f688d0305c23ad1f00f9703c41d825c522381a476b70be7a3f0acae54c1fdd1bfc0d93d5bccb80116e6a207c53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h639ff2ce1f21524b8540c0381be76c44dc7de98b0dfc3169a7f32570bf1559302e5b3d2cd4795759efea503af347b306a7c52e00cf477f4d66321bf4a72eb2f882f207ccb97fb471ff6b3d23493789e27cf502bd776b2a8fbab5d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11feefe3db2c08e66367fa8af5592d66e3dd342c442a7287ebfa9b885e41e12b9e200090bdfbd600aa5b7514beab1daa7b701d68928b6dbaa54cdaf1dbff25d6125e6c05b73525f71103a13750d7fd2e78a66cf5cc9e68fcdcd1f8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb3f621deba88c46545d0f8c882566d8f7b20fba125e71c39e5f8420023685099133f2448b230f7dcb91425b6e6017ad7f693b36190246ce7f6a4c51cdbc71e8e55c07a1e82e9d8a28f0ea9f141fef4c30bf36ff8fec9347582a8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c587c6082bd994f717281725000786e262bceb8cc6e83dcef528f851d85576992798423b779b8d0a9c4a3e4de72c6d870f1e8d5b5f2c59c8b5392f6a22f0d8352452d01aa8c59808353cc443d15ee46c80c7b3673a14a75cbbeeb;
        #1
        $finish();
    end
endmodule
