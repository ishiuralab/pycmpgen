module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71,
        output wire [0:0] dst72);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    reg [485:0] src32;
    reg [485:0] src33;
    reg [485:0] src34;
    reg [485:0] src35;
    reg [485:0] src36;
    reg [485:0] src37;
    reg [485:0] src38;
    reg [485:0] src39;
    reg [485:0] src40;
    reg [485:0] src41;
    reg [485:0] src42;
    reg [485:0] src43;
    reg [485:0] src44;
    reg [485:0] src45;
    reg [485:0] src46;
    reg [485:0] src47;
    reg [485:0] src48;
    reg [485:0] src49;
    reg [485:0] src50;
    reg [485:0] src51;
    reg [485:0] src52;
    reg [485:0] src53;
    reg [485:0] src54;
    reg [485:0] src55;
    reg [485:0] src56;
    reg [485:0] src57;
    reg [485:0] src58;
    reg [485:0] src59;
    reg [485:0] src60;
    reg [485:0] src61;
    reg [485:0] src62;
    reg [485:0] src63;
    compressor2_1_486_64 compressor2_1_486_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71),
            .dst72(dst72));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
        src12 <= 486'h0;
        src13 <= 486'h0;
        src14 <= 486'h0;
        src15 <= 486'h0;
        src16 <= 486'h0;
        src17 <= 486'h0;
        src18 <= 486'h0;
        src19 <= 486'h0;
        src20 <= 486'h0;
        src21 <= 486'h0;
        src22 <= 486'h0;
        src23 <= 486'h0;
        src24 <= 486'h0;
        src25 <= 486'h0;
        src26 <= 486'h0;
        src27 <= 486'h0;
        src28 <= 486'h0;
        src29 <= 486'h0;
        src30 <= 486'h0;
        src31 <= 486'h0;
        src32 <= 486'h0;
        src33 <= 486'h0;
        src34 <= 486'h0;
        src35 <= 486'h0;
        src36 <= 486'h0;
        src37 <= 486'h0;
        src38 <= 486'h0;
        src39 <= 486'h0;
        src40 <= 486'h0;
        src41 <= 486'h0;
        src42 <= 486'h0;
        src43 <= 486'h0;
        src44 <= 486'h0;
        src45 <= 486'h0;
        src46 <= 486'h0;
        src47 <= 486'h0;
        src48 <= 486'h0;
        src49 <= 486'h0;
        src50 <= 486'h0;
        src51 <= 486'h0;
        src52 <= 486'h0;
        src53 <= 486'h0;
        src54 <= 486'h0;
        src55 <= 486'h0;
        src56 <= 486'h0;
        src57 <= 486'h0;
        src58 <= 486'h0;
        src59 <= 486'h0;
        src60 <= 486'h0;
        src61 <= 486'h0;
        src62 <= 486'h0;
        src63 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor2_1_486_64(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    input [485:0]src12,
    input [485:0]src13,
    input [485:0]src14,
    input [485:0]src15,
    input [485:0]src16,
    input [485:0]src17,
    input [485:0]src18,
    input [485:0]src19,
    input [485:0]src20,
    input [485:0]src21,
    input [485:0]src22,
    input [485:0]src23,
    input [485:0]src24,
    input [485:0]src25,
    input [485:0]src26,
    input [485:0]src27,
    input [485:0]src28,
    input [485:0]src29,
    input [485:0]src30,
    input [485:0]src31,
    input [485:0]src32,
    input [485:0]src33,
    input [485:0]src34,
    input [485:0]src35,
    input [485:0]src36,
    input [485:0]src37,
    input [485:0]src38,
    input [485:0]src39,
    input [485:0]src40,
    input [485:0]src41,
    input [485:0]src42,
    input [485:0]src43,
    input [485:0]src44,
    input [485:0]src45,
    input [485:0]src46,
    input [485:0]src47,
    input [485:0]src48,
    input [485:0]src49,
    input [485:0]src50,
    input [485:0]src51,
    input [485:0]src52,
    input [485:0]src53,
    input [485:0]src54,
    input [485:0]src55,
    input [485:0]src56,
    input [485:0]src57,
    input [485:0]src58,
    input [485:0]src59,
    input [485:0]src60,
    input [485:0]src61,
    input [485:0]src62,
    input [485:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71,
    output dst72);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [0:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [0:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [1:0] comp_out70;
    wire [1:0] comp_out71;
    wire [1:0] comp_out72;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71),
        .dst72(comp_out72)
    );
    rowadder2_1_73 rowadder2_1inst(
        .src0({comp_out72[0], comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out72[1], comp_out71[1], comp_out70[1], comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], 1'h0, comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], 1'h0, comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], 1'h0}),
        .dst0({dst72, dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      input wire [485:0] src12,
      input wire [485:0] src13,
      input wire [485:0] src14,
      input wire [485:0] src15,
      input wire [485:0] src16,
      input wire [485:0] src17,
      input wire [485:0] src18,
      input wire [485:0] src19,
      input wire [485:0] src20,
      input wire [485:0] src21,
      input wire [485:0] src22,
      input wire [485:0] src23,
      input wire [485:0] src24,
      input wire [485:0] src25,
      input wire [485:0] src26,
      input wire [485:0] src27,
      input wire [485:0] src28,
      input wire [485:0] src29,
      input wire [485:0] src30,
      input wire [485:0] src31,
      input wire [485:0] src32,
      input wire [485:0] src33,
      input wire [485:0] src34,
      input wire [485:0] src35,
      input wire [485:0] src36,
      input wire [485:0] src37,
      input wire [485:0] src38,
      input wire [485:0] src39,
      input wire [485:0] src40,
      input wire [485:0] src41,
      input wire [485:0] src42,
      input wire [485:0] src43,
      input wire [485:0] src44,
      input wire [485:0] src45,
      input wire [485:0] src46,
      input wire [485:0] src47,
      input wire [485:0] src48,
      input wire [485:0] src49,
      input wire [485:0] src50,
      input wire [485:0] src51,
      input wire [485:0] src52,
      input wire [485:0] src53,
      input wire [485:0] src54,
      input wire [485:0] src55,
      input wire [485:0] src56,
      input wire [485:0] src57,
      input wire [485:0] src58,
      input wire [485:0] src59,
      input wire [485:0] src60,
      input wire [485:0] src61,
      input wire [485:0] src62,
      input wire [485:0] src63,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [0:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [0:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [1:0] dst70,
      output wire [1:0] dst71,
      output wire [1:0] dst72);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [485:0] stage0_12;
   wire [485:0] stage0_13;
   wire [485:0] stage0_14;
   wire [485:0] stage0_15;
   wire [485:0] stage0_16;
   wire [485:0] stage0_17;
   wire [485:0] stage0_18;
   wire [485:0] stage0_19;
   wire [485:0] stage0_20;
   wire [485:0] stage0_21;
   wire [485:0] stage0_22;
   wire [485:0] stage0_23;
   wire [485:0] stage0_24;
   wire [485:0] stage0_25;
   wire [485:0] stage0_26;
   wire [485:0] stage0_27;
   wire [485:0] stage0_28;
   wire [485:0] stage0_29;
   wire [485:0] stage0_30;
   wire [485:0] stage0_31;
   wire [485:0] stage0_32;
   wire [485:0] stage0_33;
   wire [485:0] stage0_34;
   wire [485:0] stage0_35;
   wire [485:0] stage0_36;
   wire [485:0] stage0_37;
   wire [485:0] stage0_38;
   wire [485:0] stage0_39;
   wire [485:0] stage0_40;
   wire [485:0] stage0_41;
   wire [485:0] stage0_42;
   wire [485:0] stage0_43;
   wire [485:0] stage0_44;
   wire [485:0] stage0_45;
   wire [485:0] stage0_46;
   wire [485:0] stage0_47;
   wire [485:0] stage0_48;
   wire [485:0] stage0_49;
   wire [485:0] stage0_50;
   wire [485:0] stage0_51;
   wire [485:0] stage0_52;
   wire [485:0] stage0_53;
   wire [485:0] stage0_54;
   wire [485:0] stage0_55;
   wire [485:0] stage0_56;
   wire [485:0] stage0_57;
   wire [485:0] stage0_58;
   wire [485:0] stage0_59;
   wire [485:0] stage0_60;
   wire [485:0] stage0_61;
   wire [485:0] stage0_62;
   wire [485:0] stage0_63;
   wire [124:0] stage1_0;
   wire [175:0] stage1_1;
   wire [157:0] stage1_2;
   wire [214:0] stage1_3;
   wire [227:0] stage1_4;
   wire [197:0] stage1_5;
   wire [213:0] stage1_6;
   wire [220:0] stage1_7;
   wire [205:0] stage1_8;
   wire [213:0] stage1_9;
   wire [284:0] stage1_10;
   wire [276:0] stage1_11;
   wire [188:0] stage1_12;
   wire [304:0] stage1_13;
   wire [218:0] stage1_14;
   wire [170:0] stage1_15;
   wire [221:0] stage1_16;
   wire [228:0] stage1_17;
   wire [208:0] stage1_18;
   wire [275:0] stage1_19;
   wire [267:0] stage1_20;
   wire [189:0] stage1_21;
   wire [170:0] stage1_22;
   wire [286:0] stage1_23;
   wire [213:0] stage1_24;
   wire [183:0] stage1_25;
   wire [250:0] stage1_26;
   wire [205:0] stage1_27;
   wire [223:0] stage1_28;
   wire [228:0] stage1_29;
   wire [191:0] stage1_30;
   wire [217:0] stage1_31;
   wire [216:0] stage1_32;
   wire [258:0] stage1_33;
   wire [189:0] stage1_34;
   wire [216:0] stage1_35;
   wire [201:0] stage1_36;
   wire [307:0] stage1_37;
   wire [264:0] stage1_38;
   wire [212:0] stage1_39;
   wire [303:0] stage1_40;
   wire [170:0] stage1_41;
   wire [173:0] stage1_42;
   wire [253:0] stage1_43;
   wire [255:0] stage1_44;
   wire [211:0] stage1_45;
   wire [297:0] stage1_46;
   wire [235:0] stage1_47;
   wire [197:0] stage1_48;
   wire [172:0] stage1_49;
   wire [189:0] stage1_50;
   wire [274:0] stage1_51;
   wire [198:0] stage1_52;
   wire [168:0] stage1_53;
   wire [230:0] stage1_54;
   wire [266:0] stage1_55;
   wire [186:0] stage1_56;
   wire [188:0] stage1_57;
   wire [219:0] stage1_58;
   wire [205:0] stage1_59;
   wire [214:0] stage1_60;
   wire [218:0] stage1_61;
   wire [192:0] stage1_62;
   wire [307:0] stage1_63;
   wire [123:0] stage1_64;
   wire [53:0] stage1_65;
   wire [37:0] stage2_0;
   wire [53:0] stage2_1;
   wire [62:0] stage2_2;
   wire [113:0] stage2_3;
   wire [111:0] stage2_4;
   wire [151:0] stage2_5;
   wire [91:0] stage2_6;
   wire [72:0] stage2_7;
   wire [159:0] stage2_8;
   wire [142:0] stage2_9;
   wire [163:0] stage2_10;
   wire [138:0] stage2_11;
   wire [106:0] stage2_12;
   wire [77:0] stage2_13;
   wire [107:0] stage2_14;
   wire [140:0] stage2_15;
   wire [82:0] stage2_16;
   wire [86:0] stage2_17;
   wire [118:0] stage2_18;
   wire [112:0] stage2_19;
   wire [92:0] stage2_20;
   wire [127:0] stage2_21;
   wire [107:0] stage2_22;
   wire [75:0] stage2_23;
   wire [101:0] stage2_24;
   wire [95:0] stage2_25;
   wire [84:0] stage2_26;
   wire [105:0] stage2_27;
   wire [91:0] stage2_28;
   wire [86:0] stage2_29;
   wire [116:0] stage2_30;
   wire [98:0] stage2_31;
   wire [105:0] stage2_32;
   wire [75:0] stage2_33;
   wire [131:0] stage2_34;
   wire [132:0] stage2_35;
   wire [74:0] stage2_36;
   wire [89:0] stage2_37;
   wire [139:0] stage2_38;
   wire [136:0] stage2_39;
   wire [112:0] stage2_40;
   wire [105:0] stage2_41;
   wire [85:0] stage2_42;
   wire [78:0] stage2_43;
   wire [118:0] stage2_44;
   wire [117:0] stage2_45;
   wire [87:0] stage2_46;
   wire [103:0] stage2_47;
   wire [129:0] stage2_48;
   wire [95:0] stage2_49;
   wire [85:0] stage2_50;
   wire [87:0] stage2_51;
   wire [104:0] stage2_52;
   wire [114:0] stage2_53;
   wire [99:0] stage2_54;
   wire [105:0] stage2_55;
   wire [114:0] stage2_56;
   wire [65:0] stage2_57;
   wire [85:0] stage2_58;
   wire [109:0] stage2_59;
   wire [84:0] stage2_60;
   wire [74:0] stage2_61;
   wire [104:0] stage2_62;
   wire [98:0] stage2_63;
   wire [141:0] stage2_64;
   wire [55:0] stage2_65;
   wire [41:0] stage2_66;
   wire [20:0] stage3_0;
   wire [21:0] stage3_1;
   wire [42:0] stage3_2;
   wire [28:0] stage3_3;
   wire [111:0] stage3_4;
   wire [52:0] stage3_5;
   wire [77:0] stage3_6;
   wire [50:0] stage3_7;
   wire [34:0] stage3_8;
   wire [53:0] stage3_9;
   wire [99:0] stage3_10;
   wire [57:0] stage3_11;
   wire [67:0] stage3_12;
   wire [56:0] stage3_13;
   wire [31:0] stage3_14;
   wire [47:0] stage3_15;
   wire [50:0] stage3_16;
   wire [35:0] stage3_17;
   wire [59:0] stage3_18;
   wire [47:0] stage3_19;
   wire [82:0] stage3_20;
   wire [38:0] stage3_21;
   wire [72:0] stage3_22;
   wire [42:0] stage3_23;
   wire [28:0] stage3_24;
   wire [32:0] stage3_25;
   wire [48:0] stage3_26;
   wire [48:0] stage3_27;
   wire [56:0] stage3_28;
   wire [47:0] stage3_29;
   wire [41:0] stage3_30;
   wire [37:0] stage3_31;
   wire [53:0] stage3_32;
   wire [45:0] stage3_33;
   wire [41:0] stage3_34;
   wire [56:0] stage3_35;
   wire [45:0] stage3_36;
   wire [52:0] stage3_37;
   wire [59:0] stage3_38;
   wire [57:0] stage3_39;
   wire [51:0] stage3_40;
   wire [42:0] stage3_41;
   wire [49:0] stage3_42;
   wire [45:0] stage3_43;
   wire [40:0] stage3_44;
   wire [43:0] stage3_45;
   wire [57:0] stage3_46;
   wire [43:0] stage3_47;
   wire [41:0] stage3_48;
   wire [41:0] stage3_49;
   wire [46:0] stage3_50;
   wire [62:0] stage3_51;
   wire [62:0] stage3_52;
   wire [74:0] stage3_53;
   wire [38:0] stage3_54;
   wire [66:0] stage3_55;
   wire [31:0] stage3_56;
   wire [53:0] stage3_57;
   wire [61:0] stage3_58;
   wire [49:0] stage3_59;
   wire [41:0] stage3_60;
   wire [52:0] stage3_61;
   wire [33:0] stage3_62;
   wire [47:0] stage3_63;
   wire [50:0] stage3_64;
   wire [37:0] stage3_65;
   wire [37:0] stage3_66;
   wire [13:0] stage3_67;
   wire [5:0] stage3_68;
   wire [8:0] stage4_0;
   wire [6:0] stage4_1;
   wire [10:0] stage4_2;
   wire [16:0] stage4_3;
   wire [30:0] stage4_4;
   wire [35:0] stage4_5;
   wire [23:0] stage4_6;
   wire [38:0] stage4_7;
   wire [27:0] stage4_8;
   wire [13:0] stage4_9;
   wire [41:0] stage4_10;
   wire [28:0] stage4_11;
   wire [23:0] stage4_12;
   wire [31:0] stage4_13;
   wire [29:0] stage4_14;
   wire [14:0] stage4_15;
   wire [26:0] stage4_16;
   wire [17:0] stage4_17;
   wire [20:0] stage4_18;
   wire [28:0] stage4_19;
   wire [33:0] stage4_20;
   wire [36:0] stage4_21;
   wire [17:0] stage4_22;
   wire [20:0] stage4_23;
   wire [21:0] stage4_24;
   wire [20:0] stage4_25;
   wire [18:0] stage4_26;
   wire [26:0] stage4_27;
   wire [18:0] stage4_28;
   wire [21:0] stage4_29;
   wire [32:0] stage4_30;
   wire [14:0] stage4_31;
   wire [29:0] stage4_32;
   wire [28:0] stage4_33;
   wire [18:0] stage4_34;
   wire [35:0] stage4_35;
   wire [35:0] stage4_36;
   wire [17:0] stage4_37;
   wire [19:0] stage4_38;
   wire [23:0] stage4_39;
   wire [27:0] stage4_40;
   wire [19:0] stage4_41;
   wire [37:0] stage4_42;
   wire [13:0] stage4_43;
   wire [24:0] stage4_44;
   wire [28:0] stage4_45;
   wire [16:0] stage4_46;
   wire [20:0] stage4_47;
   wire [22:0] stage4_48;
   wire [12:0] stage4_49;
   wire [21:0] stage4_50;
   wire [35:0] stage4_51;
   wire [18:0] stage4_52;
   wire [43:0] stage4_53;
   wire [25:0] stage4_54;
   wire [38:0] stage4_55;
   wire [13:0] stage4_56;
   wire [25:0] stage4_57;
   wire [23:0] stage4_58;
   wire [20:0] stage4_59;
   wire [21:0] stage4_60;
   wire [31:0] stage4_61;
   wire [16:0] stage4_62;
   wire [13:0] stage4_63;
   wire [33:0] stage4_64;
   wire [35:0] stage4_65;
   wire [10:0] stage4_66;
   wire [10:0] stage4_67;
   wire [13:0] stage4_68;
   wire [1:0] stage4_69;
   wire [4:0] stage5_0;
   wire [1:0] stage5_1;
   wire [4:0] stage5_2;
   wire [7:0] stage5_3;
   wire [10:0] stage5_4;
   wire [15:0] stage5_5;
   wire [9:0] stage5_6;
   wire [10:0] stage5_7;
   wire [18:0] stage5_8;
   wire [10:0] stage5_9;
   wire [20:0] stage5_10;
   wire [13:0] stage5_11;
   wire [10:0] stage5_12;
   wire [14:0] stage5_13;
   wire [15:0] stage5_14;
   wire [11:0] stage5_15;
   wire [7:0] stage5_16;
   wire [6:0] stage5_17;
   wire [11:0] stage5_18;
   wire [15:0] stage5_19;
   wire [13:0] stage5_20;
   wire [10:0] stage5_21;
   wire [13:0] stage5_22;
   wire [9:0] stage5_23;
   wire [8:0] stage5_24;
   wire [9:0] stage5_25;
   wire [14:0] stage5_26;
   wire [5:0] stage5_27;
   wire [9:0] stage5_28;
   wire [14:0] stage5_29;
   wire [8:0] stage5_30;
   wire [9:0] stage5_31;
   wire [19:0] stage5_32;
   wire [11:0] stage5_33;
   wire [13:0] stage5_34;
   wire [13:0] stage5_35;
   wire [12:0] stage5_36;
   wire [10:0] stage5_37;
   wire [9:0] stage5_38;
   wire [9:0] stage5_39;
   wire [10:0] stage5_40;
   wire [8:0] stage5_41;
   wire [18:0] stage5_42;
   wire [10:0] stage5_43;
   wire [12:0] stage5_44;
   wire [14:0] stage5_45;
   wire [11:0] stage5_46;
   wire [11:0] stage5_47;
   wire [13:0] stage5_48;
   wire [5:0] stage5_49;
   wire [11:0] stage5_50;
   wire [18:0] stage5_51;
   wire [9:0] stage5_52;
   wire [12:0] stage5_53;
   wire [16:0] stage5_54;
   wire [21:0] stage5_55;
   wire [8:0] stage5_56;
   wire [13:0] stage5_57;
   wire [15:0] stage5_58;
   wire [7:0] stage5_59;
   wire [14:0] stage5_60;
   wire [15:0] stage5_61;
   wire [11:0] stage5_62;
   wire [8:0] stage5_63;
   wire [14:0] stage5_64;
   wire [17:0] stage5_65;
   wire [7:0] stage5_66;
   wire [10:0] stage5_67;
   wire [13:0] stage5_68;
   wire [2:0] stage5_69;
   wire [0:0] stage5_70;
   wire [4:0] stage6_0;
   wire [1:0] stage6_1;
   wire [4:0] stage6_2;
   wire [1:0] stage6_3;
   wire [5:0] stage6_4;
   wire [3:0] stage6_5;
   wire [7:0] stage6_6;
   wire [4:0] stage6_7;
   wire [5:0] stage6_8;
   wire [9:0] stage6_9;
   wire [4:0] stage6_10;
   wire [6:0] stage6_11;
   wire [6:0] stage6_12;
   wire [9:0] stage6_13;
   wire [6:0] stage6_14;
   wire [5:0] stage6_15;
   wire [4:0] stage6_16;
   wire [4:0] stage6_17;
   wire [5:0] stage6_18;
   wire [4:0] stage6_19;
   wire [5:0] stage6_20;
   wire [5:0] stage6_21;
   wire [5:0] stage6_22;
   wire [6:0] stage6_23;
   wire [6:0] stage6_24;
   wire [2:0] stage6_25;
   wire [7:0] stage6_26;
   wire [4:0] stage6_27;
   wire [5:0] stage6_28;
   wire [5:0] stage6_29;
   wire [4:0] stage6_30;
   wire [5:0] stage6_31;
   wire [5:0] stage6_32;
   wire [5:0] stage6_33;
   wire [8:0] stage6_34;
   wire [4:0] stage6_35;
   wire [5:0] stage6_36;
   wire [5:0] stage6_37;
   wire [4:0] stage6_38;
   wire [3:0] stage6_39;
   wire [5:0] stage6_40;
   wire [7:0] stage6_41;
   wire [6:0] stage6_42;
   wire [6:0] stage6_43;
   wire [4:0] stage6_44;
   wire [8:0] stage6_45;
   wire [4:0] stage6_46;
   wire [6:0] stage6_47;
   wire [4:0] stage6_48;
   wire [5:0] stage6_49;
   wire [2:0] stage6_50;
   wire [7:0] stage6_51;
   wire [6:0] stage6_52;
   wire [4:0] stage6_53;
   wire [5:0] stage6_54;
   wire [9:0] stage6_55;
   wire [9:0] stage6_56;
   wire [6:0] stage6_57;
   wire [5:0] stage6_58;
   wire [4:0] stage6_59;
   wire [4:0] stage6_60;
   wire [8:0] stage6_61;
   wire [5:0] stage6_62;
   wire [4:0] stage6_63;
   wire [8:0] stage6_64;
   wire [4:0] stage6_65;
   wire [4:0] stage6_66;
   wire [4:0] stage6_67;
   wire [16:0] stage6_68;
   wire [4:0] stage6_69;
   wire [0:0] stage6_70;
   wire [4:0] stage7_0;
   wire [1:0] stage7_1;
   wire [4:0] stage7_2;
   wire [1:0] stage7_3;
   wire [0:0] stage7_4;
   wire [1:0] stage7_5;
   wire [2:0] stage7_6;
   wire [2:0] stage7_7;
   wire [4:0] stage7_8;
   wire [5:0] stage7_9;
   wire [1:0] stage7_10;
   wire [3:0] stage7_11;
   wire [1:0] stage7_12;
   wire [5:0] stage7_13;
   wire [2:0] stage7_14;
   wire [5:0] stage7_15;
   wire [2:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [6:0] stage7_19;
   wire [2:0] stage7_20;
   wire [5:0] stage7_21;
   wire [6:0] stage7_22;
   wire [0:0] stage7_23;
   wire [3:0] stage7_24;
   wire [1:0] stage7_25;
   wire [5:0] stage7_26;
   wire [4:0] stage7_27;
   wire [0:0] stage7_28;
   wire [4:0] stage7_29;
   wire [6:0] stage7_30;
   wire [1:0] stage7_31;
   wire [5:0] stage7_32;
   wire [0:0] stage7_33;
   wire [5:0] stage7_34;
   wire [5:0] stage7_35;
   wire [0:0] stage7_36;
   wire [1:0] stage7_37;
   wire [6:0] stage7_38;
   wire [0:0] stage7_39;
   wire [6:0] stage7_40;
   wire [4:0] stage7_41;
   wire [2:0] stage7_42;
   wire [3:0] stage7_43;
   wire [1:0] stage7_44;
   wire [4:0] stage7_45;
   wire [2:0] stage7_46;
   wire [7:0] stage7_47;
   wire [0:0] stage7_48;
   wire [1:0] stage7_49;
   wire [2:0] stage7_50;
   wire [3:0] stage7_51;
   wire [3:0] stage7_52;
   wire [5:0] stage7_53;
   wire [0:0] stage7_54;
   wire [6:0] stage7_55;
   wire [6:0] stage7_56;
   wire [1:0] stage7_57;
   wire [1:0] stage7_58;
   wire [6:0] stage7_59;
   wire [5:0] stage7_60;
   wire [1:0] stage7_61;
   wire [1:0] stage7_62;
   wire [2:0] stage7_63;
   wire [3:0] stage7_64;
   wire [2:0] stage7_65;
   wire [5:0] stage7_66;
   wire [0:0] stage7_67;
   wire [4:0] stage7_68;
   wire [4:0] stage7_69;
   wire [2:0] stage7_70;
   wire [1:0] stage7_71;
   wire [0:0] stage8_0;
   wire [1:0] stage8_1;
   wire [1:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [0:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [1:0] stage8_39;
   wire [1:0] stage8_40;
   wire [1:0] stage8_41;
   wire [1:0] stage8_42;
   wire [1:0] stage8_43;
   wire [1:0] stage8_44;
   wire [1:0] stage8_45;
   wire [0:0] stage8_46;
   wire [1:0] stage8_47;
   wire [1:0] stage8_48;
   wire [1:0] stage8_49;
   wire [1:0] stage8_50;
   wire [1:0] stage8_51;
   wire [1:0] stage8_52;
   wire [1:0] stage8_53;
   wire [1:0] stage8_54;
   wire [1:0] stage8_55;
   wire [1:0] stage8_56;
   wire [1:0] stage8_57;
   wire [1:0] stage8_58;
   wire [1:0] stage8_59;
   wire [1:0] stage8_60;
   wire [1:0] stage8_61;
   wire [1:0] stage8_62;
   wire [1:0] stage8_63;
   wire [1:0] stage8_64;
   wire [1:0] stage8_65;
   wire [1:0] stage8_66;
   wire [1:0] stage8_67;
   wire [1:0] stage8_68;
   wire [1:0] stage8_69;
   wire [1:0] stage8_70;
   wire [1:0] stage8_71;
   wire [1:0] stage8_72;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;
   assign dst41 = stage8_41;
   assign dst42 = stage8_42;
   assign dst43 = stage8_43;
   assign dst44 = stage8_44;
   assign dst45 = stage8_45;
   assign dst46 = stage8_46;
   assign dst47 = stage8_47;
   assign dst48 = stage8_48;
   assign dst49 = stage8_49;
   assign dst50 = stage8_50;
   assign dst51 = stage8_51;
   assign dst52 = stage8_52;
   assign dst53 = stage8_53;
   assign dst54 = stage8_54;
   assign dst55 = stage8_55;
   assign dst56 = stage8_56;
   assign dst57 = stage8_57;
   assign dst58 = stage8_58;
   assign dst59 = stage8_59;
   assign dst60 = stage8_60;
   assign dst61 = stage8_61;
   assign dst62 = stage8_62;
   assign dst63 = stage8_63;
   assign dst64 = stage8_64;
   assign dst65 = stage8_65;
   assign dst66 = stage8_66;
   assign dst67 = stage8_67;
   assign dst68 = stage8_68;
   assign dst69 = stage8_69;
   assign dst70 = stage8_70;
   assign dst71 = stage8_71;
   assign dst72 = stage8_72;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[2]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_1[3]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[4]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[5]},
      {stage0_2[5]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[6]},
      {stage0_2[6]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc117_4 gpc7 (
      {stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[7]},
      {stage0_2[7]},
      {stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc117_4 gpc8 (
      {stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[8]},
      {stage0_2[8]},
      {stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc117_4 gpc9 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[9]},
      {stage0_2[9]},
      {stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc117_4 gpc10 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_1[10]},
      {stage0_2[10]},
      {stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc117_4 gpc11 (
      {stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[11]},
      {stage0_2[11]},
      {stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc117_4 gpc12 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[12]},
      {stage0_2[12]},
      {stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_2[13]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_2[14]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_2[15]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_2[16]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_2[17]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_2[18]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54]},
      {stage0_2[19]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60]},
      {stage0_2[20]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66]},
      {stage0_2[21]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72]},
      {stage0_2[22]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78]},
      {stage0_2[23]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84]},
      {stage0_2[24]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90]},
      {stage0_2[25]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96]},
      {stage0_2[26]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102]},
      {stage0_2[27]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108]},
      {stage0_2[28]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114]},
      {stage0_2[29]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120]},
      {stage0_2[30]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126]},
      {stage0_2[31]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132]},
      {stage0_2[32]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138]},
      {stage0_2[33]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144]},
      {stage0_2[34]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150]},
      {stage0_2[35]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156]},
      {stage0_2[36]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162]},
      {stage0_2[37]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168]},
      {stage0_2[38]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174]},
      {stage0_2[39]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180]},
      {stage0_2[40]},
      {stage0_3[27]},
      {stage1_4[27],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186]},
      {stage0_2[41]},
      {stage0_3[28]},
      {stage1_4[28],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[29],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[30],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[31],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[32],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[33],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213]},
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77]},
      {stage1_4[34],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219]},
      {stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83]},
      {stage1_4[35],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225]},
      {stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89]},
      {stage1_4[36],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231]},
      {stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95]},
      {stage1_4[37],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage1_4[38],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243]},
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107]},
      {stage1_4[39],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249]},
      {stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113]},
      {stage1_4[40],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255]},
      {stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119]},
      {stage1_4[41],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[256], stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261]},
      {stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage1_4[42],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[262], stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267]},
      {stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage1_4[43],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273]},
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137]},
      {stage1_4[44],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279]},
      {stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143]},
      {stage1_4[45],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[280], stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285]},
      {stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage1_4[46],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[286], stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291]},
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155]},
      {stage1_4[47],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[292], stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297]},
      {stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage1_4[48],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303]},
      {stage0_2[162], stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167]},
      {stage1_4[49],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309]},
      {stage0_2[168], stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173]},
      {stage1_4[50],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[310], stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315]},
      {stage0_2[174], stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179]},
      {stage1_4[51],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[316], stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321]},
      {stage0_2[180], stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185]},
      {stage1_4[52],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[322], stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327]},
      {stage0_2[186], stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191]},
      {stage1_4[53],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333]},
      {stage0_2[192], stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197]},
      {stage1_4[54],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339]},
      {stage0_2[198], stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203]},
      {stage1_4[55],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[340], stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345]},
      {stage0_2[204], stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209]},
      {stage1_4[56],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[346], stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351]},
      {stage0_2[210], stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215]},
      {stage1_4[57],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[352], stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357]},
      {stage0_2[216], stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221]},
      {stage1_4[58],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363]},
      {stage0_2[222], stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227]},
      {stage1_4[59],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369]},
      {stage0_2[228], stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233]},
      {stage1_4[60],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[370], stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375]},
      {stage0_2[234], stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239]},
      {stage1_4[61],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[376], stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381]},
      {stage0_2[240], stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage1_4[62],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[382], stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387]},
      {stage0_2[246], stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251]},
      {stage1_4[63],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393]},
      {stage0_2[252], stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257]},
      {stage1_4[64],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399]},
      {stage0_2[258], stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263]},
      {stage1_4[65],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[400], stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405]},
      {stage0_2[264], stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269]},
      {stage1_4[66],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[406], stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411]},
      {stage0_2[270], stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275]},
      {stage1_4[67],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[412], stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417]},
      {stage0_2[276], stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281]},
      {stage1_4[68],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423]},
      {stage0_2[282], stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287]},
      {stage1_4[69],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[424], stage0_0[425], stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429]},
      {stage0_2[288], stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293]},
      {stage1_4[70],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[430], stage0_0[431], stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435]},
      {stage0_2[294], stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299]},
      {stage1_4[71],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[436], stage0_0[437], stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441]},
      {stage0_2[300], stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305]},
      {stage1_4[72],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_0[442], stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447]},
      {stage0_2[306], stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311]},
      {stage1_4[73],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192]},
      {stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage1_5[0],stage1_4[74],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198]},
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40]},
      {stage1_5[1],stage1_4[75],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204]},
      {stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46]},
      {stage1_5[2],stage1_4[76],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210]},
      {stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52]},
      {stage1_5[3],stage1_4[77],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216]},
      {stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58]},
      {stage1_5[4],stage1_4[78],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222]},
      {stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64]},
      {stage1_5[5],stage1_4[79],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228]},
      {stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70]},
      {stage1_5[6],stage1_4[80],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234]},
      {stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76]},
      {stage1_5[7],stage1_4[81],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240]},
      {stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82]},
      {stage1_5[8],stage1_4[82],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246]},
      {stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88]},
      {stage1_5[9],stage1_4[83],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252]},
      {stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94]},
      {stage1_5[10],stage1_4[84],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258]},
      {stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100]},
      {stage1_5[11],stage1_4[85],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264]},
      {stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage1_5[12],stage1_4[86],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270]},
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112]},
      {stage1_5[13],stage1_4[87],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276]},
      {stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118]},
      {stage1_5[14],stage1_4[88],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282]},
      {stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124]},
      {stage1_5[15],stage1_4[89],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288]},
      {stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130]},
      {stage1_5[16],stage1_4[90],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294]},
      {stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136]},
      {stage1_5[17],stage1_4[91],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300]},
      {stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142]},
      {stage1_5[18],stage1_4[92],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306]},
      {stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148]},
      {stage1_5[19],stage1_4[93],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[307], stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311], stage0_1[312]},
      {stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage1_5[20],stage1_4[94],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[313], stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317], stage0_1[318]},
      {stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160]},
      {stage1_5[21],stage1_4[95],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[319], stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323], stage0_1[324]},
      {stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166]},
      {stage1_5[22],stage1_4[96],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[325], stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329], stage0_1[330]},
      {stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172]},
      {stage1_5[23],stage1_4[97],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[331], stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335], stage0_1[336]},
      {stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178]},
      {stage1_5[24],stage1_4[98],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[337], stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341], stage0_1[342]},
      {stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184]},
      {stage1_5[25],stage1_4[99],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[343], stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347], stage0_1[348]},
      {stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190]},
      {stage1_5[26],stage1_4[100],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[349], stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353], stage0_1[354]},
      {stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage1_5[27],stage1_4[101],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[355], stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359], stage0_1[360]},
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202]},
      {stage1_5[28],stage1_4[102],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[361], stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365], stage0_1[366]},
      {stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208]},
      {stage1_5[29],stage1_4[103],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371], stage0_1[372]},
      {stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214]},
      {stage1_5[30],stage1_4[104],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378]},
      {stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220]},
      {stage1_5[31],stage1_4[105],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384]},
      {stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage1_5[32],stage1_4[106],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390]},
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232]},
      {stage1_5[33],stage1_4[107],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396]},
      {stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238]},
      {stage1_5[34],stage1_4[108],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402]},
      {stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244]},
      {stage1_5[35],stage1_4[109],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408]},
      {stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250]},
      {stage1_5[36],stage1_4[110],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414]},
      {stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256]},
      {stage1_5[37],stage1_4[111],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420]},
      {stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262]},
      {stage1_5[38],stage1_4[112],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426]},
      {stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268]},
      {stage1_5[39],stage1_4[113],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432]},
      {stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274]},
      {stage1_5[40],stage1_4[114],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438]},
      {stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280]},
      {stage1_5[41],stage1_4[115],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_2[312], stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[42],stage1_4[116],stage1_3[129],stage1_2[129]}
   );
   gpc606_5 gpc130 (
      {stage0_2[318], stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[43],stage1_4[117],stage1_3[130],stage1_2[130]}
   );
   gpc606_5 gpc131 (
      {stage0_2[324], stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[44],stage1_4[118],stage1_3[131],stage1_2[131]}
   );
   gpc606_5 gpc132 (
      {stage0_2[330], stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[45],stage1_4[119],stage1_3[132],stage1_2[132]}
   );
   gpc606_5 gpc133 (
      {stage0_2[336], stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[46],stage1_4[120],stage1_3[133],stage1_2[133]}
   );
   gpc606_5 gpc134 (
      {stage0_2[342], stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[47],stage1_4[121],stage1_3[134],stage1_2[134]}
   );
   gpc606_5 gpc135 (
      {stage0_2[348], stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[48],stage1_4[122],stage1_3[135],stage1_2[135]}
   );
   gpc606_5 gpc136 (
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[49],stage1_4[123],stage1_3[136],stage1_2[136]}
   );
   gpc606_5 gpc137 (
      {stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[50],stage1_4[124],stage1_3[137],stage1_2[137]}
   );
   gpc606_5 gpc138 (
      {stage0_2[366], stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[51],stage1_4[125],stage1_3[138],stage1_2[138]}
   );
   gpc606_5 gpc139 (
      {stage0_2[372], stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[52],stage1_4[126],stage1_3[139],stage1_2[139]}
   );
   gpc606_5 gpc140 (
      {stage0_2[378], stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[53],stage1_4[127],stage1_3[140],stage1_2[140]}
   );
   gpc606_5 gpc141 (
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[54],stage1_4[128],stage1_3[141],stage1_2[141]}
   );
   gpc606_5 gpc142 (
      {stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394], stage0_2[395]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[55],stage1_4[129],stage1_3[142],stage1_2[142]}
   );
   gpc606_5 gpc143 (
      {stage0_2[396], stage0_2[397], stage0_2[398], stage0_2[399], stage0_2[400], stage0_2[401]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[56],stage1_4[130],stage1_3[143],stage1_2[143]}
   );
   gpc606_5 gpc144 (
      {stage0_2[402], stage0_2[403], stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[57],stage1_4[131],stage1_3[144],stage1_2[144]}
   );
   gpc606_5 gpc145 (
      {stage0_2[408], stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[58],stage1_4[132],stage1_3[145],stage1_2[145]}
   );
   gpc606_5 gpc146 (
      {stage0_2[414], stage0_2[415], stage0_2[416], stage0_2[417], stage0_2[418], stage0_2[419]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[59],stage1_4[133],stage1_3[146],stage1_2[146]}
   );
   gpc606_5 gpc147 (
      {stage0_2[420], stage0_2[421], stage0_2[422], stage0_2[423], stage0_2[424], stage0_2[425]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[60],stage1_4[134],stage1_3[147],stage1_2[147]}
   );
   gpc606_5 gpc148 (
      {stage0_2[426], stage0_2[427], stage0_2[428], stage0_2[429], stage0_2[430], stage0_2[431]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[61],stage1_4[135],stage1_3[148],stage1_2[148]}
   );
   gpc606_5 gpc149 (
      {stage0_2[432], stage0_2[433], stage0_2[434], stage0_2[435], stage0_2[436], stage0_2[437]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[62],stage1_4[136],stage1_3[149],stage1_2[149]}
   );
   gpc606_5 gpc150 (
      {stage0_2[438], stage0_2[439], stage0_2[440], stage0_2[441], stage0_2[442], stage0_2[443]},
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage1_6[21],stage1_5[63],stage1_4[137],stage1_3[150],stage1_2[150]}
   );
   gpc606_5 gpc151 (
      {stage0_2[444], stage0_2[445], stage0_2[446], stage0_2[447], stage0_2[448], stage0_2[449]},
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage1_6[22],stage1_5[64],stage1_4[138],stage1_3[151],stage1_2[151]}
   );
   gpc606_5 gpc152 (
      {stage0_2[450], stage0_2[451], stage0_2[452], stage0_2[453], stage0_2[454], stage0_2[455]},
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage1_6[23],stage1_5[65],stage1_4[139],stage1_3[152],stage1_2[152]}
   );
   gpc606_5 gpc153 (
      {stage0_2[456], stage0_2[457], stage0_2[458], stage0_2[459], stage0_2[460], stage0_2[461]},
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage1_6[24],stage1_5[66],stage1_4[140],stage1_3[153],stage1_2[153]}
   );
   gpc606_5 gpc154 (
      {stage0_2[462], stage0_2[463], stage0_2[464], stage0_2[465], stage0_2[466], stage0_2[467]},
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage1_6[25],stage1_5[67],stage1_4[141],stage1_3[154],stage1_2[154]}
   );
   gpc606_5 gpc155 (
      {stage0_2[468], stage0_2[469], stage0_2[470], stage0_2[471], stage0_2[472], stage0_2[473]},
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage1_6[26],stage1_5[68],stage1_4[142],stage1_3[155],stage1_2[155]}
   );
   gpc606_5 gpc156 (
      {stage0_2[474], stage0_2[475], stage0_2[476], stage0_2[477], stage0_2[478], stage0_2[479]},
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage1_6[27],stage1_5[69],stage1_4[143],stage1_3[156],stage1_2[156]}
   );
   gpc606_5 gpc157 (
      {stage0_2[480], stage0_2[481], stage0_2[482], stage0_2[483], stage0_2[484], stage0_2[485]},
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage1_6[28],stage1_5[70],stage1_4[144],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285]},
      {stage0_4[174]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[29],stage1_5[71],stage1_4[145],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[286], stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290]},
      {stage0_4[175]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[30],stage1_5[72],stage1_4[146],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295]},
      {stage0_4[176]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[31],stage1_5[73],stage1_4[147],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[296], stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300]},
      {stage0_4[177]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[32],stage1_5[74],stage1_4[148],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[301], stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305]},
      {stage0_4[178]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[33],stage1_5[75],stage1_4[149],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[306], stage0_3[307], stage0_3[308], stage0_3[309], stage0_3[310]},
      {stage0_4[179]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[34],stage1_5[76],stage1_4[150],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[311], stage0_3[312], stage0_3[313], stage0_3[314], stage0_3[315]},
      {stage0_4[180]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[35],stage1_5[77],stage1_4[151],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[316], stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320]},
      {stage0_4[181]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[36],stage1_5[78],stage1_4[152],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[321], stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325]},
      {stage0_4[182]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[37],stage1_5[79],stage1_4[153],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[326], stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330]},
      {stage0_4[183]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[38],stage1_5[80],stage1_4[154],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[331], stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335]},
      {stage0_4[184]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[39],stage1_5[81],stage1_4[155],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[336], stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340]},
      {stage0_4[185]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[40],stage1_5[82],stage1_4[156],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[341], stage0_3[342], stage0_3[343], stage0_3[344], stage0_3[345]},
      {stage0_4[186]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[41],stage1_5[83],stage1_4[157],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[346], stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350]},
      {stage0_4[187]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[42],stage1_5[84],stage1_4[158],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[351], stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355]},
      {stage0_4[188]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[43],stage1_5[85],stage1_4[159],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[356], stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360]},
      {stage0_4[189]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[44],stage1_5[86],stage1_4[160],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[361], stage0_3[362], stage0_3[363], stage0_3[364], stage0_3[365]},
      {stage0_4[190]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[45],stage1_5[87],stage1_4[161],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[366], stage0_3[367], stage0_3[368], stage0_3[369], stage0_3[370]},
      {stage0_4[191]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[46],stage1_5[88],stage1_4[162],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[371], stage0_3[372], stage0_3[373], stage0_3[374], stage0_3[375]},
      {stage0_4[192]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[47],stage1_5[89],stage1_4[163],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage0_4[193]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[48],stage1_5[90],stage1_4[164],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385]},
      {stage0_4[194]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[49],stage1_5[91],stage1_4[165],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[386], stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390]},
      {stage0_4[195]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[50],stage1_5[92],stage1_4[166],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[391], stage0_3[392], stage0_3[393], stage0_3[394], stage0_3[395]},
      {stage0_4[196]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[51],stage1_5[93],stage1_4[167],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[396], stage0_3[397], stage0_3[398], stage0_3[399], stage0_3[400]},
      {stage0_4[197]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[52],stage1_5[94],stage1_4[168],stage1_3[181]}
   );
   gpc615_5 gpc182 (
      {stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404], stage0_3[405]},
      {stage0_4[198]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[53],stage1_5[95],stage1_4[169],stage1_3[182]}
   );
   gpc615_5 gpc183 (
      {stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage0_4[199]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[54],stage1_5[96],stage1_4[170],stage1_3[183]}
   );
   gpc615_5 gpc184 (
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415]},
      {stage0_4[200]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[55],stage1_5[97],stage1_4[171],stage1_3[184]}
   );
   gpc615_5 gpc185 (
      {stage0_3[416], stage0_3[417], stage0_3[418], stage0_3[419], stage0_3[420]},
      {stage0_4[201]},
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage1_7[27],stage1_6[56],stage1_5[98],stage1_4[172],stage1_3[185]}
   );
   gpc615_5 gpc186 (
      {stage0_3[421], stage0_3[422], stage0_3[423], stage0_3[424], stage0_3[425]},
      {stage0_4[202]},
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage1_7[28],stage1_6[57],stage1_5[99],stage1_4[173],stage1_3[186]}
   );
   gpc615_5 gpc187 (
      {stage0_3[426], stage0_3[427], stage0_3[428], stage0_3[429], stage0_3[430]},
      {stage0_4[203]},
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage1_7[29],stage1_6[58],stage1_5[100],stage1_4[174],stage1_3[187]}
   );
   gpc615_5 gpc188 (
      {stage0_3[431], stage0_3[432], stage0_3[433], stage0_3[434], stage0_3[435]},
      {stage0_4[204]},
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage1_7[30],stage1_6[59],stage1_5[101],stage1_4[175],stage1_3[188]}
   );
   gpc615_5 gpc189 (
      {stage0_3[436], stage0_3[437], stage0_3[438], stage0_3[439], stage0_3[440]},
      {stage0_4[205]},
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage1_7[31],stage1_6[60],stage1_5[102],stage1_4[176],stage1_3[189]}
   );
   gpc615_5 gpc190 (
      {stage0_3[441], stage0_3[442], stage0_3[443], stage0_3[444], stage0_3[445]},
      {stage0_4[206]},
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage1_7[32],stage1_6[61],stage1_5[103],stage1_4[177],stage1_3[190]}
   );
   gpc615_5 gpc191 (
      {stage0_3[446], stage0_3[447], stage0_3[448], stage0_3[449], stage0_3[450]},
      {stage0_4[207]},
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage1_7[33],stage1_6[62],stage1_5[104],stage1_4[178],stage1_3[191]}
   );
   gpc615_5 gpc192 (
      {stage0_3[451], stage0_3[452], stage0_3[453], stage0_3[454], stage0_3[455]},
      {stage0_4[208]},
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage1_7[34],stage1_6[63],stage1_5[105],stage1_4[179],stage1_3[192]}
   );
   gpc615_5 gpc193 (
      {stage0_3[456], stage0_3[457], stage0_3[458], stage0_3[459], stage0_3[460]},
      {stage0_4[209]},
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage1_7[35],stage1_6[64],stage1_5[106],stage1_4[180],stage1_3[193]}
   );
   gpc615_5 gpc194 (
      {stage0_3[461], stage0_3[462], stage0_3[463], stage0_3[464], stage0_3[465]},
      {stage0_4[210]},
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage1_7[36],stage1_6[65],stage1_5[107],stage1_4[181],stage1_3[194]}
   );
   gpc606_5 gpc195 (
      {stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[37],stage1_6[66],stage1_5[108],stage1_4[182]}
   );
   gpc606_5 gpc196 (
      {stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[38],stage1_6[67],stage1_5[109],stage1_4[183]}
   );
   gpc606_5 gpc197 (
      {stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[39],stage1_6[68],stage1_5[110],stage1_4[184]}
   );
   gpc606_5 gpc198 (
      {stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[40],stage1_6[69],stage1_5[111],stage1_4[185]}
   );
   gpc606_5 gpc199 (
      {stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[41],stage1_6[70],stage1_5[112],stage1_4[186]}
   );
   gpc606_5 gpc200 (
      {stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[42],stage1_6[71],stage1_5[113],stage1_4[187]}
   );
   gpc606_5 gpc201 (
      {stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[43],stage1_6[72],stage1_5[114],stage1_4[188]}
   );
   gpc606_5 gpc202 (
      {stage0_4[253], stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[44],stage1_6[73],stage1_5[115],stage1_4[189]}
   );
   gpc606_5 gpc203 (
      {stage0_4[259], stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[45],stage1_6[74],stage1_5[116],stage1_4[190]}
   );
   gpc606_5 gpc204 (
      {stage0_4[265], stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[46],stage1_6[75],stage1_5[117],stage1_4[191]}
   );
   gpc606_5 gpc205 (
      {stage0_4[271], stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[47],stage1_6[76],stage1_5[118],stage1_4[192]}
   );
   gpc606_5 gpc206 (
      {stage0_4[277], stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[48],stage1_6[77],stage1_5[119],stage1_4[193]}
   );
   gpc606_5 gpc207 (
      {stage0_4[283], stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[49],stage1_6[78],stage1_5[120],stage1_4[194]}
   );
   gpc606_5 gpc208 (
      {stage0_4[289], stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[50],stage1_6[79],stage1_5[121],stage1_4[195]}
   );
   gpc606_5 gpc209 (
      {stage0_4[295], stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[51],stage1_6[80],stage1_5[122],stage1_4[196]}
   );
   gpc606_5 gpc210 (
      {stage0_4[301], stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[52],stage1_6[81],stage1_5[123],stage1_4[197]}
   );
   gpc606_5 gpc211 (
      {stage0_4[307], stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[53],stage1_6[82],stage1_5[124],stage1_4[198]}
   );
   gpc606_5 gpc212 (
      {stage0_4[313], stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[54],stage1_6[83],stage1_5[125],stage1_4[199]}
   );
   gpc606_5 gpc213 (
      {stage0_4[319], stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[55],stage1_6[84],stage1_5[126],stage1_4[200]}
   );
   gpc606_5 gpc214 (
      {stage0_4[325], stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[56],stage1_6[85],stage1_5[127],stage1_4[201]}
   );
   gpc606_5 gpc215 (
      {stage0_4[331], stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[57],stage1_6[86],stage1_5[128],stage1_4[202]}
   );
   gpc606_5 gpc216 (
      {stage0_4[337], stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[58],stage1_6[87],stage1_5[129],stage1_4[203]}
   );
   gpc606_5 gpc217 (
      {stage0_4[343], stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[59],stage1_6[88],stage1_5[130],stage1_4[204]}
   );
   gpc606_5 gpc218 (
      {stage0_4[349], stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[60],stage1_6[89],stage1_5[131],stage1_4[205]}
   );
   gpc606_5 gpc219 (
      {stage0_4[355], stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[61],stage1_6[90],stage1_5[132],stage1_4[206]}
   );
   gpc606_5 gpc220 (
      {stage0_4[361], stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[62],stage1_6[91],stage1_5[133],stage1_4[207]}
   );
   gpc606_5 gpc221 (
      {stage0_4[367], stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[63],stage1_6[92],stage1_5[134],stage1_4[208]}
   );
   gpc606_5 gpc222 (
      {stage0_4[373], stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[64],stage1_6[93],stage1_5[135],stage1_4[209]}
   );
   gpc606_5 gpc223 (
      {stage0_4[379], stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[65],stage1_6[94],stage1_5[136],stage1_4[210]}
   );
   gpc606_5 gpc224 (
      {stage0_4[385], stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[66],stage1_6[95],stage1_5[137],stage1_4[211]}
   );
   gpc606_5 gpc225 (
      {stage0_4[391], stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[67],stage1_6[96],stage1_5[138],stage1_4[212]}
   );
   gpc606_5 gpc226 (
      {stage0_4[397], stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[68],stage1_6[97],stage1_5[139],stage1_4[213]}
   );
   gpc606_5 gpc227 (
      {stage0_4[403], stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[69],stage1_6[98],stage1_5[140],stage1_4[214]}
   );
   gpc606_5 gpc228 (
      {stage0_4[409], stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[70],stage1_6[99],stage1_5[141],stage1_4[215]}
   );
   gpc606_5 gpc229 (
      {stage0_4[415], stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[71],stage1_6[100],stage1_5[142],stage1_4[216]}
   );
   gpc606_5 gpc230 (
      {stage0_4[421], stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[72],stage1_6[101],stage1_5[143],stage1_4[217]}
   );
   gpc606_5 gpc231 (
      {stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[73],stage1_6[102],stage1_5[144],stage1_4[218]}
   );
   gpc606_5 gpc232 (
      {stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[74],stage1_6[103],stage1_5[145],stage1_4[219]}
   );
   gpc606_5 gpc233 (
      {stage0_4[439], stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[75],stage1_6[104],stage1_5[146],stage1_4[220]}
   );
   gpc606_5 gpc234 (
      {stage0_4[445], stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[76],stage1_6[105],stage1_5[147],stage1_4[221]}
   );
   gpc606_5 gpc235 (
      {stage0_4[451], stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[77],stage1_6[106],stage1_5[148],stage1_4[222]}
   );
   gpc606_5 gpc236 (
      {stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461], stage0_4[462]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[78],stage1_6[107],stage1_5[149],stage1_4[223]}
   );
   gpc606_5 gpc237 (
      {stage0_4[463], stage0_4[464], stage0_4[465], stage0_4[466], stage0_4[467], stage0_4[468]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[79],stage1_6[108],stage1_5[150],stage1_4[224]}
   );
   gpc606_5 gpc238 (
      {stage0_4[469], stage0_4[470], stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[80],stage1_6[109],stage1_5[151],stage1_4[225]}
   );
   gpc606_5 gpc239 (
      {stage0_4[475], stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[81],stage1_6[110],stage1_5[152],stage1_4[226]}
   );
   gpc606_5 gpc240 (
      {stage0_4[481], stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], 1'b0},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[82],stage1_6[111],stage1_5[153],stage1_4[227]}
   );
   gpc606_5 gpc241 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[46],stage1_7[83],stage1_6[112],stage1_5[154]}
   );
   gpc606_5 gpc242 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[47],stage1_7[84],stage1_6[113],stage1_5[155]}
   );
   gpc606_5 gpc243 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[48],stage1_7[85],stage1_6[114],stage1_5[156]}
   );
   gpc606_5 gpc244 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[49],stage1_7[86],stage1_6[115],stage1_5[157]}
   );
   gpc606_5 gpc245 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[50],stage1_7[87],stage1_6[116],stage1_5[158]}
   );
   gpc606_5 gpc246 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[51],stage1_7[88],stage1_6[117],stage1_5[159]}
   );
   gpc606_5 gpc247 (
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[52],stage1_7[89],stage1_6[118],stage1_5[160]}
   );
   gpc606_5 gpc248 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[53],stage1_7[90],stage1_6[119],stage1_5[161]}
   );
   gpc606_5 gpc249 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[54],stage1_7[91],stage1_6[120],stage1_5[162]}
   );
   gpc606_5 gpc250 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[55],stage1_7[92],stage1_6[121],stage1_5[163]}
   );
   gpc606_5 gpc251 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[56],stage1_7[93],stage1_6[122],stage1_5[164]}
   );
   gpc606_5 gpc252 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[57],stage1_7[94],stage1_6[123],stage1_5[165]}
   );
   gpc606_5 gpc253 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[58],stage1_7[95],stage1_6[124],stage1_5[166]}
   );
   gpc606_5 gpc254 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[59],stage1_7[96],stage1_6[125],stage1_5[167]}
   );
   gpc606_5 gpc255 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[60],stage1_7[97],stage1_6[126],stage1_5[168]}
   );
   gpc606_5 gpc256 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[61],stage1_7[98],stage1_6[127],stage1_5[169]}
   );
   gpc606_5 gpc257 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[62],stage1_7[99],stage1_6[128],stage1_5[170]}
   );
   gpc606_5 gpc258 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[63],stage1_7[100],stage1_6[129],stage1_5[171]}
   );
   gpc606_5 gpc259 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[64],stage1_7[101],stage1_6[130],stage1_5[172]}
   );
   gpc606_5 gpc260 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[65],stage1_7[102],stage1_6[131],stage1_5[173]}
   );
   gpc606_5 gpc261 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[66],stage1_7[103],stage1_6[132],stage1_5[174]}
   );
   gpc606_5 gpc262 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[67],stage1_7[104],stage1_6[133],stage1_5[175]}
   );
   gpc606_5 gpc263 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[68],stage1_7[105],stage1_6[134],stage1_5[176]}
   );
   gpc606_5 gpc264 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[69],stage1_7[106],stage1_6[135],stage1_5[177]}
   );
   gpc606_5 gpc265 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[70],stage1_7[107],stage1_6[136],stage1_5[178]}
   );
   gpc606_5 gpc266 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[71],stage1_7[108],stage1_6[137],stage1_5[179]}
   );
   gpc606_5 gpc267 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[72],stage1_7[109],stage1_6[138],stage1_5[180]}
   );
   gpc606_5 gpc268 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[73],stage1_7[110],stage1_6[139],stage1_5[181]}
   );
   gpc606_5 gpc269 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[74],stage1_7[111],stage1_6[140],stage1_5[182]}
   );
   gpc606_5 gpc270 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[75],stage1_7[112],stage1_6[141],stage1_5[183]}
   );
   gpc606_5 gpc271 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[76],stage1_7[113],stage1_6[142],stage1_5[184]}
   );
   gpc606_5 gpc272 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[77],stage1_7[114],stage1_6[143],stage1_5[185]}
   );
   gpc606_5 gpc273 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[78],stage1_7[115],stage1_6[144],stage1_5[186]}
   );
   gpc606_5 gpc274 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[79],stage1_7[116],stage1_6[145],stage1_5[187]}
   );
   gpc606_5 gpc275 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[80],stage1_7[117],stage1_6[146],stage1_5[188]}
   );
   gpc606_5 gpc276 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[81],stage1_7[118],stage1_6[147],stage1_5[189]}
   );
   gpc606_5 gpc277 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[82],stage1_7[119],stage1_6[148],stage1_5[190]}
   );
   gpc606_5 gpc278 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[83],stage1_7[120],stage1_6[149],stage1_5[191]}
   );
   gpc606_5 gpc279 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[84],stage1_7[121],stage1_6[150],stage1_5[192]}
   );
   gpc606_5 gpc280 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[85],stage1_7[122],stage1_6[151],stage1_5[193]}
   );
   gpc606_5 gpc281 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[86],stage1_7[123],stage1_6[152],stage1_5[194]}
   );
   gpc606_5 gpc282 (
      {stage0_5[468], stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[87],stage1_7[124],stage1_6[153],stage1_5[195]}
   );
   gpc606_5 gpc283 (
      {stage0_5[474], stage0_5[475], stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[88],stage1_7[125],stage1_6[154],stage1_5[196]}
   );
   gpc606_5 gpc284 (
      {stage0_5[480], stage0_5[481], stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[89],stage1_7[126],stage1_6[155],stage1_5[197]}
   );
   gpc615_5 gpc285 (
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280]},
      {stage0_7[264]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[44],stage1_8[90],stage1_7[127],stage1_6[156]}
   );
   gpc615_5 gpc286 (
      {stage0_6[281], stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285]},
      {stage0_7[265]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[45],stage1_8[91],stage1_7[128],stage1_6[157]}
   );
   gpc615_5 gpc287 (
      {stage0_6[286], stage0_6[287], stage0_6[288], stage0_6[289], stage0_6[290]},
      {stage0_7[266]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[46],stage1_8[92],stage1_7[129],stage1_6[158]}
   );
   gpc615_5 gpc288 (
      {stage0_6[291], stage0_6[292], stage0_6[293], stage0_6[294], stage0_6[295]},
      {stage0_7[267]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[47],stage1_8[93],stage1_7[130],stage1_6[159]}
   );
   gpc615_5 gpc289 (
      {stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299], stage0_6[300]},
      {stage0_7[268]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[48],stage1_8[94],stage1_7[131],stage1_6[160]}
   );
   gpc615_5 gpc290 (
      {stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage0_7[269]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[49],stage1_8[95],stage1_7[132],stage1_6[161]}
   );
   gpc615_5 gpc291 (
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310]},
      {stage0_7[270]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[50],stage1_8[96],stage1_7[133],stage1_6[162]}
   );
   gpc615_5 gpc292 (
      {stage0_6[311], stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315]},
      {stage0_7[271]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[51],stage1_8[97],stage1_7[134],stage1_6[163]}
   );
   gpc615_5 gpc293 (
      {stage0_6[316], stage0_6[317], stage0_6[318], stage0_6[319], stage0_6[320]},
      {stage0_7[272]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[52],stage1_8[98],stage1_7[135],stage1_6[164]}
   );
   gpc615_5 gpc294 (
      {stage0_6[321], stage0_6[322], stage0_6[323], stage0_6[324], stage0_6[325]},
      {stage0_7[273]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[53],stage1_8[99],stage1_7[136],stage1_6[165]}
   );
   gpc615_5 gpc295 (
      {stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329], stage0_6[330]},
      {stage0_7[274]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[54],stage1_8[100],stage1_7[137],stage1_6[166]}
   );
   gpc615_5 gpc296 (
      {stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage0_7[275]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[55],stage1_8[101],stage1_7[138],stage1_6[167]}
   );
   gpc615_5 gpc297 (
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340]},
      {stage0_7[276]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[56],stage1_8[102],stage1_7[139],stage1_6[168]}
   );
   gpc615_5 gpc298 (
      {stage0_6[341], stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345]},
      {stage0_7[277]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[57],stage1_8[103],stage1_7[140],stage1_6[169]}
   );
   gpc615_5 gpc299 (
      {stage0_6[346], stage0_6[347], stage0_6[348], stage0_6[349], stage0_6[350]},
      {stage0_7[278]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[58],stage1_8[104],stage1_7[141],stage1_6[170]}
   );
   gpc615_5 gpc300 (
      {stage0_6[351], stage0_6[352], stage0_6[353], stage0_6[354], stage0_6[355]},
      {stage0_7[279]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[59],stage1_8[105],stage1_7[142],stage1_6[171]}
   );
   gpc615_5 gpc301 (
      {stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359], stage0_6[360]},
      {stage0_7[280]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[60],stage1_8[106],stage1_7[143],stage1_6[172]}
   );
   gpc615_5 gpc302 (
      {stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage0_7[281]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[61],stage1_8[107],stage1_7[144],stage1_6[173]}
   );
   gpc615_5 gpc303 (
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370]},
      {stage0_7[282]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[62],stage1_8[108],stage1_7[145],stage1_6[174]}
   );
   gpc615_5 gpc304 (
      {stage0_6[371], stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375]},
      {stage0_7[283]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[63],stage1_8[109],stage1_7[146],stage1_6[175]}
   );
   gpc615_5 gpc305 (
      {stage0_6[376], stage0_6[377], stage0_6[378], stage0_6[379], stage0_6[380]},
      {stage0_7[284]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[64],stage1_8[110],stage1_7[147],stage1_6[176]}
   );
   gpc615_5 gpc306 (
      {stage0_6[381], stage0_6[382], stage0_6[383], stage0_6[384], stage0_6[385]},
      {stage0_7[285]},
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage1_10[21],stage1_9[65],stage1_8[111],stage1_7[148],stage1_6[177]}
   );
   gpc615_5 gpc307 (
      {stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389], stage0_6[390]},
      {stage0_7[286]},
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage1_10[22],stage1_9[66],stage1_8[112],stage1_7[149],stage1_6[178]}
   );
   gpc615_5 gpc308 (
      {stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage0_7[287]},
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage1_10[23],stage1_9[67],stage1_8[113],stage1_7[150],stage1_6[179]}
   );
   gpc615_5 gpc309 (
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400]},
      {stage0_7[288]},
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage1_10[24],stage1_9[68],stage1_8[114],stage1_7[151],stage1_6[180]}
   );
   gpc615_5 gpc310 (
      {stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405]},
      {stage0_7[289]},
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage1_10[25],stage1_9[69],stage1_8[115],stage1_7[152],stage1_6[181]}
   );
   gpc615_5 gpc311 (
      {stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409], stage0_6[410]},
      {stage0_7[290]},
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage1_10[26],stage1_9[70],stage1_8[116],stage1_7[153],stage1_6[182]}
   );
   gpc615_5 gpc312 (
      {stage0_6[411], stage0_6[412], stage0_6[413], stage0_6[414], stage0_6[415]},
      {stage0_7[291]},
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage1_10[27],stage1_9[71],stage1_8[117],stage1_7[154],stage1_6[183]}
   );
   gpc615_5 gpc313 (
      {stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419], stage0_6[420]},
      {stage0_7[292]},
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage1_10[28],stage1_9[72],stage1_8[118],stage1_7[155],stage1_6[184]}
   );
   gpc615_5 gpc314 (
      {stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage0_7[293]},
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage1_10[29],stage1_9[73],stage1_8[119],stage1_7[156],stage1_6[185]}
   );
   gpc615_5 gpc315 (
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430]},
      {stage0_7[294]},
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage1_10[30],stage1_9[74],stage1_8[120],stage1_7[157],stage1_6[186]}
   );
   gpc615_5 gpc316 (
      {stage0_6[431], stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435]},
      {stage0_7[295]},
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage1_10[31],stage1_9[75],stage1_8[121],stage1_7[158],stage1_6[187]}
   );
   gpc615_5 gpc317 (
      {stage0_6[436], stage0_6[437], stage0_6[438], stage0_6[439], stage0_6[440]},
      {stage0_7[296]},
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage1_10[32],stage1_9[76],stage1_8[122],stage1_7[159],stage1_6[188]}
   );
   gpc615_5 gpc318 (
      {stage0_6[441], stage0_6[442], stage0_6[443], stage0_6[444], stage0_6[445]},
      {stage0_7[297]},
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage1_10[33],stage1_9[77],stage1_8[123],stage1_7[160],stage1_6[189]}
   );
   gpc615_5 gpc319 (
      {stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449], stage0_6[450]},
      {stage0_7[298]},
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage1_10[34],stage1_9[78],stage1_8[124],stage1_7[161],stage1_6[190]}
   );
   gpc615_5 gpc320 (
      {stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455]},
      {stage0_7[299]},
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215]},
      {stage1_10[35],stage1_9[79],stage1_8[125],stage1_7[162],stage1_6[191]}
   );
   gpc615_5 gpc321 (
      {stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459], stage0_6[460]},
      {stage0_7[300]},
      {stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221]},
      {stage1_10[36],stage1_9[80],stage1_8[126],stage1_7[163],stage1_6[192]}
   );
   gpc615_5 gpc322 (
      {stage0_6[461], stage0_6[462], stage0_6[463], stage0_6[464], stage0_6[465]},
      {stage0_7[301]},
      {stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage1_10[37],stage1_9[81],stage1_8[127],stage1_7[164],stage1_6[193]}
   );
   gpc615_5 gpc323 (
      {stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305], stage0_7[306]},
      {stage0_8[228]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[38],stage1_9[82],stage1_8[128],stage1_7[165]}
   );
   gpc615_5 gpc324 (
      {stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage0_8[229]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[39],stage1_9[83],stage1_8[129],stage1_7[166]}
   );
   gpc615_5 gpc325 (
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316]},
      {stage0_8[230]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[40],stage1_9[84],stage1_8[130],stage1_7[167]}
   );
   gpc615_5 gpc326 (
      {stage0_7[317], stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321]},
      {stage0_8[231]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[41],stage1_9[85],stage1_8[131],stage1_7[168]}
   );
   gpc615_5 gpc327 (
      {stage0_7[322], stage0_7[323], stage0_7[324], stage0_7[325], stage0_7[326]},
      {stage0_8[232]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[42],stage1_9[86],stage1_8[132],stage1_7[169]}
   );
   gpc615_5 gpc328 (
      {stage0_7[327], stage0_7[328], stage0_7[329], stage0_7[330], stage0_7[331]},
      {stage0_8[233]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[43],stage1_9[87],stage1_8[133],stage1_7[170]}
   );
   gpc615_5 gpc329 (
      {stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335], stage0_7[336]},
      {stage0_8[234]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[44],stage1_9[88],stage1_8[134],stage1_7[171]}
   );
   gpc615_5 gpc330 (
      {stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340], stage0_7[341]},
      {stage0_8[235]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[45],stage1_9[89],stage1_8[135],stage1_7[172]}
   );
   gpc615_5 gpc331 (
      {stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345], stage0_7[346]},
      {stage0_8[236]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[46],stage1_9[90],stage1_8[136],stage1_7[173]}
   );
   gpc615_5 gpc332 (
      {stage0_7[347], stage0_7[348], stage0_7[349], stage0_7[350], stage0_7[351]},
      {stage0_8[237]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[47],stage1_9[91],stage1_8[137],stage1_7[174]}
   );
   gpc615_5 gpc333 (
      {stage0_7[352], stage0_7[353], stage0_7[354], stage0_7[355], stage0_7[356]},
      {stage0_8[238]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[48],stage1_9[92],stage1_8[138],stage1_7[175]}
   );
   gpc615_5 gpc334 (
      {stage0_7[357], stage0_7[358], stage0_7[359], stage0_7[360], stage0_7[361]},
      {stage0_8[239]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[49],stage1_9[93],stage1_8[139],stage1_7[176]}
   );
   gpc615_5 gpc335 (
      {stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365], stage0_7[366]},
      {stage0_8[240]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[50],stage1_9[94],stage1_8[140],stage1_7[177]}
   );
   gpc615_5 gpc336 (
      {stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370], stage0_7[371]},
      {stage0_8[241]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[51],stage1_9[95],stage1_8[141],stage1_7[178]}
   );
   gpc615_5 gpc337 (
      {stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375], stage0_7[376]},
      {stage0_8[242]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[52],stage1_9[96],stage1_8[142],stage1_7[179]}
   );
   gpc615_5 gpc338 (
      {stage0_7[377], stage0_7[378], stage0_7[379], stage0_7[380], stage0_7[381]},
      {stage0_8[243]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[53],stage1_9[97],stage1_8[143],stage1_7[180]}
   );
   gpc615_5 gpc339 (
      {stage0_7[382], stage0_7[383], stage0_7[384], stage0_7[385], stage0_7[386]},
      {stage0_8[244]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[54],stage1_9[98],stage1_8[144],stage1_7[181]}
   );
   gpc615_5 gpc340 (
      {stage0_7[387], stage0_7[388], stage0_7[389], stage0_7[390], stage0_7[391]},
      {stage0_8[245]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[55],stage1_9[99],stage1_8[145],stage1_7[182]}
   );
   gpc615_5 gpc341 (
      {stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395], stage0_7[396]},
      {stage0_8[246]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[56],stage1_9[100],stage1_8[146],stage1_7[183]}
   );
   gpc615_5 gpc342 (
      {stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400], stage0_7[401]},
      {stage0_8[247]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[57],stage1_9[101],stage1_8[147],stage1_7[184]}
   );
   gpc615_5 gpc343 (
      {stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406]},
      {stage0_8[248]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[58],stage1_9[102],stage1_8[148],stage1_7[185]}
   );
   gpc615_5 gpc344 (
      {stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411]},
      {stage0_8[249]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[59],stage1_9[103],stage1_8[149],stage1_7[186]}
   );
   gpc615_5 gpc345 (
      {stage0_7[412], stage0_7[413], stage0_7[414], stage0_7[415], stage0_7[416]},
      {stage0_8[250]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[60],stage1_9[104],stage1_8[150],stage1_7[187]}
   );
   gpc615_5 gpc346 (
      {stage0_7[417], stage0_7[418], stage0_7[419], stage0_7[420], stage0_7[421]},
      {stage0_8[251]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[61],stage1_9[105],stage1_8[151],stage1_7[188]}
   );
   gpc615_5 gpc347 (
      {stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425], stage0_7[426]},
      {stage0_8[252]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[62],stage1_9[106],stage1_8[152],stage1_7[189]}
   );
   gpc615_5 gpc348 (
      {stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430], stage0_7[431]},
      {stage0_8[253]},
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage1_11[25],stage1_10[63],stage1_9[107],stage1_8[153],stage1_7[190]}
   );
   gpc615_5 gpc349 (
      {stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436]},
      {stage0_8[254]},
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage1_11[26],stage1_10[64],stage1_9[108],stage1_8[154],stage1_7[191]}
   );
   gpc615_5 gpc350 (
      {stage0_7[437], stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441]},
      {stage0_8[255]},
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage1_11[27],stage1_10[65],stage1_9[109],stage1_8[155],stage1_7[192]}
   );
   gpc615_5 gpc351 (
      {stage0_7[442], stage0_7[443], stage0_7[444], stage0_7[445], stage0_7[446]},
      {stage0_8[256]},
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage1_11[28],stage1_10[66],stage1_9[110],stage1_8[156],stage1_7[193]}
   );
   gpc615_5 gpc352 (
      {stage0_7[447], stage0_7[448], stage0_7[449], stage0_7[450], stage0_7[451]},
      {stage0_8[257]},
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage1_11[29],stage1_10[67],stage1_9[111],stage1_8[157],stage1_7[194]}
   );
   gpc615_5 gpc353 (
      {stage0_7[452], stage0_7[453], stage0_7[454], stage0_7[455], stage0_7[456]},
      {stage0_8[258]},
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage1_11[30],stage1_10[68],stage1_9[112],stage1_8[158],stage1_7[195]}
   );
   gpc615_5 gpc354 (
      {stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460], stage0_7[461]},
      {stage0_8[259]},
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage1_11[31],stage1_10[69],stage1_9[113],stage1_8[159],stage1_7[196]}
   );
   gpc606_5 gpc355 (
      {stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264], stage0_8[265]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[32],stage1_10[70],stage1_9[114],stage1_8[160]}
   );
   gpc606_5 gpc356 (
      {stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270], stage0_8[271]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[33],stage1_10[71],stage1_9[115],stage1_8[161]}
   );
   gpc606_5 gpc357 (
      {stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276], stage0_8[277]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[34],stage1_10[72],stage1_9[116],stage1_8[162]}
   );
   gpc606_5 gpc358 (
      {stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282], stage0_8[283]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[35],stage1_10[73],stage1_9[117],stage1_8[163]}
   );
   gpc606_5 gpc359 (
      {stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288], stage0_8[289]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[36],stage1_10[74],stage1_9[118],stage1_8[164]}
   );
   gpc606_5 gpc360 (
      {stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294], stage0_8[295]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[37],stage1_10[75],stage1_9[119],stage1_8[165]}
   );
   gpc606_5 gpc361 (
      {stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300], stage0_8[301]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[38],stage1_10[76],stage1_9[120],stage1_8[166]}
   );
   gpc606_5 gpc362 (
      {stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306], stage0_8[307]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[39],stage1_10[77],stage1_9[121],stage1_8[167]}
   );
   gpc606_5 gpc363 (
      {stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312], stage0_8[313]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[40],stage1_10[78],stage1_9[122],stage1_8[168]}
   );
   gpc606_5 gpc364 (
      {stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318], stage0_8[319]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[41],stage1_10[79],stage1_9[123],stage1_8[169]}
   );
   gpc606_5 gpc365 (
      {stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324], stage0_8[325]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[42],stage1_10[80],stage1_9[124],stage1_8[170]}
   );
   gpc606_5 gpc366 (
      {stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330], stage0_8[331]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[43],stage1_10[81],stage1_9[125],stage1_8[171]}
   );
   gpc606_5 gpc367 (
      {stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336], stage0_8[337]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[44],stage1_10[82],stage1_9[126],stage1_8[172]}
   );
   gpc606_5 gpc368 (
      {stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342], stage0_8[343]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[45],stage1_10[83],stage1_9[127],stage1_8[173]}
   );
   gpc606_5 gpc369 (
      {stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348], stage0_8[349]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[46],stage1_10[84],stage1_9[128],stage1_8[174]}
   );
   gpc606_5 gpc370 (
      {stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354], stage0_8[355]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[47],stage1_10[85],stage1_9[129],stage1_8[175]}
   );
   gpc606_5 gpc371 (
      {stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360], stage0_8[361]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[48],stage1_10[86],stage1_9[130],stage1_8[176]}
   );
   gpc606_5 gpc372 (
      {stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366], stage0_8[367]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[49],stage1_10[87],stage1_9[131],stage1_8[177]}
   );
   gpc606_5 gpc373 (
      {stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372], stage0_8[373]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[50],stage1_10[88],stage1_9[132],stage1_8[178]}
   );
   gpc606_5 gpc374 (
      {stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378], stage0_8[379]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[51],stage1_10[89],stage1_9[133],stage1_8[179]}
   );
   gpc606_5 gpc375 (
      {stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384], stage0_8[385]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[52],stage1_10[90],stage1_9[134],stage1_8[180]}
   );
   gpc606_5 gpc376 (
      {stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390], stage0_8[391]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[53],stage1_10[91],stage1_9[135],stage1_8[181]}
   );
   gpc606_5 gpc377 (
      {stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396], stage0_8[397]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[54],stage1_10[92],stage1_9[136],stage1_8[182]}
   );
   gpc606_5 gpc378 (
      {stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402], stage0_8[403]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[55],stage1_10[93],stage1_9[137],stage1_8[183]}
   );
   gpc606_5 gpc379 (
      {stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408], stage0_8[409]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[56],stage1_10[94],stage1_9[138],stage1_8[184]}
   );
   gpc606_5 gpc380 (
      {stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414], stage0_8[415]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[57],stage1_10[95],stage1_9[139],stage1_8[185]}
   );
   gpc606_5 gpc381 (
      {stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420], stage0_8[421]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[58],stage1_10[96],stage1_9[140],stage1_8[186]}
   );
   gpc606_5 gpc382 (
      {stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426], stage0_8[427]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[59],stage1_10[97],stage1_9[141],stage1_8[187]}
   );
   gpc606_5 gpc383 (
      {stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432], stage0_8[433]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[60],stage1_10[98],stage1_9[142],stage1_8[188]}
   );
   gpc606_5 gpc384 (
      {stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438], stage0_8[439]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[61],stage1_10[99],stage1_9[143],stage1_8[189]}
   );
   gpc606_5 gpc385 (
      {stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444], stage0_8[445]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[62],stage1_10[100],stage1_9[144],stage1_8[190]}
   );
   gpc606_5 gpc386 (
      {stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450], stage0_8[451]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[63],stage1_10[101],stage1_9[145],stage1_8[191]}
   );
   gpc606_5 gpc387 (
      {stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456], stage0_8[457]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[64],stage1_10[102],stage1_9[146],stage1_8[192]}
   );
   gpc606_5 gpc388 (
      {stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462], stage0_8[463]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[65],stage1_10[103],stage1_9[147],stage1_8[193]}
   );
   gpc606_5 gpc389 (
      {stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468], stage0_8[469]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[66],stage1_10[104],stage1_9[148],stage1_8[194]}
   );
   gpc606_5 gpc390 (
      {stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474], stage0_8[475]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[67],stage1_10[105],stage1_9[149],stage1_8[195]}
   );
   gpc606_5 gpc391 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[36],stage1_11[68],stage1_10[106],stage1_9[150]}
   );
   gpc606_5 gpc392 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[37],stage1_11[69],stage1_10[107],stage1_9[151]}
   );
   gpc606_5 gpc393 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[38],stage1_11[70],stage1_10[108],stage1_9[152]}
   );
   gpc606_5 gpc394 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[39],stage1_11[71],stage1_10[109],stage1_9[153]}
   );
   gpc606_5 gpc395 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[40],stage1_11[72],stage1_10[110],stage1_9[154]}
   );
   gpc606_5 gpc396 (
      {stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[41],stage1_11[73],stage1_10[111],stage1_9[155]}
   );
   gpc606_5 gpc397 (
      {stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[42],stage1_11[74],stage1_10[112],stage1_9[156]}
   );
   gpc606_5 gpc398 (
      {stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[43],stage1_11[75],stage1_10[113],stage1_9[157]}
   );
   gpc606_5 gpc399 (
      {stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[44],stage1_11[76],stage1_10[114],stage1_9[158]}
   );
   gpc606_5 gpc400 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[45],stage1_11[77],stage1_10[115],stage1_9[159]}
   );
   gpc606_5 gpc401 (
      {stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[46],stage1_11[78],stage1_10[116],stage1_9[160]}
   );
   gpc606_5 gpc402 (
      {stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[47],stage1_11[79],stage1_10[117],stage1_9[161]}
   );
   gpc606_5 gpc403 (
      {stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[48],stage1_11[80],stage1_10[118],stage1_9[162]}
   );
   gpc606_5 gpc404 (
      {stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[49],stage1_11[81],stage1_10[119],stage1_9[163]}
   );
   gpc606_5 gpc405 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[50],stage1_11[82],stage1_10[120],stage1_9[164]}
   );
   gpc606_5 gpc406 (
      {stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[51],stage1_11[83],stage1_10[121],stage1_9[165]}
   );
   gpc606_5 gpc407 (
      {stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[52],stage1_11[84],stage1_10[122],stage1_9[166]}
   );
   gpc606_5 gpc408 (
      {stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[53],stage1_11[85],stage1_10[123],stage1_9[167]}
   );
   gpc606_5 gpc409 (
      {stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[54],stage1_11[86],stage1_10[124],stage1_9[168]}
   );
   gpc606_5 gpc410 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[55],stage1_11[87],stage1_10[125],stage1_9[169]}
   );
   gpc606_5 gpc411 (
      {stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315], stage0_9[316], stage0_9[317]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[56],stage1_11[88],stage1_10[126],stage1_9[170]}
   );
   gpc606_5 gpc412 (
      {stage0_9[318], stage0_9[319], stage0_9[320], stage0_9[321], stage0_9[322], stage0_9[323]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[57],stage1_11[89],stage1_10[127],stage1_9[171]}
   );
   gpc606_5 gpc413 (
      {stage0_9[324], stage0_9[325], stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[58],stage1_11[90],stage1_10[128],stage1_9[172]}
   );
   gpc606_5 gpc414 (
      {stage0_9[330], stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[59],stage1_11[91],stage1_10[129],stage1_9[173]}
   );
   gpc606_5 gpc415 (
      {stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340], stage0_9[341]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[60],stage1_11[92],stage1_10[130],stage1_9[174]}
   );
   gpc606_5 gpc416 (
      {stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345], stage0_9[346], stage0_9[347]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[61],stage1_11[93],stage1_10[131],stage1_9[175]}
   );
   gpc606_5 gpc417 (
      {stage0_9[348], stage0_9[349], stage0_9[350], stage0_9[351], stage0_9[352], stage0_9[353]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[62],stage1_11[94],stage1_10[132],stage1_9[176]}
   );
   gpc606_5 gpc418 (
      {stage0_9[354], stage0_9[355], stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[63],stage1_11[95],stage1_10[133],stage1_9[177]}
   );
   gpc606_5 gpc419 (
      {stage0_9[360], stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[64],stage1_11[96],stage1_10[134],stage1_9[178]}
   );
   gpc606_5 gpc420 (
      {stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370], stage0_9[371]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[65],stage1_11[97],stage1_10[135],stage1_9[179]}
   );
   gpc606_5 gpc421 (
      {stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375], stage0_9[376], stage0_9[377]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[66],stage1_11[98],stage1_10[136],stage1_9[180]}
   );
   gpc606_5 gpc422 (
      {stage0_9[378], stage0_9[379], stage0_9[380], stage0_9[381], stage0_9[382], stage0_9[383]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[67],stage1_11[99],stage1_10[137],stage1_9[181]}
   );
   gpc606_5 gpc423 (
      {stage0_9[384], stage0_9[385], stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[68],stage1_11[100],stage1_10[138],stage1_9[182]}
   );
   gpc606_5 gpc424 (
      {stage0_9[390], stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[69],stage1_11[101],stage1_10[139],stage1_9[183]}
   );
   gpc606_5 gpc425 (
      {stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400], stage0_9[401]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[70],stage1_11[102],stage1_10[140],stage1_9[184]}
   );
   gpc606_5 gpc426 (
      {stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[71],stage1_11[103],stage1_10[141],stage1_9[185]}
   );
   gpc606_5 gpc427 (
      {stage0_9[408], stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[72],stage1_11[104],stage1_10[142],stage1_9[186]}
   );
   gpc606_5 gpc428 (
      {stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[73],stage1_11[105],stage1_10[143],stage1_9[187]}
   );
   gpc606_5 gpc429 (
      {stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[74],stage1_11[106],stage1_10[144],stage1_9[188]}
   );
   gpc606_5 gpc430 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430], stage0_9[431]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[75],stage1_11[107],stage1_10[145],stage1_9[189]}
   );
   gpc606_5 gpc431 (
      {stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435], stage0_9[436], stage0_9[437]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[76],stage1_11[108],stage1_10[146],stage1_9[190]}
   );
   gpc606_5 gpc432 (
      {stage0_9[438], stage0_9[439], stage0_9[440], stage0_9[441], stage0_9[442], stage0_9[443]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[77],stage1_11[109],stage1_10[147],stage1_9[191]}
   );
   gpc606_5 gpc433 (
      {stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[78],stage1_11[110],stage1_10[148],stage1_9[192]}
   );
   gpc606_5 gpc434 (
      {stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[79],stage1_11[111],stage1_10[149],stage1_9[193]}
   );
   gpc606_5 gpc435 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460], stage0_9[461]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[80],stage1_11[112],stage1_10[150],stage1_9[194]}
   );
   gpc606_5 gpc436 (
      {stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465], stage0_9[466], stage0_9[467]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[81],stage1_11[113],stage1_10[151],stage1_9[195]}
   );
   gpc2135_5 gpc437 (
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220]},
      {stage0_11[276], stage0_11[277], stage0_11[278]},
      {stage0_12[0]},
      {stage0_13[0], stage0_13[1]},
      {stage1_14[0],stage1_13[46],stage1_12[82],stage1_11[114],stage1_10[152]}
   );
   gpc2135_5 gpc438 (
      {stage0_10[221], stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225]},
      {stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage0_12[1]},
      {stage0_13[2], stage0_13[3]},
      {stage1_14[1],stage1_13[47],stage1_12[83],stage1_11[115],stage1_10[153]}
   );
   gpc2135_5 gpc439 (
      {stage0_10[226], stage0_10[227], stage0_10[228], stage0_10[229], stage0_10[230]},
      {stage0_11[282], stage0_11[283], stage0_11[284]},
      {stage0_12[2]},
      {stage0_13[4], stage0_13[5]},
      {stage1_14[2],stage1_13[48],stage1_12[84],stage1_11[116],stage1_10[154]}
   );
   gpc2135_5 gpc440 (
      {stage0_10[231], stage0_10[232], stage0_10[233], stage0_10[234], stage0_10[235]},
      {stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage0_12[3]},
      {stage0_13[6], stage0_13[7]},
      {stage1_14[3],stage1_13[49],stage1_12[85],stage1_11[117],stage1_10[155]}
   );
   gpc606_5 gpc441 (
      {stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239], stage0_10[240], stage0_10[241]},
      {stage0_12[4], stage0_12[5], stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9]},
      {stage1_14[4],stage1_13[50],stage1_12[86],stage1_11[118],stage1_10[156]}
   );
   gpc606_5 gpc442 (
      {stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245], stage0_10[246], stage0_10[247]},
      {stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15]},
      {stage1_14[5],stage1_13[51],stage1_12[87],stage1_11[119],stage1_10[157]}
   );
   gpc606_5 gpc443 (
      {stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251], stage0_10[252], stage0_10[253]},
      {stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21]},
      {stage1_14[6],stage1_13[52],stage1_12[88],stage1_11[120],stage1_10[158]}
   );
   gpc606_5 gpc444 (
      {stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257], stage0_10[258], stage0_10[259]},
      {stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27]},
      {stage1_14[7],stage1_13[53],stage1_12[89],stage1_11[121],stage1_10[159]}
   );
   gpc606_5 gpc445 (
      {stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263], stage0_10[264], stage0_10[265]},
      {stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33]},
      {stage1_14[8],stage1_13[54],stage1_12[90],stage1_11[122],stage1_10[160]}
   );
   gpc606_5 gpc446 (
      {stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269], stage0_10[270], stage0_10[271]},
      {stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39]},
      {stage1_14[9],stage1_13[55],stage1_12[91],stage1_11[123],stage1_10[161]}
   );
   gpc606_5 gpc447 (
      {stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275], stage0_10[276], stage0_10[277]},
      {stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45]},
      {stage1_14[10],stage1_13[56],stage1_12[92],stage1_11[124],stage1_10[162]}
   );
   gpc606_5 gpc448 (
      {stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281], stage0_10[282], stage0_10[283]},
      {stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51]},
      {stage1_14[11],stage1_13[57],stage1_12[93],stage1_11[125],stage1_10[163]}
   );
   gpc606_5 gpc449 (
      {stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287], stage0_10[288], stage0_10[289]},
      {stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57]},
      {stage1_14[12],stage1_13[58],stage1_12[94],stage1_11[126],stage1_10[164]}
   );
   gpc606_5 gpc450 (
      {stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293], stage0_10[294], stage0_10[295]},
      {stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63]},
      {stage1_14[13],stage1_13[59],stage1_12[95],stage1_11[127],stage1_10[165]}
   );
   gpc606_5 gpc451 (
      {stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299], stage0_10[300], stage0_10[301]},
      {stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69]},
      {stage1_14[14],stage1_13[60],stage1_12[96],stage1_11[128],stage1_10[166]}
   );
   gpc606_5 gpc452 (
      {stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305], stage0_10[306], stage0_10[307]},
      {stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75]},
      {stage1_14[15],stage1_13[61],stage1_12[97],stage1_11[129],stage1_10[167]}
   );
   gpc606_5 gpc453 (
      {stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311], stage0_10[312], stage0_10[313]},
      {stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81]},
      {stage1_14[16],stage1_13[62],stage1_12[98],stage1_11[130],stage1_10[168]}
   );
   gpc615_5 gpc454 (
      {stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317], stage0_10[318]},
      {stage0_11[288]},
      {stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87]},
      {stage1_14[17],stage1_13[63],stage1_12[99],stage1_11[131],stage1_10[169]}
   );
   gpc615_5 gpc455 (
      {stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage0_11[289]},
      {stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93]},
      {stage1_14[18],stage1_13[64],stage1_12[100],stage1_11[132],stage1_10[170]}
   );
   gpc615_5 gpc456 (
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328]},
      {stage0_11[290]},
      {stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99]},
      {stage1_14[19],stage1_13[65],stage1_12[101],stage1_11[133],stage1_10[171]}
   );
   gpc615_5 gpc457 (
      {stage0_10[329], stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333]},
      {stage0_11[291]},
      {stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105]},
      {stage1_14[20],stage1_13[66],stage1_12[102],stage1_11[134],stage1_10[172]}
   );
   gpc615_5 gpc458 (
      {stage0_10[334], stage0_10[335], stage0_10[336], stage0_10[337], stage0_10[338]},
      {stage0_11[292]},
      {stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111]},
      {stage1_14[21],stage1_13[67],stage1_12[103],stage1_11[135],stage1_10[173]}
   );
   gpc615_5 gpc459 (
      {stage0_10[339], stage0_10[340], stage0_10[341], stage0_10[342], stage0_10[343]},
      {stage0_11[293]},
      {stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117]},
      {stage1_14[22],stage1_13[68],stage1_12[104],stage1_11[136],stage1_10[174]}
   );
   gpc615_5 gpc460 (
      {stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347], stage0_10[348]},
      {stage0_11[294]},
      {stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123]},
      {stage1_14[23],stage1_13[69],stage1_12[105],stage1_11[137],stage1_10[175]}
   );
   gpc615_5 gpc461 (
      {stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage0_11[295]},
      {stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129]},
      {stage1_14[24],stage1_13[70],stage1_12[106],stage1_11[138],stage1_10[176]}
   );
   gpc615_5 gpc462 (
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358]},
      {stage0_11[296]},
      {stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135]},
      {stage1_14[25],stage1_13[71],stage1_12[107],stage1_11[139],stage1_10[177]}
   );
   gpc615_5 gpc463 (
      {stage0_10[359], stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363]},
      {stage0_11[297]},
      {stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141]},
      {stage1_14[26],stage1_13[72],stage1_12[108],stage1_11[140],stage1_10[178]}
   );
   gpc615_5 gpc464 (
      {stage0_10[364], stage0_10[365], stage0_10[366], stage0_10[367], stage0_10[368]},
      {stage0_11[298]},
      {stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147]},
      {stage1_14[27],stage1_13[73],stage1_12[109],stage1_11[141],stage1_10[179]}
   );
   gpc615_5 gpc465 (
      {stage0_10[369], stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373]},
      {stage0_11[299]},
      {stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153]},
      {stage1_14[28],stage1_13[74],stage1_12[110],stage1_11[142],stage1_10[180]}
   );
   gpc615_5 gpc466 (
      {stage0_10[374], stage0_10[375], stage0_10[376], stage0_10[377], stage0_10[378]},
      {stage0_11[300]},
      {stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159]},
      {stage1_14[29],stage1_13[75],stage1_12[111],stage1_11[143],stage1_10[181]}
   );
   gpc615_5 gpc467 (
      {stage0_10[379], stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383]},
      {stage0_11[301]},
      {stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165]},
      {stage1_14[30],stage1_13[76],stage1_12[112],stage1_11[144],stage1_10[182]}
   );
   gpc615_5 gpc468 (
      {stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305], stage0_11[306]},
      {stage0_12[166]},
      {stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12], stage0_13[13]},
      {stage1_15[0],stage1_14[31],stage1_13[77],stage1_12[113],stage1_11[145]}
   );
   gpc615_5 gpc469 (
      {stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage0_12[167]},
      {stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18], stage0_13[19]},
      {stage1_15[1],stage1_14[32],stage1_13[78],stage1_12[114],stage1_11[146]}
   );
   gpc615_5 gpc470 (
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316]},
      {stage0_12[168]},
      {stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23], stage0_13[24], stage0_13[25]},
      {stage1_15[2],stage1_14[33],stage1_13[79],stage1_12[115],stage1_11[147]}
   );
   gpc615_5 gpc471 (
      {stage0_11[317], stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321]},
      {stage0_12[169]},
      {stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30], stage0_13[31]},
      {stage1_15[3],stage1_14[34],stage1_13[80],stage1_12[116],stage1_11[148]}
   );
   gpc615_5 gpc472 (
      {stage0_11[322], stage0_11[323], stage0_11[324], stage0_11[325], stage0_11[326]},
      {stage0_12[170]},
      {stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35], stage0_13[36], stage0_13[37]},
      {stage1_15[4],stage1_14[35],stage1_13[81],stage1_12[117],stage1_11[149]}
   );
   gpc615_5 gpc473 (
      {stage0_11[327], stage0_11[328], stage0_11[329], stage0_11[330], stage0_11[331]},
      {stage0_12[171]},
      {stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41], stage0_13[42], stage0_13[43]},
      {stage1_15[5],stage1_14[36],stage1_13[82],stage1_12[118],stage1_11[150]}
   );
   gpc615_5 gpc474 (
      {stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335], stage0_11[336]},
      {stage0_12[172]},
      {stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47], stage0_13[48], stage0_13[49]},
      {stage1_15[6],stage1_14[37],stage1_13[83],stage1_12[119],stage1_11[151]}
   );
   gpc615_5 gpc475 (
      {stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage0_12[173]},
      {stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55]},
      {stage1_15[7],stage1_14[38],stage1_13[84],stage1_12[120],stage1_11[152]}
   );
   gpc615_5 gpc476 (
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346]},
      {stage0_12[174]},
      {stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage1_15[8],stage1_14[39],stage1_13[85],stage1_12[121],stage1_11[153]}
   );
   gpc615_5 gpc477 (
      {stage0_11[347], stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351]},
      {stage0_12[175]},
      {stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67]},
      {stage1_15[9],stage1_14[40],stage1_13[86],stage1_12[122],stage1_11[154]}
   );
   gpc615_5 gpc478 (
      {stage0_11[352], stage0_11[353], stage0_11[354], stage0_11[355], stage0_11[356]},
      {stage0_12[176]},
      {stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73]},
      {stage1_15[10],stage1_14[41],stage1_13[87],stage1_12[123],stage1_11[155]}
   );
   gpc615_5 gpc479 (
      {stage0_11[357], stage0_11[358], stage0_11[359], stage0_11[360], stage0_11[361]},
      {stage0_12[177]},
      {stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77], stage0_13[78], stage0_13[79]},
      {stage1_15[11],stage1_14[42],stage1_13[88],stage1_12[124],stage1_11[156]}
   );
   gpc615_5 gpc480 (
      {stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365], stage0_11[366]},
      {stage0_12[178]},
      {stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85]},
      {stage1_15[12],stage1_14[43],stage1_13[89],stage1_12[125],stage1_11[157]}
   );
   gpc615_5 gpc481 (
      {stage0_12[179], stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183]},
      {stage0_13[86]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[13],stage1_14[44],stage1_13[90],stage1_12[126]}
   );
   gpc615_5 gpc482 (
      {stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188]},
      {stage0_13[87]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[14],stage1_14[45],stage1_13[91],stage1_12[127]}
   );
   gpc615_5 gpc483 (
      {stage0_12[189], stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193]},
      {stage0_13[88]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[15],stage1_14[46],stage1_13[92],stage1_12[128]}
   );
   gpc615_5 gpc484 (
      {stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198]},
      {stage0_13[89]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[16],stage1_14[47],stage1_13[93],stage1_12[129]}
   );
   gpc615_5 gpc485 (
      {stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage0_13[90]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[17],stage1_14[48],stage1_13[94],stage1_12[130]}
   );
   gpc615_5 gpc486 (
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208]},
      {stage0_13[91]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[18],stage1_14[49],stage1_13[95],stage1_12[131]}
   );
   gpc615_5 gpc487 (
      {stage0_12[209], stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213]},
      {stage0_13[92]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[19],stage1_14[50],stage1_13[96],stage1_12[132]}
   );
   gpc615_5 gpc488 (
      {stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218]},
      {stage0_13[93]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[20],stage1_14[51],stage1_13[97],stage1_12[133]}
   );
   gpc615_5 gpc489 (
      {stage0_12[219], stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223]},
      {stage0_13[94]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[21],stage1_14[52],stage1_13[98],stage1_12[134]}
   );
   gpc615_5 gpc490 (
      {stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227], stage0_12[228]},
      {stage0_13[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[22],stage1_14[53],stage1_13[99],stage1_12[135]}
   );
   gpc615_5 gpc491 (
      {stage0_12[229], stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233]},
      {stage0_13[96]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[23],stage1_14[54],stage1_13[100],stage1_12[136]}
   );
   gpc615_5 gpc492 (
      {stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238]},
      {stage0_13[97]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[24],stage1_14[55],stage1_13[101],stage1_12[137]}
   );
   gpc615_5 gpc493 (
      {stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243]},
      {stage0_13[98]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[25],stage1_14[56],stage1_13[102],stage1_12[138]}
   );
   gpc615_5 gpc494 (
      {stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248]},
      {stage0_13[99]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[26],stage1_14[57],stage1_13[103],stage1_12[139]}
   );
   gpc615_5 gpc495 (
      {stage0_12[249], stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253]},
      {stage0_13[100]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[27],stage1_14[58],stage1_13[104],stage1_12[140]}
   );
   gpc615_5 gpc496 (
      {stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257], stage0_12[258]},
      {stage0_13[101]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[28],stage1_14[59],stage1_13[105],stage1_12[141]}
   );
   gpc615_5 gpc497 (
      {stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263]},
      {stage0_13[102]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[29],stage1_14[60],stage1_13[106],stage1_12[142]}
   );
   gpc615_5 gpc498 (
      {stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268]},
      {stage0_13[103]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[30],stage1_14[61],stage1_13[107],stage1_12[143]}
   );
   gpc615_5 gpc499 (
      {stage0_12[269], stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273]},
      {stage0_13[104]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[31],stage1_14[62],stage1_13[108],stage1_12[144]}
   );
   gpc615_5 gpc500 (
      {stage0_12[274], stage0_12[275], stage0_12[276], stage0_12[277], stage0_12[278]},
      {stage0_13[105]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[32],stage1_14[63],stage1_13[109],stage1_12[145]}
   );
   gpc615_5 gpc501 (
      {stage0_12[279], stage0_12[280], stage0_12[281], stage0_12[282], stage0_12[283]},
      {stage0_13[106]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[33],stage1_14[64],stage1_13[110],stage1_12[146]}
   );
   gpc615_5 gpc502 (
      {stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287], stage0_12[288]},
      {stage0_13[107]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[34],stage1_14[65],stage1_13[111],stage1_12[147]}
   );
   gpc615_5 gpc503 (
      {stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293]},
      {stage0_13[108]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[35],stage1_14[66],stage1_13[112],stage1_12[148]}
   );
   gpc615_5 gpc504 (
      {stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298]},
      {stage0_13[109]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[36],stage1_14[67],stage1_13[113],stage1_12[149]}
   );
   gpc615_5 gpc505 (
      {stage0_12[299], stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303]},
      {stage0_13[110]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[37],stage1_14[68],stage1_13[114],stage1_12[150]}
   );
   gpc615_5 gpc506 (
      {stage0_12[304], stage0_12[305], stage0_12[306], stage0_12[307], stage0_12[308]},
      {stage0_13[111]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[38],stage1_14[69],stage1_13[115],stage1_12[151]}
   );
   gpc615_5 gpc507 (
      {stage0_12[309], stage0_12[310], stage0_12[311], stage0_12[312], stage0_12[313]},
      {stage0_13[112]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[39],stage1_14[70],stage1_13[116],stage1_12[152]}
   );
   gpc615_5 gpc508 (
      {stage0_12[314], stage0_12[315], stage0_12[316], stage0_12[317], stage0_12[318]},
      {stage0_13[113]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[40],stage1_14[71],stage1_13[117],stage1_12[153]}
   );
   gpc615_5 gpc509 (
      {stage0_12[319], stage0_12[320], stage0_12[321], stage0_12[322], stage0_12[323]},
      {stage0_13[114]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[41],stage1_14[72],stage1_13[118],stage1_12[154]}
   );
   gpc615_5 gpc510 (
      {stage0_12[324], stage0_12[325], stage0_12[326], stage0_12[327], stage0_12[328]},
      {stage0_13[115]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[42],stage1_14[73],stage1_13[119],stage1_12[155]}
   );
   gpc615_5 gpc511 (
      {stage0_12[329], stage0_12[330], stage0_12[331], stage0_12[332], stage0_12[333]},
      {stage0_13[116]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[43],stage1_14[74],stage1_13[120],stage1_12[156]}
   );
   gpc615_5 gpc512 (
      {stage0_12[334], stage0_12[335], stage0_12[336], stage0_12[337], stage0_12[338]},
      {stage0_13[117]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[44],stage1_14[75],stage1_13[121],stage1_12[157]}
   );
   gpc615_5 gpc513 (
      {stage0_12[339], stage0_12[340], stage0_12[341], stage0_12[342], stage0_12[343]},
      {stage0_13[118]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[45],stage1_14[76],stage1_13[122],stage1_12[158]}
   );
   gpc615_5 gpc514 (
      {stage0_12[344], stage0_12[345], stage0_12[346], stage0_12[347], stage0_12[348]},
      {stage0_13[119]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[46],stage1_14[77],stage1_13[123],stage1_12[159]}
   );
   gpc615_5 gpc515 (
      {stage0_12[349], stage0_12[350], stage0_12[351], stage0_12[352], stage0_12[353]},
      {stage0_13[120]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[47],stage1_14[78],stage1_13[124],stage1_12[160]}
   );
   gpc615_5 gpc516 (
      {stage0_12[354], stage0_12[355], stage0_12[356], stage0_12[357], stage0_12[358]},
      {stage0_13[121]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[48],stage1_14[79],stage1_13[125],stage1_12[161]}
   );
   gpc615_5 gpc517 (
      {stage0_12[359], stage0_12[360], stage0_12[361], stage0_12[362], stage0_12[363]},
      {stage0_13[122]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[49],stage1_14[80],stage1_13[126],stage1_12[162]}
   );
   gpc615_5 gpc518 (
      {stage0_12[364], stage0_12[365], stage0_12[366], stage0_12[367], stage0_12[368]},
      {stage0_13[123]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[50],stage1_14[81],stage1_13[127],stage1_12[163]}
   );
   gpc615_5 gpc519 (
      {stage0_12[369], stage0_12[370], stage0_12[371], stage0_12[372], stage0_12[373]},
      {stage0_13[124]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[51],stage1_14[82],stage1_13[128],stage1_12[164]}
   );
   gpc615_5 gpc520 (
      {stage0_12[374], stage0_12[375], stage0_12[376], stage0_12[377], stage0_12[378]},
      {stage0_13[125]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[52],stage1_14[83],stage1_13[129],stage1_12[165]}
   );
   gpc615_5 gpc521 (
      {stage0_12[379], stage0_12[380], stage0_12[381], stage0_12[382], stage0_12[383]},
      {stage0_13[126]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[53],stage1_14[84],stage1_13[130],stage1_12[166]}
   );
   gpc615_5 gpc522 (
      {stage0_12[384], stage0_12[385], stage0_12[386], stage0_12[387], stage0_12[388]},
      {stage0_13[127]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[54],stage1_14[85],stage1_13[131],stage1_12[167]}
   );
   gpc615_5 gpc523 (
      {stage0_12[389], stage0_12[390], stage0_12[391], stage0_12[392], stage0_12[393]},
      {stage0_13[128]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[55],stage1_14[86],stage1_13[132],stage1_12[168]}
   );
   gpc615_5 gpc524 (
      {stage0_12[394], stage0_12[395], stage0_12[396], stage0_12[397], stage0_12[398]},
      {stage0_13[129]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[56],stage1_14[87],stage1_13[133],stage1_12[169]}
   );
   gpc615_5 gpc525 (
      {stage0_12[399], stage0_12[400], stage0_12[401], stage0_12[402], stage0_12[403]},
      {stage0_13[130]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[57],stage1_14[88],stage1_13[134],stage1_12[170]}
   );
   gpc615_5 gpc526 (
      {stage0_12[404], stage0_12[405], stage0_12[406], stage0_12[407], stage0_12[408]},
      {stage0_13[131]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[58],stage1_14[89],stage1_13[135],stage1_12[171]}
   );
   gpc615_5 gpc527 (
      {stage0_12[409], stage0_12[410], stage0_12[411], stage0_12[412], stage0_12[413]},
      {stage0_13[132]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[59],stage1_14[90],stage1_13[136],stage1_12[172]}
   );
   gpc615_5 gpc528 (
      {stage0_12[414], stage0_12[415], stage0_12[416], stage0_12[417], stage0_12[418]},
      {stage0_13[133]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[60],stage1_14[91],stage1_13[137],stage1_12[173]}
   );
   gpc615_5 gpc529 (
      {stage0_12[419], stage0_12[420], stage0_12[421], stage0_12[422], stage0_12[423]},
      {stage0_13[134]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[61],stage1_14[92],stage1_13[138],stage1_12[174]}
   );
   gpc615_5 gpc530 (
      {stage0_12[424], stage0_12[425], stage0_12[426], stage0_12[427], stage0_12[428]},
      {stage0_13[135]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[62],stage1_14[93],stage1_13[139],stage1_12[175]}
   );
   gpc615_5 gpc531 (
      {stage0_12[429], stage0_12[430], stage0_12[431], stage0_12[432], stage0_12[433]},
      {stage0_13[136]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[63],stage1_14[94],stage1_13[140],stage1_12[176]}
   );
   gpc615_5 gpc532 (
      {stage0_12[434], stage0_12[435], stage0_12[436], stage0_12[437], stage0_12[438]},
      {stage0_13[137]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[64],stage1_14[95],stage1_13[141],stage1_12[177]}
   );
   gpc615_5 gpc533 (
      {stage0_12[439], stage0_12[440], stage0_12[441], stage0_12[442], stage0_12[443]},
      {stage0_13[138]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[65],stage1_14[96],stage1_13[142],stage1_12[178]}
   );
   gpc615_5 gpc534 (
      {stage0_12[444], stage0_12[445], stage0_12[446], stage0_12[447], stage0_12[448]},
      {stage0_13[139]},
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage1_16[53],stage1_15[66],stage1_14[97],stage1_13[143],stage1_12[179]}
   );
   gpc615_5 gpc535 (
      {stage0_12[449], stage0_12[450], stage0_12[451], stage0_12[452], stage0_12[453]},
      {stage0_13[140]},
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage1_16[54],stage1_15[67],stage1_14[98],stage1_13[144],stage1_12[180]}
   );
   gpc615_5 gpc536 (
      {stage0_12[454], stage0_12[455], stage0_12[456], stage0_12[457], stage0_12[458]},
      {stage0_13[141]},
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage1_16[55],stage1_15[68],stage1_14[99],stage1_13[145],stage1_12[181]}
   );
   gpc615_5 gpc537 (
      {stage0_12[459], stage0_12[460], stage0_12[461], stage0_12[462], stage0_12[463]},
      {stage0_13[142]},
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage1_16[56],stage1_15[69],stage1_14[100],stage1_13[146],stage1_12[182]}
   );
   gpc615_5 gpc538 (
      {stage0_12[464], stage0_12[465], stage0_12[466], stage0_12[467], stage0_12[468]},
      {stage0_13[143]},
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage1_16[57],stage1_15[70],stage1_14[101],stage1_13[147],stage1_12[183]}
   );
   gpc615_5 gpc539 (
      {stage0_12[469], stage0_12[470], stage0_12[471], stage0_12[472], stage0_12[473]},
      {stage0_13[144]},
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage1_16[58],stage1_15[71],stage1_14[102],stage1_13[148],stage1_12[184]}
   );
   gpc615_5 gpc540 (
      {stage0_12[474], stage0_12[475], stage0_12[476], stage0_12[477], stage0_12[478]},
      {stage0_13[145]},
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage1_16[59],stage1_15[72],stage1_14[103],stage1_13[149],stage1_12[185]}
   );
   gpc615_5 gpc541 (
      {stage0_12[479], stage0_12[480], stage0_12[481], stage0_12[482], stage0_12[483]},
      {stage0_13[146]},
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage1_16[60],stage1_15[73],stage1_14[104],stage1_13[150],stage1_12[186]}
   );
   gpc606_5 gpc542 (
      {stage0_13[147], stage0_13[148], stage0_13[149], stage0_13[150], stage0_13[151], stage0_13[152]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[61],stage1_15[74],stage1_14[105],stage1_13[151]}
   );
   gpc606_5 gpc543 (
      {stage0_13[153], stage0_13[154], stage0_13[155], stage0_13[156], stage0_13[157], stage0_13[158]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[62],stage1_15[75],stage1_14[106],stage1_13[152]}
   );
   gpc606_5 gpc544 (
      {stage0_13[159], stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[63],stage1_15[76],stage1_14[107],stage1_13[153]}
   );
   gpc606_5 gpc545 (
      {stage0_13[165], stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[64],stage1_15[77],stage1_14[108],stage1_13[154]}
   );
   gpc606_5 gpc546 (
      {stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175], stage0_13[176]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[65],stage1_15[78],stage1_14[109],stage1_13[155]}
   );
   gpc606_5 gpc547 (
      {stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181], stage0_13[182]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[66],stage1_15[79],stage1_14[110],stage1_13[156]}
   );
   gpc606_5 gpc548 (
      {stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[67],stage1_15[80],stage1_14[111],stage1_13[157]}
   );
   gpc606_5 gpc549 (
      {stage0_13[189], stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[68],stage1_15[81],stage1_14[112],stage1_13[158]}
   );
   gpc606_5 gpc550 (
      {stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[69],stage1_15[82],stage1_14[113],stage1_13[159]}
   );
   gpc615_5 gpc551 (
      {stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205]},
      {stage0_14[366]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[70],stage1_15[83],stage1_14[114],stage1_13[160]}
   );
   gpc615_5 gpc552 (
      {stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210]},
      {stage0_14[367]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[71],stage1_15[84],stage1_14[115],stage1_13[161]}
   );
   gpc615_5 gpc553 (
      {stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage0_14[368]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[72],stage1_15[85],stage1_14[116],stage1_13[162]}
   );
   gpc615_5 gpc554 (
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220]},
      {stage0_14[369]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[73],stage1_15[86],stage1_14[117],stage1_13[163]}
   );
   gpc615_5 gpc555 (
      {stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225]},
      {stage0_14[370]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[74],stage1_15[87],stage1_14[118],stage1_13[164]}
   );
   gpc615_5 gpc556 (
      {stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_14[371]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[75],stage1_15[88],stage1_14[119],stage1_13[165]}
   );
   gpc615_5 gpc557 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_14[372]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[76],stage1_15[89],stage1_14[120],stage1_13[166]}
   );
   gpc615_5 gpc558 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240]},
      {stage0_14[373]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[77],stage1_15[90],stage1_14[121],stage1_13[167]}
   );
   gpc615_5 gpc559 (
      {stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_14[374]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[78],stage1_15[91],stage1_14[122],stage1_13[168]}
   );
   gpc615_5 gpc560 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250]},
      {stage0_14[375]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[79],stage1_15[92],stage1_14[123],stage1_13[169]}
   );
   gpc615_5 gpc561 (
      {stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255]},
      {stage0_14[376]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[80],stage1_15[93],stage1_14[124],stage1_13[170]}
   );
   gpc615_5 gpc562 (
      {stage0_13[256], stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260]},
      {stage0_14[377]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[81],stage1_15[94],stage1_14[125],stage1_13[171]}
   );
   gpc615_5 gpc563 (
      {stage0_13[261], stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265]},
      {stage0_14[378]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[82],stage1_15[95],stage1_14[126],stage1_13[172]}
   );
   gpc615_5 gpc564 (
      {stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270]},
      {stage0_14[379]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[83],stage1_15[96],stage1_14[127],stage1_13[173]}
   );
   gpc615_5 gpc565 (
      {stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage0_14[380]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[84],stage1_15[97],stage1_14[128],stage1_13[174]}
   );
   gpc615_5 gpc566 (
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280]},
      {stage0_14[381]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[85],stage1_15[98],stage1_14[129],stage1_13[175]}
   );
   gpc615_5 gpc567 (
      {stage0_13[281], stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285]},
      {stage0_14[382]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[86],stage1_15[99],stage1_14[130],stage1_13[176]}
   );
   gpc615_5 gpc568 (
      {stage0_13[286], stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290]},
      {stage0_14[383]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[87],stage1_15[100],stage1_14[131],stage1_13[177]}
   );
   gpc615_5 gpc569 (
      {stage0_13[291], stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295]},
      {stage0_14[384]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[88],stage1_15[101],stage1_14[132],stage1_13[178]}
   );
   gpc615_5 gpc570 (
      {stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300]},
      {stage0_14[385]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[89],stage1_15[102],stage1_14[133],stage1_13[179]}
   );
   gpc615_5 gpc571 (
      {stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_14[386]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[90],stage1_15[103],stage1_14[134],stage1_13[180]}
   );
   gpc615_5 gpc572 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310]},
      {stage0_14[387]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[91],stage1_15[104],stage1_14[135],stage1_13[181]}
   );
   gpc615_5 gpc573 (
      {stage0_13[311], stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315]},
      {stage0_14[388]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[92],stage1_15[105],stage1_14[136],stage1_13[182]}
   );
   gpc615_5 gpc574 (
      {stage0_13[316], stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320]},
      {stage0_14[389]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[93],stage1_15[106],stage1_14[137],stage1_13[183]}
   );
   gpc615_5 gpc575 (
      {stage0_13[321], stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325]},
      {stage0_14[390]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[94],stage1_15[107],stage1_14[138],stage1_13[184]}
   );
   gpc615_5 gpc576 (
      {stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330]},
      {stage0_14[391]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[95],stage1_15[108],stage1_14[139],stage1_13[185]}
   );
   gpc615_5 gpc577 (
      {stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_14[392]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[96],stage1_15[109],stage1_14[140],stage1_13[186]}
   );
   gpc615_5 gpc578 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340]},
      {stage0_14[393]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[97],stage1_15[110],stage1_14[141],stage1_13[187]}
   );
   gpc615_5 gpc579 (
      {stage0_13[341], stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345]},
      {stage0_14[394]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[98],stage1_15[111],stage1_14[142],stage1_13[188]}
   );
   gpc615_5 gpc580 (
      {stage0_13[346], stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350]},
      {stage0_14[395]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[99],stage1_15[112],stage1_14[143],stage1_13[189]}
   );
   gpc615_5 gpc581 (
      {stage0_13[351], stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355]},
      {stage0_14[396]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[100],stage1_15[113],stage1_14[144],stage1_13[190]}
   );
   gpc615_5 gpc582 (
      {stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360]},
      {stage0_14[397]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[101],stage1_15[114],stage1_14[145],stage1_13[191]}
   );
   gpc615_5 gpc583 (
      {stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_14[398]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[102],stage1_15[115],stage1_14[146],stage1_13[192]}
   );
   gpc615_5 gpc584 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370]},
      {stage0_14[399]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[103],stage1_15[116],stage1_14[147],stage1_13[193]}
   );
   gpc615_5 gpc585 (
      {stage0_13[371], stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375]},
      {stage0_14[400]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[104],stage1_15[117],stage1_14[148],stage1_13[194]}
   );
   gpc606_5 gpc586 (
      {stage0_14[401], stage0_14[402], stage0_14[403], stage0_14[404], stage0_14[405], stage0_14[406]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[44],stage1_16[105],stage1_15[118],stage1_14[149]}
   );
   gpc606_5 gpc587 (
      {stage0_14[407], stage0_14[408], stage0_14[409], stage0_14[410], stage0_14[411], stage0_14[412]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[45],stage1_16[106],stage1_15[119],stage1_14[150]}
   );
   gpc606_5 gpc588 (
      {stage0_14[413], stage0_14[414], stage0_14[415], stage0_14[416], stage0_14[417], stage0_14[418]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[46],stage1_16[107],stage1_15[120],stage1_14[151]}
   );
   gpc615_5 gpc589 (
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268]},
      {stage0_16[18]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[3],stage1_17[47],stage1_16[108],stage1_15[121]}
   );
   gpc615_5 gpc590 (
      {stage0_15[269], stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273]},
      {stage0_16[19]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[4],stage1_17[48],stage1_16[109],stage1_15[122]}
   );
   gpc615_5 gpc591 (
      {stage0_15[274], stage0_15[275], stage0_15[276], stage0_15[277], stage0_15[278]},
      {stage0_16[20]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[5],stage1_17[49],stage1_16[110],stage1_15[123]}
   );
   gpc615_5 gpc592 (
      {stage0_15[279], stage0_15[280], stage0_15[281], stage0_15[282], stage0_15[283]},
      {stage0_16[21]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[6],stage1_17[50],stage1_16[111],stage1_15[124]}
   );
   gpc615_5 gpc593 (
      {stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287], stage0_15[288]},
      {stage0_16[22]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[7],stage1_17[51],stage1_16[112],stage1_15[125]}
   );
   gpc615_5 gpc594 (
      {stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage0_16[23]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[8],stage1_17[52],stage1_16[113],stage1_15[126]}
   );
   gpc615_5 gpc595 (
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298]},
      {stage0_16[24]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[9],stage1_17[53],stage1_16[114],stage1_15[127]}
   );
   gpc615_5 gpc596 (
      {stage0_15[299], stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303]},
      {stage0_16[25]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[10],stage1_17[54],stage1_16[115],stage1_15[128]}
   );
   gpc615_5 gpc597 (
      {stage0_15[304], stage0_15[305], stage0_15[306], stage0_15[307], stage0_15[308]},
      {stage0_16[26]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[11],stage1_17[55],stage1_16[116],stage1_15[129]}
   );
   gpc615_5 gpc598 (
      {stage0_15[309], stage0_15[310], stage0_15[311], stage0_15[312], stage0_15[313]},
      {stage0_16[27]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[12],stage1_17[56],stage1_16[117],stage1_15[130]}
   );
   gpc615_5 gpc599 (
      {stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317], stage0_15[318]},
      {stage0_16[28]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[13],stage1_17[57],stage1_16[118],stage1_15[131]}
   );
   gpc615_5 gpc600 (
      {stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage0_16[29]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[14],stage1_17[58],stage1_16[119],stage1_15[132]}
   );
   gpc615_5 gpc601 (
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328]},
      {stage0_16[30]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[15],stage1_17[59],stage1_16[120],stage1_15[133]}
   );
   gpc615_5 gpc602 (
      {stage0_15[329], stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333]},
      {stage0_16[31]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[16],stage1_17[60],stage1_16[121],stage1_15[134]}
   );
   gpc615_5 gpc603 (
      {stage0_15[334], stage0_15[335], stage0_15[336], stage0_15[337], stage0_15[338]},
      {stage0_16[32]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[17],stage1_17[61],stage1_16[122],stage1_15[135]}
   );
   gpc615_5 gpc604 (
      {stage0_15[339], stage0_15[340], stage0_15[341], stage0_15[342], stage0_15[343]},
      {stage0_16[33]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[18],stage1_17[62],stage1_16[123],stage1_15[136]}
   );
   gpc615_5 gpc605 (
      {stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347], stage0_15[348]},
      {stage0_16[34]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[19],stage1_17[63],stage1_16[124],stage1_15[137]}
   );
   gpc615_5 gpc606 (
      {stage0_15[349], stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353]},
      {stage0_16[35]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[20],stage1_17[64],stage1_16[125],stage1_15[138]}
   );
   gpc615_5 gpc607 (
      {stage0_15[354], stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358]},
      {stage0_16[36]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[21],stage1_17[65],stage1_16[126],stage1_15[139]}
   );
   gpc615_5 gpc608 (
      {stage0_15[359], stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363]},
      {stage0_16[37]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[22],stage1_17[66],stage1_16[127],stage1_15[140]}
   );
   gpc615_5 gpc609 (
      {stage0_15[364], stage0_15[365], stage0_15[366], stage0_15[367], stage0_15[368]},
      {stage0_16[38]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[23],stage1_17[67],stage1_16[128],stage1_15[141]}
   );
   gpc615_5 gpc610 (
      {stage0_15[369], stage0_15[370], stage0_15[371], stage0_15[372], stage0_15[373]},
      {stage0_16[39]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[24],stage1_17[68],stage1_16[129],stage1_15[142]}
   );
   gpc615_5 gpc611 (
      {stage0_15[374], stage0_15[375], stage0_15[376], stage0_15[377], stage0_15[378]},
      {stage0_16[40]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[25],stage1_17[69],stage1_16[130],stage1_15[143]}
   );
   gpc615_5 gpc612 (
      {stage0_15[379], stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383]},
      {stage0_16[41]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[26],stage1_17[70],stage1_16[131],stage1_15[144]}
   );
   gpc615_5 gpc613 (
      {stage0_15[384], stage0_15[385], stage0_15[386], stage0_15[387], stage0_15[388]},
      {stage0_16[42]},
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage1_19[24],stage1_18[27],stage1_17[71],stage1_16[132],stage1_15[145]}
   );
   gpc615_5 gpc614 (
      {stage0_15[389], stage0_15[390], stage0_15[391], stage0_15[392], stage0_15[393]},
      {stage0_16[43]},
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage1_19[25],stage1_18[28],stage1_17[72],stage1_16[133],stage1_15[146]}
   );
   gpc615_5 gpc615 (
      {stage0_15[394], stage0_15[395], stage0_15[396], stage0_15[397], stage0_15[398]},
      {stage0_16[44]},
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage1_19[26],stage1_18[29],stage1_17[73],stage1_16[134],stage1_15[147]}
   );
   gpc615_5 gpc616 (
      {stage0_15[399], stage0_15[400], stage0_15[401], stage0_15[402], stage0_15[403]},
      {stage0_16[45]},
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage1_19[27],stage1_18[30],stage1_17[74],stage1_16[135],stage1_15[148]}
   );
   gpc615_5 gpc617 (
      {stage0_15[404], stage0_15[405], stage0_15[406], stage0_15[407], stage0_15[408]},
      {stage0_16[46]},
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage1_19[28],stage1_18[31],stage1_17[75],stage1_16[136],stage1_15[149]}
   );
   gpc615_5 gpc618 (
      {stage0_15[409], stage0_15[410], stage0_15[411], stage0_15[412], stage0_15[413]},
      {stage0_16[47]},
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage1_19[29],stage1_18[32],stage1_17[76],stage1_16[137],stage1_15[150]}
   );
   gpc615_5 gpc619 (
      {stage0_15[414], stage0_15[415], stage0_15[416], stage0_15[417], stage0_15[418]},
      {stage0_16[48]},
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage1_19[30],stage1_18[33],stage1_17[77],stage1_16[138],stage1_15[151]}
   );
   gpc615_5 gpc620 (
      {stage0_15[419], stage0_15[420], stage0_15[421], stage0_15[422], stage0_15[423]},
      {stage0_16[49]},
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage1_19[31],stage1_18[34],stage1_17[78],stage1_16[139],stage1_15[152]}
   );
   gpc615_5 gpc621 (
      {stage0_15[424], stage0_15[425], stage0_15[426], stage0_15[427], stage0_15[428]},
      {stage0_16[50]},
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage1_19[32],stage1_18[35],stage1_17[79],stage1_16[140],stage1_15[153]}
   );
   gpc615_5 gpc622 (
      {stage0_15[429], stage0_15[430], stage0_15[431], stage0_15[432], stage0_15[433]},
      {stage0_16[51]},
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage1_19[33],stage1_18[36],stage1_17[80],stage1_16[141],stage1_15[154]}
   );
   gpc615_5 gpc623 (
      {stage0_15[434], stage0_15[435], stage0_15[436], stage0_15[437], stage0_15[438]},
      {stage0_16[52]},
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage1_19[34],stage1_18[37],stage1_17[81],stage1_16[142],stage1_15[155]}
   );
   gpc615_5 gpc624 (
      {stage0_15[439], stage0_15[440], stage0_15[441], stage0_15[442], stage0_15[443]},
      {stage0_16[53]},
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage1_19[35],stage1_18[38],stage1_17[82],stage1_16[143],stage1_15[156]}
   );
   gpc615_5 gpc625 (
      {stage0_15[444], stage0_15[445], stage0_15[446], stage0_15[447], stage0_15[448]},
      {stage0_16[54]},
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage1_19[36],stage1_18[39],stage1_17[83],stage1_16[144],stage1_15[157]}
   );
   gpc615_5 gpc626 (
      {stage0_15[449], stage0_15[450], stage0_15[451], stage0_15[452], stage0_15[453]},
      {stage0_16[55]},
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage1_19[37],stage1_18[40],stage1_17[84],stage1_16[145],stage1_15[158]}
   );
   gpc615_5 gpc627 (
      {stage0_15[454], stage0_15[455], stage0_15[456], stage0_15[457], stage0_15[458]},
      {stage0_16[56]},
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage1_19[38],stage1_18[41],stage1_17[85],stage1_16[146],stage1_15[159]}
   );
   gpc615_5 gpc628 (
      {stage0_15[459], stage0_15[460], stage0_15[461], stage0_15[462], stage0_15[463]},
      {stage0_16[57]},
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage1_19[39],stage1_18[42],stage1_17[86],stage1_16[147],stage1_15[160]}
   );
   gpc615_5 gpc629 (
      {stage0_15[464], stage0_15[465], stage0_15[466], stage0_15[467], stage0_15[468]},
      {stage0_16[58]},
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage1_19[40],stage1_18[43],stage1_17[87],stage1_16[148],stage1_15[161]}
   );
   gpc615_5 gpc630 (
      {stage0_15[469], stage0_15[470], stage0_15[471], stage0_15[472], stage0_15[473]},
      {stage0_16[59]},
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage1_19[41],stage1_18[44],stage1_17[88],stage1_16[149],stage1_15[162]}
   );
   gpc615_5 gpc631 (
      {stage0_15[474], stage0_15[475], stage0_15[476], stage0_15[477], stage0_15[478]},
      {stage0_16[60]},
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage1_19[42],stage1_18[45],stage1_17[89],stage1_16[150],stage1_15[163]}
   );
   gpc606_5 gpc632 (
      {stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65], stage0_16[66]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[43],stage1_18[46],stage1_17[90],stage1_16[151]}
   );
   gpc606_5 gpc633 (
      {stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71], stage0_16[72]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[44],stage1_18[47],stage1_17[91],stage1_16[152]}
   );
   gpc606_5 gpc634 (
      {stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[45],stage1_18[48],stage1_17[92],stage1_16[153]}
   );
   gpc606_5 gpc635 (
      {stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[46],stage1_18[49],stage1_17[93],stage1_16[154]}
   );
   gpc606_5 gpc636 (
      {stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[47],stage1_18[50],stage1_17[94],stage1_16[155]}
   );
   gpc606_5 gpc637 (
      {stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[48],stage1_18[51],stage1_17[95],stage1_16[156]}
   );
   gpc606_5 gpc638 (
      {stage0_16[97], stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[49],stage1_18[52],stage1_17[96],stage1_16[157]}
   );
   gpc606_5 gpc639 (
      {stage0_16[103], stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[50],stage1_18[53],stage1_17[97],stage1_16[158]}
   );
   gpc606_5 gpc640 (
      {stage0_16[109], stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[51],stage1_18[54],stage1_17[98],stage1_16[159]}
   );
   gpc606_5 gpc641 (
      {stage0_16[115], stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[52],stage1_18[55],stage1_17[99],stage1_16[160]}
   );
   gpc606_5 gpc642 (
      {stage0_16[121], stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[53],stage1_18[56],stage1_17[100],stage1_16[161]}
   );
   gpc606_5 gpc643 (
      {stage0_16[127], stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[54],stage1_18[57],stage1_17[101],stage1_16[162]}
   );
   gpc606_5 gpc644 (
      {stage0_16[133], stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[55],stage1_18[58],stage1_17[102],stage1_16[163]}
   );
   gpc606_5 gpc645 (
      {stage0_16[139], stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[56],stage1_18[59],stage1_17[103],stage1_16[164]}
   );
   gpc606_5 gpc646 (
      {stage0_16[145], stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[57],stage1_18[60],stage1_17[104],stage1_16[165]}
   );
   gpc606_5 gpc647 (
      {stage0_16[151], stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[58],stage1_18[61],stage1_17[105],stage1_16[166]}
   );
   gpc606_5 gpc648 (
      {stage0_16[157], stage0_16[158], stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[59],stage1_18[62],stage1_17[106],stage1_16[167]}
   );
   gpc606_5 gpc649 (
      {stage0_16[163], stage0_16[164], stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[60],stage1_18[63],stage1_17[107],stage1_16[168]}
   );
   gpc606_5 gpc650 (
      {stage0_16[169], stage0_16[170], stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[61],stage1_18[64],stage1_17[108],stage1_16[169]}
   );
   gpc606_5 gpc651 (
      {stage0_16[175], stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[62],stage1_18[65],stage1_17[109],stage1_16[170]}
   );
   gpc606_5 gpc652 (
      {stage0_16[181], stage0_16[182], stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[63],stage1_18[66],stage1_17[110],stage1_16[171]}
   );
   gpc606_5 gpc653 (
      {stage0_16[187], stage0_16[188], stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[64],stage1_18[67],stage1_17[111],stage1_16[172]}
   );
   gpc606_5 gpc654 (
      {stage0_16[193], stage0_16[194], stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[65],stage1_18[68],stage1_17[112],stage1_16[173]}
   );
   gpc606_5 gpc655 (
      {stage0_16[199], stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[66],stage1_18[69],stage1_17[113],stage1_16[174]}
   );
   gpc606_5 gpc656 (
      {stage0_16[205], stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[67],stage1_18[70],stage1_17[114],stage1_16[175]}
   );
   gpc606_5 gpc657 (
      {stage0_16[211], stage0_16[212], stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[68],stage1_18[71],stage1_17[115],stage1_16[176]}
   );
   gpc606_5 gpc658 (
      {stage0_16[217], stage0_16[218], stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[69],stage1_18[72],stage1_17[116],stage1_16[177]}
   );
   gpc606_5 gpc659 (
      {stage0_16[223], stage0_16[224], stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[70],stage1_18[73],stage1_17[117],stage1_16[178]}
   );
   gpc606_5 gpc660 (
      {stage0_16[229], stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[71],stage1_18[74],stage1_17[118],stage1_16[179]}
   );
   gpc606_5 gpc661 (
      {stage0_16[235], stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[72],stage1_18[75],stage1_17[119],stage1_16[180]}
   );
   gpc606_5 gpc662 (
      {stage0_16[241], stage0_16[242], stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[73],stage1_18[76],stage1_17[120],stage1_16[181]}
   );
   gpc606_5 gpc663 (
      {stage0_16[247], stage0_16[248], stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[74],stage1_18[77],stage1_17[121],stage1_16[182]}
   );
   gpc606_5 gpc664 (
      {stage0_16[253], stage0_16[254], stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[75],stage1_18[78],stage1_17[122],stage1_16[183]}
   );
   gpc606_5 gpc665 (
      {stage0_16[259], stage0_16[260], stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[76],stage1_18[79],stage1_17[123],stage1_16[184]}
   );
   gpc606_5 gpc666 (
      {stage0_16[265], stage0_16[266], stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[77],stage1_18[80],stage1_17[124],stage1_16[185]}
   );
   gpc606_5 gpc667 (
      {stage0_16[271], stage0_16[272], stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[78],stage1_18[81],stage1_17[125],stage1_16[186]}
   );
   gpc606_5 gpc668 (
      {stage0_16[277], stage0_16[278], stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[79],stage1_18[82],stage1_17[126],stage1_16[187]}
   );
   gpc606_5 gpc669 (
      {stage0_16[283], stage0_16[284], stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[80],stage1_18[83],stage1_17[127],stage1_16[188]}
   );
   gpc606_5 gpc670 (
      {stage0_16[289], stage0_16[290], stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[81],stage1_18[84],stage1_17[128],stage1_16[189]}
   );
   gpc606_5 gpc671 (
      {stage0_16[295], stage0_16[296], stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[82],stage1_18[85],stage1_17[129],stage1_16[190]}
   );
   gpc606_5 gpc672 (
      {stage0_16[301], stage0_16[302], stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[83],stage1_18[86],stage1_17[130],stage1_16[191]}
   );
   gpc606_5 gpc673 (
      {stage0_16[307], stage0_16[308], stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[84],stage1_18[87],stage1_17[131],stage1_16[192]}
   );
   gpc606_5 gpc674 (
      {stage0_16[313], stage0_16[314], stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[85],stage1_18[88],stage1_17[132],stage1_16[193]}
   );
   gpc606_5 gpc675 (
      {stage0_16[319], stage0_16[320], stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[86],stage1_18[89],stage1_17[133],stage1_16[194]}
   );
   gpc606_5 gpc676 (
      {stage0_16[325], stage0_16[326], stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[87],stage1_18[90],stage1_17[134],stage1_16[195]}
   );
   gpc606_5 gpc677 (
      {stage0_16[331], stage0_16[332], stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[88],stage1_18[91],stage1_17[135],stage1_16[196]}
   );
   gpc606_5 gpc678 (
      {stage0_16[337], stage0_16[338], stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[89],stage1_18[92],stage1_17[136],stage1_16[197]}
   );
   gpc606_5 gpc679 (
      {stage0_16[343], stage0_16[344], stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[90],stage1_18[93],stage1_17[137],stage1_16[198]}
   );
   gpc606_5 gpc680 (
      {stage0_16[349], stage0_16[350], stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354]},
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage1_20[48],stage1_19[91],stage1_18[94],stage1_17[138],stage1_16[199]}
   );
   gpc606_5 gpc681 (
      {stage0_16[355], stage0_16[356], stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360]},
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage1_20[49],stage1_19[92],stage1_18[95],stage1_17[139],stage1_16[200]}
   );
   gpc606_5 gpc682 (
      {stage0_16[361], stage0_16[362], stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366]},
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage1_20[50],stage1_19[93],stage1_18[96],stage1_17[140],stage1_16[201]}
   );
   gpc606_5 gpc683 (
      {stage0_16[367], stage0_16[368], stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372]},
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage1_20[51],stage1_19[94],stage1_18[97],stage1_17[141],stage1_16[202]}
   );
   gpc606_5 gpc684 (
      {stage0_16[373], stage0_16[374], stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378]},
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316], stage0_18[317]},
      {stage1_20[52],stage1_19[95],stage1_18[98],stage1_17[142],stage1_16[203]}
   );
   gpc606_5 gpc685 (
      {stage0_16[379], stage0_16[380], stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384]},
      {stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321], stage0_18[322], stage0_18[323]},
      {stage1_20[53],stage1_19[96],stage1_18[99],stage1_17[143],stage1_16[204]}
   );
   gpc606_5 gpc686 (
      {stage0_16[385], stage0_16[386], stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390]},
      {stage0_18[324], stage0_18[325], stage0_18[326], stage0_18[327], stage0_18[328], stage0_18[329]},
      {stage1_20[54],stage1_19[97],stage1_18[100],stage1_17[144],stage1_16[205]}
   );
   gpc606_5 gpc687 (
      {stage0_16[391], stage0_16[392], stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396]},
      {stage0_18[330], stage0_18[331], stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335]},
      {stage1_20[55],stage1_19[98],stage1_18[101],stage1_17[145],stage1_16[206]}
   );
   gpc606_5 gpc688 (
      {stage0_16[397], stage0_16[398], stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402]},
      {stage0_18[336], stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340], stage0_18[341]},
      {stage1_20[56],stage1_19[99],stage1_18[102],stage1_17[146],stage1_16[207]}
   );
   gpc606_5 gpc689 (
      {stage0_16[403], stage0_16[404], stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408]},
      {stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345], stage0_18[346], stage0_18[347]},
      {stage1_20[57],stage1_19[100],stage1_18[103],stage1_17[147],stage1_16[208]}
   );
   gpc606_5 gpc690 (
      {stage0_16[409], stage0_16[410], stage0_16[411], stage0_16[412], stage0_16[413], stage0_16[414]},
      {stage0_18[348], stage0_18[349], stage0_18[350], stage0_18[351], stage0_18[352], stage0_18[353]},
      {stage1_20[58],stage1_19[101],stage1_18[104],stage1_17[148],stage1_16[209]}
   );
   gpc606_5 gpc691 (
      {stage0_16[415], stage0_16[416], stage0_16[417], stage0_16[418], stage0_16[419], stage0_16[420]},
      {stage0_18[354], stage0_18[355], stage0_18[356], stage0_18[357], stage0_18[358], stage0_18[359]},
      {stage1_20[59],stage1_19[102],stage1_18[105],stage1_17[149],stage1_16[210]}
   );
   gpc606_5 gpc692 (
      {stage0_16[421], stage0_16[422], stage0_16[423], stage0_16[424], stage0_16[425], stage0_16[426]},
      {stage0_18[360], stage0_18[361], stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365]},
      {stage1_20[60],stage1_19[103],stage1_18[106],stage1_17[150],stage1_16[211]}
   );
   gpc606_5 gpc693 (
      {stage0_16[427], stage0_16[428], stage0_16[429], stage0_16[430], stage0_16[431], stage0_16[432]},
      {stage0_18[366], stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370], stage0_18[371]},
      {stage1_20[61],stage1_19[104],stage1_18[107],stage1_17[151],stage1_16[212]}
   );
   gpc606_5 gpc694 (
      {stage0_16[433], stage0_16[434], stage0_16[435], stage0_16[436], stage0_16[437], stage0_16[438]},
      {stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375], stage0_18[376], stage0_18[377]},
      {stage1_20[62],stage1_19[105],stage1_18[108],stage1_17[152],stage1_16[213]}
   );
   gpc606_5 gpc695 (
      {stage0_16[439], stage0_16[440], stage0_16[441], stage0_16[442], stage0_16[443], stage0_16[444]},
      {stage0_18[378], stage0_18[379], stage0_18[380], stage0_18[381], stage0_18[382], stage0_18[383]},
      {stage1_20[63],stage1_19[106],stage1_18[109],stage1_17[153],stage1_16[214]}
   );
   gpc606_5 gpc696 (
      {stage0_16[445], stage0_16[446], stage0_16[447], stage0_16[448], stage0_16[449], stage0_16[450]},
      {stage0_18[384], stage0_18[385], stage0_18[386], stage0_18[387], stage0_18[388], stage0_18[389]},
      {stage1_20[64],stage1_19[107],stage1_18[110],stage1_17[154],stage1_16[215]}
   );
   gpc606_5 gpc697 (
      {stage0_16[451], stage0_16[452], stage0_16[453], stage0_16[454], stage0_16[455], stage0_16[456]},
      {stage0_18[390], stage0_18[391], stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395]},
      {stage1_20[65],stage1_19[108],stage1_18[111],stage1_17[155],stage1_16[216]}
   );
   gpc606_5 gpc698 (
      {stage0_16[457], stage0_16[458], stage0_16[459], stage0_16[460], stage0_16[461], stage0_16[462]},
      {stage0_18[396], stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400], stage0_18[401]},
      {stage1_20[66],stage1_19[109],stage1_18[112],stage1_17[156],stage1_16[217]}
   );
   gpc606_5 gpc699 (
      {stage0_16[463], stage0_16[464], stage0_16[465], stage0_16[466], stage0_16[467], stage0_16[468]},
      {stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405], stage0_18[406], stage0_18[407]},
      {stage1_20[67],stage1_19[110],stage1_18[113],stage1_17[157],stage1_16[218]}
   );
   gpc606_5 gpc700 (
      {stage0_16[469], stage0_16[470], stage0_16[471], stage0_16[472], stage0_16[473], stage0_16[474]},
      {stage0_18[408], stage0_18[409], stage0_18[410], stage0_18[411], stage0_18[412], stage0_18[413]},
      {stage1_20[68],stage1_19[111],stage1_18[114],stage1_17[158],stage1_16[219]}
   );
   gpc606_5 gpc701 (
      {stage0_16[475], stage0_16[476], stage0_16[477], stage0_16[478], stage0_16[479], stage0_16[480]},
      {stage0_18[414], stage0_18[415], stage0_18[416], stage0_18[417], stage0_18[418], stage0_18[419]},
      {stage1_20[69],stage1_19[112],stage1_18[115],stage1_17[159],stage1_16[220]}
   );
   gpc606_5 gpc702 (
      {stage0_16[481], stage0_16[482], stage0_16[483], stage0_16[484], stage0_16[485], 1'b0},
      {stage0_18[420], stage0_18[421], stage0_18[422], stage0_18[423], stage0_18[424], stage0_18[425]},
      {stage1_20[70],stage1_19[113],stage1_18[116],stage1_17[160],stage1_16[221]}
   );
   gpc606_5 gpc703 (
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[71],stage1_19[114],stage1_18[117],stage1_17[161]}
   );
   gpc606_5 gpc704 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[72],stage1_19[115],stage1_18[118],stage1_17[162]}
   );
   gpc606_5 gpc705 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[73],stage1_19[116],stage1_18[119],stage1_17[163]}
   );
   gpc606_5 gpc706 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[74],stage1_19[117],stage1_18[120],stage1_17[164]}
   );
   gpc606_5 gpc707 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[75],stage1_19[118],stage1_18[121],stage1_17[165]}
   );
   gpc606_5 gpc708 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[76],stage1_19[119],stage1_18[122],stage1_17[166]}
   );
   gpc606_5 gpc709 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[77],stage1_19[120],stage1_18[123],stage1_17[167]}
   );
   gpc606_5 gpc710 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[78],stage1_19[121],stage1_18[124],stage1_17[168]}
   );
   gpc606_5 gpc711 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[79],stage1_19[122],stage1_18[125],stage1_17[169]}
   );
   gpc606_5 gpc712 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[80],stage1_19[123],stage1_18[126],stage1_17[170]}
   );
   gpc606_5 gpc713 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[81],stage1_19[124],stage1_18[127],stage1_17[171]}
   );
   gpc606_5 gpc714 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[82],stage1_19[125],stage1_18[128],stage1_17[172]}
   );
   gpc606_5 gpc715 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[83],stage1_19[126],stage1_18[129],stage1_17[173]}
   );
   gpc606_5 gpc716 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[84],stage1_19[127],stage1_18[130],stage1_17[174]}
   );
   gpc606_5 gpc717 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[85],stage1_19[128],stage1_18[131],stage1_17[175]}
   );
   gpc606_5 gpc718 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[86],stage1_19[129],stage1_18[132],stage1_17[176]}
   );
   gpc606_5 gpc719 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[87],stage1_19[130],stage1_18[133],stage1_17[177]}
   );
   gpc606_5 gpc720 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[88],stage1_19[131],stage1_18[134],stage1_17[178]}
   );
   gpc606_5 gpc721 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[89],stage1_19[132],stage1_18[135],stage1_17[179]}
   );
   gpc606_5 gpc722 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[90],stage1_19[133],stage1_18[136],stage1_17[180]}
   );
   gpc606_5 gpc723 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[91],stage1_19[134],stage1_18[137],stage1_17[181]}
   );
   gpc606_5 gpc724 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[92],stage1_19[135],stage1_18[138],stage1_17[182]}
   );
   gpc606_5 gpc725 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[93],stage1_19[136],stage1_18[139],stage1_17[183]}
   );
   gpc606_5 gpc726 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[94],stage1_19[137],stage1_18[140],stage1_17[184]}
   );
   gpc606_5 gpc727 (
      {stage0_17[402], stage0_17[403], stage0_17[404], stage0_17[405], stage0_17[406], stage0_17[407]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[95],stage1_19[138],stage1_18[141],stage1_17[185]}
   );
   gpc606_5 gpc728 (
      {stage0_17[408], stage0_17[409], stage0_17[410], stage0_17[411], stage0_17[412], stage0_17[413]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[96],stage1_19[139],stage1_18[142],stage1_17[186]}
   );
   gpc606_5 gpc729 (
      {stage0_17[414], stage0_17[415], stage0_17[416], stage0_17[417], stage0_17[418], stage0_17[419]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[97],stage1_19[140],stage1_18[143],stage1_17[187]}
   );
   gpc606_5 gpc730 (
      {stage0_17[420], stage0_17[421], stage0_17[422], stage0_17[423], stage0_17[424], stage0_17[425]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[98],stage1_19[141],stage1_18[144],stage1_17[188]}
   );
   gpc606_5 gpc731 (
      {stage0_17[426], stage0_17[427], stage0_17[428], stage0_17[429], stage0_17[430], stage0_17[431]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[99],stage1_19[142],stage1_18[145],stage1_17[189]}
   );
   gpc606_5 gpc732 (
      {stage0_17[432], stage0_17[433], stage0_17[434], stage0_17[435], stage0_17[436], stage0_17[437]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[100],stage1_19[143],stage1_18[146],stage1_17[190]}
   );
   gpc606_5 gpc733 (
      {stage0_17[438], stage0_17[439], stage0_17[440], stage0_17[441], stage0_17[442], stage0_17[443]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[101],stage1_19[144],stage1_18[147],stage1_17[191]}
   );
   gpc606_5 gpc734 (
      {stage0_17[444], stage0_17[445], stage0_17[446], stage0_17[447], stage0_17[448], stage0_17[449]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[102],stage1_19[145],stage1_18[148],stage1_17[192]}
   );
   gpc615_5 gpc735 (
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196]},
      {stage0_20[0]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[0],stage1_21[32],stage1_20[103],stage1_19[146]}
   );
   gpc615_5 gpc736 (
      {stage0_19[197], stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201]},
      {stage0_20[1]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[1],stage1_21[33],stage1_20[104],stage1_19[147]}
   );
   gpc615_5 gpc737 (
      {stage0_19[202], stage0_19[203], stage0_19[204], stage0_19[205], stage0_19[206]},
      {stage0_20[2]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[2],stage1_21[34],stage1_20[105],stage1_19[148]}
   );
   gpc615_5 gpc738 (
      {stage0_19[207], stage0_19[208], stage0_19[209], stage0_19[210], stage0_19[211]},
      {stage0_20[3]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[3],stage1_21[35],stage1_20[106],stage1_19[149]}
   );
   gpc615_5 gpc739 (
      {stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215], stage0_19[216]},
      {stage0_20[4]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[4],stage1_21[36],stage1_20[107],stage1_19[150]}
   );
   gpc615_5 gpc740 (
      {stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage0_20[5]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[5],stage1_21[37],stage1_20[108],stage1_19[151]}
   );
   gpc615_5 gpc741 (
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226]},
      {stage0_20[6]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[6],stage1_21[38],stage1_20[109],stage1_19[152]}
   );
   gpc615_5 gpc742 (
      {stage0_19[227], stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231]},
      {stage0_20[7]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[7],stage1_21[39],stage1_20[110],stage1_19[153]}
   );
   gpc615_5 gpc743 (
      {stage0_19[232], stage0_19[233], stage0_19[234], stage0_19[235], stage0_19[236]},
      {stage0_20[8]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[8],stage1_21[40],stage1_20[111],stage1_19[154]}
   );
   gpc615_5 gpc744 (
      {stage0_19[237], stage0_19[238], stage0_19[239], stage0_19[240], stage0_19[241]},
      {stage0_20[9]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[9],stage1_21[41],stage1_20[112],stage1_19[155]}
   );
   gpc615_5 gpc745 (
      {stage0_19[242], stage0_19[243], stage0_19[244], stage0_19[245], stage0_19[246]},
      {stage0_20[10]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[10],stage1_21[42],stage1_20[113],stage1_19[156]}
   );
   gpc615_5 gpc746 (
      {stage0_19[247], stage0_19[248], stage0_19[249], stage0_19[250], stage0_19[251]},
      {stage0_20[11]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[11],stage1_21[43],stage1_20[114],stage1_19[157]}
   );
   gpc615_5 gpc747 (
      {stage0_19[252], stage0_19[253], stage0_19[254], stage0_19[255], stage0_19[256]},
      {stage0_20[12]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[12],stage1_21[44],stage1_20[115],stage1_19[158]}
   );
   gpc615_5 gpc748 (
      {stage0_19[257], stage0_19[258], stage0_19[259], stage0_19[260], stage0_19[261]},
      {stage0_20[13]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[13],stage1_21[45],stage1_20[116],stage1_19[159]}
   );
   gpc615_5 gpc749 (
      {stage0_19[262], stage0_19[263], stage0_19[264], stage0_19[265], stage0_19[266]},
      {stage0_20[14]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage1_23[14],stage1_22[14],stage1_21[46],stage1_20[117],stage1_19[160]}
   );
   gpc615_5 gpc750 (
      {stage0_19[267], stage0_19[268], stage0_19[269], stage0_19[270], stage0_19[271]},
      {stage0_20[15]},
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage1_23[15],stage1_22[15],stage1_21[47],stage1_20[118],stage1_19[161]}
   );
   gpc615_5 gpc751 (
      {stage0_19[272], stage0_19[273], stage0_19[274], stage0_19[275], stage0_19[276]},
      {stage0_20[16]},
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage1_23[16],stage1_22[16],stage1_21[48],stage1_20[119],stage1_19[162]}
   );
   gpc615_5 gpc752 (
      {stage0_19[277], stage0_19[278], stage0_19[279], stage0_19[280], stage0_19[281]},
      {stage0_20[17]},
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage1_23[17],stage1_22[17],stage1_21[49],stage1_20[120],stage1_19[163]}
   );
   gpc615_5 gpc753 (
      {stage0_19[282], stage0_19[283], stage0_19[284], stage0_19[285], stage0_19[286]},
      {stage0_20[18]},
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage1_23[18],stage1_22[18],stage1_21[50],stage1_20[121],stage1_19[164]}
   );
   gpc615_5 gpc754 (
      {stage0_19[287], stage0_19[288], stage0_19[289], stage0_19[290], stage0_19[291]},
      {stage0_20[19]},
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage1_23[19],stage1_22[19],stage1_21[51],stage1_20[122],stage1_19[165]}
   );
   gpc615_5 gpc755 (
      {stage0_19[292], stage0_19[293], stage0_19[294], stage0_19[295], stage0_19[296]},
      {stage0_20[20]},
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage1_23[20],stage1_22[20],stage1_21[52],stage1_20[123],stage1_19[166]}
   );
   gpc615_5 gpc756 (
      {stage0_19[297], stage0_19[298], stage0_19[299], stage0_19[300], stage0_19[301]},
      {stage0_20[21]},
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage1_23[21],stage1_22[21],stage1_21[53],stage1_20[124],stage1_19[167]}
   );
   gpc615_5 gpc757 (
      {stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305], stage0_19[306]},
      {stage0_20[22]},
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage1_23[22],stage1_22[22],stage1_21[54],stage1_20[125],stage1_19[168]}
   );
   gpc615_5 gpc758 (
      {stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage0_20[23]},
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage1_23[23],stage1_22[23],stage1_21[55],stage1_20[126],stage1_19[169]}
   );
   gpc615_5 gpc759 (
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316]},
      {stage0_20[24]},
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage1_23[24],stage1_22[24],stage1_21[56],stage1_20[127],stage1_19[170]}
   );
   gpc615_5 gpc760 (
      {stage0_19[317], stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321]},
      {stage0_20[25]},
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage1_23[25],stage1_22[25],stage1_21[57],stage1_20[128],stage1_19[171]}
   );
   gpc615_5 gpc761 (
      {stage0_19[322], stage0_19[323], stage0_19[324], stage0_19[325], stage0_19[326]},
      {stage0_20[26]},
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage1_23[26],stage1_22[26],stage1_21[58],stage1_20[129],stage1_19[172]}
   );
   gpc615_5 gpc762 (
      {stage0_19[327], stage0_19[328], stage0_19[329], stage0_19[330], stage0_19[331]},
      {stage0_20[27]},
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage1_23[27],stage1_22[27],stage1_21[59],stage1_20[130],stage1_19[173]}
   );
   gpc615_5 gpc763 (
      {stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335], stage0_19[336]},
      {stage0_20[28]},
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage1_23[28],stage1_22[28],stage1_21[60],stage1_20[131],stage1_19[174]}
   );
   gpc615_5 gpc764 (
      {stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage0_20[29]},
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage1_23[29],stage1_22[29],stage1_21[61],stage1_20[132],stage1_19[175]}
   );
   gpc615_5 gpc765 (
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346]},
      {stage0_20[30]},
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage1_23[30],stage1_22[30],stage1_21[62],stage1_20[133],stage1_19[176]}
   );
   gpc615_5 gpc766 (
      {stage0_19[347], stage0_19[348], stage0_19[349], stage0_19[350], stage0_19[351]},
      {stage0_20[31]},
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage1_23[31],stage1_22[31],stage1_21[63],stage1_20[134],stage1_19[177]}
   );
   gpc615_5 gpc767 (
      {stage0_19[352], stage0_19[353], stage0_19[354], stage0_19[355], stage0_19[356]},
      {stage0_20[32]},
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage1_23[32],stage1_22[32],stage1_21[64],stage1_20[135],stage1_19[178]}
   );
   gpc615_5 gpc768 (
      {stage0_19[357], stage0_19[358], stage0_19[359], stage0_19[360], stage0_19[361]},
      {stage0_20[33]},
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage1_23[33],stage1_22[33],stage1_21[65],stage1_20[136],stage1_19[179]}
   );
   gpc615_5 gpc769 (
      {stage0_19[362], stage0_19[363], stage0_19[364], stage0_19[365], stage0_19[366]},
      {stage0_20[34]},
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage1_23[34],stage1_22[34],stage1_21[66],stage1_20[137],stage1_19[180]}
   );
   gpc615_5 gpc770 (
      {stage0_19[367], stage0_19[368], stage0_19[369], stage0_19[370], stage0_19[371]},
      {stage0_20[35]},
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage1_23[35],stage1_22[35],stage1_21[67],stage1_20[138],stage1_19[181]}
   );
   gpc615_5 gpc771 (
      {stage0_19[372], stage0_19[373], stage0_19[374], stage0_19[375], stage0_19[376]},
      {stage0_20[36]},
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage1_23[36],stage1_22[36],stage1_21[68],stage1_20[139],stage1_19[182]}
   );
   gpc615_5 gpc772 (
      {stage0_19[377], stage0_19[378], stage0_19[379], stage0_19[380], stage0_19[381]},
      {stage0_20[37]},
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage1_23[37],stage1_22[37],stage1_21[69],stage1_20[140],stage1_19[183]}
   );
   gpc615_5 gpc773 (
      {stage0_19[382], stage0_19[383], stage0_19[384], stage0_19[385], stage0_19[386]},
      {stage0_20[38]},
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage1_23[38],stage1_22[38],stage1_21[70],stage1_20[141],stage1_19[184]}
   );
   gpc615_5 gpc774 (
      {stage0_19[387], stage0_19[388], stage0_19[389], stage0_19[390], stage0_19[391]},
      {stage0_20[39]},
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage1_23[39],stage1_22[39],stage1_21[71],stage1_20[142],stage1_19[185]}
   );
   gpc615_5 gpc775 (
      {stage0_19[392], stage0_19[393], stage0_19[394], stage0_19[395], stage0_19[396]},
      {stage0_20[40]},
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage1_23[40],stage1_22[40],stage1_21[72],stage1_20[143],stage1_19[186]}
   );
   gpc1343_5 gpc776 (
      {stage0_20[41], stage0_20[42], stage0_20[43]},
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249]},
      {stage0_22[0], stage0_22[1], stage0_22[2]},
      {stage0_23[0]},
      {stage1_24[0],stage1_23[41],stage1_22[41],stage1_21[73],stage1_20[144]}
   );
   gpc1163_5 gpc777 (
      {stage0_20[44], stage0_20[45], stage0_20[46]},
      {stage0_21[250], stage0_21[251], stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255]},
      {stage0_22[3]},
      {stage0_23[1]},
      {stage1_24[1],stage1_23[42],stage1_22[42],stage1_21[74],stage1_20[145]}
   );
   gpc1163_5 gpc778 (
      {stage0_20[47], stage0_20[48], stage0_20[49]},
      {stage0_21[256], stage0_21[257], stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261]},
      {stage0_22[4]},
      {stage0_23[2]},
      {stage1_24[2],stage1_23[43],stage1_22[43],stage1_21[75],stage1_20[146]}
   );
   gpc1163_5 gpc779 (
      {stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[262], stage0_21[263], stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267]},
      {stage0_22[5]},
      {stage0_23[3]},
      {stage1_24[3],stage1_23[44],stage1_22[44],stage1_21[76],stage1_20[147]}
   );
   gpc1163_5 gpc780 (
      {stage0_20[53], stage0_20[54], stage0_20[55]},
      {stage0_21[268], stage0_21[269], stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273]},
      {stage0_22[6]},
      {stage0_23[4]},
      {stage1_24[4],stage1_23[45],stage1_22[45],stage1_21[77],stage1_20[148]}
   );
   gpc1163_5 gpc781 (
      {stage0_20[56], stage0_20[57], stage0_20[58]},
      {stage0_21[274], stage0_21[275], stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279]},
      {stage0_22[7]},
      {stage0_23[5]},
      {stage1_24[5],stage1_23[46],stage1_22[46],stage1_21[78],stage1_20[149]}
   );
   gpc1163_5 gpc782 (
      {stage0_20[59], stage0_20[60], stage0_20[61]},
      {stage0_21[280], stage0_21[281], stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285]},
      {stage0_22[8]},
      {stage0_23[6]},
      {stage1_24[6],stage1_23[47],stage1_22[47],stage1_21[79],stage1_20[150]}
   );
   gpc606_5 gpc783 (
      {stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65], stage0_20[66], stage0_20[67]},
      {stage0_22[9], stage0_22[10], stage0_22[11], stage0_22[12], stage0_22[13], stage0_22[14]},
      {stage1_24[7],stage1_23[48],stage1_22[48],stage1_21[80],stage1_20[151]}
   );
   gpc606_5 gpc784 (
      {stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73]},
      {stage0_22[15], stage0_22[16], stage0_22[17], stage0_22[18], stage0_22[19], stage0_22[20]},
      {stage1_24[8],stage1_23[49],stage1_22[49],stage1_21[81],stage1_20[152]}
   );
   gpc606_5 gpc785 (
      {stage0_20[74], stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79]},
      {stage0_22[21], stage0_22[22], stage0_22[23], stage0_22[24], stage0_22[25], stage0_22[26]},
      {stage1_24[9],stage1_23[50],stage1_22[50],stage1_21[82],stage1_20[153]}
   );
   gpc606_5 gpc786 (
      {stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85]},
      {stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30], stage0_22[31], stage0_22[32]},
      {stage1_24[10],stage1_23[51],stage1_22[51],stage1_21[83],stage1_20[154]}
   );
   gpc606_5 gpc787 (
      {stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91]},
      {stage0_22[33], stage0_22[34], stage0_22[35], stage0_22[36], stage0_22[37], stage0_22[38]},
      {stage1_24[11],stage1_23[52],stage1_22[52],stage1_21[84],stage1_20[155]}
   );
   gpc606_5 gpc788 (
      {stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97]},
      {stage0_22[39], stage0_22[40], stage0_22[41], stage0_22[42], stage0_22[43], stage0_22[44]},
      {stage1_24[12],stage1_23[53],stage1_22[53],stage1_21[85],stage1_20[156]}
   );
   gpc606_5 gpc789 (
      {stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103]},
      {stage0_22[45], stage0_22[46], stage0_22[47], stage0_22[48], stage0_22[49], stage0_22[50]},
      {stage1_24[13],stage1_23[54],stage1_22[54],stage1_21[86],stage1_20[157]}
   );
   gpc606_5 gpc790 (
      {stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109]},
      {stage0_22[51], stage0_22[52], stage0_22[53], stage0_22[54], stage0_22[55], stage0_22[56]},
      {stage1_24[14],stage1_23[55],stage1_22[55],stage1_21[87],stage1_20[158]}
   );
   gpc606_5 gpc791 (
      {stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115]},
      {stage0_22[57], stage0_22[58], stage0_22[59], stage0_22[60], stage0_22[61], stage0_22[62]},
      {stage1_24[15],stage1_23[56],stage1_22[56],stage1_21[88],stage1_20[159]}
   );
   gpc606_5 gpc792 (
      {stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119], stage0_20[120], stage0_20[121]},
      {stage0_22[63], stage0_22[64], stage0_22[65], stage0_22[66], stage0_22[67], stage0_22[68]},
      {stage1_24[16],stage1_23[57],stage1_22[57],stage1_21[89],stage1_20[160]}
   );
   gpc606_5 gpc793 (
      {stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125], stage0_20[126], stage0_20[127]},
      {stage0_22[69], stage0_22[70], stage0_22[71], stage0_22[72], stage0_22[73], stage0_22[74]},
      {stage1_24[17],stage1_23[58],stage1_22[58],stage1_21[90],stage1_20[161]}
   );
   gpc606_5 gpc794 (
      {stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131], stage0_20[132], stage0_20[133]},
      {stage0_22[75], stage0_22[76], stage0_22[77], stage0_22[78], stage0_22[79], stage0_22[80]},
      {stage1_24[18],stage1_23[59],stage1_22[59],stage1_21[91],stage1_20[162]}
   );
   gpc606_5 gpc795 (
      {stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137], stage0_20[138], stage0_20[139]},
      {stage0_22[81], stage0_22[82], stage0_22[83], stage0_22[84], stage0_22[85], stage0_22[86]},
      {stage1_24[19],stage1_23[60],stage1_22[60],stage1_21[92],stage1_20[163]}
   );
   gpc606_5 gpc796 (
      {stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143], stage0_20[144], stage0_20[145]},
      {stage0_22[87], stage0_22[88], stage0_22[89], stage0_22[90], stage0_22[91], stage0_22[92]},
      {stage1_24[20],stage1_23[61],stage1_22[61],stage1_21[93],stage1_20[164]}
   );
   gpc606_5 gpc797 (
      {stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149], stage0_20[150], stage0_20[151]},
      {stage0_22[93], stage0_22[94], stage0_22[95], stage0_22[96], stage0_22[97], stage0_22[98]},
      {stage1_24[21],stage1_23[62],stage1_22[62],stage1_21[94],stage1_20[165]}
   );
   gpc606_5 gpc798 (
      {stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155], stage0_20[156], stage0_20[157]},
      {stage0_22[99], stage0_22[100], stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104]},
      {stage1_24[22],stage1_23[63],stage1_22[63],stage1_21[95],stage1_20[166]}
   );
   gpc606_5 gpc799 (
      {stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161], stage0_20[162], stage0_20[163]},
      {stage0_22[105], stage0_22[106], stage0_22[107], stage0_22[108], stage0_22[109], stage0_22[110]},
      {stage1_24[23],stage1_23[64],stage1_22[64],stage1_21[96],stage1_20[167]}
   );
   gpc606_5 gpc800 (
      {stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167], stage0_20[168], stage0_20[169]},
      {stage0_22[111], stage0_22[112], stage0_22[113], stage0_22[114], stage0_22[115], stage0_22[116]},
      {stage1_24[24],stage1_23[65],stage1_22[65],stage1_21[97],stage1_20[168]}
   );
   gpc606_5 gpc801 (
      {stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173], stage0_20[174], stage0_20[175]},
      {stage0_22[117], stage0_22[118], stage0_22[119], stage0_22[120], stage0_22[121], stage0_22[122]},
      {stage1_24[25],stage1_23[66],stage1_22[66],stage1_21[98],stage1_20[169]}
   );
   gpc606_5 gpc802 (
      {stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179], stage0_20[180], stage0_20[181]},
      {stage0_22[123], stage0_22[124], stage0_22[125], stage0_22[126], stage0_22[127], stage0_22[128]},
      {stage1_24[26],stage1_23[67],stage1_22[67],stage1_21[99],stage1_20[170]}
   );
   gpc606_5 gpc803 (
      {stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185], stage0_20[186], stage0_20[187]},
      {stage0_22[129], stage0_22[130], stage0_22[131], stage0_22[132], stage0_22[133], stage0_22[134]},
      {stage1_24[27],stage1_23[68],stage1_22[68],stage1_21[100],stage1_20[171]}
   );
   gpc606_5 gpc804 (
      {stage0_20[188], stage0_20[189], stage0_20[190], stage0_20[191], stage0_20[192], stage0_20[193]},
      {stage0_22[135], stage0_22[136], stage0_22[137], stage0_22[138], stage0_22[139], stage0_22[140]},
      {stage1_24[28],stage1_23[69],stage1_22[69],stage1_21[101],stage1_20[172]}
   );
   gpc606_5 gpc805 (
      {stage0_20[194], stage0_20[195], stage0_20[196], stage0_20[197], stage0_20[198], stage0_20[199]},
      {stage0_22[141], stage0_22[142], stage0_22[143], stage0_22[144], stage0_22[145], stage0_22[146]},
      {stage1_24[29],stage1_23[70],stage1_22[70],stage1_21[102],stage1_20[173]}
   );
   gpc606_5 gpc806 (
      {stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203], stage0_20[204], stage0_20[205]},
      {stage0_22[147], stage0_22[148], stage0_22[149], stage0_22[150], stage0_22[151], stage0_22[152]},
      {stage1_24[30],stage1_23[71],stage1_22[71],stage1_21[103],stage1_20[174]}
   );
   gpc606_5 gpc807 (
      {stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209], stage0_20[210], stage0_20[211]},
      {stage0_22[153], stage0_22[154], stage0_22[155], stage0_22[156], stage0_22[157], stage0_22[158]},
      {stage1_24[31],stage1_23[72],stage1_22[72],stage1_21[104],stage1_20[175]}
   );
   gpc606_5 gpc808 (
      {stage0_20[212], stage0_20[213], stage0_20[214], stage0_20[215], stage0_20[216], stage0_20[217]},
      {stage0_22[159], stage0_22[160], stage0_22[161], stage0_22[162], stage0_22[163], stage0_22[164]},
      {stage1_24[32],stage1_23[73],stage1_22[73],stage1_21[105],stage1_20[176]}
   );
   gpc606_5 gpc809 (
      {stage0_20[218], stage0_20[219], stage0_20[220], stage0_20[221], stage0_20[222], stage0_20[223]},
      {stage0_22[165], stage0_22[166], stage0_22[167], stage0_22[168], stage0_22[169], stage0_22[170]},
      {stage1_24[33],stage1_23[74],stage1_22[74],stage1_21[106],stage1_20[177]}
   );
   gpc606_5 gpc810 (
      {stage0_20[224], stage0_20[225], stage0_20[226], stage0_20[227], stage0_20[228], stage0_20[229]},
      {stage0_22[171], stage0_22[172], stage0_22[173], stage0_22[174], stage0_22[175], stage0_22[176]},
      {stage1_24[34],stage1_23[75],stage1_22[75],stage1_21[107],stage1_20[178]}
   );
   gpc606_5 gpc811 (
      {stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233], stage0_20[234], stage0_20[235]},
      {stage0_22[177], stage0_22[178], stage0_22[179], stage0_22[180], stage0_22[181], stage0_22[182]},
      {stage1_24[35],stage1_23[76],stage1_22[76],stage1_21[108],stage1_20[179]}
   );
   gpc606_5 gpc812 (
      {stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239], stage0_20[240], stage0_20[241]},
      {stage0_22[183], stage0_22[184], stage0_22[185], stage0_22[186], stage0_22[187], stage0_22[188]},
      {stage1_24[36],stage1_23[77],stage1_22[77],stage1_21[109],stage1_20[180]}
   );
   gpc606_5 gpc813 (
      {stage0_20[242], stage0_20[243], stage0_20[244], stage0_20[245], stage0_20[246], stage0_20[247]},
      {stage0_22[189], stage0_22[190], stage0_22[191], stage0_22[192], stage0_22[193], stage0_22[194]},
      {stage1_24[37],stage1_23[78],stage1_22[78],stage1_21[110],stage1_20[181]}
   );
   gpc606_5 gpc814 (
      {stage0_20[248], stage0_20[249], stage0_20[250], stage0_20[251], stage0_20[252], stage0_20[253]},
      {stage0_22[195], stage0_22[196], stage0_22[197], stage0_22[198], stage0_22[199], stage0_22[200]},
      {stage1_24[38],stage1_23[79],stage1_22[79],stage1_21[111],stage1_20[182]}
   );
   gpc606_5 gpc815 (
      {stage0_20[254], stage0_20[255], stage0_20[256], stage0_20[257], stage0_20[258], stage0_20[259]},
      {stage0_22[201], stage0_22[202], stage0_22[203], stage0_22[204], stage0_22[205], stage0_22[206]},
      {stage1_24[39],stage1_23[80],stage1_22[80],stage1_21[112],stage1_20[183]}
   );
   gpc606_5 gpc816 (
      {stage0_20[260], stage0_20[261], stage0_20[262], stage0_20[263], stage0_20[264], stage0_20[265]},
      {stage0_22[207], stage0_22[208], stage0_22[209], stage0_22[210], stage0_22[211], stage0_22[212]},
      {stage1_24[40],stage1_23[81],stage1_22[81],stage1_21[113],stage1_20[184]}
   );
   gpc606_5 gpc817 (
      {stage0_20[266], stage0_20[267], stage0_20[268], stage0_20[269], stage0_20[270], stage0_20[271]},
      {stage0_22[213], stage0_22[214], stage0_22[215], stage0_22[216], stage0_22[217], stage0_22[218]},
      {stage1_24[41],stage1_23[82],stage1_22[82],stage1_21[114],stage1_20[185]}
   );
   gpc606_5 gpc818 (
      {stage0_20[272], stage0_20[273], stage0_20[274], stage0_20[275], stage0_20[276], stage0_20[277]},
      {stage0_22[219], stage0_22[220], stage0_22[221], stage0_22[222], stage0_22[223], stage0_22[224]},
      {stage1_24[42],stage1_23[83],stage1_22[83],stage1_21[115],stage1_20[186]}
   );
   gpc606_5 gpc819 (
      {stage0_20[278], stage0_20[279], stage0_20[280], stage0_20[281], stage0_20[282], stage0_20[283]},
      {stage0_22[225], stage0_22[226], stage0_22[227], stage0_22[228], stage0_22[229], stage0_22[230]},
      {stage1_24[43],stage1_23[84],stage1_22[84],stage1_21[116],stage1_20[187]}
   );
   gpc606_5 gpc820 (
      {stage0_20[284], stage0_20[285], stage0_20[286], stage0_20[287], stage0_20[288], stage0_20[289]},
      {stage0_22[231], stage0_22[232], stage0_22[233], stage0_22[234], stage0_22[235], stage0_22[236]},
      {stage1_24[44],stage1_23[85],stage1_22[85],stage1_21[117],stage1_20[188]}
   );
   gpc606_5 gpc821 (
      {stage0_20[290], stage0_20[291], stage0_20[292], stage0_20[293], stage0_20[294], stage0_20[295]},
      {stage0_22[237], stage0_22[238], stage0_22[239], stage0_22[240], stage0_22[241], stage0_22[242]},
      {stage1_24[45],stage1_23[86],stage1_22[86],stage1_21[118],stage1_20[189]}
   );
   gpc606_5 gpc822 (
      {stage0_20[296], stage0_20[297], stage0_20[298], stage0_20[299], stage0_20[300], stage0_20[301]},
      {stage0_22[243], stage0_22[244], stage0_22[245], stage0_22[246], stage0_22[247], stage0_22[248]},
      {stage1_24[46],stage1_23[87],stage1_22[87],stage1_21[119],stage1_20[190]}
   );
   gpc606_5 gpc823 (
      {stage0_20[302], stage0_20[303], stage0_20[304], stage0_20[305], stage0_20[306], stage0_20[307]},
      {stage0_22[249], stage0_22[250], stage0_22[251], stage0_22[252], stage0_22[253], stage0_22[254]},
      {stage1_24[47],stage1_23[88],stage1_22[88],stage1_21[120],stage1_20[191]}
   );
   gpc606_5 gpc824 (
      {stage0_20[308], stage0_20[309], stage0_20[310], stage0_20[311], stage0_20[312], stage0_20[313]},
      {stage0_22[255], stage0_22[256], stage0_22[257], stage0_22[258], stage0_22[259], stage0_22[260]},
      {stage1_24[48],stage1_23[89],stage1_22[89],stage1_21[121],stage1_20[192]}
   );
   gpc606_5 gpc825 (
      {stage0_20[314], stage0_20[315], stage0_20[316], stage0_20[317], stage0_20[318], stage0_20[319]},
      {stage0_22[261], stage0_22[262], stage0_22[263], stage0_22[264], stage0_22[265], stage0_22[266]},
      {stage1_24[49],stage1_23[90],stage1_22[90],stage1_21[122],stage1_20[193]}
   );
   gpc606_5 gpc826 (
      {stage0_20[320], stage0_20[321], stage0_20[322], stage0_20[323], stage0_20[324], stage0_20[325]},
      {stage0_22[267], stage0_22[268], stage0_22[269], stage0_22[270], stage0_22[271], stage0_22[272]},
      {stage1_24[50],stage1_23[91],stage1_22[91],stage1_21[123],stage1_20[194]}
   );
   gpc606_5 gpc827 (
      {stage0_20[326], stage0_20[327], stage0_20[328], stage0_20[329], stage0_20[330], stage0_20[331]},
      {stage0_22[273], stage0_22[274], stage0_22[275], stage0_22[276], stage0_22[277], stage0_22[278]},
      {stage1_24[51],stage1_23[92],stage1_22[92],stage1_21[124],stage1_20[195]}
   );
   gpc606_5 gpc828 (
      {stage0_20[332], stage0_20[333], stage0_20[334], stage0_20[335], stage0_20[336], stage0_20[337]},
      {stage0_22[279], stage0_22[280], stage0_22[281], stage0_22[282], stage0_22[283], stage0_22[284]},
      {stage1_24[52],stage1_23[93],stage1_22[93],stage1_21[125],stage1_20[196]}
   );
   gpc606_5 gpc829 (
      {stage0_20[338], stage0_20[339], stage0_20[340], stage0_20[341], stage0_20[342], stage0_20[343]},
      {stage0_22[285], stage0_22[286], stage0_22[287], stage0_22[288], stage0_22[289], stage0_22[290]},
      {stage1_24[53],stage1_23[94],stage1_22[94],stage1_21[126],stage1_20[197]}
   );
   gpc606_5 gpc830 (
      {stage0_20[344], stage0_20[345], stage0_20[346], stage0_20[347], stage0_20[348], stage0_20[349]},
      {stage0_22[291], stage0_22[292], stage0_22[293], stage0_22[294], stage0_22[295], stage0_22[296]},
      {stage1_24[54],stage1_23[95],stage1_22[95],stage1_21[127],stage1_20[198]}
   );
   gpc606_5 gpc831 (
      {stage0_20[350], stage0_20[351], stage0_20[352], stage0_20[353], stage0_20[354], stage0_20[355]},
      {stage0_22[297], stage0_22[298], stage0_22[299], stage0_22[300], stage0_22[301], stage0_22[302]},
      {stage1_24[55],stage1_23[96],stage1_22[96],stage1_21[128],stage1_20[199]}
   );
   gpc606_5 gpc832 (
      {stage0_20[356], stage0_20[357], stage0_20[358], stage0_20[359], stage0_20[360], stage0_20[361]},
      {stage0_22[303], stage0_22[304], stage0_22[305], stage0_22[306], stage0_22[307], stage0_22[308]},
      {stage1_24[56],stage1_23[97],stage1_22[97],stage1_21[129],stage1_20[200]}
   );
   gpc606_5 gpc833 (
      {stage0_20[362], stage0_20[363], stage0_20[364], stage0_20[365], stage0_20[366], stage0_20[367]},
      {stage0_22[309], stage0_22[310], stage0_22[311], stage0_22[312], stage0_22[313], stage0_22[314]},
      {stage1_24[57],stage1_23[98],stage1_22[98],stage1_21[130],stage1_20[201]}
   );
   gpc606_5 gpc834 (
      {stage0_20[368], stage0_20[369], stage0_20[370], stage0_20[371], stage0_20[372], stage0_20[373]},
      {stage0_22[315], stage0_22[316], stage0_22[317], stage0_22[318], stage0_22[319], stage0_22[320]},
      {stage1_24[58],stage1_23[99],stage1_22[99],stage1_21[131],stage1_20[202]}
   );
   gpc606_5 gpc835 (
      {stage0_20[374], stage0_20[375], stage0_20[376], stage0_20[377], stage0_20[378], stage0_20[379]},
      {stage0_22[321], stage0_22[322], stage0_22[323], stage0_22[324], stage0_22[325], stage0_22[326]},
      {stage1_24[59],stage1_23[100],stage1_22[100],stage1_21[132],stage1_20[203]}
   );
   gpc606_5 gpc836 (
      {stage0_20[380], stage0_20[381], stage0_20[382], stage0_20[383], stage0_20[384], stage0_20[385]},
      {stage0_22[327], stage0_22[328], stage0_22[329], stage0_22[330], stage0_22[331], stage0_22[332]},
      {stage1_24[60],stage1_23[101],stage1_22[101],stage1_21[133],stage1_20[204]}
   );
   gpc606_5 gpc837 (
      {stage0_20[386], stage0_20[387], stage0_20[388], stage0_20[389], stage0_20[390], stage0_20[391]},
      {stage0_22[333], stage0_22[334], stage0_22[335], stage0_22[336], stage0_22[337], stage0_22[338]},
      {stage1_24[61],stage1_23[102],stage1_22[102],stage1_21[134],stage1_20[205]}
   );
   gpc615_5 gpc838 (
      {stage0_20[392], stage0_20[393], stage0_20[394], stage0_20[395], stage0_20[396]},
      {stage0_21[286]},
      {stage0_22[339], stage0_22[340], stage0_22[341], stage0_22[342], stage0_22[343], stage0_22[344]},
      {stage1_24[62],stage1_23[103],stage1_22[103],stage1_21[135],stage1_20[206]}
   );
   gpc615_5 gpc839 (
      {stage0_20[397], stage0_20[398], stage0_20[399], stage0_20[400], stage0_20[401]},
      {stage0_21[287]},
      {stage0_22[345], stage0_22[346], stage0_22[347], stage0_22[348], stage0_22[349], stage0_22[350]},
      {stage1_24[63],stage1_23[104],stage1_22[104],stage1_21[136],stage1_20[207]}
   );
   gpc615_5 gpc840 (
      {stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405], stage0_20[406]},
      {stage0_21[288]},
      {stage0_22[351], stage0_22[352], stage0_22[353], stage0_22[354], stage0_22[355], stage0_22[356]},
      {stage1_24[64],stage1_23[105],stage1_22[105],stage1_21[137],stage1_20[208]}
   );
   gpc615_5 gpc841 (
      {stage0_20[407], stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411]},
      {stage0_21[289]},
      {stage0_22[357], stage0_22[358], stage0_22[359], stage0_22[360], stage0_22[361], stage0_22[362]},
      {stage1_24[65],stage1_23[106],stage1_22[106],stage1_21[138],stage1_20[209]}
   );
   gpc615_5 gpc842 (
      {stage0_20[412], stage0_20[413], stage0_20[414], stage0_20[415], stage0_20[416]},
      {stage0_21[290]},
      {stage0_22[363], stage0_22[364], stage0_22[365], stage0_22[366], stage0_22[367], stage0_22[368]},
      {stage1_24[66],stage1_23[107],stage1_22[107],stage1_21[139],stage1_20[210]}
   );
   gpc615_5 gpc843 (
      {stage0_20[417], stage0_20[418], stage0_20[419], stage0_20[420], stage0_20[421]},
      {stage0_21[291]},
      {stage0_22[369], stage0_22[370], stage0_22[371], stage0_22[372], stage0_22[373], stage0_22[374]},
      {stage1_24[67],stage1_23[108],stage1_22[108],stage1_21[140],stage1_20[211]}
   );
   gpc615_5 gpc844 (
      {stage0_20[422], stage0_20[423], stage0_20[424], stage0_20[425], stage0_20[426]},
      {stage0_21[292]},
      {stage0_22[375], stage0_22[376], stage0_22[377], stage0_22[378], stage0_22[379], stage0_22[380]},
      {stage1_24[68],stage1_23[109],stage1_22[109],stage1_21[141],stage1_20[212]}
   );
   gpc615_5 gpc845 (
      {stage0_20[427], stage0_20[428], stage0_20[429], stage0_20[430], stage0_20[431]},
      {stage0_21[293]},
      {stage0_22[381], stage0_22[382], stage0_22[383], stage0_22[384], stage0_22[385], stage0_22[386]},
      {stage1_24[69],stage1_23[110],stage1_22[110],stage1_21[142],stage1_20[213]}
   );
   gpc606_5 gpc846 (
      {stage0_21[294], stage0_21[295], stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299]},
      {stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11], stage0_23[12]},
      {stage1_25[0],stage1_24[70],stage1_23[111],stage1_22[111],stage1_21[143]}
   );
   gpc606_5 gpc847 (
      {stage0_21[300], stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17], stage0_23[18]},
      {stage1_25[1],stage1_24[71],stage1_23[112],stage1_22[112],stage1_21[144]}
   );
   gpc606_5 gpc848 (
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310], stage0_21[311]},
      {stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23], stage0_23[24]},
      {stage1_25[2],stage1_24[72],stage1_23[113],stage1_22[113],stage1_21[145]}
   );
   gpc606_5 gpc849 (
      {stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315], stage0_21[316], stage0_21[317]},
      {stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29], stage0_23[30]},
      {stage1_25[3],stage1_24[73],stage1_23[114],stage1_22[114],stage1_21[146]}
   );
   gpc606_5 gpc850 (
      {stage0_21[318], stage0_21[319], stage0_21[320], stage0_21[321], stage0_21[322], stage0_21[323]},
      {stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35], stage0_23[36]},
      {stage1_25[4],stage1_24[74],stage1_23[115],stage1_22[115],stage1_21[147]}
   );
   gpc606_5 gpc851 (
      {stage0_21[324], stage0_21[325], stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329]},
      {stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41], stage0_23[42]},
      {stage1_25[5],stage1_24[75],stage1_23[116],stage1_22[116],stage1_21[148]}
   );
   gpc606_5 gpc852 (
      {stage0_21[330], stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47], stage0_23[48]},
      {stage1_25[6],stage1_24[76],stage1_23[117],stage1_22[117],stage1_21[149]}
   );
   gpc606_5 gpc853 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340], stage0_21[341]},
      {stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53], stage0_23[54]},
      {stage1_25[7],stage1_24[77],stage1_23[118],stage1_22[118],stage1_21[150]}
   );
   gpc606_5 gpc854 (
      {stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345], stage0_21[346], stage0_21[347]},
      {stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59], stage0_23[60]},
      {stage1_25[8],stage1_24[78],stage1_23[119],stage1_22[119],stage1_21[151]}
   );
   gpc606_5 gpc855 (
      {stage0_21[348], stage0_21[349], stage0_21[350], stage0_21[351], stage0_21[352], stage0_21[353]},
      {stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65], stage0_23[66]},
      {stage1_25[9],stage1_24[79],stage1_23[120],stage1_22[120],stage1_21[152]}
   );
   gpc606_5 gpc856 (
      {stage0_21[354], stage0_21[355], stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359]},
      {stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71], stage0_23[72]},
      {stage1_25[10],stage1_24[80],stage1_23[121],stage1_22[121],stage1_21[153]}
   );
   gpc606_5 gpc857 (
      {stage0_21[360], stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77], stage0_23[78]},
      {stage1_25[11],stage1_24[81],stage1_23[122],stage1_22[122],stage1_21[154]}
   );
   gpc606_5 gpc858 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370], stage0_21[371]},
      {stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83], stage0_23[84]},
      {stage1_25[12],stage1_24[82],stage1_23[123],stage1_22[123],stage1_21[155]}
   );
   gpc606_5 gpc859 (
      {stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375], stage0_21[376], stage0_21[377]},
      {stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89], stage0_23[90]},
      {stage1_25[13],stage1_24[83],stage1_23[124],stage1_22[124],stage1_21[156]}
   );
   gpc606_5 gpc860 (
      {stage0_21[378], stage0_21[379], stage0_21[380], stage0_21[381], stage0_21[382], stage0_21[383]},
      {stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95], stage0_23[96]},
      {stage1_25[14],stage1_24[84],stage1_23[125],stage1_22[125],stage1_21[157]}
   );
   gpc606_5 gpc861 (
      {stage0_21[384], stage0_21[385], stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389]},
      {stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101], stage0_23[102]},
      {stage1_25[15],stage1_24[85],stage1_23[126],stage1_22[126],stage1_21[158]}
   );
   gpc606_5 gpc862 (
      {stage0_21[390], stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107], stage0_23[108]},
      {stage1_25[16],stage1_24[86],stage1_23[127],stage1_22[127],stage1_21[159]}
   );
   gpc606_5 gpc863 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400], stage0_21[401]},
      {stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113], stage0_23[114]},
      {stage1_25[17],stage1_24[87],stage1_23[128],stage1_22[128],stage1_21[160]}
   );
   gpc606_5 gpc864 (
      {stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405], stage0_21[406], stage0_21[407]},
      {stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120]},
      {stage1_25[18],stage1_24[88],stage1_23[129],stage1_22[129],stage1_21[161]}
   );
   gpc606_5 gpc865 (
      {stage0_21[408], stage0_21[409], stage0_21[410], stage0_21[411], stage0_21[412], stage0_21[413]},
      {stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125], stage0_23[126]},
      {stage1_25[19],stage1_24[89],stage1_23[130],stage1_22[130],stage1_21[162]}
   );
   gpc606_5 gpc866 (
      {stage0_21[414], stage0_21[415], stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419]},
      {stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131], stage0_23[132]},
      {stage1_25[20],stage1_24[90],stage1_23[131],stage1_22[131],stage1_21[163]}
   );
   gpc606_5 gpc867 (
      {stage0_21[420], stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137], stage0_23[138]},
      {stage1_25[21],stage1_24[91],stage1_23[132],stage1_22[132],stage1_21[164]}
   );
   gpc606_5 gpc868 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430], stage0_21[431]},
      {stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143], stage0_23[144]},
      {stage1_25[22],stage1_24[92],stage1_23[133],stage1_22[133],stage1_21[165]}
   );
   gpc606_5 gpc869 (
      {stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435], stage0_21[436], stage0_21[437]},
      {stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149], stage0_23[150]},
      {stage1_25[23],stage1_24[93],stage1_23[134],stage1_22[134],stage1_21[166]}
   );
   gpc606_5 gpc870 (
      {stage0_21[438], stage0_21[439], stage0_21[440], stage0_21[441], stage0_21[442], stage0_21[443]},
      {stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155], stage0_23[156]},
      {stage1_25[24],stage1_24[94],stage1_23[135],stage1_22[135],stage1_21[167]}
   );
   gpc606_5 gpc871 (
      {stage0_21[444], stage0_21[445], stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449]},
      {stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161], stage0_23[162]},
      {stage1_25[25],stage1_24[95],stage1_23[136],stage1_22[136],stage1_21[168]}
   );
   gpc606_5 gpc872 (
      {stage0_21[450], stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167], stage0_23[168]},
      {stage1_25[26],stage1_24[96],stage1_23[137],stage1_22[137],stage1_21[169]}
   );
   gpc606_5 gpc873 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460], stage0_21[461]},
      {stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173], stage0_23[174]},
      {stage1_25[27],stage1_24[97],stage1_23[138],stage1_22[138],stage1_21[170]}
   );
   gpc606_5 gpc874 (
      {stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465], stage0_21[466], stage0_21[467]},
      {stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179], stage0_23[180]},
      {stage1_25[28],stage1_24[98],stage1_23[139],stage1_22[139],stage1_21[171]}
   );
   gpc615_5 gpc875 (
      {stage0_22[387], stage0_22[388], stage0_22[389], stage0_22[390], stage0_22[391]},
      {stage0_23[181]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[29],stage1_24[99],stage1_23[140],stage1_22[140]}
   );
   gpc615_5 gpc876 (
      {stage0_22[392], stage0_22[393], stage0_22[394], stage0_22[395], stage0_22[396]},
      {stage0_23[182]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[30],stage1_24[100],stage1_23[141],stage1_22[141]}
   );
   gpc615_5 gpc877 (
      {stage0_22[397], stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401]},
      {stage0_23[183]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[31],stage1_24[101],stage1_23[142],stage1_22[142]}
   );
   gpc615_5 gpc878 (
      {stage0_22[402], stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406]},
      {stage0_23[184]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[32],stage1_24[102],stage1_23[143],stage1_22[143]}
   );
   gpc615_5 gpc879 (
      {stage0_22[407], stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411]},
      {stage0_23[185]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[33],stage1_24[103],stage1_23[144],stage1_22[144]}
   );
   gpc615_5 gpc880 (
      {stage0_22[412], stage0_22[413], stage0_22[414], stage0_22[415], stage0_22[416]},
      {stage0_23[186]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[34],stage1_24[104],stage1_23[145],stage1_22[145]}
   );
   gpc615_5 gpc881 (
      {stage0_22[417], stage0_22[418], stage0_22[419], stage0_22[420], stage0_22[421]},
      {stage0_23[187]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[35],stage1_24[105],stage1_23[146],stage1_22[146]}
   );
   gpc615_5 gpc882 (
      {stage0_22[422], stage0_22[423], stage0_22[424], stage0_22[425], stage0_22[426]},
      {stage0_23[188]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[36],stage1_24[106],stage1_23[147],stage1_22[147]}
   );
   gpc615_5 gpc883 (
      {stage0_22[427], stage0_22[428], stage0_22[429], stage0_22[430], stage0_22[431]},
      {stage0_23[189]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[37],stage1_24[107],stage1_23[148],stage1_22[148]}
   );
   gpc615_5 gpc884 (
      {stage0_22[432], stage0_22[433], stage0_22[434], stage0_22[435], stage0_22[436]},
      {stage0_23[190]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[38],stage1_24[108],stage1_23[149],stage1_22[149]}
   );
   gpc615_5 gpc885 (
      {stage0_22[437], stage0_22[438], stage0_22[439], stage0_22[440], stage0_22[441]},
      {stage0_23[191]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[39],stage1_24[109],stage1_23[150],stage1_22[150]}
   );
   gpc615_5 gpc886 (
      {stage0_22[442], stage0_22[443], stage0_22[444], stage0_22[445], stage0_22[446]},
      {stage0_23[192]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[40],stage1_24[110],stage1_23[151],stage1_22[151]}
   );
   gpc615_5 gpc887 (
      {stage0_22[447], stage0_22[448], stage0_22[449], stage0_22[450], stage0_22[451]},
      {stage0_23[193]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[41],stage1_24[111],stage1_23[152],stage1_22[152]}
   );
   gpc615_5 gpc888 (
      {stage0_22[452], stage0_22[453], stage0_22[454], stage0_22[455], stage0_22[456]},
      {stage0_23[194]},
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage1_26[13],stage1_25[42],stage1_24[112],stage1_23[153],stage1_22[153]}
   );
   gpc615_5 gpc889 (
      {stage0_22[457], stage0_22[458], stage0_22[459], stage0_22[460], stage0_22[461]},
      {stage0_23[195]},
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage1_26[14],stage1_25[43],stage1_24[113],stage1_23[154],stage1_22[154]}
   );
   gpc615_5 gpc890 (
      {stage0_22[462], stage0_22[463], stage0_22[464], stage0_22[465], stage0_22[466]},
      {stage0_23[196]},
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage1_26[15],stage1_25[44],stage1_24[114],stage1_23[155],stage1_22[155]}
   );
   gpc615_5 gpc891 (
      {stage0_22[467], stage0_22[468], stage0_22[469], stage0_22[470], stage0_22[471]},
      {stage0_23[197]},
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage1_26[16],stage1_25[45],stage1_24[115],stage1_23[156],stage1_22[156]}
   );
   gpc615_5 gpc892 (
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202]},
      {stage0_24[102]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[17],stage1_25[46],stage1_24[116],stage1_23[157]}
   );
   gpc615_5 gpc893 (
      {stage0_23[203], stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207]},
      {stage0_24[103]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[18],stage1_25[47],stage1_24[117],stage1_23[158]}
   );
   gpc615_5 gpc894 (
      {stage0_23[208], stage0_23[209], stage0_23[210], stage0_23[211], stage0_23[212]},
      {stage0_24[104]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[19],stage1_25[48],stage1_24[118],stage1_23[159]}
   );
   gpc615_5 gpc895 (
      {stage0_23[213], stage0_23[214], stage0_23[215], stage0_23[216], stage0_23[217]},
      {stage0_24[105]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[20],stage1_25[49],stage1_24[119],stage1_23[160]}
   );
   gpc615_5 gpc896 (
      {stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221], stage0_23[222]},
      {stage0_24[106]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[21],stage1_25[50],stage1_24[120],stage1_23[161]}
   );
   gpc615_5 gpc897 (
      {stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage0_24[107]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[22],stage1_25[51],stage1_24[121],stage1_23[162]}
   );
   gpc615_5 gpc898 (
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232]},
      {stage0_24[108]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[23],stage1_25[52],stage1_24[122],stage1_23[163]}
   );
   gpc615_5 gpc899 (
      {stage0_23[233], stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237]},
      {stage0_24[109]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[24],stage1_25[53],stage1_24[123],stage1_23[164]}
   );
   gpc615_5 gpc900 (
      {stage0_23[238], stage0_23[239], stage0_23[240], stage0_23[241], stage0_23[242]},
      {stage0_24[110]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[25],stage1_25[54],stage1_24[124],stage1_23[165]}
   );
   gpc615_5 gpc901 (
      {stage0_23[243], stage0_23[244], stage0_23[245], stage0_23[246], stage0_23[247]},
      {stage0_24[111]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[26],stage1_25[55],stage1_24[125],stage1_23[166]}
   );
   gpc615_5 gpc902 (
      {stage0_23[248], stage0_23[249], stage0_23[250], stage0_23[251], stage0_23[252]},
      {stage0_24[112]},
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage1_27[10],stage1_26[27],stage1_25[56],stage1_24[126],stage1_23[167]}
   );
   gpc615_5 gpc903 (
      {stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256], stage0_23[257]},
      {stage0_24[113]},
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage1_27[11],stage1_26[28],stage1_25[57],stage1_24[127],stage1_23[168]}
   );
   gpc615_5 gpc904 (
      {stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262]},
      {stage0_24[114]},
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage1_27[12],stage1_26[29],stage1_25[58],stage1_24[128],stage1_23[169]}
   );
   gpc615_5 gpc905 (
      {stage0_23[263], stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267]},
      {stage0_24[115]},
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage1_27[13],stage1_26[30],stage1_25[59],stage1_24[129],stage1_23[170]}
   );
   gpc615_5 gpc906 (
      {stage0_23[268], stage0_23[269], stage0_23[270], stage0_23[271], stage0_23[272]},
      {stage0_24[116]},
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage1_27[14],stage1_26[31],stage1_25[60],stage1_24[130],stage1_23[171]}
   );
   gpc615_5 gpc907 (
      {stage0_23[273], stage0_23[274], stage0_23[275], stage0_23[276], stage0_23[277]},
      {stage0_24[117]},
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage1_27[15],stage1_26[32],stage1_25[61],stage1_24[131],stage1_23[172]}
   );
   gpc615_5 gpc908 (
      {stage0_23[278], stage0_23[279], stage0_23[280], stage0_23[281], stage0_23[282]},
      {stage0_24[118]},
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage1_27[16],stage1_26[33],stage1_25[62],stage1_24[132],stage1_23[173]}
   );
   gpc615_5 gpc909 (
      {stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286], stage0_23[287]},
      {stage0_24[119]},
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage1_27[17],stage1_26[34],stage1_25[63],stage1_24[133],stage1_23[174]}
   );
   gpc615_5 gpc910 (
      {stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292]},
      {stage0_24[120]},
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage1_27[18],stage1_26[35],stage1_25[64],stage1_24[134],stage1_23[175]}
   );
   gpc615_5 gpc911 (
      {stage0_23[293], stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297]},
      {stage0_24[121]},
      {stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119]},
      {stage1_27[19],stage1_26[36],stage1_25[65],stage1_24[135],stage1_23[176]}
   );
   gpc615_5 gpc912 (
      {stage0_23[298], stage0_23[299], stage0_23[300], stage0_23[301], stage0_23[302]},
      {stage0_24[122]},
      {stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125]},
      {stage1_27[20],stage1_26[37],stage1_25[66],stage1_24[136],stage1_23[177]}
   );
   gpc615_5 gpc913 (
      {stage0_23[303], stage0_23[304], stage0_23[305], stage0_23[306], stage0_23[307]},
      {stage0_24[123]},
      {stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131]},
      {stage1_27[21],stage1_26[38],stage1_25[67],stage1_24[137],stage1_23[178]}
   );
   gpc615_5 gpc914 (
      {stage0_23[308], stage0_23[309], stage0_23[310], stage0_23[311], stage0_23[312]},
      {stage0_24[124]},
      {stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage1_27[22],stage1_26[39],stage1_25[68],stage1_24[138],stage1_23[179]}
   );
   gpc615_5 gpc915 (
      {stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316], stage0_23[317]},
      {stage0_24[125]},
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143]},
      {stage1_27[23],stage1_26[40],stage1_25[69],stage1_24[139],stage1_23[180]}
   );
   gpc615_5 gpc916 (
      {stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322]},
      {stage0_24[126]},
      {stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149]},
      {stage1_27[24],stage1_26[41],stage1_25[70],stage1_24[140],stage1_23[181]}
   );
   gpc615_5 gpc917 (
      {stage0_23[323], stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327]},
      {stage0_24[127]},
      {stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155]},
      {stage1_27[25],stage1_26[42],stage1_25[71],stage1_24[141],stage1_23[182]}
   );
   gpc615_5 gpc918 (
      {stage0_23[328], stage0_23[329], stage0_23[330], stage0_23[331], stage0_23[332]},
      {stage0_24[128]},
      {stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161]},
      {stage1_27[26],stage1_26[43],stage1_25[72],stage1_24[142],stage1_23[183]}
   );
   gpc615_5 gpc919 (
      {stage0_23[333], stage0_23[334], stage0_23[335], stage0_23[336], stage0_23[337]},
      {stage0_24[129]},
      {stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167]},
      {stage1_27[27],stage1_26[44],stage1_25[73],stage1_24[143],stage1_23[184]}
   );
   gpc615_5 gpc920 (
      {stage0_23[338], stage0_23[339], stage0_23[340], stage0_23[341], stage0_23[342]},
      {stage0_24[130]},
      {stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173]},
      {stage1_27[28],stage1_26[45],stage1_25[74],stage1_24[144],stage1_23[185]}
   );
   gpc615_5 gpc921 (
      {stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346], stage0_23[347]},
      {stage0_24[131]},
      {stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179]},
      {stage1_27[29],stage1_26[46],stage1_25[75],stage1_24[145],stage1_23[186]}
   );
   gpc615_5 gpc922 (
      {stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352]},
      {stage0_24[132]},
      {stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185]},
      {stage1_27[30],stage1_26[47],stage1_25[76],stage1_24[146],stage1_23[187]}
   );
   gpc615_5 gpc923 (
      {stage0_23[353], stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357]},
      {stage0_24[133]},
      {stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191]},
      {stage1_27[31],stage1_26[48],stage1_25[77],stage1_24[147],stage1_23[188]}
   );
   gpc615_5 gpc924 (
      {stage0_23[358], stage0_23[359], stage0_23[360], stage0_23[361], stage0_23[362]},
      {stage0_24[134]},
      {stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197]},
      {stage1_27[32],stage1_26[49],stage1_25[78],stage1_24[148],stage1_23[189]}
   );
   gpc615_5 gpc925 (
      {stage0_23[363], stage0_23[364], stage0_23[365], stage0_23[366], stage0_23[367]},
      {stage0_24[135]},
      {stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203]},
      {stage1_27[33],stage1_26[50],stage1_25[79],stage1_24[149],stage1_23[190]}
   );
   gpc615_5 gpc926 (
      {stage0_23[368], stage0_23[369], stage0_23[370], stage0_23[371], stage0_23[372]},
      {stage0_24[136]},
      {stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209]},
      {stage1_27[34],stage1_26[51],stage1_25[80],stage1_24[150],stage1_23[191]}
   );
   gpc615_5 gpc927 (
      {stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376], stage0_23[377]},
      {stage0_24[137]},
      {stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215]},
      {stage1_27[35],stage1_26[52],stage1_25[81],stage1_24[151],stage1_23[192]}
   );
   gpc615_5 gpc928 (
      {stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382]},
      {stage0_24[138]},
      {stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221]},
      {stage1_27[36],stage1_26[53],stage1_25[82],stage1_24[152],stage1_23[193]}
   );
   gpc615_5 gpc929 (
      {stage0_23[383], stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387]},
      {stage0_24[139]},
      {stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225], stage0_25[226], stage0_25[227]},
      {stage1_27[37],stage1_26[54],stage1_25[83],stage1_24[153],stage1_23[194]}
   );
   gpc615_5 gpc930 (
      {stage0_23[388], stage0_23[389], stage0_23[390], stage0_23[391], stage0_23[392]},
      {stage0_24[140]},
      {stage0_25[228], stage0_25[229], stage0_25[230], stage0_25[231], stage0_25[232], stage0_25[233]},
      {stage1_27[38],stage1_26[55],stage1_25[84],stage1_24[154],stage1_23[195]}
   );
   gpc623_5 gpc931 (
      {stage0_23[393], stage0_23[394], stage0_23[395]},
      {stage0_24[141], stage0_24[142]},
      {stage0_25[234], stage0_25[235], stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239]},
      {stage1_27[39],stage1_26[56],stage1_25[85],stage1_24[155],stage1_23[196]}
   );
   gpc606_5 gpc932 (
      {stage0_24[143], stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[40],stage1_26[57],stage1_25[86],stage1_24[156]}
   );
   gpc606_5 gpc933 (
      {stage0_24[149], stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[41],stage1_26[58],stage1_25[87],stage1_24[157]}
   );
   gpc606_5 gpc934 (
      {stage0_24[155], stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[42],stage1_26[59],stage1_25[88],stage1_24[158]}
   );
   gpc606_5 gpc935 (
      {stage0_24[161], stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165], stage0_24[166]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[43],stage1_26[60],stage1_25[89],stage1_24[159]}
   );
   gpc606_5 gpc936 (
      {stage0_24[167], stage0_24[168], stage0_24[169], stage0_24[170], stage0_24[171], stage0_24[172]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[44],stage1_26[61],stage1_25[90],stage1_24[160]}
   );
   gpc606_5 gpc937 (
      {stage0_24[173], stage0_24[174], stage0_24[175], stage0_24[176], stage0_24[177], stage0_24[178]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[45],stage1_26[62],stage1_25[91],stage1_24[161]}
   );
   gpc606_5 gpc938 (
      {stage0_24[179], stage0_24[180], stage0_24[181], stage0_24[182], stage0_24[183], stage0_24[184]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[46],stage1_26[63],stage1_25[92],stage1_24[162]}
   );
   gpc606_5 gpc939 (
      {stage0_24[185], stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189], stage0_24[190]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[47],stage1_26[64],stage1_25[93],stage1_24[163]}
   );
   gpc606_5 gpc940 (
      {stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195], stage0_24[196]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[48],stage1_26[65],stage1_25[94],stage1_24[164]}
   );
   gpc606_5 gpc941 (
      {stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200], stage0_24[201], stage0_24[202]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[49],stage1_26[66],stage1_25[95],stage1_24[165]}
   );
   gpc606_5 gpc942 (
      {stage0_24[203], stage0_24[204], stage0_24[205], stage0_24[206], stage0_24[207], stage0_24[208]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[50],stage1_26[67],stage1_25[96],stage1_24[166]}
   );
   gpc606_5 gpc943 (
      {stage0_24[209], stage0_24[210], stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[51],stage1_26[68],stage1_25[97],stage1_24[167]}
   );
   gpc606_5 gpc944 (
      {stage0_24[215], stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[52],stage1_26[69],stage1_25[98],stage1_24[168]}
   );
   gpc606_5 gpc945 (
      {stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225], stage0_24[226]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[53],stage1_26[70],stage1_25[99],stage1_24[169]}
   );
   gpc606_5 gpc946 (
      {stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230], stage0_24[231], stage0_24[232]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[54],stage1_26[71],stage1_25[100],stage1_24[170]}
   );
   gpc606_5 gpc947 (
      {stage0_24[233], stage0_24[234], stage0_24[235], stage0_24[236], stage0_24[237], stage0_24[238]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[55],stage1_26[72],stage1_25[101],stage1_24[171]}
   );
   gpc606_5 gpc948 (
      {stage0_24[239], stage0_24[240], stage0_24[241], stage0_24[242], stage0_24[243], stage0_24[244]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[56],stage1_26[73],stage1_25[102],stage1_24[172]}
   );
   gpc606_5 gpc949 (
      {stage0_24[245], stage0_24[246], stage0_24[247], stage0_24[248], stage0_24[249], stage0_24[250]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[57],stage1_26[74],stage1_25[103],stage1_24[173]}
   );
   gpc606_5 gpc950 (
      {stage0_24[251], stage0_24[252], stage0_24[253], stage0_24[254], stage0_24[255], stage0_24[256]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[58],stage1_26[75],stage1_25[104],stage1_24[174]}
   );
   gpc606_5 gpc951 (
      {stage0_24[257], stage0_24[258], stage0_24[259], stage0_24[260], stage0_24[261], stage0_24[262]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[59],stage1_26[76],stage1_25[105],stage1_24[175]}
   );
   gpc606_5 gpc952 (
      {stage0_24[263], stage0_24[264], stage0_24[265], stage0_24[266], stage0_24[267], stage0_24[268]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[60],stage1_26[77],stage1_25[106],stage1_24[176]}
   );
   gpc606_5 gpc953 (
      {stage0_24[269], stage0_24[270], stage0_24[271], stage0_24[272], stage0_24[273], stage0_24[274]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[61],stage1_26[78],stage1_25[107],stage1_24[177]}
   );
   gpc606_5 gpc954 (
      {stage0_24[275], stage0_24[276], stage0_24[277], stage0_24[278], stage0_24[279], stage0_24[280]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[62],stage1_26[79],stage1_25[108],stage1_24[178]}
   );
   gpc606_5 gpc955 (
      {stage0_24[281], stage0_24[282], stage0_24[283], stage0_24[284], stage0_24[285], stage0_24[286]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[63],stage1_26[80],stage1_25[109],stage1_24[179]}
   );
   gpc606_5 gpc956 (
      {stage0_24[287], stage0_24[288], stage0_24[289], stage0_24[290], stage0_24[291], stage0_24[292]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[64],stage1_26[81],stage1_25[110],stage1_24[180]}
   );
   gpc606_5 gpc957 (
      {stage0_24[293], stage0_24[294], stage0_24[295], stage0_24[296], stage0_24[297], stage0_24[298]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[65],stage1_26[82],stage1_25[111],stage1_24[181]}
   );
   gpc606_5 gpc958 (
      {stage0_24[299], stage0_24[300], stage0_24[301], stage0_24[302], stage0_24[303], stage0_24[304]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[66],stage1_26[83],stage1_25[112],stage1_24[182]}
   );
   gpc606_5 gpc959 (
      {stage0_24[305], stage0_24[306], stage0_24[307], stage0_24[308], stage0_24[309], stage0_24[310]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[67],stage1_26[84],stage1_25[113],stage1_24[183]}
   );
   gpc606_5 gpc960 (
      {stage0_24[311], stage0_24[312], stage0_24[313], stage0_24[314], stage0_24[315], stage0_24[316]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[68],stage1_26[85],stage1_25[114],stage1_24[184]}
   );
   gpc606_5 gpc961 (
      {stage0_24[317], stage0_24[318], stage0_24[319], stage0_24[320], stage0_24[321], stage0_24[322]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[69],stage1_26[86],stage1_25[115],stage1_24[185]}
   );
   gpc606_5 gpc962 (
      {stage0_24[323], stage0_24[324], stage0_24[325], stage0_24[326], stage0_24[327], stage0_24[328]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[70],stage1_26[87],stage1_25[116],stage1_24[186]}
   );
   gpc606_5 gpc963 (
      {stage0_24[329], stage0_24[330], stage0_24[331], stage0_24[332], stage0_24[333], stage0_24[334]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[71],stage1_26[88],stage1_25[117],stage1_24[187]}
   );
   gpc606_5 gpc964 (
      {stage0_24[335], stage0_24[336], stage0_24[337], stage0_24[338], stage0_24[339], stage0_24[340]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[72],stage1_26[89],stage1_25[118],stage1_24[188]}
   );
   gpc606_5 gpc965 (
      {stage0_24[341], stage0_24[342], stage0_24[343], stage0_24[344], stage0_24[345], stage0_24[346]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[73],stage1_26[90],stage1_25[119],stage1_24[189]}
   );
   gpc606_5 gpc966 (
      {stage0_24[347], stage0_24[348], stage0_24[349], stage0_24[350], stage0_24[351], stage0_24[352]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[74],stage1_26[91],stage1_25[120],stage1_24[190]}
   );
   gpc606_5 gpc967 (
      {stage0_24[353], stage0_24[354], stage0_24[355], stage0_24[356], stage0_24[357], stage0_24[358]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[75],stage1_26[92],stage1_25[121],stage1_24[191]}
   );
   gpc606_5 gpc968 (
      {stage0_24[359], stage0_24[360], stage0_24[361], stage0_24[362], stage0_24[363], stage0_24[364]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[76],stage1_26[93],stage1_25[122],stage1_24[192]}
   );
   gpc606_5 gpc969 (
      {stage0_24[365], stage0_24[366], stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[77],stage1_26[94],stage1_25[123],stage1_24[193]}
   );
   gpc606_5 gpc970 (
      {stage0_24[371], stage0_24[372], stage0_24[373], stage0_24[374], stage0_24[375], stage0_24[376]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[78],stage1_26[95],stage1_25[124],stage1_24[194]}
   );
   gpc606_5 gpc971 (
      {stage0_24[377], stage0_24[378], stage0_24[379], stage0_24[380], stage0_24[381], stage0_24[382]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[79],stage1_26[96],stage1_25[125],stage1_24[195]}
   );
   gpc606_5 gpc972 (
      {stage0_24[383], stage0_24[384], stage0_24[385], stage0_24[386], stage0_24[387], stage0_24[388]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[80],stage1_26[97],stage1_25[126],stage1_24[196]}
   );
   gpc606_5 gpc973 (
      {stage0_24[389], stage0_24[390], stage0_24[391], stage0_24[392], stage0_24[393], stage0_24[394]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[81],stage1_26[98],stage1_25[127],stage1_24[197]}
   );
   gpc606_5 gpc974 (
      {stage0_24[395], stage0_24[396], stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[82],stage1_26[99],stage1_25[128],stage1_24[198]}
   );
   gpc606_5 gpc975 (
      {stage0_24[401], stage0_24[402], stage0_24[403], stage0_24[404], stage0_24[405], stage0_24[406]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[83],stage1_26[100],stage1_25[129],stage1_24[199]}
   );
   gpc606_5 gpc976 (
      {stage0_24[407], stage0_24[408], stage0_24[409], stage0_24[410], stage0_24[411], stage0_24[412]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[84],stage1_26[101],stage1_25[130],stage1_24[200]}
   );
   gpc606_5 gpc977 (
      {stage0_24[413], stage0_24[414], stage0_24[415], stage0_24[416], stage0_24[417], stage0_24[418]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[85],stage1_26[102],stage1_25[131],stage1_24[201]}
   );
   gpc606_5 gpc978 (
      {stage0_24[419], stage0_24[420], stage0_24[421], stage0_24[422], stage0_24[423], stage0_24[424]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[86],stage1_26[103],stage1_25[132],stage1_24[202]}
   );
   gpc606_5 gpc979 (
      {stage0_24[425], stage0_24[426], stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[87],stage1_26[104],stage1_25[133],stage1_24[203]}
   );
   gpc606_5 gpc980 (
      {stage0_24[431], stage0_24[432], stage0_24[433], stage0_24[434], stage0_24[435], stage0_24[436]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[88],stage1_26[105],stage1_25[134],stage1_24[204]}
   );
   gpc606_5 gpc981 (
      {stage0_24[437], stage0_24[438], stage0_24[439], stage0_24[440], stage0_24[441], stage0_24[442]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[89],stage1_26[106],stage1_25[135],stage1_24[205]}
   );
   gpc606_5 gpc982 (
      {stage0_24[443], stage0_24[444], stage0_24[445], stage0_24[446], stage0_24[447], stage0_24[448]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[90],stage1_26[107],stage1_25[136],stage1_24[206]}
   );
   gpc606_5 gpc983 (
      {stage0_24[449], stage0_24[450], stage0_24[451], stage0_24[452], stage0_24[453], stage0_24[454]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[91],stage1_26[108],stage1_25[137],stage1_24[207]}
   );
   gpc606_5 gpc984 (
      {stage0_24[455], stage0_24[456], stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[92],stage1_26[109],stage1_25[138],stage1_24[208]}
   );
   gpc606_5 gpc985 (
      {stage0_24[461], stage0_24[462], stage0_24[463], stage0_24[464], stage0_24[465], stage0_24[466]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[93],stage1_26[110],stage1_25[139],stage1_24[209]}
   );
   gpc606_5 gpc986 (
      {stage0_24[467], stage0_24[468], stage0_24[469], stage0_24[470], stage0_24[471], stage0_24[472]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[94],stage1_26[111],stage1_25[140],stage1_24[210]}
   );
   gpc606_5 gpc987 (
      {stage0_24[473], stage0_24[474], stage0_24[475], stage0_24[476], stage0_24[477], stage0_24[478]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[95],stage1_26[112],stage1_25[141],stage1_24[211]}
   );
   gpc606_5 gpc988 (
      {stage0_24[479], stage0_24[480], stage0_24[481], stage0_24[482], stage0_24[483], stage0_24[484]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[96],stage1_26[113],stage1_25[142],stage1_24[212]}
   );
   gpc606_5 gpc989 (
      {stage0_25[240], stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[57],stage1_27[97],stage1_26[114],stage1_25[143]}
   );
   gpc606_5 gpc990 (
      {stage0_25[246], stage0_25[247], stage0_25[248], stage0_25[249], stage0_25[250], stage0_25[251]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[58],stage1_27[98],stage1_26[115],stage1_25[144]}
   );
   gpc606_5 gpc991 (
      {stage0_25[252], stage0_25[253], stage0_25[254], stage0_25[255], stage0_25[256], stage0_25[257]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[59],stage1_27[99],stage1_26[116],stage1_25[145]}
   );
   gpc606_5 gpc992 (
      {stage0_25[258], stage0_25[259], stage0_25[260], stage0_25[261], stage0_25[262], stage0_25[263]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[60],stage1_27[100],stage1_26[117],stage1_25[146]}
   );
   gpc606_5 gpc993 (
      {stage0_25[264], stage0_25[265], stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[61],stage1_27[101],stage1_26[118],stage1_25[147]}
   );
   gpc606_5 gpc994 (
      {stage0_25[270], stage0_25[271], stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[62],stage1_27[102],stage1_26[119],stage1_25[148]}
   );
   gpc606_5 gpc995 (
      {stage0_25[276], stage0_25[277], stage0_25[278], stage0_25[279], stage0_25[280], stage0_25[281]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[63],stage1_27[103],stage1_26[120],stage1_25[149]}
   );
   gpc606_5 gpc996 (
      {stage0_25[282], stage0_25[283], stage0_25[284], stage0_25[285], stage0_25[286], stage0_25[287]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[64],stage1_27[104],stage1_26[121],stage1_25[150]}
   );
   gpc606_5 gpc997 (
      {stage0_25[288], stage0_25[289], stage0_25[290], stage0_25[291], stage0_25[292], stage0_25[293]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[65],stage1_27[105],stage1_26[122],stage1_25[151]}
   );
   gpc606_5 gpc998 (
      {stage0_25[294], stage0_25[295], stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[66],stage1_27[106],stage1_26[123],stage1_25[152]}
   );
   gpc606_5 gpc999 (
      {stage0_25[300], stage0_25[301], stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[67],stage1_27[107],stage1_26[124],stage1_25[153]}
   );
   gpc606_5 gpc1000 (
      {stage0_25[306], stage0_25[307], stage0_25[308], stage0_25[309], stage0_25[310], stage0_25[311]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[68],stage1_27[108],stage1_26[125],stage1_25[154]}
   );
   gpc606_5 gpc1001 (
      {stage0_25[312], stage0_25[313], stage0_25[314], stage0_25[315], stage0_25[316], stage0_25[317]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[69],stage1_27[109],stage1_26[126],stage1_25[155]}
   );
   gpc606_5 gpc1002 (
      {stage0_25[318], stage0_25[319], stage0_25[320], stage0_25[321], stage0_25[322], stage0_25[323]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[70],stage1_27[110],stage1_26[127],stage1_25[156]}
   );
   gpc606_5 gpc1003 (
      {stage0_25[324], stage0_25[325], stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[71],stage1_27[111],stage1_26[128],stage1_25[157]}
   );
   gpc606_5 gpc1004 (
      {stage0_25[330], stage0_25[331], stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[72],stage1_27[112],stage1_26[129],stage1_25[158]}
   );
   gpc606_5 gpc1005 (
      {stage0_25[336], stage0_25[337], stage0_25[338], stage0_25[339], stage0_25[340], stage0_25[341]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[73],stage1_27[113],stage1_26[130],stage1_25[159]}
   );
   gpc606_5 gpc1006 (
      {stage0_25[342], stage0_25[343], stage0_25[344], stage0_25[345], stage0_25[346], stage0_25[347]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[74],stage1_27[114],stage1_26[131],stage1_25[160]}
   );
   gpc606_5 gpc1007 (
      {stage0_25[348], stage0_25[349], stage0_25[350], stage0_25[351], stage0_25[352], stage0_25[353]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[75],stage1_27[115],stage1_26[132],stage1_25[161]}
   );
   gpc606_5 gpc1008 (
      {stage0_25[354], stage0_25[355], stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[76],stage1_27[116],stage1_26[133],stage1_25[162]}
   );
   gpc606_5 gpc1009 (
      {stage0_25[360], stage0_25[361], stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[77],stage1_27[117],stage1_26[134],stage1_25[163]}
   );
   gpc606_5 gpc1010 (
      {stage0_25[366], stage0_25[367], stage0_25[368], stage0_25[369], stage0_25[370], stage0_25[371]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[78],stage1_27[118],stage1_26[135],stage1_25[164]}
   );
   gpc606_5 gpc1011 (
      {stage0_25[372], stage0_25[373], stage0_25[374], stage0_25[375], stage0_25[376], stage0_25[377]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[79],stage1_27[119],stage1_26[136],stage1_25[165]}
   );
   gpc606_5 gpc1012 (
      {stage0_25[378], stage0_25[379], stage0_25[380], stage0_25[381], stage0_25[382], stage0_25[383]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[80],stage1_27[120],stage1_26[137],stage1_25[166]}
   );
   gpc606_5 gpc1013 (
      {stage0_25[384], stage0_25[385], stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[81],stage1_27[121],stage1_26[138],stage1_25[167]}
   );
   gpc606_5 gpc1014 (
      {stage0_25[390], stage0_25[391], stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[82],stage1_27[122],stage1_26[139],stage1_25[168]}
   );
   gpc606_5 gpc1015 (
      {stage0_25[396], stage0_25[397], stage0_25[398], stage0_25[399], stage0_25[400], stage0_25[401]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[83],stage1_27[123],stage1_26[140],stage1_25[169]}
   );
   gpc606_5 gpc1016 (
      {stage0_25[402], stage0_25[403], stage0_25[404], stage0_25[405], stage0_25[406], stage0_25[407]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[84],stage1_27[124],stage1_26[141],stage1_25[170]}
   );
   gpc606_5 gpc1017 (
      {stage0_25[408], stage0_25[409], stage0_25[410], stage0_25[411], stage0_25[412], stage0_25[413]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[85],stage1_27[125],stage1_26[142],stage1_25[171]}
   );
   gpc606_5 gpc1018 (
      {stage0_25[414], stage0_25[415], stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[86],stage1_27[126],stage1_26[143],stage1_25[172]}
   );
   gpc606_5 gpc1019 (
      {stage0_25[420], stage0_25[421], stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[87],stage1_27[127],stage1_26[144],stage1_25[173]}
   );
   gpc606_5 gpc1020 (
      {stage0_25[426], stage0_25[427], stage0_25[428], stage0_25[429], stage0_25[430], stage0_25[431]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[88],stage1_27[128],stage1_26[145],stage1_25[174]}
   );
   gpc606_5 gpc1021 (
      {stage0_25[432], stage0_25[433], stage0_25[434], stage0_25[435], stage0_25[436], stage0_25[437]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[89],stage1_27[129],stage1_26[146],stage1_25[175]}
   );
   gpc606_5 gpc1022 (
      {stage0_25[438], stage0_25[439], stage0_25[440], stage0_25[441], stage0_25[442], stage0_25[443]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[90],stage1_27[130],stage1_26[147],stage1_25[176]}
   );
   gpc606_5 gpc1023 (
      {stage0_25[444], stage0_25[445], stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[91],stage1_27[131],stage1_26[148],stage1_25[177]}
   );
   gpc606_5 gpc1024 (
      {stage0_25[450], stage0_25[451], stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[92],stage1_27[132],stage1_26[149],stage1_25[178]}
   );
   gpc606_5 gpc1025 (
      {stage0_25[456], stage0_25[457], stage0_25[458], stage0_25[459], stage0_25[460], stage0_25[461]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[93],stage1_27[133],stage1_26[150],stage1_25[179]}
   );
   gpc606_5 gpc1026 (
      {stage0_25[462], stage0_25[463], stage0_25[464], stage0_25[465], stage0_25[466], stage0_25[467]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[94],stage1_27[134],stage1_26[151],stage1_25[180]}
   );
   gpc606_5 gpc1027 (
      {stage0_25[468], stage0_25[469], stage0_25[470], stage0_25[471], stage0_25[472], stage0_25[473]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[95],stage1_27[135],stage1_26[152],stage1_25[181]}
   );
   gpc606_5 gpc1028 (
      {stage0_25[474], stage0_25[475], stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[96],stage1_27[136],stage1_26[153],stage1_25[182]}
   );
   gpc606_5 gpc1029 (
      {stage0_25[480], stage0_25[481], stage0_25[482], stage0_25[483], stage0_25[484], stage0_25[485]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[97],stage1_27[137],stage1_26[154],stage1_25[183]}
   );
   gpc615_5 gpc1030 (
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346]},
      {stage0_27[246]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[41],stage1_28[98],stage1_27[138],stage1_26[155]}
   );
   gpc615_5 gpc1031 (
      {stage0_26[347], stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351]},
      {stage0_27[247]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[42],stage1_28[99],stage1_27[139],stage1_26[156]}
   );
   gpc615_5 gpc1032 (
      {stage0_26[352], stage0_26[353], stage0_26[354], stage0_26[355], stage0_26[356]},
      {stage0_27[248]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[43],stage1_28[100],stage1_27[140],stage1_26[157]}
   );
   gpc615_5 gpc1033 (
      {stage0_26[357], stage0_26[358], stage0_26[359], stage0_26[360], stage0_26[361]},
      {stage0_27[249]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[44],stage1_28[101],stage1_27[141],stage1_26[158]}
   );
   gpc615_5 gpc1034 (
      {stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365], stage0_26[366]},
      {stage0_27[250]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[45],stage1_28[102],stage1_27[142],stage1_26[159]}
   );
   gpc615_5 gpc1035 (
      {stage0_26[367], stage0_26[368], stage0_26[369], stage0_26[370], stage0_26[371]},
      {stage0_27[251]},
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage1_30[5],stage1_29[46],stage1_28[103],stage1_27[143],stage1_26[160]}
   );
   gpc615_5 gpc1036 (
      {stage0_26[372], stage0_26[373], stage0_26[374], stage0_26[375], stage0_26[376]},
      {stage0_27[252]},
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage1_30[6],stage1_29[47],stage1_28[104],stage1_27[144],stage1_26[161]}
   );
   gpc615_5 gpc1037 (
      {stage0_26[377], stage0_26[378], stage0_26[379], stage0_26[380], stage0_26[381]},
      {stage0_27[253]},
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage1_30[7],stage1_29[48],stage1_28[105],stage1_27[145],stage1_26[162]}
   );
   gpc615_5 gpc1038 (
      {stage0_26[382], stage0_26[383], stage0_26[384], stage0_26[385], stage0_26[386]},
      {stage0_27[254]},
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage1_30[8],stage1_29[49],stage1_28[106],stage1_27[146],stage1_26[163]}
   );
   gpc615_5 gpc1039 (
      {stage0_26[387], stage0_26[388], stage0_26[389], stage0_26[390], stage0_26[391]},
      {stage0_27[255]},
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage1_30[9],stage1_29[50],stage1_28[107],stage1_27[147],stage1_26[164]}
   );
   gpc615_5 gpc1040 (
      {stage0_26[392], stage0_26[393], stage0_26[394], stage0_26[395], stage0_26[396]},
      {stage0_27[256]},
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage1_30[10],stage1_29[51],stage1_28[108],stage1_27[148],stage1_26[165]}
   );
   gpc615_5 gpc1041 (
      {stage0_26[397], stage0_26[398], stage0_26[399], stage0_26[400], stage0_26[401]},
      {stage0_27[257]},
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage1_30[11],stage1_29[52],stage1_28[109],stage1_27[149],stage1_26[166]}
   );
   gpc615_5 gpc1042 (
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262]},
      {stage0_28[72]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[12],stage1_29[53],stage1_28[110],stage1_27[150]}
   );
   gpc615_5 gpc1043 (
      {stage0_27[263], stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267]},
      {stage0_28[73]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[13],stage1_29[54],stage1_28[111],stage1_27[151]}
   );
   gpc615_5 gpc1044 (
      {stage0_27[268], stage0_27[269], stage0_27[270], stage0_27[271], stage0_27[272]},
      {stage0_28[74]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[14],stage1_29[55],stage1_28[112],stage1_27[152]}
   );
   gpc615_5 gpc1045 (
      {stage0_27[273], stage0_27[274], stage0_27[275], stage0_27[276], stage0_27[277]},
      {stage0_28[75]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[15],stage1_29[56],stage1_28[113],stage1_27[153]}
   );
   gpc615_5 gpc1046 (
      {stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281], stage0_27[282]},
      {stage0_28[76]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[16],stage1_29[57],stage1_28[114],stage1_27[154]}
   );
   gpc615_5 gpc1047 (
      {stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage0_28[77]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[17],stage1_29[58],stage1_28[115],stage1_27[155]}
   );
   gpc615_5 gpc1048 (
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292]},
      {stage0_28[78]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[18],stage1_29[59],stage1_28[116],stage1_27[156]}
   );
   gpc615_5 gpc1049 (
      {stage0_27[293], stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297]},
      {stage0_28[79]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[19],stage1_29[60],stage1_28[117],stage1_27[157]}
   );
   gpc615_5 gpc1050 (
      {stage0_27[298], stage0_27[299], stage0_27[300], stage0_27[301], stage0_27[302]},
      {stage0_28[80]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[20],stage1_29[61],stage1_28[118],stage1_27[158]}
   );
   gpc615_5 gpc1051 (
      {stage0_27[303], stage0_27[304], stage0_27[305], stage0_27[306], stage0_27[307]},
      {stage0_28[81]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[21],stage1_29[62],stage1_28[119],stage1_27[159]}
   );
   gpc615_5 gpc1052 (
      {stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311], stage0_27[312]},
      {stage0_28[82]},
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage1_31[10],stage1_30[22],stage1_29[63],stage1_28[120],stage1_27[160]}
   );
   gpc615_5 gpc1053 (
      {stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage0_28[83]},
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage1_31[11],stage1_30[23],stage1_29[64],stage1_28[121],stage1_27[161]}
   );
   gpc615_5 gpc1054 (
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322]},
      {stage0_28[84]},
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage1_31[12],stage1_30[24],stage1_29[65],stage1_28[122],stage1_27[162]}
   );
   gpc615_5 gpc1055 (
      {stage0_27[323], stage0_27[324], stage0_27[325], stage0_27[326], stage0_27[327]},
      {stage0_28[85]},
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage1_31[13],stage1_30[25],stage1_29[66],stage1_28[123],stage1_27[163]}
   );
   gpc615_5 gpc1056 (
      {stage0_27[328], stage0_27[329], stage0_27[330], stage0_27[331], stage0_27[332]},
      {stage0_28[86]},
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage1_31[14],stage1_30[26],stage1_29[67],stage1_28[124],stage1_27[164]}
   );
   gpc615_5 gpc1057 (
      {stage0_27[333], stage0_27[334], stage0_27[335], stage0_27[336], stage0_27[337]},
      {stage0_28[87]},
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage1_31[15],stage1_30[27],stage1_29[68],stage1_28[125],stage1_27[165]}
   );
   gpc615_5 gpc1058 (
      {stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341], stage0_27[342]},
      {stage0_28[88]},
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage1_31[16],stage1_30[28],stage1_29[69],stage1_28[126],stage1_27[166]}
   );
   gpc615_5 gpc1059 (
      {stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage0_28[89]},
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage1_31[17],stage1_30[29],stage1_29[70],stage1_28[127],stage1_27[167]}
   );
   gpc615_5 gpc1060 (
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352]},
      {stage0_28[90]},
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage1_31[18],stage1_30[30],stage1_29[71],stage1_28[128],stage1_27[168]}
   );
   gpc615_5 gpc1061 (
      {stage0_27[353], stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357]},
      {stage0_28[91]},
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage1_31[19],stage1_30[31],stage1_29[72],stage1_28[129],stage1_27[169]}
   );
   gpc615_5 gpc1062 (
      {stage0_27[358], stage0_27[359], stage0_27[360], stage0_27[361], stage0_27[362]},
      {stage0_28[92]},
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage1_31[20],stage1_30[32],stage1_29[73],stage1_28[130],stage1_27[170]}
   );
   gpc615_5 gpc1063 (
      {stage0_27[363], stage0_27[364], stage0_27[365], stage0_27[366], stage0_27[367]},
      {stage0_28[93]},
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage1_31[21],stage1_30[33],stage1_29[74],stage1_28[131],stage1_27[171]}
   );
   gpc615_5 gpc1064 (
      {stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371], stage0_27[372]},
      {stage0_28[94]},
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage1_31[22],stage1_30[34],stage1_29[75],stage1_28[132],stage1_27[172]}
   );
   gpc615_5 gpc1065 (
      {stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage0_28[95]},
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage1_31[23],stage1_30[35],stage1_29[76],stage1_28[133],stage1_27[173]}
   );
   gpc615_5 gpc1066 (
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382]},
      {stage0_28[96]},
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage1_31[24],stage1_30[36],stage1_29[77],stage1_28[134],stage1_27[174]}
   );
   gpc615_5 gpc1067 (
      {stage0_27[383], stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387]},
      {stage0_28[97]},
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage1_31[25],stage1_30[37],stage1_29[78],stage1_28[135],stage1_27[175]}
   );
   gpc615_5 gpc1068 (
      {stage0_27[388], stage0_27[389], stage0_27[390], stage0_27[391], stage0_27[392]},
      {stage0_28[98]},
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage1_31[26],stage1_30[38],stage1_29[79],stage1_28[136],stage1_27[176]}
   );
   gpc615_5 gpc1069 (
      {stage0_27[393], stage0_27[394], stage0_27[395], stage0_27[396], stage0_27[397]},
      {stage0_28[99]},
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage1_31[27],stage1_30[39],stage1_29[80],stage1_28[137],stage1_27[177]}
   );
   gpc615_5 gpc1070 (
      {stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401], stage0_27[402]},
      {stage0_28[100]},
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage1_31[28],stage1_30[40],stage1_29[81],stage1_28[138],stage1_27[178]}
   );
   gpc615_5 gpc1071 (
      {stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage0_28[101]},
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage1_31[29],stage1_30[41],stage1_29[82],stage1_28[139],stage1_27[179]}
   );
   gpc615_5 gpc1072 (
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412]},
      {stage0_28[102]},
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage1_31[30],stage1_30[42],stage1_29[83],stage1_28[140],stage1_27[180]}
   );
   gpc615_5 gpc1073 (
      {stage0_27[413], stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417]},
      {stage0_28[103]},
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191]},
      {stage1_31[31],stage1_30[43],stage1_29[84],stage1_28[141],stage1_27[181]}
   );
   gpc615_5 gpc1074 (
      {stage0_27[418], stage0_27[419], stage0_27[420], stage0_27[421], stage0_27[422]},
      {stage0_28[104]},
      {stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197]},
      {stage1_31[32],stage1_30[44],stage1_29[85],stage1_28[142],stage1_27[182]}
   );
   gpc615_5 gpc1075 (
      {stage0_27[423], stage0_27[424], stage0_27[425], stage0_27[426], stage0_27[427]},
      {stage0_28[105]},
      {stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203]},
      {stage1_31[33],stage1_30[45],stage1_29[86],stage1_28[143],stage1_27[183]}
   );
   gpc615_5 gpc1076 (
      {stage0_27[428], stage0_27[429], stage0_27[430], stage0_27[431], stage0_27[432]},
      {stage0_28[106]},
      {stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209]},
      {stage1_31[34],stage1_30[46],stage1_29[87],stage1_28[144],stage1_27[184]}
   );
   gpc615_5 gpc1077 (
      {stage0_27[433], stage0_27[434], stage0_27[435], stage0_27[436], stage0_27[437]},
      {stage0_28[107]},
      {stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage1_31[35],stage1_30[47],stage1_29[88],stage1_28[145],stage1_27[185]}
   );
   gpc615_5 gpc1078 (
      {stage0_27[438], stage0_27[439], stage0_27[440], stage0_27[441], stage0_27[442]},
      {stage0_28[108]},
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221]},
      {stage1_31[36],stage1_30[48],stage1_29[89],stage1_28[146],stage1_27[186]}
   );
   gpc615_5 gpc1079 (
      {stage0_27[443], stage0_27[444], stage0_27[445], stage0_27[446], stage0_27[447]},
      {stage0_28[109]},
      {stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227]},
      {stage1_31[37],stage1_30[49],stage1_29[90],stage1_28[147],stage1_27[187]}
   );
   gpc615_5 gpc1080 (
      {stage0_27[448], stage0_27[449], stage0_27[450], stage0_27[451], stage0_27[452]},
      {stage0_28[110]},
      {stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233]},
      {stage1_31[38],stage1_30[50],stage1_29[91],stage1_28[148],stage1_27[188]}
   );
   gpc615_5 gpc1081 (
      {stage0_27[453], stage0_27[454], stage0_27[455], stage0_27[456], stage0_27[457]},
      {stage0_28[111]},
      {stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239]},
      {stage1_31[39],stage1_30[51],stage1_29[92],stage1_28[149],stage1_27[189]}
   );
   gpc615_5 gpc1082 (
      {stage0_27[458], stage0_27[459], stage0_27[460], stage0_27[461], stage0_27[462]},
      {stage0_28[112]},
      {stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage1_31[40],stage1_30[52],stage1_29[93],stage1_28[150],stage1_27[190]}
   );
   gpc615_5 gpc1083 (
      {stage0_27[463], stage0_27[464], stage0_27[465], stage0_27[466], stage0_27[467]},
      {stage0_28[113]},
      {stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250], stage0_29[251]},
      {stage1_31[41],stage1_30[53],stage1_29[94],stage1_28[151],stage1_27[191]}
   );
   gpc615_5 gpc1084 (
      {stage0_27[468], stage0_27[469], stage0_27[470], stage0_27[471], stage0_27[472]},
      {stage0_28[114]},
      {stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255], stage0_29[256], stage0_29[257]},
      {stage1_31[42],stage1_30[54],stage1_29[95],stage1_28[152],stage1_27[192]}
   );
   gpc606_5 gpc1085 (
      {stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[43],stage1_30[55],stage1_29[96],stage1_28[153]}
   );
   gpc606_5 gpc1086 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[44],stage1_30[56],stage1_29[97],stage1_28[154]}
   );
   gpc606_5 gpc1087 (
      {stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[45],stage1_30[57],stage1_29[98],stage1_28[155]}
   );
   gpc606_5 gpc1088 (
      {stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[46],stage1_30[58],stage1_29[99],stage1_28[156]}
   );
   gpc606_5 gpc1089 (
      {stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[47],stage1_30[59],stage1_29[100],stage1_28[157]}
   );
   gpc606_5 gpc1090 (
      {stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[48],stage1_30[60],stage1_29[101],stage1_28[158]}
   );
   gpc606_5 gpc1091 (
      {stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[49],stage1_30[61],stage1_29[102],stage1_28[159]}
   );
   gpc606_5 gpc1092 (
      {stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[50],stage1_30[62],stage1_29[103],stage1_28[160]}
   );
   gpc606_5 gpc1093 (
      {stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[51],stage1_30[63],stage1_29[104],stage1_28[161]}
   );
   gpc606_5 gpc1094 (
      {stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[52],stage1_30[64],stage1_29[105],stage1_28[162]}
   );
   gpc606_5 gpc1095 (
      {stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[53],stage1_30[65],stage1_29[106],stage1_28[163]}
   );
   gpc606_5 gpc1096 (
      {stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[54],stage1_30[66],stage1_29[107],stage1_28[164]}
   );
   gpc606_5 gpc1097 (
      {stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[55],stage1_30[67],stage1_29[108],stage1_28[165]}
   );
   gpc606_5 gpc1098 (
      {stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[56],stage1_30[68],stage1_29[109],stage1_28[166]}
   );
   gpc606_5 gpc1099 (
      {stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[57],stage1_30[69],stage1_29[110],stage1_28[167]}
   );
   gpc606_5 gpc1100 (
      {stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[58],stage1_30[70],stage1_29[111],stage1_28[168]}
   );
   gpc606_5 gpc1101 (
      {stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[59],stage1_30[71],stage1_29[112],stage1_28[169]}
   );
   gpc606_5 gpc1102 (
      {stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[60],stage1_30[72],stage1_29[113],stage1_28[170]}
   );
   gpc606_5 gpc1103 (
      {stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[61],stage1_30[73],stage1_29[114],stage1_28[171]}
   );
   gpc606_5 gpc1104 (
      {stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[62],stage1_30[74],stage1_29[115],stage1_28[172]}
   );
   gpc606_5 gpc1105 (
      {stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239], stage0_28[240]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[63],stage1_30[75],stage1_29[116],stage1_28[173]}
   );
   gpc606_5 gpc1106 (
      {stage0_28[241], stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245], stage0_28[246]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[64],stage1_30[76],stage1_29[117],stage1_28[174]}
   );
   gpc606_5 gpc1107 (
      {stage0_28[247], stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251], stage0_28[252]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[65],stage1_30[77],stage1_29[118],stage1_28[175]}
   );
   gpc606_5 gpc1108 (
      {stage0_28[253], stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257], stage0_28[258]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[66],stage1_30[78],stage1_29[119],stage1_28[176]}
   );
   gpc606_5 gpc1109 (
      {stage0_28[259], stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263], stage0_28[264]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[67],stage1_30[79],stage1_29[120],stage1_28[177]}
   );
   gpc606_5 gpc1110 (
      {stage0_28[265], stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269], stage0_28[270]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[68],stage1_30[80],stage1_29[121],stage1_28[178]}
   );
   gpc606_5 gpc1111 (
      {stage0_28[271], stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275], stage0_28[276]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[69],stage1_30[81],stage1_29[122],stage1_28[179]}
   );
   gpc606_5 gpc1112 (
      {stage0_28[277], stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281], stage0_28[282]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[70],stage1_30[82],stage1_29[123],stage1_28[180]}
   );
   gpc606_5 gpc1113 (
      {stage0_28[283], stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287], stage0_28[288]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[71],stage1_30[83],stage1_29[124],stage1_28[181]}
   );
   gpc606_5 gpc1114 (
      {stage0_28[289], stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293], stage0_28[294]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[72],stage1_30[84],stage1_29[125],stage1_28[182]}
   );
   gpc606_5 gpc1115 (
      {stage0_28[295], stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299], stage0_28[300]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[73],stage1_30[85],stage1_29[126],stage1_28[183]}
   );
   gpc606_5 gpc1116 (
      {stage0_28[301], stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305], stage0_28[306]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[74],stage1_30[86],stage1_29[127],stage1_28[184]}
   );
   gpc606_5 gpc1117 (
      {stage0_28[307], stage0_28[308], stage0_28[309], stage0_28[310], stage0_28[311], stage0_28[312]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[75],stage1_30[87],stage1_29[128],stage1_28[185]}
   );
   gpc606_5 gpc1118 (
      {stage0_28[313], stage0_28[314], stage0_28[315], stage0_28[316], stage0_28[317], stage0_28[318]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[76],stage1_30[88],stage1_29[129],stage1_28[186]}
   );
   gpc606_5 gpc1119 (
      {stage0_28[319], stage0_28[320], stage0_28[321], stage0_28[322], stage0_28[323], stage0_28[324]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[77],stage1_30[89],stage1_29[130],stage1_28[187]}
   );
   gpc606_5 gpc1120 (
      {stage0_28[325], stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329], stage0_28[330]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[78],stage1_30[90],stage1_29[131],stage1_28[188]}
   );
   gpc606_5 gpc1121 (
      {stage0_28[331], stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335], stage0_28[336]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[79],stage1_30[91],stage1_29[132],stage1_28[189]}
   );
   gpc606_5 gpc1122 (
      {stage0_28[337], stage0_28[338], stage0_28[339], stage0_28[340], stage0_28[341], stage0_28[342]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[80],stage1_30[92],stage1_29[133],stage1_28[190]}
   );
   gpc606_5 gpc1123 (
      {stage0_28[343], stage0_28[344], stage0_28[345], stage0_28[346], stage0_28[347], stage0_28[348]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[81],stage1_30[93],stage1_29[134],stage1_28[191]}
   );
   gpc606_5 gpc1124 (
      {stage0_28[349], stage0_28[350], stage0_28[351], stage0_28[352], stage0_28[353], stage0_28[354]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[82],stage1_30[94],stage1_29[135],stage1_28[192]}
   );
   gpc606_5 gpc1125 (
      {stage0_28[355], stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359], stage0_28[360]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[83],stage1_30[95],stage1_29[136],stage1_28[193]}
   );
   gpc606_5 gpc1126 (
      {stage0_28[361], stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365], stage0_28[366]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[84],stage1_30[96],stage1_29[137],stage1_28[194]}
   );
   gpc606_5 gpc1127 (
      {stage0_28[367], stage0_28[368], stage0_28[369], stage0_28[370], stage0_28[371], stage0_28[372]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[85],stage1_30[97],stage1_29[138],stage1_28[195]}
   );
   gpc606_5 gpc1128 (
      {stage0_28[373], stage0_28[374], stage0_28[375], stage0_28[376], stage0_28[377], stage0_28[378]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[86],stage1_30[98],stage1_29[139],stage1_28[196]}
   );
   gpc606_5 gpc1129 (
      {stage0_28[379], stage0_28[380], stage0_28[381], stage0_28[382], stage0_28[383], stage0_28[384]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[87],stage1_30[99],stage1_29[140],stage1_28[197]}
   );
   gpc606_5 gpc1130 (
      {stage0_28[385], stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389], stage0_28[390]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[88],stage1_30[100],stage1_29[141],stage1_28[198]}
   );
   gpc606_5 gpc1131 (
      {stage0_28[391], stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395], stage0_28[396]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[89],stage1_30[101],stage1_29[142],stage1_28[199]}
   );
   gpc606_5 gpc1132 (
      {stage0_28[397], stage0_28[398], stage0_28[399], stage0_28[400], stage0_28[401], stage0_28[402]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[90],stage1_30[102],stage1_29[143],stage1_28[200]}
   );
   gpc606_5 gpc1133 (
      {stage0_28[403], stage0_28[404], stage0_28[405], stage0_28[406], stage0_28[407], stage0_28[408]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[91],stage1_30[103],stage1_29[144],stage1_28[201]}
   );
   gpc606_5 gpc1134 (
      {stage0_28[409], stage0_28[410], stage0_28[411], stage0_28[412], stage0_28[413], stage0_28[414]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[92],stage1_30[104],stage1_29[145],stage1_28[202]}
   );
   gpc606_5 gpc1135 (
      {stage0_28[415], stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419], stage0_28[420]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[93],stage1_30[105],stage1_29[146],stage1_28[203]}
   );
   gpc606_5 gpc1136 (
      {stage0_28[421], stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425], stage0_28[426]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[94],stage1_30[106],stage1_29[147],stage1_28[204]}
   );
   gpc606_5 gpc1137 (
      {stage0_28[427], stage0_28[428], stage0_28[429], stage0_28[430], stage0_28[431], stage0_28[432]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[95],stage1_30[107],stage1_29[148],stage1_28[205]}
   );
   gpc606_5 gpc1138 (
      {stage0_28[433], stage0_28[434], stage0_28[435], stage0_28[436], stage0_28[437], stage0_28[438]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[96],stage1_30[108],stage1_29[149],stage1_28[206]}
   );
   gpc606_5 gpc1139 (
      {stage0_28[439], stage0_28[440], stage0_28[441], stage0_28[442], stage0_28[443], stage0_28[444]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[97],stage1_30[109],stage1_29[150],stage1_28[207]}
   );
   gpc606_5 gpc1140 (
      {stage0_28[445], stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449], stage0_28[450]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[98],stage1_30[110],stage1_29[151],stage1_28[208]}
   );
   gpc606_5 gpc1141 (
      {stage0_28[451], stage0_28[452], stage0_28[453], stage0_28[454], stage0_28[455], stage0_28[456]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[99],stage1_30[111],stage1_29[152],stage1_28[209]}
   );
   gpc606_5 gpc1142 (
      {stage0_28[457], stage0_28[458], stage0_28[459], stage0_28[460], stage0_28[461], stage0_28[462]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[100],stage1_30[112],stage1_29[153],stage1_28[210]}
   );
   gpc606_5 gpc1143 (
      {stage0_28[463], stage0_28[464], stage0_28[465], stage0_28[466], stage0_28[467], stage0_28[468]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[101],stage1_30[113],stage1_29[154],stage1_28[211]}
   );
   gpc606_5 gpc1144 (
      {stage0_28[469], stage0_28[470], stage0_28[471], stage0_28[472], stage0_28[473], stage0_28[474]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[102],stage1_30[114],stage1_29[155],stage1_28[212]}
   );
   gpc606_5 gpc1145 (
      {stage0_29[258], stage0_29[259], stage0_29[260], stage0_29[261], stage0_29[262], stage0_29[263]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[60],stage1_31[103],stage1_30[115],stage1_29[156]}
   );
   gpc606_5 gpc1146 (
      {stage0_29[264], stage0_29[265], stage0_29[266], stage0_29[267], stage0_29[268], stage0_29[269]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[61],stage1_31[104],stage1_30[116],stage1_29[157]}
   );
   gpc606_5 gpc1147 (
      {stage0_29[270], stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274], stage0_29[275]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[62],stage1_31[105],stage1_30[117],stage1_29[158]}
   );
   gpc606_5 gpc1148 (
      {stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280], stage0_29[281]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[63],stage1_31[106],stage1_30[118],stage1_29[159]}
   );
   gpc606_5 gpc1149 (
      {stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285], stage0_29[286], stage0_29[287]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[64],stage1_31[107],stage1_30[119],stage1_29[160]}
   );
   gpc606_5 gpc1150 (
      {stage0_29[288], stage0_29[289], stage0_29[290], stage0_29[291], stage0_29[292], stage0_29[293]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[65],stage1_31[108],stage1_30[120],stage1_29[161]}
   );
   gpc606_5 gpc1151 (
      {stage0_29[294], stage0_29[295], stage0_29[296], stage0_29[297], stage0_29[298], stage0_29[299]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[66],stage1_31[109],stage1_30[121],stage1_29[162]}
   );
   gpc606_5 gpc1152 (
      {stage0_29[300], stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304], stage0_29[305]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[67],stage1_31[110],stage1_30[122],stage1_29[163]}
   );
   gpc606_5 gpc1153 (
      {stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310], stage0_29[311]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[68],stage1_31[111],stage1_30[123],stage1_29[164]}
   );
   gpc606_5 gpc1154 (
      {stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315], stage0_29[316], stage0_29[317]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[69],stage1_31[112],stage1_30[124],stage1_29[165]}
   );
   gpc606_5 gpc1155 (
      {stage0_29[318], stage0_29[319], stage0_29[320], stage0_29[321], stage0_29[322], stage0_29[323]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[70],stage1_31[113],stage1_30[125],stage1_29[166]}
   );
   gpc606_5 gpc1156 (
      {stage0_29[324], stage0_29[325], stage0_29[326], stage0_29[327], stage0_29[328], stage0_29[329]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[71],stage1_31[114],stage1_30[126],stage1_29[167]}
   );
   gpc606_5 gpc1157 (
      {stage0_29[330], stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334], stage0_29[335]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[72],stage1_31[115],stage1_30[127],stage1_29[168]}
   );
   gpc606_5 gpc1158 (
      {stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340], stage0_29[341]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[73],stage1_31[116],stage1_30[128],stage1_29[169]}
   );
   gpc606_5 gpc1159 (
      {stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345], stage0_29[346], stage0_29[347]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[74],stage1_31[117],stage1_30[129],stage1_29[170]}
   );
   gpc606_5 gpc1160 (
      {stage0_29[348], stage0_29[349], stage0_29[350], stage0_29[351], stage0_29[352], stage0_29[353]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[75],stage1_31[118],stage1_30[130],stage1_29[171]}
   );
   gpc606_5 gpc1161 (
      {stage0_29[354], stage0_29[355], stage0_29[356], stage0_29[357], stage0_29[358], stage0_29[359]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[76],stage1_31[119],stage1_30[131],stage1_29[172]}
   );
   gpc606_5 gpc1162 (
      {stage0_29[360], stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364], stage0_29[365]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[77],stage1_31[120],stage1_30[132],stage1_29[173]}
   );
   gpc606_5 gpc1163 (
      {stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370], stage0_29[371]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[78],stage1_31[121],stage1_30[133],stage1_29[174]}
   );
   gpc606_5 gpc1164 (
      {stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375], stage0_29[376], stage0_29[377]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[79],stage1_31[122],stage1_30[134],stage1_29[175]}
   );
   gpc606_5 gpc1165 (
      {stage0_29[378], stage0_29[379], stage0_29[380], stage0_29[381], stage0_29[382], stage0_29[383]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[80],stage1_31[123],stage1_30[135],stage1_29[176]}
   );
   gpc606_5 gpc1166 (
      {stage0_29[384], stage0_29[385], stage0_29[386], stage0_29[387], stage0_29[388], stage0_29[389]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[81],stage1_31[124],stage1_30[136],stage1_29[177]}
   );
   gpc606_5 gpc1167 (
      {stage0_29[390], stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394], stage0_29[395]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[82],stage1_31[125],stage1_30[137],stage1_29[178]}
   );
   gpc606_5 gpc1168 (
      {stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400], stage0_29[401]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[83],stage1_31[126],stage1_30[138],stage1_29[179]}
   );
   gpc606_5 gpc1169 (
      {stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405], stage0_29[406], stage0_29[407]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[84],stage1_31[127],stage1_30[139],stage1_29[180]}
   );
   gpc606_5 gpc1170 (
      {stage0_29[408], stage0_29[409], stage0_29[410], stage0_29[411], stage0_29[412], stage0_29[413]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[85],stage1_31[128],stage1_30[140],stage1_29[181]}
   );
   gpc606_5 gpc1171 (
      {stage0_29[414], stage0_29[415], stage0_29[416], stage0_29[417], stage0_29[418], stage0_29[419]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[86],stage1_31[129],stage1_30[141],stage1_29[182]}
   );
   gpc606_5 gpc1172 (
      {stage0_29[420], stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424], stage0_29[425]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[87],stage1_31[130],stage1_30[142],stage1_29[183]}
   );
   gpc606_5 gpc1173 (
      {stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430], stage0_29[431]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[88],stage1_31[131],stage1_30[143],stage1_29[184]}
   );
   gpc606_5 gpc1174 (
      {stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435], stage0_29[436], stage0_29[437]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[89],stage1_31[132],stage1_30[144],stage1_29[185]}
   );
   gpc606_5 gpc1175 (
      {stage0_29[438], stage0_29[439], stage0_29[440], stage0_29[441], stage0_29[442], stage0_29[443]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[90],stage1_31[133],stage1_30[145],stage1_29[186]}
   );
   gpc615_5 gpc1176 (
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364]},
      {stage0_31[186]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[31],stage1_32[91],stage1_31[134],stage1_30[146]}
   );
   gpc615_5 gpc1177 (
      {stage0_30[365], stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369]},
      {stage0_31[187]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[32],stage1_32[92],stage1_31[135],stage1_30[147]}
   );
   gpc615_5 gpc1178 (
      {stage0_30[370], stage0_30[371], stage0_30[372], stage0_30[373], stage0_30[374]},
      {stage0_31[188]},
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage1_34[2],stage1_33[33],stage1_32[93],stage1_31[136],stage1_30[148]}
   );
   gpc615_5 gpc1179 (
      {stage0_30[375], stage0_30[376], stage0_30[377], stage0_30[378], stage0_30[379]},
      {stage0_31[189]},
      {stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21], stage0_32[22], stage0_32[23]},
      {stage1_34[3],stage1_33[34],stage1_32[94],stage1_31[137],stage1_30[149]}
   );
   gpc615_5 gpc1180 (
      {stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383], stage0_30[384]},
      {stage0_31[190]},
      {stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27], stage0_32[28], stage0_32[29]},
      {stage1_34[4],stage1_33[35],stage1_32[95],stage1_31[138],stage1_30[150]}
   );
   gpc615_5 gpc1181 (
      {stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage0_31[191]},
      {stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33], stage0_32[34], stage0_32[35]},
      {stage1_34[5],stage1_33[36],stage1_32[96],stage1_31[139],stage1_30[151]}
   );
   gpc615_5 gpc1182 (
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394]},
      {stage0_31[192]},
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage1_34[6],stage1_33[37],stage1_32[97],stage1_31[140],stage1_30[152]}
   );
   gpc615_5 gpc1183 (
      {stage0_30[395], stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399]},
      {stage0_31[193]},
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage1_34[7],stage1_33[38],stage1_32[98],stage1_31[141],stage1_30[153]}
   );
   gpc615_5 gpc1184 (
      {stage0_30[400], stage0_30[401], stage0_30[402], stage0_30[403], stage0_30[404]},
      {stage0_31[194]},
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52], stage0_32[53]},
      {stage1_34[8],stage1_33[39],stage1_32[99],stage1_31[142],stage1_30[154]}
   );
   gpc615_5 gpc1185 (
      {stage0_30[405], stage0_30[406], stage0_30[407], stage0_30[408], stage0_30[409]},
      {stage0_31[195]},
      {stage0_32[54], stage0_32[55], stage0_32[56], stage0_32[57], stage0_32[58], stage0_32[59]},
      {stage1_34[9],stage1_33[40],stage1_32[100],stage1_31[143],stage1_30[155]}
   );
   gpc615_5 gpc1186 (
      {stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413], stage0_30[414]},
      {stage0_31[196]},
      {stage0_32[60], stage0_32[61], stage0_32[62], stage0_32[63], stage0_32[64], stage0_32[65]},
      {stage1_34[10],stage1_33[41],stage1_32[101],stage1_31[144],stage1_30[156]}
   );
   gpc615_5 gpc1187 (
      {stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage0_31[197]},
      {stage0_32[66], stage0_32[67], stage0_32[68], stage0_32[69], stage0_32[70], stage0_32[71]},
      {stage1_34[11],stage1_33[42],stage1_32[102],stage1_31[145],stage1_30[157]}
   );
   gpc615_5 gpc1188 (
      {stage0_30[420], stage0_30[421], stage0_30[422], stage0_30[423], stage0_30[424]},
      {stage0_31[198]},
      {stage0_32[72], stage0_32[73], stage0_32[74], stage0_32[75], stage0_32[76], stage0_32[77]},
      {stage1_34[12],stage1_33[43],stage1_32[103],stage1_31[146],stage1_30[158]}
   );
   gpc615_5 gpc1189 (
      {stage0_30[425], stage0_30[426], stage0_30[427], stage0_30[428], stage0_30[429]},
      {stage0_31[199]},
      {stage0_32[78], stage0_32[79], stage0_32[80], stage0_32[81], stage0_32[82], stage0_32[83]},
      {stage1_34[13],stage1_33[44],stage1_32[104],stage1_31[147],stage1_30[159]}
   );
   gpc615_5 gpc1190 (
      {stage0_30[430], stage0_30[431], stage0_30[432], stage0_30[433], stage0_30[434]},
      {stage0_31[200]},
      {stage0_32[84], stage0_32[85], stage0_32[86], stage0_32[87], stage0_32[88], stage0_32[89]},
      {stage1_34[14],stage1_33[45],stage1_32[105],stage1_31[148],stage1_30[160]}
   );
   gpc615_5 gpc1191 (
      {stage0_30[435], stage0_30[436], stage0_30[437], stage0_30[438], stage0_30[439]},
      {stage0_31[201]},
      {stage0_32[90], stage0_32[91], stage0_32[92], stage0_32[93], stage0_32[94], stage0_32[95]},
      {stage1_34[15],stage1_33[46],stage1_32[106],stage1_31[149],stage1_30[161]}
   );
   gpc615_5 gpc1192 (
      {stage0_30[440], stage0_30[441], stage0_30[442], stage0_30[443], stage0_30[444]},
      {stage0_31[202]},
      {stage0_32[96], stage0_32[97], stage0_32[98], stage0_32[99], stage0_32[100], stage0_32[101]},
      {stage1_34[16],stage1_33[47],stage1_32[107],stage1_31[150],stage1_30[162]}
   );
   gpc615_5 gpc1193 (
      {stage0_30[445], stage0_30[446], stage0_30[447], stage0_30[448], stage0_30[449]},
      {stage0_31[203]},
      {stage0_32[102], stage0_32[103], stage0_32[104], stage0_32[105], stage0_32[106], stage0_32[107]},
      {stage1_34[17],stage1_33[48],stage1_32[108],stage1_31[151],stage1_30[163]}
   );
   gpc615_5 gpc1194 (
      {stage0_30[450], stage0_30[451], stage0_30[452], stage0_30[453], stage0_30[454]},
      {stage0_31[204]},
      {stage0_32[108], stage0_32[109], stage0_32[110], stage0_32[111], stage0_32[112], stage0_32[113]},
      {stage1_34[18],stage1_33[49],stage1_32[109],stage1_31[152],stage1_30[164]}
   );
   gpc615_5 gpc1195 (
      {stage0_30[455], stage0_30[456], stage0_30[457], stage0_30[458], stage0_30[459]},
      {stage0_31[205]},
      {stage0_32[114], stage0_32[115], stage0_32[116], stage0_32[117], stage0_32[118], stage0_32[119]},
      {stage1_34[19],stage1_33[50],stage1_32[110],stage1_31[153],stage1_30[165]}
   );
   gpc615_5 gpc1196 (
      {stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209], stage0_31[210]},
      {stage0_32[120]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[20],stage1_33[51],stage1_32[111],stage1_31[154]}
   );
   gpc615_5 gpc1197 (
      {stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage0_32[121]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[21],stage1_33[52],stage1_32[112],stage1_31[155]}
   );
   gpc615_5 gpc1198 (
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220]},
      {stage0_32[122]},
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage1_35[2],stage1_34[22],stage1_33[53],stage1_32[113],stage1_31[156]}
   );
   gpc615_5 gpc1199 (
      {stage0_31[221], stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225]},
      {stage0_32[123]},
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage1_35[3],stage1_34[23],stage1_33[54],stage1_32[114],stage1_31[157]}
   );
   gpc615_5 gpc1200 (
      {stage0_31[226], stage0_31[227], stage0_31[228], stage0_31[229], stage0_31[230]},
      {stage0_32[124]},
      {stage0_33[24], stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29]},
      {stage1_35[4],stage1_34[24],stage1_33[55],stage1_32[115],stage1_31[158]}
   );
   gpc615_5 gpc1201 (
      {stage0_31[231], stage0_31[232], stage0_31[233], stage0_31[234], stage0_31[235]},
      {stage0_32[125]},
      {stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35]},
      {stage1_35[5],stage1_34[25],stage1_33[56],stage1_32[116],stage1_31[159]}
   );
   gpc615_5 gpc1202 (
      {stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239], stage0_31[240]},
      {stage0_32[126]},
      {stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41]},
      {stage1_35[6],stage1_34[26],stage1_33[57],stage1_32[117],stage1_31[160]}
   );
   gpc615_5 gpc1203 (
      {stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage0_32[127]},
      {stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47]},
      {stage1_35[7],stage1_34[27],stage1_33[58],stage1_32[118],stage1_31[161]}
   );
   gpc615_5 gpc1204 (
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250]},
      {stage0_32[128]},
      {stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53]},
      {stage1_35[8],stage1_34[28],stage1_33[59],stage1_32[119],stage1_31[162]}
   );
   gpc615_5 gpc1205 (
      {stage0_31[251], stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255]},
      {stage0_32[129]},
      {stage0_33[54], stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59]},
      {stage1_35[9],stage1_34[29],stage1_33[60],stage1_32[120],stage1_31[163]}
   );
   gpc615_5 gpc1206 (
      {stage0_31[256], stage0_31[257], stage0_31[258], stage0_31[259], stage0_31[260]},
      {stage0_32[130]},
      {stage0_33[60], stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65]},
      {stage1_35[10],stage1_34[30],stage1_33[61],stage1_32[121],stage1_31[164]}
   );
   gpc615_5 gpc1207 (
      {stage0_31[261], stage0_31[262], stage0_31[263], stage0_31[264], stage0_31[265]},
      {stage0_32[131]},
      {stage0_33[66], stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71]},
      {stage1_35[11],stage1_34[31],stage1_33[62],stage1_32[122],stage1_31[165]}
   );
   gpc615_5 gpc1208 (
      {stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269], stage0_31[270]},
      {stage0_32[132]},
      {stage0_33[72], stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77]},
      {stage1_35[12],stage1_34[32],stage1_33[63],stage1_32[123],stage1_31[166]}
   );
   gpc615_5 gpc1209 (
      {stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage0_32[133]},
      {stage0_33[78], stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83]},
      {stage1_35[13],stage1_34[33],stage1_33[64],stage1_32[124],stage1_31[167]}
   );
   gpc615_5 gpc1210 (
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280]},
      {stage0_32[134]},
      {stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88], stage0_33[89]},
      {stage1_35[14],stage1_34[34],stage1_33[65],stage1_32[125],stage1_31[168]}
   );
   gpc615_5 gpc1211 (
      {stage0_31[281], stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285]},
      {stage0_32[135]},
      {stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93], stage0_33[94], stage0_33[95]},
      {stage1_35[15],stage1_34[35],stage1_33[66],stage1_32[126],stage1_31[169]}
   );
   gpc615_5 gpc1212 (
      {stage0_31[286], stage0_31[287], stage0_31[288], stage0_31[289], stage0_31[290]},
      {stage0_32[136]},
      {stage0_33[96], stage0_33[97], stage0_33[98], stage0_33[99], stage0_33[100], stage0_33[101]},
      {stage1_35[16],stage1_34[36],stage1_33[67],stage1_32[127],stage1_31[170]}
   );
   gpc615_5 gpc1213 (
      {stage0_31[291], stage0_31[292], stage0_31[293], stage0_31[294], stage0_31[295]},
      {stage0_32[137]},
      {stage0_33[102], stage0_33[103], stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107]},
      {stage1_35[17],stage1_34[37],stage1_33[68],stage1_32[128],stage1_31[171]}
   );
   gpc615_5 gpc1214 (
      {stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299], stage0_31[300]},
      {stage0_32[138]},
      {stage0_33[108], stage0_33[109], stage0_33[110], stage0_33[111], stage0_33[112], stage0_33[113]},
      {stage1_35[18],stage1_34[38],stage1_33[69],stage1_32[129],stage1_31[172]}
   );
   gpc615_5 gpc1215 (
      {stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage0_32[139]},
      {stage0_33[114], stage0_33[115], stage0_33[116], stage0_33[117], stage0_33[118], stage0_33[119]},
      {stage1_35[19],stage1_34[39],stage1_33[70],stage1_32[130],stage1_31[173]}
   );
   gpc615_5 gpc1216 (
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310]},
      {stage0_32[140]},
      {stage0_33[120], stage0_33[121], stage0_33[122], stage0_33[123], stage0_33[124], stage0_33[125]},
      {stage1_35[20],stage1_34[40],stage1_33[71],stage1_32[131],stage1_31[174]}
   );
   gpc615_5 gpc1217 (
      {stage0_31[311], stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315]},
      {stage0_32[141]},
      {stage0_33[126], stage0_33[127], stage0_33[128], stage0_33[129], stage0_33[130], stage0_33[131]},
      {stage1_35[21],stage1_34[41],stage1_33[72],stage1_32[132],stage1_31[175]}
   );
   gpc615_5 gpc1218 (
      {stage0_31[316], stage0_31[317], stage0_31[318], stage0_31[319], stage0_31[320]},
      {stage0_32[142]},
      {stage0_33[132], stage0_33[133], stage0_33[134], stage0_33[135], stage0_33[136], stage0_33[137]},
      {stage1_35[22],stage1_34[42],stage1_33[73],stage1_32[133],stage1_31[176]}
   );
   gpc615_5 gpc1219 (
      {stage0_31[321], stage0_31[322], stage0_31[323], stage0_31[324], stage0_31[325]},
      {stage0_32[143]},
      {stage0_33[138], stage0_33[139], stage0_33[140], stage0_33[141], stage0_33[142], stage0_33[143]},
      {stage1_35[23],stage1_34[43],stage1_33[74],stage1_32[134],stage1_31[177]}
   );
   gpc615_5 gpc1220 (
      {stage0_31[326], stage0_31[327], stage0_31[328], stage0_31[329], stage0_31[330]},
      {stage0_32[144]},
      {stage0_33[144], stage0_33[145], stage0_33[146], stage0_33[147], stage0_33[148], stage0_33[149]},
      {stage1_35[24],stage1_34[44],stage1_33[75],stage1_32[135],stage1_31[178]}
   );
   gpc615_5 gpc1221 (
      {stage0_31[331], stage0_31[332], stage0_31[333], stage0_31[334], stage0_31[335]},
      {stage0_32[145]},
      {stage0_33[150], stage0_33[151], stage0_33[152], stage0_33[153], stage0_33[154], stage0_33[155]},
      {stage1_35[25],stage1_34[45],stage1_33[76],stage1_32[136],stage1_31[179]}
   );
   gpc615_5 gpc1222 (
      {stage0_31[336], stage0_31[337], stage0_31[338], stage0_31[339], stage0_31[340]},
      {stage0_32[146]},
      {stage0_33[156], stage0_33[157], stage0_33[158], stage0_33[159], stage0_33[160], stage0_33[161]},
      {stage1_35[26],stage1_34[46],stage1_33[77],stage1_32[137],stage1_31[180]}
   );
   gpc615_5 gpc1223 (
      {stage0_31[341], stage0_31[342], stage0_31[343], stage0_31[344], stage0_31[345]},
      {stage0_32[147]},
      {stage0_33[162], stage0_33[163], stage0_33[164], stage0_33[165], stage0_33[166], stage0_33[167]},
      {stage1_35[27],stage1_34[47],stage1_33[78],stage1_32[138],stage1_31[181]}
   );
   gpc615_5 gpc1224 (
      {stage0_31[346], stage0_31[347], stage0_31[348], stage0_31[349], stage0_31[350]},
      {stage0_32[148]},
      {stage0_33[168], stage0_33[169], stage0_33[170], stage0_33[171], stage0_33[172], stage0_33[173]},
      {stage1_35[28],stage1_34[48],stage1_33[79],stage1_32[139],stage1_31[182]}
   );
   gpc615_5 gpc1225 (
      {stage0_31[351], stage0_31[352], stage0_31[353], stage0_31[354], stage0_31[355]},
      {stage0_32[149]},
      {stage0_33[174], stage0_33[175], stage0_33[176], stage0_33[177], stage0_33[178], stage0_33[179]},
      {stage1_35[29],stage1_34[49],stage1_33[80],stage1_32[140],stage1_31[183]}
   );
   gpc615_5 gpc1226 (
      {stage0_31[356], stage0_31[357], stage0_31[358], stage0_31[359], stage0_31[360]},
      {stage0_32[150]},
      {stage0_33[180], stage0_33[181], stage0_33[182], stage0_33[183], stage0_33[184], stage0_33[185]},
      {stage1_35[30],stage1_34[50],stage1_33[81],stage1_32[141],stage1_31[184]}
   );
   gpc615_5 gpc1227 (
      {stage0_31[361], stage0_31[362], stage0_31[363], stage0_31[364], stage0_31[365]},
      {stage0_32[151]},
      {stage0_33[186], stage0_33[187], stage0_33[188], stage0_33[189], stage0_33[190], stage0_33[191]},
      {stage1_35[31],stage1_34[51],stage1_33[82],stage1_32[142],stage1_31[185]}
   );
   gpc615_5 gpc1228 (
      {stage0_31[366], stage0_31[367], stage0_31[368], stage0_31[369], stage0_31[370]},
      {stage0_32[152]},
      {stage0_33[192], stage0_33[193], stage0_33[194], stage0_33[195], stage0_33[196], stage0_33[197]},
      {stage1_35[32],stage1_34[52],stage1_33[83],stage1_32[143],stage1_31[186]}
   );
   gpc615_5 gpc1229 (
      {stage0_31[371], stage0_31[372], stage0_31[373], stage0_31[374], stage0_31[375]},
      {stage0_32[153]},
      {stage0_33[198], stage0_33[199], stage0_33[200], stage0_33[201], stage0_33[202], stage0_33[203]},
      {stage1_35[33],stage1_34[53],stage1_33[84],stage1_32[144],stage1_31[187]}
   );
   gpc615_5 gpc1230 (
      {stage0_31[376], stage0_31[377], stage0_31[378], stage0_31[379], stage0_31[380]},
      {stage0_32[154]},
      {stage0_33[204], stage0_33[205], stage0_33[206], stage0_33[207], stage0_33[208], stage0_33[209]},
      {stage1_35[34],stage1_34[54],stage1_33[85],stage1_32[145],stage1_31[188]}
   );
   gpc615_5 gpc1231 (
      {stage0_31[381], stage0_31[382], stage0_31[383], stage0_31[384], stage0_31[385]},
      {stage0_32[155]},
      {stage0_33[210], stage0_33[211], stage0_33[212], stage0_33[213], stage0_33[214], stage0_33[215]},
      {stage1_35[35],stage1_34[55],stage1_33[86],stage1_32[146],stage1_31[189]}
   );
   gpc615_5 gpc1232 (
      {stage0_31[386], stage0_31[387], stage0_31[388], stage0_31[389], stage0_31[390]},
      {stage0_32[156]},
      {stage0_33[216], stage0_33[217], stage0_33[218], stage0_33[219], stage0_33[220], stage0_33[221]},
      {stage1_35[36],stage1_34[56],stage1_33[87],stage1_32[147],stage1_31[190]}
   );
   gpc615_5 gpc1233 (
      {stage0_31[391], stage0_31[392], stage0_31[393], stage0_31[394], stage0_31[395]},
      {stage0_32[157]},
      {stage0_33[222], stage0_33[223], stage0_33[224], stage0_33[225], stage0_33[226], stage0_33[227]},
      {stage1_35[37],stage1_34[57],stage1_33[88],stage1_32[148],stage1_31[191]}
   );
   gpc615_5 gpc1234 (
      {stage0_31[396], stage0_31[397], stage0_31[398], stage0_31[399], stage0_31[400]},
      {stage0_32[158]},
      {stage0_33[228], stage0_33[229], stage0_33[230], stage0_33[231], stage0_33[232], stage0_33[233]},
      {stage1_35[38],stage1_34[58],stage1_33[89],stage1_32[149],stage1_31[192]}
   );
   gpc615_5 gpc1235 (
      {stage0_31[401], stage0_31[402], stage0_31[403], stage0_31[404], stage0_31[405]},
      {stage0_32[159]},
      {stage0_33[234], stage0_33[235], stage0_33[236], stage0_33[237], stage0_33[238], stage0_33[239]},
      {stage1_35[39],stage1_34[59],stage1_33[90],stage1_32[150],stage1_31[193]}
   );
   gpc615_5 gpc1236 (
      {stage0_31[406], stage0_31[407], stage0_31[408], stage0_31[409], stage0_31[410]},
      {stage0_32[160]},
      {stage0_33[240], stage0_33[241], stage0_33[242], stage0_33[243], stage0_33[244], stage0_33[245]},
      {stage1_35[40],stage1_34[60],stage1_33[91],stage1_32[151],stage1_31[194]}
   );
   gpc615_5 gpc1237 (
      {stage0_31[411], stage0_31[412], stage0_31[413], stage0_31[414], stage0_31[415]},
      {stage0_32[161]},
      {stage0_33[246], stage0_33[247], stage0_33[248], stage0_33[249], stage0_33[250], stage0_33[251]},
      {stage1_35[41],stage1_34[61],stage1_33[92],stage1_32[152],stage1_31[195]}
   );
   gpc615_5 gpc1238 (
      {stage0_31[416], stage0_31[417], stage0_31[418], stage0_31[419], stage0_31[420]},
      {stage0_32[162]},
      {stage0_33[252], stage0_33[253], stage0_33[254], stage0_33[255], stage0_33[256], stage0_33[257]},
      {stage1_35[42],stage1_34[62],stage1_33[93],stage1_32[153],stage1_31[196]}
   );
   gpc615_5 gpc1239 (
      {stage0_31[421], stage0_31[422], stage0_31[423], stage0_31[424], stage0_31[425]},
      {stage0_32[163]},
      {stage0_33[258], stage0_33[259], stage0_33[260], stage0_33[261], stage0_33[262], stage0_33[263]},
      {stage1_35[43],stage1_34[63],stage1_33[94],stage1_32[154],stage1_31[197]}
   );
   gpc615_5 gpc1240 (
      {stage0_31[426], stage0_31[427], stage0_31[428], stage0_31[429], stage0_31[430]},
      {stage0_32[164]},
      {stage0_33[264], stage0_33[265], stage0_33[266], stage0_33[267], stage0_33[268], stage0_33[269]},
      {stage1_35[44],stage1_34[64],stage1_33[95],stage1_32[155],stage1_31[198]}
   );
   gpc615_5 gpc1241 (
      {stage0_31[431], stage0_31[432], stage0_31[433], stage0_31[434], stage0_31[435]},
      {stage0_32[165]},
      {stage0_33[270], stage0_33[271], stage0_33[272], stage0_33[273], stage0_33[274], stage0_33[275]},
      {stage1_35[45],stage1_34[65],stage1_33[96],stage1_32[156],stage1_31[199]}
   );
   gpc615_5 gpc1242 (
      {stage0_31[436], stage0_31[437], stage0_31[438], stage0_31[439], stage0_31[440]},
      {stage0_32[166]},
      {stage0_33[276], stage0_33[277], stage0_33[278], stage0_33[279], stage0_33[280], stage0_33[281]},
      {stage1_35[46],stage1_34[66],stage1_33[97],stage1_32[157],stage1_31[200]}
   );
   gpc615_5 gpc1243 (
      {stage0_31[441], stage0_31[442], stage0_31[443], stage0_31[444], stage0_31[445]},
      {stage0_32[167]},
      {stage0_33[282], stage0_33[283], stage0_33[284], stage0_33[285], stage0_33[286], stage0_33[287]},
      {stage1_35[47],stage1_34[67],stage1_33[98],stage1_32[158],stage1_31[201]}
   );
   gpc615_5 gpc1244 (
      {stage0_31[446], stage0_31[447], stage0_31[448], stage0_31[449], stage0_31[450]},
      {stage0_32[168]},
      {stage0_33[288], stage0_33[289], stage0_33[290], stage0_33[291], stage0_33[292], stage0_33[293]},
      {stage1_35[48],stage1_34[68],stage1_33[99],stage1_32[159],stage1_31[202]}
   );
   gpc615_5 gpc1245 (
      {stage0_31[451], stage0_31[452], stage0_31[453], stage0_31[454], stage0_31[455]},
      {stage0_32[169]},
      {stage0_33[294], stage0_33[295], stage0_33[296], stage0_33[297], stage0_33[298], stage0_33[299]},
      {stage1_35[49],stage1_34[69],stage1_33[100],stage1_32[160],stage1_31[203]}
   );
   gpc615_5 gpc1246 (
      {stage0_31[456], stage0_31[457], stage0_31[458], stage0_31[459], stage0_31[460]},
      {stage0_32[170]},
      {stage0_33[300], stage0_33[301], stage0_33[302], stage0_33[303], stage0_33[304], stage0_33[305]},
      {stage1_35[50],stage1_34[70],stage1_33[101],stage1_32[161],stage1_31[204]}
   );
   gpc615_5 gpc1247 (
      {stage0_31[461], stage0_31[462], stage0_31[463], stage0_31[464], stage0_31[465]},
      {stage0_32[171]},
      {stage0_33[306], stage0_33[307], stage0_33[308], stage0_33[309], stage0_33[310], stage0_33[311]},
      {stage1_35[51],stage1_34[71],stage1_33[102],stage1_32[162],stage1_31[205]}
   );
   gpc615_5 gpc1248 (
      {stage0_31[466], stage0_31[467], stage0_31[468], stage0_31[469], stage0_31[470]},
      {stage0_32[172]},
      {stage0_33[312], stage0_33[313], stage0_33[314], stage0_33[315], stage0_33[316], stage0_33[317]},
      {stage1_35[52],stage1_34[72],stage1_33[103],stage1_32[163],stage1_31[206]}
   );
   gpc615_5 gpc1249 (
      {stage0_31[471], stage0_31[472], stage0_31[473], stage0_31[474], stage0_31[475]},
      {stage0_32[173]},
      {stage0_33[318], stage0_33[319], stage0_33[320], stage0_33[321], stage0_33[322], stage0_33[323]},
      {stage1_35[53],stage1_34[73],stage1_33[104],stage1_32[164],stage1_31[207]}
   );
   gpc606_5 gpc1250 (
      {stage0_32[174], stage0_32[175], stage0_32[176], stage0_32[177], stage0_32[178], stage0_32[179]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[54],stage1_34[74],stage1_33[105],stage1_32[165]}
   );
   gpc606_5 gpc1251 (
      {stage0_32[180], stage0_32[181], stage0_32[182], stage0_32[183], stage0_32[184], stage0_32[185]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[55],stage1_34[75],stage1_33[106],stage1_32[166]}
   );
   gpc606_5 gpc1252 (
      {stage0_32[186], stage0_32[187], stage0_32[188], stage0_32[189], stage0_32[190], stage0_32[191]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[56],stage1_34[76],stage1_33[107],stage1_32[167]}
   );
   gpc606_5 gpc1253 (
      {stage0_32[192], stage0_32[193], stage0_32[194], stage0_32[195], stage0_32[196], stage0_32[197]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[57],stage1_34[77],stage1_33[108],stage1_32[168]}
   );
   gpc606_5 gpc1254 (
      {stage0_32[198], stage0_32[199], stage0_32[200], stage0_32[201], stage0_32[202], stage0_32[203]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[58],stage1_34[78],stage1_33[109],stage1_32[169]}
   );
   gpc606_5 gpc1255 (
      {stage0_32[204], stage0_32[205], stage0_32[206], stage0_32[207], stage0_32[208], stage0_32[209]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[59],stage1_34[79],stage1_33[110],stage1_32[170]}
   );
   gpc606_5 gpc1256 (
      {stage0_32[210], stage0_32[211], stage0_32[212], stage0_32[213], stage0_32[214], stage0_32[215]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[60],stage1_34[80],stage1_33[111],stage1_32[171]}
   );
   gpc606_5 gpc1257 (
      {stage0_32[216], stage0_32[217], stage0_32[218], stage0_32[219], stage0_32[220], stage0_32[221]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[61],stage1_34[81],stage1_33[112],stage1_32[172]}
   );
   gpc606_5 gpc1258 (
      {stage0_32[222], stage0_32[223], stage0_32[224], stage0_32[225], stage0_32[226], stage0_32[227]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[62],stage1_34[82],stage1_33[113],stage1_32[173]}
   );
   gpc606_5 gpc1259 (
      {stage0_32[228], stage0_32[229], stage0_32[230], stage0_32[231], stage0_32[232], stage0_32[233]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[63],stage1_34[83],stage1_33[114],stage1_32[174]}
   );
   gpc606_5 gpc1260 (
      {stage0_32[234], stage0_32[235], stage0_32[236], stage0_32[237], stage0_32[238], stage0_32[239]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[64],stage1_34[84],stage1_33[115],stage1_32[175]}
   );
   gpc606_5 gpc1261 (
      {stage0_32[240], stage0_32[241], stage0_32[242], stage0_32[243], stage0_32[244], stage0_32[245]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[65],stage1_34[85],stage1_33[116],stage1_32[176]}
   );
   gpc606_5 gpc1262 (
      {stage0_32[246], stage0_32[247], stage0_32[248], stage0_32[249], stage0_32[250], stage0_32[251]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[66],stage1_34[86],stage1_33[117],stage1_32[177]}
   );
   gpc606_5 gpc1263 (
      {stage0_32[252], stage0_32[253], stage0_32[254], stage0_32[255], stage0_32[256], stage0_32[257]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[67],stage1_34[87],stage1_33[118],stage1_32[178]}
   );
   gpc606_5 gpc1264 (
      {stage0_32[258], stage0_32[259], stage0_32[260], stage0_32[261], stage0_32[262], stage0_32[263]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[68],stage1_34[88],stage1_33[119],stage1_32[179]}
   );
   gpc606_5 gpc1265 (
      {stage0_32[264], stage0_32[265], stage0_32[266], stage0_32[267], stage0_32[268], stage0_32[269]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[69],stage1_34[89],stage1_33[120],stage1_32[180]}
   );
   gpc606_5 gpc1266 (
      {stage0_32[270], stage0_32[271], stage0_32[272], stage0_32[273], stage0_32[274], stage0_32[275]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[70],stage1_34[90],stage1_33[121],stage1_32[181]}
   );
   gpc606_5 gpc1267 (
      {stage0_32[276], stage0_32[277], stage0_32[278], stage0_32[279], stage0_32[280], stage0_32[281]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[71],stage1_34[91],stage1_33[122],stage1_32[182]}
   );
   gpc606_5 gpc1268 (
      {stage0_32[282], stage0_32[283], stage0_32[284], stage0_32[285], stage0_32[286], stage0_32[287]},
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112], stage0_34[113]},
      {stage1_36[18],stage1_35[72],stage1_34[92],stage1_33[123],stage1_32[183]}
   );
   gpc606_5 gpc1269 (
      {stage0_32[288], stage0_32[289], stage0_32[290], stage0_32[291], stage0_32[292], stage0_32[293]},
      {stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117], stage0_34[118], stage0_34[119]},
      {stage1_36[19],stage1_35[73],stage1_34[93],stage1_33[124],stage1_32[184]}
   );
   gpc606_5 gpc1270 (
      {stage0_32[294], stage0_32[295], stage0_32[296], stage0_32[297], stage0_32[298], stage0_32[299]},
      {stage0_34[120], stage0_34[121], stage0_34[122], stage0_34[123], stage0_34[124], stage0_34[125]},
      {stage1_36[20],stage1_35[74],stage1_34[94],stage1_33[125],stage1_32[185]}
   );
   gpc606_5 gpc1271 (
      {stage0_32[300], stage0_32[301], stage0_32[302], stage0_32[303], stage0_32[304], stage0_32[305]},
      {stage0_34[126], stage0_34[127], stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131]},
      {stage1_36[21],stage1_35[75],stage1_34[95],stage1_33[126],stage1_32[186]}
   );
   gpc606_5 gpc1272 (
      {stage0_32[306], stage0_32[307], stage0_32[308], stage0_32[309], stage0_32[310], stage0_32[311]},
      {stage0_34[132], stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage1_36[22],stage1_35[76],stage1_34[96],stage1_33[127],stage1_32[187]}
   );
   gpc606_5 gpc1273 (
      {stage0_32[312], stage0_32[313], stage0_32[314], stage0_32[315], stage0_32[316], stage0_32[317]},
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142], stage0_34[143]},
      {stage1_36[23],stage1_35[77],stage1_34[97],stage1_33[128],stage1_32[188]}
   );
   gpc606_5 gpc1274 (
      {stage0_32[318], stage0_32[319], stage0_32[320], stage0_32[321], stage0_32[322], stage0_32[323]},
      {stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147], stage0_34[148], stage0_34[149]},
      {stage1_36[24],stage1_35[78],stage1_34[98],stage1_33[129],stage1_32[189]}
   );
   gpc606_5 gpc1275 (
      {stage0_32[324], stage0_32[325], stage0_32[326], stage0_32[327], stage0_32[328], stage0_32[329]},
      {stage0_34[150], stage0_34[151], stage0_34[152], stage0_34[153], stage0_34[154], stage0_34[155]},
      {stage1_36[25],stage1_35[79],stage1_34[99],stage1_33[130],stage1_32[190]}
   );
   gpc606_5 gpc1276 (
      {stage0_32[330], stage0_32[331], stage0_32[332], stage0_32[333], stage0_32[334], stage0_32[335]},
      {stage0_34[156], stage0_34[157], stage0_34[158], stage0_34[159], stage0_34[160], stage0_34[161]},
      {stage1_36[26],stage1_35[80],stage1_34[100],stage1_33[131],stage1_32[191]}
   );
   gpc606_5 gpc1277 (
      {stage0_32[336], stage0_32[337], stage0_32[338], stage0_32[339], stage0_32[340], stage0_32[341]},
      {stage0_34[162], stage0_34[163], stage0_34[164], stage0_34[165], stage0_34[166], stage0_34[167]},
      {stage1_36[27],stage1_35[81],stage1_34[101],stage1_33[132],stage1_32[192]}
   );
   gpc606_5 gpc1278 (
      {stage0_32[342], stage0_32[343], stage0_32[344], stage0_32[345], stage0_32[346], stage0_32[347]},
      {stage0_34[168], stage0_34[169], stage0_34[170], stage0_34[171], stage0_34[172], stage0_34[173]},
      {stage1_36[28],stage1_35[82],stage1_34[102],stage1_33[133],stage1_32[193]}
   );
   gpc606_5 gpc1279 (
      {stage0_32[348], stage0_32[349], stage0_32[350], stage0_32[351], stage0_32[352], stage0_32[353]},
      {stage0_34[174], stage0_34[175], stage0_34[176], stage0_34[177], stage0_34[178], stage0_34[179]},
      {stage1_36[29],stage1_35[83],stage1_34[103],stage1_33[134],stage1_32[194]}
   );
   gpc606_5 gpc1280 (
      {stage0_32[354], stage0_32[355], stage0_32[356], stage0_32[357], stage0_32[358], stage0_32[359]},
      {stage0_34[180], stage0_34[181], stage0_34[182], stage0_34[183], stage0_34[184], stage0_34[185]},
      {stage1_36[30],stage1_35[84],stage1_34[104],stage1_33[135],stage1_32[195]}
   );
   gpc606_5 gpc1281 (
      {stage0_32[360], stage0_32[361], stage0_32[362], stage0_32[363], stage0_32[364], stage0_32[365]},
      {stage0_34[186], stage0_34[187], stage0_34[188], stage0_34[189], stage0_34[190], stage0_34[191]},
      {stage1_36[31],stage1_35[85],stage1_34[105],stage1_33[136],stage1_32[196]}
   );
   gpc606_5 gpc1282 (
      {stage0_32[366], stage0_32[367], stage0_32[368], stage0_32[369], stage0_32[370], stage0_32[371]},
      {stage0_34[192], stage0_34[193], stage0_34[194], stage0_34[195], stage0_34[196], stage0_34[197]},
      {stage1_36[32],stage1_35[86],stage1_34[106],stage1_33[137],stage1_32[197]}
   );
   gpc606_5 gpc1283 (
      {stage0_32[372], stage0_32[373], stage0_32[374], stage0_32[375], stage0_32[376], stage0_32[377]},
      {stage0_34[198], stage0_34[199], stage0_34[200], stage0_34[201], stage0_34[202], stage0_34[203]},
      {stage1_36[33],stage1_35[87],stage1_34[107],stage1_33[138],stage1_32[198]}
   );
   gpc606_5 gpc1284 (
      {stage0_32[378], stage0_32[379], stage0_32[380], stage0_32[381], stage0_32[382], stage0_32[383]},
      {stage0_34[204], stage0_34[205], stage0_34[206], stage0_34[207], stage0_34[208], stage0_34[209]},
      {stage1_36[34],stage1_35[88],stage1_34[108],stage1_33[139],stage1_32[199]}
   );
   gpc606_5 gpc1285 (
      {stage0_32[384], stage0_32[385], stage0_32[386], stage0_32[387], stage0_32[388], stage0_32[389]},
      {stage0_34[210], stage0_34[211], stage0_34[212], stage0_34[213], stage0_34[214], stage0_34[215]},
      {stage1_36[35],stage1_35[89],stage1_34[109],stage1_33[140],stage1_32[200]}
   );
   gpc606_5 gpc1286 (
      {stage0_32[390], stage0_32[391], stage0_32[392], stage0_32[393], stage0_32[394], stage0_32[395]},
      {stage0_34[216], stage0_34[217], stage0_34[218], stage0_34[219], stage0_34[220], stage0_34[221]},
      {stage1_36[36],stage1_35[90],stage1_34[110],stage1_33[141],stage1_32[201]}
   );
   gpc606_5 gpc1287 (
      {stage0_32[396], stage0_32[397], stage0_32[398], stage0_32[399], stage0_32[400], stage0_32[401]},
      {stage0_34[222], stage0_34[223], stage0_34[224], stage0_34[225], stage0_34[226], stage0_34[227]},
      {stage1_36[37],stage1_35[91],stage1_34[111],stage1_33[142],stage1_32[202]}
   );
   gpc606_5 gpc1288 (
      {stage0_32[402], stage0_32[403], stage0_32[404], stage0_32[405], stage0_32[406], stage0_32[407]},
      {stage0_34[228], stage0_34[229], stage0_34[230], stage0_34[231], stage0_34[232], stage0_34[233]},
      {stage1_36[38],stage1_35[92],stage1_34[112],stage1_33[143],stage1_32[203]}
   );
   gpc606_5 gpc1289 (
      {stage0_32[408], stage0_32[409], stage0_32[410], stage0_32[411], stage0_32[412], stage0_32[413]},
      {stage0_34[234], stage0_34[235], stage0_34[236], stage0_34[237], stage0_34[238], stage0_34[239]},
      {stage1_36[39],stage1_35[93],stage1_34[113],stage1_33[144],stage1_32[204]}
   );
   gpc606_5 gpc1290 (
      {stage0_32[414], stage0_32[415], stage0_32[416], stage0_32[417], stage0_32[418], stage0_32[419]},
      {stage0_34[240], stage0_34[241], stage0_34[242], stage0_34[243], stage0_34[244], stage0_34[245]},
      {stage1_36[40],stage1_35[94],stage1_34[114],stage1_33[145],stage1_32[205]}
   );
   gpc606_5 gpc1291 (
      {stage0_32[420], stage0_32[421], stage0_32[422], stage0_32[423], stage0_32[424], stage0_32[425]},
      {stage0_34[246], stage0_34[247], stage0_34[248], stage0_34[249], stage0_34[250], stage0_34[251]},
      {stage1_36[41],stage1_35[95],stage1_34[115],stage1_33[146],stage1_32[206]}
   );
   gpc606_5 gpc1292 (
      {stage0_32[426], stage0_32[427], stage0_32[428], stage0_32[429], stage0_32[430], stage0_32[431]},
      {stage0_34[252], stage0_34[253], stage0_34[254], stage0_34[255], stage0_34[256], stage0_34[257]},
      {stage1_36[42],stage1_35[96],stage1_34[116],stage1_33[147],stage1_32[207]}
   );
   gpc606_5 gpc1293 (
      {stage0_32[432], stage0_32[433], stage0_32[434], stage0_32[435], stage0_32[436], stage0_32[437]},
      {stage0_34[258], stage0_34[259], stage0_34[260], stage0_34[261], stage0_34[262], stage0_34[263]},
      {stage1_36[43],stage1_35[97],stage1_34[117],stage1_33[148],stage1_32[208]}
   );
   gpc606_5 gpc1294 (
      {stage0_32[438], stage0_32[439], stage0_32[440], stage0_32[441], stage0_32[442], stage0_32[443]},
      {stage0_34[264], stage0_34[265], stage0_34[266], stage0_34[267], stage0_34[268], stage0_34[269]},
      {stage1_36[44],stage1_35[98],stage1_34[118],stage1_33[149],stage1_32[209]}
   );
   gpc606_5 gpc1295 (
      {stage0_32[444], stage0_32[445], stage0_32[446], stage0_32[447], stage0_32[448], stage0_32[449]},
      {stage0_34[270], stage0_34[271], stage0_34[272], stage0_34[273], stage0_34[274], stage0_34[275]},
      {stage1_36[45],stage1_35[99],stage1_34[119],stage1_33[150],stage1_32[210]}
   );
   gpc606_5 gpc1296 (
      {stage0_32[450], stage0_32[451], stage0_32[452], stage0_32[453], stage0_32[454], stage0_32[455]},
      {stage0_34[276], stage0_34[277], stage0_34[278], stage0_34[279], stage0_34[280], stage0_34[281]},
      {stage1_36[46],stage1_35[100],stage1_34[120],stage1_33[151],stage1_32[211]}
   );
   gpc606_5 gpc1297 (
      {stage0_32[456], stage0_32[457], stage0_32[458], stage0_32[459], stage0_32[460], stage0_32[461]},
      {stage0_34[282], stage0_34[283], stage0_34[284], stage0_34[285], stage0_34[286], stage0_34[287]},
      {stage1_36[47],stage1_35[101],stage1_34[121],stage1_33[152],stage1_32[212]}
   );
   gpc606_5 gpc1298 (
      {stage0_32[462], stage0_32[463], stage0_32[464], stage0_32[465], stage0_32[466], stage0_32[467]},
      {stage0_34[288], stage0_34[289], stage0_34[290], stage0_34[291], stage0_34[292], stage0_34[293]},
      {stage1_36[48],stage1_35[102],stage1_34[122],stage1_33[153],stage1_32[213]}
   );
   gpc606_5 gpc1299 (
      {stage0_32[468], stage0_32[469], stage0_32[470], stage0_32[471], stage0_32[472], stage0_32[473]},
      {stage0_34[294], stage0_34[295], stage0_34[296], stage0_34[297], stage0_34[298], stage0_34[299]},
      {stage1_36[49],stage1_35[103],stage1_34[123],stage1_33[154],stage1_32[214]}
   );
   gpc606_5 gpc1300 (
      {stage0_32[474], stage0_32[475], stage0_32[476], stage0_32[477], stage0_32[478], stage0_32[479]},
      {stage0_34[300], stage0_34[301], stage0_34[302], stage0_34[303], stage0_34[304], stage0_34[305]},
      {stage1_36[50],stage1_35[104],stage1_34[124],stage1_33[155],stage1_32[215]}
   );
   gpc606_5 gpc1301 (
      {stage0_32[480], stage0_32[481], stage0_32[482], stage0_32[483], stage0_32[484], stage0_32[485]},
      {stage0_34[306], stage0_34[307], stage0_34[308], stage0_34[309], stage0_34[310], stage0_34[311]},
      {stage1_36[51],stage1_35[105],stage1_34[125],stage1_33[156],stage1_32[216]}
   );
   gpc606_5 gpc1302 (
      {stage0_33[324], stage0_33[325], stage0_33[326], stage0_33[327], stage0_33[328], stage0_33[329]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[52],stage1_35[106],stage1_34[126],stage1_33[157]}
   );
   gpc606_5 gpc1303 (
      {stage0_33[330], stage0_33[331], stage0_33[332], stage0_33[333], stage0_33[334], stage0_33[335]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[53],stage1_35[107],stage1_34[127],stage1_33[158]}
   );
   gpc606_5 gpc1304 (
      {stage0_33[336], stage0_33[337], stage0_33[338], stage0_33[339], stage0_33[340], stage0_33[341]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[54],stage1_35[108],stage1_34[128],stage1_33[159]}
   );
   gpc606_5 gpc1305 (
      {stage0_33[342], stage0_33[343], stage0_33[344], stage0_33[345], stage0_33[346], stage0_33[347]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[55],stage1_35[109],stage1_34[129],stage1_33[160]}
   );
   gpc606_5 gpc1306 (
      {stage0_33[348], stage0_33[349], stage0_33[350], stage0_33[351], stage0_33[352], stage0_33[353]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[56],stage1_35[110],stage1_34[130],stage1_33[161]}
   );
   gpc606_5 gpc1307 (
      {stage0_33[354], stage0_33[355], stage0_33[356], stage0_33[357], stage0_33[358], stage0_33[359]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[57],stage1_35[111],stage1_34[131],stage1_33[162]}
   );
   gpc606_5 gpc1308 (
      {stage0_33[360], stage0_33[361], stage0_33[362], stage0_33[363], stage0_33[364], stage0_33[365]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[58],stage1_35[112],stage1_34[132],stage1_33[163]}
   );
   gpc606_5 gpc1309 (
      {stage0_33[366], stage0_33[367], stage0_33[368], stage0_33[369], stage0_33[370], stage0_33[371]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[59],stage1_35[113],stage1_34[133],stage1_33[164]}
   );
   gpc606_5 gpc1310 (
      {stage0_33[372], stage0_33[373], stage0_33[374], stage0_33[375], stage0_33[376], stage0_33[377]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[60],stage1_35[114],stage1_34[134],stage1_33[165]}
   );
   gpc606_5 gpc1311 (
      {stage0_33[378], stage0_33[379], stage0_33[380], stage0_33[381], stage0_33[382], stage0_33[383]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[61],stage1_35[115],stage1_34[135],stage1_33[166]}
   );
   gpc606_5 gpc1312 (
      {stage0_33[384], stage0_33[385], stage0_33[386], stage0_33[387], stage0_33[388], stage0_33[389]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[62],stage1_35[116],stage1_34[136],stage1_33[167]}
   );
   gpc606_5 gpc1313 (
      {stage0_33[390], stage0_33[391], stage0_33[392], stage0_33[393], stage0_33[394], stage0_33[395]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[63],stage1_35[117],stage1_34[137],stage1_33[168]}
   );
   gpc1163_5 gpc1314 (
      {stage0_34[312], stage0_34[313], stage0_34[314]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage0_36[0]},
      {stage0_37[0]},
      {stage1_38[0],stage1_37[12],stage1_36[64],stage1_35[118],stage1_34[138]}
   );
   gpc1163_5 gpc1315 (
      {stage0_34[315], stage0_34[316], stage0_34[317]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage0_36[1]},
      {stage0_37[1]},
      {stage1_38[1],stage1_37[13],stage1_36[65],stage1_35[119],stage1_34[139]}
   );
   gpc1163_5 gpc1316 (
      {stage0_34[318], stage0_34[319], stage0_34[320]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage0_36[2]},
      {stage0_37[2]},
      {stage1_38[2],stage1_37[14],stage1_36[66],stage1_35[120],stage1_34[140]}
   );
   gpc1163_5 gpc1317 (
      {stage0_34[321], stage0_34[322], stage0_34[323]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage0_36[3]},
      {stage0_37[3]},
      {stage1_38[3],stage1_37[15],stage1_36[67],stage1_35[121],stage1_34[141]}
   );
   gpc1163_5 gpc1318 (
      {stage0_34[324], stage0_34[325], stage0_34[326]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage0_36[4]},
      {stage0_37[4]},
      {stage1_38[4],stage1_37[16],stage1_36[68],stage1_35[122],stage1_34[142]}
   );
   gpc1163_5 gpc1319 (
      {stage0_34[327], stage0_34[328], stage0_34[329]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage0_36[5]},
      {stage0_37[5]},
      {stage1_38[5],stage1_37[17],stage1_36[69],stage1_35[123],stage1_34[143]}
   );
   gpc1163_5 gpc1320 (
      {stage0_34[330], stage0_34[331], stage0_34[332]},
      {stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111], stage0_35[112], stage0_35[113]},
      {stage0_36[6]},
      {stage0_37[6]},
      {stage1_38[6],stage1_37[18],stage1_36[70],stage1_35[124],stage1_34[144]}
   );
   gpc1163_5 gpc1321 (
      {stage0_34[333], stage0_34[334], stage0_34[335]},
      {stage0_35[114], stage0_35[115], stage0_35[116], stage0_35[117], stage0_35[118], stage0_35[119]},
      {stage0_36[7]},
      {stage0_37[7]},
      {stage1_38[7],stage1_37[19],stage1_36[71],stage1_35[125],stage1_34[145]}
   );
   gpc1163_5 gpc1322 (
      {stage0_34[336], stage0_34[337], stage0_34[338]},
      {stage0_35[120], stage0_35[121], stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125]},
      {stage0_36[8]},
      {stage0_37[8]},
      {stage1_38[8],stage1_37[20],stage1_36[72],stage1_35[126],stage1_34[146]}
   );
   gpc1163_5 gpc1323 (
      {stage0_34[339], stage0_34[340], stage0_34[341]},
      {stage0_35[126], stage0_35[127], stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131]},
      {stage0_36[9]},
      {stage0_37[9]},
      {stage1_38[9],stage1_37[21],stage1_36[73],stage1_35[127],stage1_34[147]}
   );
   gpc1163_5 gpc1324 (
      {stage0_34[342], stage0_34[343], stage0_34[344]},
      {stage0_35[132], stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage0_36[10]},
      {stage0_37[10]},
      {stage1_38[10],stage1_37[22],stage1_36[74],stage1_35[128],stage1_34[148]}
   );
   gpc1163_5 gpc1325 (
      {stage0_34[345], stage0_34[346], stage0_34[347]},
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142], stage0_35[143]},
      {stage0_36[11]},
      {stage0_37[11]},
      {stage1_38[11],stage1_37[23],stage1_36[75],stage1_35[129],stage1_34[149]}
   );
   gpc1163_5 gpc1326 (
      {stage0_34[348], stage0_34[349], stage0_34[350]},
      {stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147], stage0_35[148], stage0_35[149]},
      {stage0_36[12]},
      {stage0_37[12]},
      {stage1_38[12],stage1_37[24],stage1_36[76],stage1_35[130],stage1_34[150]}
   );
   gpc1163_5 gpc1327 (
      {stage0_34[351], stage0_34[352], stage0_34[353]},
      {stage0_35[150], stage0_35[151], stage0_35[152], stage0_35[153], stage0_35[154], stage0_35[155]},
      {stage0_36[13]},
      {stage0_37[13]},
      {stage1_38[13],stage1_37[25],stage1_36[77],stage1_35[131],stage1_34[151]}
   );
   gpc1163_5 gpc1328 (
      {stage0_34[354], stage0_34[355], stage0_34[356]},
      {stage0_35[156], stage0_35[157], stage0_35[158], stage0_35[159], stage0_35[160], stage0_35[161]},
      {stage0_36[14]},
      {stage0_37[14]},
      {stage1_38[14],stage1_37[26],stage1_36[78],stage1_35[132],stage1_34[152]}
   );
   gpc1163_5 gpc1329 (
      {stage0_34[357], stage0_34[358], stage0_34[359]},
      {stage0_35[162], stage0_35[163], stage0_35[164], stage0_35[165], stage0_35[166], stage0_35[167]},
      {stage0_36[15]},
      {stage0_37[15]},
      {stage1_38[15],stage1_37[27],stage1_36[79],stage1_35[133],stage1_34[153]}
   );
   gpc1163_5 gpc1330 (
      {stage0_34[360], stage0_34[361], stage0_34[362]},
      {stage0_35[168], stage0_35[169], stage0_35[170], stage0_35[171], stage0_35[172], stage0_35[173]},
      {stage0_36[16]},
      {stage0_37[16]},
      {stage1_38[16],stage1_37[28],stage1_36[80],stage1_35[134],stage1_34[154]}
   );
   gpc1163_5 gpc1331 (
      {stage0_34[363], stage0_34[364], stage0_34[365]},
      {stage0_35[174], stage0_35[175], stage0_35[176], stage0_35[177], stage0_35[178], stage0_35[179]},
      {stage0_36[17]},
      {stage0_37[17]},
      {stage1_38[17],stage1_37[29],stage1_36[81],stage1_35[135],stage1_34[155]}
   );
   gpc1163_5 gpc1332 (
      {stage0_34[366], stage0_34[367], stage0_34[368]},
      {stage0_35[180], stage0_35[181], stage0_35[182], stage0_35[183], stage0_35[184], stage0_35[185]},
      {stage0_36[18]},
      {stage0_37[18]},
      {stage1_38[18],stage1_37[30],stage1_36[82],stage1_35[136],stage1_34[156]}
   );
   gpc1163_5 gpc1333 (
      {stage0_34[369], stage0_34[370], stage0_34[371]},
      {stage0_35[186], stage0_35[187], stage0_35[188], stage0_35[189], stage0_35[190], stage0_35[191]},
      {stage0_36[19]},
      {stage0_37[19]},
      {stage1_38[19],stage1_37[31],stage1_36[83],stage1_35[137],stage1_34[157]}
   );
   gpc1163_5 gpc1334 (
      {stage0_34[372], stage0_34[373], stage0_34[374]},
      {stage0_35[192], stage0_35[193], stage0_35[194], stage0_35[195], stage0_35[196], stage0_35[197]},
      {stage0_36[20]},
      {stage0_37[20]},
      {stage1_38[20],stage1_37[32],stage1_36[84],stage1_35[138],stage1_34[158]}
   );
   gpc1163_5 gpc1335 (
      {stage0_34[375], stage0_34[376], stage0_34[377]},
      {stage0_35[198], stage0_35[199], stage0_35[200], stage0_35[201], stage0_35[202], stage0_35[203]},
      {stage0_36[21]},
      {stage0_37[21]},
      {stage1_38[21],stage1_37[33],stage1_36[85],stage1_35[139],stage1_34[159]}
   );
   gpc1163_5 gpc1336 (
      {stage0_34[378], stage0_34[379], stage0_34[380]},
      {stage0_35[204], stage0_35[205], stage0_35[206], stage0_35[207], stage0_35[208], stage0_35[209]},
      {stage0_36[22]},
      {stage0_37[22]},
      {stage1_38[22],stage1_37[34],stage1_36[86],stage1_35[140],stage1_34[160]}
   );
   gpc1163_5 gpc1337 (
      {stage0_34[381], stage0_34[382], stage0_34[383]},
      {stage0_35[210], stage0_35[211], stage0_35[212], stage0_35[213], stage0_35[214], stage0_35[215]},
      {stage0_36[23]},
      {stage0_37[23]},
      {stage1_38[23],stage1_37[35],stage1_36[87],stage1_35[141],stage1_34[161]}
   );
   gpc1163_5 gpc1338 (
      {stage0_34[384], stage0_34[385], stage0_34[386]},
      {stage0_35[216], stage0_35[217], stage0_35[218], stage0_35[219], stage0_35[220], stage0_35[221]},
      {stage0_36[24]},
      {stage0_37[24]},
      {stage1_38[24],stage1_37[36],stage1_36[88],stage1_35[142],stage1_34[162]}
   );
   gpc1163_5 gpc1339 (
      {stage0_34[387], stage0_34[388], stage0_34[389]},
      {stage0_35[222], stage0_35[223], stage0_35[224], stage0_35[225], stage0_35[226], stage0_35[227]},
      {stage0_36[25]},
      {stage0_37[25]},
      {stage1_38[25],stage1_37[37],stage1_36[89],stage1_35[143],stage1_34[163]}
   );
   gpc1163_5 gpc1340 (
      {stage0_34[390], stage0_34[391], stage0_34[392]},
      {stage0_35[228], stage0_35[229], stage0_35[230], stage0_35[231], stage0_35[232], stage0_35[233]},
      {stage0_36[26]},
      {stage0_37[26]},
      {stage1_38[26],stage1_37[38],stage1_36[90],stage1_35[144],stage1_34[164]}
   );
   gpc1163_5 gpc1341 (
      {stage0_34[393], stage0_34[394], stage0_34[395]},
      {stage0_35[234], stage0_35[235], stage0_35[236], stage0_35[237], stage0_35[238], stage0_35[239]},
      {stage0_36[27]},
      {stage0_37[27]},
      {stage1_38[27],stage1_37[39],stage1_36[91],stage1_35[145],stage1_34[165]}
   );
   gpc1163_5 gpc1342 (
      {stage0_34[396], stage0_34[397], stage0_34[398]},
      {stage0_35[240], stage0_35[241], stage0_35[242], stage0_35[243], stage0_35[244], stage0_35[245]},
      {stage0_36[28]},
      {stage0_37[28]},
      {stage1_38[28],stage1_37[40],stage1_36[92],stage1_35[146],stage1_34[166]}
   );
   gpc1163_5 gpc1343 (
      {stage0_34[399], stage0_34[400], stage0_34[401]},
      {stage0_35[246], stage0_35[247], stage0_35[248], stage0_35[249], stage0_35[250], stage0_35[251]},
      {stage0_36[29]},
      {stage0_37[29]},
      {stage1_38[29],stage1_37[41],stage1_36[93],stage1_35[147],stage1_34[167]}
   );
   gpc1163_5 gpc1344 (
      {stage0_34[402], stage0_34[403], stage0_34[404]},
      {stage0_35[252], stage0_35[253], stage0_35[254], stage0_35[255], stage0_35[256], stage0_35[257]},
      {stage0_36[30]},
      {stage0_37[30]},
      {stage1_38[30],stage1_37[42],stage1_36[94],stage1_35[148],stage1_34[168]}
   );
   gpc1163_5 gpc1345 (
      {stage0_34[405], stage0_34[406], stage0_34[407]},
      {stage0_35[258], stage0_35[259], stage0_35[260], stage0_35[261], stage0_35[262], stage0_35[263]},
      {stage0_36[31]},
      {stage0_37[31]},
      {stage1_38[31],stage1_37[43],stage1_36[95],stage1_35[149],stage1_34[169]}
   );
   gpc1163_5 gpc1346 (
      {stage0_34[408], stage0_34[409], stage0_34[410]},
      {stage0_35[264], stage0_35[265], stage0_35[266], stage0_35[267], stage0_35[268], stage0_35[269]},
      {stage0_36[32]},
      {stage0_37[32]},
      {stage1_38[32],stage1_37[44],stage1_36[96],stage1_35[150],stage1_34[170]}
   );
   gpc1163_5 gpc1347 (
      {stage0_34[411], stage0_34[412], stage0_34[413]},
      {stage0_35[270], stage0_35[271], stage0_35[272], stage0_35[273], stage0_35[274], stage0_35[275]},
      {stage0_36[33]},
      {stage0_37[33]},
      {stage1_38[33],stage1_37[45],stage1_36[97],stage1_35[151],stage1_34[171]}
   );
   gpc1163_5 gpc1348 (
      {stage0_34[414], stage0_34[415], stage0_34[416]},
      {stage0_35[276], stage0_35[277], stage0_35[278], stage0_35[279], stage0_35[280], stage0_35[281]},
      {stage0_36[34]},
      {stage0_37[34]},
      {stage1_38[34],stage1_37[46],stage1_36[98],stage1_35[152],stage1_34[172]}
   );
   gpc1163_5 gpc1349 (
      {stage0_34[417], stage0_34[418], stage0_34[419]},
      {stage0_35[282], stage0_35[283], stage0_35[284], stage0_35[285], stage0_35[286], stage0_35[287]},
      {stage0_36[35]},
      {stage0_37[35]},
      {stage1_38[35],stage1_37[47],stage1_36[99],stage1_35[153],stage1_34[173]}
   );
   gpc1163_5 gpc1350 (
      {stage0_34[420], stage0_34[421], stage0_34[422]},
      {stage0_35[288], stage0_35[289], stage0_35[290], stage0_35[291], stage0_35[292], stage0_35[293]},
      {stage0_36[36]},
      {stage0_37[36]},
      {stage1_38[36],stage1_37[48],stage1_36[100],stage1_35[154],stage1_34[174]}
   );
   gpc1163_5 gpc1351 (
      {stage0_34[423], stage0_34[424], stage0_34[425]},
      {stage0_35[294], stage0_35[295], stage0_35[296], stage0_35[297], stage0_35[298], stage0_35[299]},
      {stage0_36[37]},
      {stage0_37[37]},
      {stage1_38[37],stage1_37[49],stage1_36[101],stage1_35[155],stage1_34[175]}
   );
   gpc1163_5 gpc1352 (
      {stage0_34[426], stage0_34[427], stage0_34[428]},
      {stage0_35[300], stage0_35[301], stage0_35[302], stage0_35[303], stage0_35[304], stage0_35[305]},
      {stage0_36[38]},
      {stage0_37[38]},
      {stage1_38[38],stage1_37[50],stage1_36[102],stage1_35[156],stage1_34[176]}
   );
   gpc1163_5 gpc1353 (
      {stage0_34[429], stage0_34[430], stage0_34[431]},
      {stage0_35[306], stage0_35[307], stage0_35[308], stage0_35[309], stage0_35[310], stage0_35[311]},
      {stage0_36[39]},
      {stage0_37[39]},
      {stage1_38[39],stage1_37[51],stage1_36[103],stage1_35[157],stage1_34[177]}
   );
   gpc1163_5 gpc1354 (
      {stage0_34[432], stage0_34[433], stage0_34[434]},
      {stage0_35[312], stage0_35[313], stage0_35[314], stage0_35[315], stage0_35[316], stage0_35[317]},
      {stage0_36[40]},
      {stage0_37[40]},
      {stage1_38[40],stage1_37[52],stage1_36[104],stage1_35[158],stage1_34[178]}
   );
   gpc1163_5 gpc1355 (
      {stage0_34[435], stage0_34[436], stage0_34[437]},
      {stage0_35[318], stage0_35[319], stage0_35[320], stage0_35[321], stage0_35[322], stage0_35[323]},
      {stage0_36[41]},
      {stage0_37[41]},
      {stage1_38[41],stage1_37[53],stage1_36[105],stage1_35[159],stage1_34[179]}
   );
   gpc1163_5 gpc1356 (
      {stage0_34[438], stage0_34[439], stage0_34[440]},
      {stage0_35[324], stage0_35[325], stage0_35[326], stage0_35[327], stage0_35[328], stage0_35[329]},
      {stage0_36[42]},
      {stage0_37[42]},
      {stage1_38[42],stage1_37[54],stage1_36[106],stage1_35[160],stage1_34[180]}
   );
   gpc615_5 gpc1357 (
      {stage0_34[441], stage0_34[442], stage0_34[443], stage0_34[444], stage0_34[445]},
      {stage0_35[330]},
      {stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47], stage0_36[48]},
      {stage1_38[43],stage1_37[55],stage1_36[107],stage1_35[161],stage1_34[181]}
   );
   gpc615_5 gpc1358 (
      {stage0_34[446], stage0_34[447], stage0_34[448], stage0_34[449], stage0_34[450]},
      {stage0_35[331]},
      {stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53], stage0_36[54]},
      {stage1_38[44],stage1_37[56],stage1_36[108],stage1_35[162],stage1_34[182]}
   );
   gpc615_5 gpc1359 (
      {stage0_34[451], stage0_34[452], stage0_34[453], stage0_34[454], stage0_34[455]},
      {stage0_35[332]},
      {stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59], stage0_36[60]},
      {stage1_38[45],stage1_37[57],stage1_36[109],stage1_35[163],stage1_34[183]}
   );
   gpc615_5 gpc1360 (
      {stage0_34[456], stage0_34[457], stage0_34[458], stage0_34[459], stage0_34[460]},
      {stage0_35[333]},
      {stage0_36[61], stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65], stage0_36[66]},
      {stage1_38[46],stage1_37[58],stage1_36[110],stage1_35[164],stage1_34[184]}
   );
   gpc615_5 gpc1361 (
      {stage0_34[461], stage0_34[462], stage0_34[463], stage0_34[464], stage0_34[465]},
      {stage0_35[334]},
      {stage0_36[67], stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71], stage0_36[72]},
      {stage1_38[47],stage1_37[59],stage1_36[111],stage1_35[165],stage1_34[185]}
   );
   gpc615_5 gpc1362 (
      {stage0_34[466], stage0_34[467], stage0_34[468], stage0_34[469], stage0_34[470]},
      {stage0_35[335]},
      {stage0_36[73], stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77], stage0_36[78]},
      {stage1_38[48],stage1_37[60],stage1_36[112],stage1_35[166],stage1_34[186]}
   );
   gpc615_5 gpc1363 (
      {stage0_34[471], stage0_34[472], stage0_34[473], stage0_34[474], stage0_34[475]},
      {stage0_35[336]},
      {stage0_36[79], stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83], stage0_36[84]},
      {stage1_38[49],stage1_37[61],stage1_36[113],stage1_35[167],stage1_34[187]}
   );
   gpc615_5 gpc1364 (
      {stage0_34[476], stage0_34[477], stage0_34[478], stage0_34[479], stage0_34[480]},
      {stage0_35[337]},
      {stage0_36[85], stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89], stage0_36[90]},
      {stage1_38[50],stage1_37[62],stage1_36[114],stage1_35[168],stage1_34[188]}
   );
   gpc615_5 gpc1365 (
      {stage0_34[481], stage0_34[482], stage0_34[483], stage0_34[484], stage0_34[485]},
      {stage0_35[338]},
      {stage0_36[91], stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95], stage0_36[96]},
      {stage1_38[51],stage1_37[63],stage1_36[115],stage1_35[169],stage1_34[189]}
   );
   gpc615_5 gpc1366 (
      {stage0_35[339], stage0_35[340], stage0_35[341], stage0_35[342], stage0_35[343]},
      {stage0_36[97]},
      {stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47], stage0_37[48]},
      {stage1_39[0],stage1_38[52],stage1_37[64],stage1_36[116],stage1_35[170]}
   );
   gpc615_5 gpc1367 (
      {stage0_35[344], stage0_35[345], stage0_35[346], stage0_35[347], stage0_35[348]},
      {stage0_36[98]},
      {stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53], stage0_37[54]},
      {stage1_39[1],stage1_38[53],stage1_37[65],stage1_36[117],stage1_35[171]}
   );
   gpc615_5 gpc1368 (
      {stage0_35[349], stage0_35[350], stage0_35[351], stage0_35[352], stage0_35[353]},
      {stage0_36[99]},
      {stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59], stage0_37[60]},
      {stage1_39[2],stage1_38[54],stage1_37[66],stage1_36[118],stage1_35[172]}
   );
   gpc615_5 gpc1369 (
      {stage0_35[354], stage0_35[355], stage0_35[356], stage0_35[357], stage0_35[358]},
      {stage0_36[100]},
      {stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65], stage0_37[66]},
      {stage1_39[3],stage1_38[55],stage1_37[67],stage1_36[119],stage1_35[173]}
   );
   gpc615_5 gpc1370 (
      {stage0_35[359], stage0_35[360], stage0_35[361], stage0_35[362], stage0_35[363]},
      {stage0_36[101]},
      {stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71], stage0_37[72]},
      {stage1_39[4],stage1_38[56],stage1_37[68],stage1_36[120],stage1_35[174]}
   );
   gpc615_5 gpc1371 (
      {stage0_35[364], stage0_35[365], stage0_35[366], stage0_35[367], stage0_35[368]},
      {stage0_36[102]},
      {stage0_37[73], stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77], stage0_37[78]},
      {stage1_39[5],stage1_38[57],stage1_37[69],stage1_36[121],stage1_35[175]}
   );
   gpc615_5 gpc1372 (
      {stage0_35[369], stage0_35[370], stage0_35[371], stage0_35[372], stage0_35[373]},
      {stage0_36[103]},
      {stage0_37[79], stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83], stage0_37[84]},
      {stage1_39[6],stage1_38[58],stage1_37[70],stage1_36[122],stage1_35[176]}
   );
   gpc615_5 gpc1373 (
      {stage0_35[374], stage0_35[375], stage0_35[376], stage0_35[377], stage0_35[378]},
      {stage0_36[104]},
      {stage0_37[85], stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89], stage0_37[90]},
      {stage1_39[7],stage1_38[59],stage1_37[71],stage1_36[123],stage1_35[177]}
   );
   gpc615_5 gpc1374 (
      {stage0_35[379], stage0_35[380], stage0_35[381], stage0_35[382], stage0_35[383]},
      {stage0_36[105]},
      {stage0_37[91], stage0_37[92], stage0_37[93], stage0_37[94], stage0_37[95], stage0_37[96]},
      {stage1_39[8],stage1_38[60],stage1_37[72],stage1_36[124],stage1_35[178]}
   );
   gpc615_5 gpc1375 (
      {stage0_35[384], stage0_35[385], stage0_35[386], stage0_35[387], stage0_35[388]},
      {stage0_36[106]},
      {stage0_37[97], stage0_37[98], stage0_37[99], stage0_37[100], stage0_37[101], stage0_37[102]},
      {stage1_39[9],stage1_38[61],stage1_37[73],stage1_36[125],stage1_35[179]}
   );
   gpc615_5 gpc1376 (
      {stage0_35[389], stage0_35[390], stage0_35[391], stage0_35[392], stage0_35[393]},
      {stage0_36[107]},
      {stage0_37[103], stage0_37[104], stage0_37[105], stage0_37[106], stage0_37[107], stage0_37[108]},
      {stage1_39[10],stage1_38[62],stage1_37[74],stage1_36[126],stage1_35[180]}
   );
   gpc615_5 gpc1377 (
      {stage0_35[394], stage0_35[395], stage0_35[396], stage0_35[397], stage0_35[398]},
      {stage0_36[108]},
      {stage0_37[109], stage0_37[110], stage0_37[111], stage0_37[112], stage0_37[113], stage0_37[114]},
      {stage1_39[11],stage1_38[63],stage1_37[75],stage1_36[127],stage1_35[181]}
   );
   gpc615_5 gpc1378 (
      {stage0_35[399], stage0_35[400], stage0_35[401], stage0_35[402], stage0_35[403]},
      {stage0_36[109]},
      {stage0_37[115], stage0_37[116], stage0_37[117], stage0_37[118], stage0_37[119], stage0_37[120]},
      {stage1_39[12],stage1_38[64],stage1_37[76],stage1_36[128],stage1_35[182]}
   );
   gpc615_5 gpc1379 (
      {stage0_35[404], stage0_35[405], stage0_35[406], stage0_35[407], stage0_35[408]},
      {stage0_36[110]},
      {stage0_37[121], stage0_37[122], stage0_37[123], stage0_37[124], stage0_37[125], stage0_37[126]},
      {stage1_39[13],stage1_38[65],stage1_37[77],stage1_36[129],stage1_35[183]}
   );
   gpc615_5 gpc1380 (
      {stage0_35[409], stage0_35[410], stage0_35[411], stage0_35[412], stage0_35[413]},
      {stage0_36[111]},
      {stage0_37[127], stage0_37[128], stage0_37[129], stage0_37[130], stage0_37[131], stage0_37[132]},
      {stage1_39[14],stage1_38[66],stage1_37[78],stage1_36[130],stage1_35[184]}
   );
   gpc615_5 gpc1381 (
      {stage0_35[414], stage0_35[415], stage0_35[416], stage0_35[417], stage0_35[418]},
      {stage0_36[112]},
      {stage0_37[133], stage0_37[134], stage0_37[135], stage0_37[136], stage0_37[137], stage0_37[138]},
      {stage1_39[15],stage1_38[67],stage1_37[79],stage1_36[131],stage1_35[185]}
   );
   gpc615_5 gpc1382 (
      {stage0_35[419], stage0_35[420], stage0_35[421], stage0_35[422], stage0_35[423]},
      {stage0_36[113]},
      {stage0_37[139], stage0_37[140], stage0_37[141], stage0_37[142], stage0_37[143], stage0_37[144]},
      {stage1_39[16],stage1_38[68],stage1_37[80],stage1_36[132],stage1_35[186]}
   );
   gpc615_5 gpc1383 (
      {stage0_35[424], stage0_35[425], stage0_35[426], stage0_35[427], stage0_35[428]},
      {stage0_36[114]},
      {stage0_37[145], stage0_37[146], stage0_37[147], stage0_37[148], stage0_37[149], stage0_37[150]},
      {stage1_39[17],stage1_38[69],stage1_37[81],stage1_36[133],stage1_35[187]}
   );
   gpc615_5 gpc1384 (
      {stage0_35[429], stage0_35[430], stage0_35[431], stage0_35[432], stage0_35[433]},
      {stage0_36[115]},
      {stage0_37[151], stage0_37[152], stage0_37[153], stage0_37[154], stage0_37[155], stage0_37[156]},
      {stage1_39[18],stage1_38[70],stage1_37[82],stage1_36[134],stage1_35[188]}
   );
   gpc615_5 gpc1385 (
      {stage0_35[434], stage0_35[435], stage0_35[436], stage0_35[437], stage0_35[438]},
      {stage0_36[116]},
      {stage0_37[157], stage0_37[158], stage0_37[159], stage0_37[160], stage0_37[161], stage0_37[162]},
      {stage1_39[19],stage1_38[71],stage1_37[83],stage1_36[135],stage1_35[189]}
   );
   gpc615_5 gpc1386 (
      {stage0_35[439], stage0_35[440], stage0_35[441], stage0_35[442], stage0_35[443]},
      {stage0_36[117]},
      {stage0_37[163], stage0_37[164], stage0_37[165], stage0_37[166], stage0_37[167], stage0_37[168]},
      {stage1_39[20],stage1_38[72],stage1_37[84],stage1_36[136],stage1_35[190]}
   );
   gpc615_5 gpc1387 (
      {stage0_35[444], stage0_35[445], stage0_35[446], stage0_35[447], stage0_35[448]},
      {stage0_36[118]},
      {stage0_37[169], stage0_37[170], stage0_37[171], stage0_37[172], stage0_37[173], stage0_37[174]},
      {stage1_39[21],stage1_38[73],stage1_37[85],stage1_36[137],stage1_35[191]}
   );
   gpc615_5 gpc1388 (
      {stage0_35[449], stage0_35[450], stage0_35[451], stage0_35[452], stage0_35[453]},
      {stage0_36[119]},
      {stage0_37[175], stage0_37[176], stage0_37[177], stage0_37[178], stage0_37[179], stage0_37[180]},
      {stage1_39[22],stage1_38[74],stage1_37[86],stage1_36[138],stage1_35[192]}
   );
   gpc615_5 gpc1389 (
      {stage0_35[454], stage0_35[455], stage0_35[456], stage0_35[457], stage0_35[458]},
      {stage0_36[120]},
      {stage0_37[181], stage0_37[182], stage0_37[183], stage0_37[184], stage0_37[185], stage0_37[186]},
      {stage1_39[23],stage1_38[75],stage1_37[87],stage1_36[139],stage1_35[193]}
   );
   gpc615_5 gpc1390 (
      {stage0_35[459], stage0_35[460], stage0_35[461], stage0_35[462], stage0_35[463]},
      {stage0_36[121]},
      {stage0_37[187], stage0_37[188], stage0_37[189], stage0_37[190], stage0_37[191], stage0_37[192]},
      {stage1_39[24],stage1_38[76],stage1_37[88],stage1_36[140],stage1_35[194]}
   );
   gpc606_5 gpc1391 (
      {stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126], stage0_36[127]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[25],stage1_38[77],stage1_37[89],stage1_36[141]}
   );
   gpc606_5 gpc1392 (
      {stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132], stage0_36[133]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[26],stage1_38[78],stage1_37[90],stage1_36[142]}
   );
   gpc606_5 gpc1393 (
      {stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138], stage0_36[139]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[27],stage1_38[79],stage1_37[91],stage1_36[143]}
   );
   gpc606_5 gpc1394 (
      {stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144], stage0_36[145]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[28],stage1_38[80],stage1_37[92],stage1_36[144]}
   );
   gpc606_5 gpc1395 (
      {stage0_36[146], stage0_36[147], stage0_36[148], stage0_36[149], stage0_36[150], stage0_36[151]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[29],stage1_38[81],stage1_37[93],stage1_36[145]}
   );
   gpc606_5 gpc1396 (
      {stage0_36[152], stage0_36[153], stage0_36[154], stage0_36[155], stage0_36[156], stage0_36[157]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[30],stage1_38[82],stage1_37[94],stage1_36[146]}
   );
   gpc606_5 gpc1397 (
      {stage0_36[158], stage0_36[159], stage0_36[160], stage0_36[161], stage0_36[162], stage0_36[163]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[31],stage1_38[83],stage1_37[95],stage1_36[147]}
   );
   gpc606_5 gpc1398 (
      {stage0_36[164], stage0_36[165], stage0_36[166], stage0_36[167], stage0_36[168], stage0_36[169]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[32],stage1_38[84],stage1_37[96],stage1_36[148]}
   );
   gpc606_5 gpc1399 (
      {stage0_36[170], stage0_36[171], stage0_36[172], stage0_36[173], stage0_36[174], stage0_36[175]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[33],stage1_38[85],stage1_37[97],stage1_36[149]}
   );
   gpc606_5 gpc1400 (
      {stage0_36[176], stage0_36[177], stage0_36[178], stage0_36[179], stage0_36[180], stage0_36[181]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[34],stage1_38[86],stage1_37[98],stage1_36[150]}
   );
   gpc606_5 gpc1401 (
      {stage0_36[182], stage0_36[183], stage0_36[184], stage0_36[185], stage0_36[186], stage0_36[187]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[35],stage1_38[87],stage1_37[99],stage1_36[151]}
   );
   gpc606_5 gpc1402 (
      {stage0_36[188], stage0_36[189], stage0_36[190], stage0_36[191], stage0_36[192], stage0_36[193]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[36],stage1_38[88],stage1_37[100],stage1_36[152]}
   );
   gpc606_5 gpc1403 (
      {stage0_36[194], stage0_36[195], stage0_36[196], stage0_36[197], stage0_36[198], stage0_36[199]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[37],stage1_38[89],stage1_37[101],stage1_36[153]}
   );
   gpc606_5 gpc1404 (
      {stage0_36[200], stage0_36[201], stage0_36[202], stage0_36[203], stage0_36[204], stage0_36[205]},
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83]},
      {stage1_40[13],stage1_39[38],stage1_38[90],stage1_37[102],stage1_36[154]}
   );
   gpc606_5 gpc1405 (
      {stage0_36[206], stage0_36[207], stage0_36[208], stage0_36[209], stage0_36[210], stage0_36[211]},
      {stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89]},
      {stage1_40[14],stage1_39[39],stage1_38[91],stage1_37[103],stage1_36[155]}
   );
   gpc606_5 gpc1406 (
      {stage0_36[212], stage0_36[213], stage0_36[214], stage0_36[215], stage0_36[216], stage0_36[217]},
      {stage0_38[90], stage0_38[91], stage0_38[92], stage0_38[93], stage0_38[94], stage0_38[95]},
      {stage1_40[15],stage1_39[40],stage1_38[92],stage1_37[104],stage1_36[156]}
   );
   gpc606_5 gpc1407 (
      {stage0_36[218], stage0_36[219], stage0_36[220], stage0_36[221], stage0_36[222], stage0_36[223]},
      {stage0_38[96], stage0_38[97], stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101]},
      {stage1_40[16],stage1_39[41],stage1_38[93],stage1_37[105],stage1_36[157]}
   );
   gpc606_5 gpc1408 (
      {stage0_36[224], stage0_36[225], stage0_36[226], stage0_36[227], stage0_36[228], stage0_36[229]},
      {stage0_38[102], stage0_38[103], stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107]},
      {stage1_40[17],stage1_39[42],stage1_38[94],stage1_37[106],stage1_36[158]}
   );
   gpc606_5 gpc1409 (
      {stage0_36[230], stage0_36[231], stage0_36[232], stage0_36[233], stage0_36[234], stage0_36[235]},
      {stage0_38[108], stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113]},
      {stage1_40[18],stage1_39[43],stage1_38[95],stage1_37[107],stage1_36[159]}
   );
   gpc606_5 gpc1410 (
      {stage0_36[236], stage0_36[237], stage0_36[238], stage0_36[239], stage0_36[240], stage0_36[241]},
      {stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118], stage0_38[119]},
      {stage1_40[19],stage1_39[44],stage1_38[96],stage1_37[108],stage1_36[160]}
   );
   gpc606_5 gpc1411 (
      {stage0_36[242], stage0_36[243], stage0_36[244], stage0_36[245], stage0_36[246], stage0_36[247]},
      {stage0_38[120], stage0_38[121], stage0_38[122], stage0_38[123], stage0_38[124], stage0_38[125]},
      {stage1_40[20],stage1_39[45],stage1_38[97],stage1_37[109],stage1_36[161]}
   );
   gpc606_5 gpc1412 (
      {stage0_36[248], stage0_36[249], stage0_36[250], stage0_36[251], stage0_36[252], stage0_36[253]},
      {stage0_38[126], stage0_38[127], stage0_38[128], stage0_38[129], stage0_38[130], stage0_38[131]},
      {stage1_40[21],stage1_39[46],stage1_38[98],stage1_37[110],stage1_36[162]}
   );
   gpc606_5 gpc1413 (
      {stage0_36[254], stage0_36[255], stage0_36[256], stage0_36[257], stage0_36[258], stage0_36[259]},
      {stage0_38[132], stage0_38[133], stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137]},
      {stage1_40[22],stage1_39[47],stage1_38[99],stage1_37[111],stage1_36[163]}
   );
   gpc606_5 gpc1414 (
      {stage0_36[260], stage0_36[261], stage0_36[262], stage0_36[263], stage0_36[264], stage0_36[265]},
      {stage0_38[138], stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142], stage0_38[143]},
      {stage1_40[23],stage1_39[48],stage1_38[100],stage1_37[112],stage1_36[164]}
   );
   gpc606_5 gpc1415 (
      {stage0_36[266], stage0_36[267], stage0_36[268], stage0_36[269], stage0_36[270], stage0_36[271]},
      {stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147], stage0_38[148], stage0_38[149]},
      {stage1_40[24],stage1_39[49],stage1_38[101],stage1_37[113],stage1_36[165]}
   );
   gpc606_5 gpc1416 (
      {stage0_36[272], stage0_36[273], stage0_36[274], stage0_36[275], stage0_36[276], stage0_36[277]},
      {stage0_38[150], stage0_38[151], stage0_38[152], stage0_38[153], stage0_38[154], stage0_38[155]},
      {stage1_40[25],stage1_39[50],stage1_38[102],stage1_37[114],stage1_36[166]}
   );
   gpc606_5 gpc1417 (
      {stage0_36[278], stage0_36[279], stage0_36[280], stage0_36[281], stage0_36[282], stage0_36[283]},
      {stage0_38[156], stage0_38[157], stage0_38[158], stage0_38[159], stage0_38[160], stage0_38[161]},
      {stage1_40[26],stage1_39[51],stage1_38[103],stage1_37[115],stage1_36[167]}
   );
   gpc606_5 gpc1418 (
      {stage0_36[284], stage0_36[285], stage0_36[286], stage0_36[287], stage0_36[288], stage0_36[289]},
      {stage0_38[162], stage0_38[163], stage0_38[164], stage0_38[165], stage0_38[166], stage0_38[167]},
      {stage1_40[27],stage1_39[52],stage1_38[104],stage1_37[116],stage1_36[168]}
   );
   gpc606_5 gpc1419 (
      {stage0_36[290], stage0_36[291], stage0_36[292], stage0_36[293], stage0_36[294], stage0_36[295]},
      {stage0_38[168], stage0_38[169], stage0_38[170], stage0_38[171], stage0_38[172], stage0_38[173]},
      {stage1_40[28],stage1_39[53],stage1_38[105],stage1_37[117],stage1_36[169]}
   );
   gpc606_5 gpc1420 (
      {stage0_36[296], stage0_36[297], stage0_36[298], stage0_36[299], stage0_36[300], stage0_36[301]},
      {stage0_38[174], stage0_38[175], stage0_38[176], stage0_38[177], stage0_38[178], stage0_38[179]},
      {stage1_40[29],stage1_39[54],stage1_38[106],stage1_37[118],stage1_36[170]}
   );
   gpc606_5 gpc1421 (
      {stage0_36[302], stage0_36[303], stage0_36[304], stage0_36[305], stage0_36[306], stage0_36[307]},
      {stage0_38[180], stage0_38[181], stage0_38[182], stage0_38[183], stage0_38[184], stage0_38[185]},
      {stage1_40[30],stage1_39[55],stage1_38[107],stage1_37[119],stage1_36[171]}
   );
   gpc606_5 gpc1422 (
      {stage0_36[308], stage0_36[309], stage0_36[310], stage0_36[311], stage0_36[312], stage0_36[313]},
      {stage0_38[186], stage0_38[187], stage0_38[188], stage0_38[189], stage0_38[190], stage0_38[191]},
      {stage1_40[31],stage1_39[56],stage1_38[108],stage1_37[120],stage1_36[172]}
   );
   gpc606_5 gpc1423 (
      {stage0_36[314], stage0_36[315], stage0_36[316], stage0_36[317], stage0_36[318], stage0_36[319]},
      {stage0_38[192], stage0_38[193], stage0_38[194], stage0_38[195], stage0_38[196], stage0_38[197]},
      {stage1_40[32],stage1_39[57],stage1_38[109],stage1_37[121],stage1_36[173]}
   );
   gpc606_5 gpc1424 (
      {stage0_36[320], stage0_36[321], stage0_36[322], stage0_36[323], stage0_36[324], stage0_36[325]},
      {stage0_38[198], stage0_38[199], stage0_38[200], stage0_38[201], stage0_38[202], stage0_38[203]},
      {stage1_40[33],stage1_39[58],stage1_38[110],stage1_37[122],stage1_36[174]}
   );
   gpc606_5 gpc1425 (
      {stage0_36[326], stage0_36[327], stage0_36[328], stage0_36[329], stage0_36[330], stage0_36[331]},
      {stage0_38[204], stage0_38[205], stage0_38[206], stage0_38[207], stage0_38[208], stage0_38[209]},
      {stage1_40[34],stage1_39[59],stage1_38[111],stage1_37[123],stage1_36[175]}
   );
   gpc606_5 gpc1426 (
      {stage0_36[332], stage0_36[333], stage0_36[334], stage0_36[335], stage0_36[336], stage0_36[337]},
      {stage0_38[210], stage0_38[211], stage0_38[212], stage0_38[213], stage0_38[214], stage0_38[215]},
      {stage1_40[35],stage1_39[60],stage1_38[112],stage1_37[124],stage1_36[176]}
   );
   gpc606_5 gpc1427 (
      {stage0_36[338], stage0_36[339], stage0_36[340], stage0_36[341], stage0_36[342], stage0_36[343]},
      {stage0_38[216], stage0_38[217], stage0_38[218], stage0_38[219], stage0_38[220], stage0_38[221]},
      {stage1_40[36],stage1_39[61],stage1_38[113],stage1_37[125],stage1_36[177]}
   );
   gpc606_5 gpc1428 (
      {stage0_36[344], stage0_36[345], stage0_36[346], stage0_36[347], stage0_36[348], stage0_36[349]},
      {stage0_38[222], stage0_38[223], stage0_38[224], stage0_38[225], stage0_38[226], stage0_38[227]},
      {stage1_40[37],stage1_39[62],stage1_38[114],stage1_37[126],stage1_36[178]}
   );
   gpc606_5 gpc1429 (
      {stage0_36[350], stage0_36[351], stage0_36[352], stage0_36[353], stage0_36[354], stage0_36[355]},
      {stage0_38[228], stage0_38[229], stage0_38[230], stage0_38[231], stage0_38[232], stage0_38[233]},
      {stage1_40[38],stage1_39[63],stage1_38[115],stage1_37[127],stage1_36[179]}
   );
   gpc606_5 gpc1430 (
      {stage0_36[356], stage0_36[357], stage0_36[358], stage0_36[359], stage0_36[360], stage0_36[361]},
      {stage0_38[234], stage0_38[235], stage0_38[236], stage0_38[237], stage0_38[238], stage0_38[239]},
      {stage1_40[39],stage1_39[64],stage1_38[116],stage1_37[128],stage1_36[180]}
   );
   gpc606_5 gpc1431 (
      {stage0_36[362], stage0_36[363], stage0_36[364], stage0_36[365], stage0_36[366], stage0_36[367]},
      {stage0_38[240], stage0_38[241], stage0_38[242], stage0_38[243], stage0_38[244], stage0_38[245]},
      {stage1_40[40],stage1_39[65],stage1_38[117],stage1_37[129],stage1_36[181]}
   );
   gpc606_5 gpc1432 (
      {stage0_36[368], stage0_36[369], stage0_36[370], stage0_36[371], stage0_36[372], stage0_36[373]},
      {stage0_38[246], stage0_38[247], stage0_38[248], stage0_38[249], stage0_38[250], stage0_38[251]},
      {stage1_40[41],stage1_39[66],stage1_38[118],stage1_37[130],stage1_36[182]}
   );
   gpc606_5 gpc1433 (
      {stage0_36[374], stage0_36[375], stage0_36[376], stage0_36[377], stage0_36[378], stage0_36[379]},
      {stage0_38[252], stage0_38[253], stage0_38[254], stage0_38[255], stage0_38[256], stage0_38[257]},
      {stage1_40[42],stage1_39[67],stage1_38[119],stage1_37[131],stage1_36[183]}
   );
   gpc606_5 gpc1434 (
      {stage0_36[380], stage0_36[381], stage0_36[382], stage0_36[383], stage0_36[384], stage0_36[385]},
      {stage0_38[258], stage0_38[259], stage0_38[260], stage0_38[261], stage0_38[262], stage0_38[263]},
      {stage1_40[43],stage1_39[68],stage1_38[120],stage1_37[132],stage1_36[184]}
   );
   gpc606_5 gpc1435 (
      {stage0_36[386], stage0_36[387], stage0_36[388], stage0_36[389], stage0_36[390], stage0_36[391]},
      {stage0_38[264], stage0_38[265], stage0_38[266], stage0_38[267], stage0_38[268], stage0_38[269]},
      {stage1_40[44],stage1_39[69],stage1_38[121],stage1_37[133],stage1_36[185]}
   );
   gpc606_5 gpc1436 (
      {stage0_36[392], stage0_36[393], stage0_36[394], stage0_36[395], stage0_36[396], stage0_36[397]},
      {stage0_38[270], stage0_38[271], stage0_38[272], stage0_38[273], stage0_38[274], stage0_38[275]},
      {stage1_40[45],stage1_39[70],stage1_38[122],stage1_37[134],stage1_36[186]}
   );
   gpc606_5 gpc1437 (
      {stage0_36[398], stage0_36[399], stage0_36[400], stage0_36[401], stage0_36[402], stage0_36[403]},
      {stage0_38[276], stage0_38[277], stage0_38[278], stage0_38[279], stage0_38[280], stage0_38[281]},
      {stage1_40[46],stage1_39[71],stage1_38[123],stage1_37[135],stage1_36[187]}
   );
   gpc606_5 gpc1438 (
      {stage0_36[404], stage0_36[405], stage0_36[406], stage0_36[407], stage0_36[408], stage0_36[409]},
      {stage0_38[282], stage0_38[283], stage0_38[284], stage0_38[285], stage0_38[286], stage0_38[287]},
      {stage1_40[47],stage1_39[72],stage1_38[124],stage1_37[136],stage1_36[188]}
   );
   gpc606_5 gpc1439 (
      {stage0_36[410], stage0_36[411], stage0_36[412], stage0_36[413], stage0_36[414], stage0_36[415]},
      {stage0_38[288], stage0_38[289], stage0_38[290], stage0_38[291], stage0_38[292], stage0_38[293]},
      {stage1_40[48],stage1_39[73],stage1_38[125],stage1_37[137],stage1_36[189]}
   );
   gpc606_5 gpc1440 (
      {stage0_36[416], stage0_36[417], stage0_36[418], stage0_36[419], stage0_36[420], stage0_36[421]},
      {stage0_38[294], stage0_38[295], stage0_38[296], stage0_38[297], stage0_38[298], stage0_38[299]},
      {stage1_40[49],stage1_39[74],stage1_38[126],stage1_37[138],stage1_36[190]}
   );
   gpc606_5 gpc1441 (
      {stage0_36[422], stage0_36[423], stage0_36[424], stage0_36[425], stage0_36[426], stage0_36[427]},
      {stage0_38[300], stage0_38[301], stage0_38[302], stage0_38[303], stage0_38[304], stage0_38[305]},
      {stage1_40[50],stage1_39[75],stage1_38[127],stage1_37[139],stage1_36[191]}
   );
   gpc606_5 gpc1442 (
      {stage0_36[428], stage0_36[429], stage0_36[430], stage0_36[431], stage0_36[432], stage0_36[433]},
      {stage0_38[306], stage0_38[307], stage0_38[308], stage0_38[309], stage0_38[310], stage0_38[311]},
      {stage1_40[51],stage1_39[76],stage1_38[128],stage1_37[140],stage1_36[192]}
   );
   gpc606_5 gpc1443 (
      {stage0_36[434], stage0_36[435], stage0_36[436], stage0_36[437], stage0_36[438], stage0_36[439]},
      {stage0_38[312], stage0_38[313], stage0_38[314], stage0_38[315], stage0_38[316], stage0_38[317]},
      {stage1_40[52],stage1_39[77],stage1_38[129],stage1_37[141],stage1_36[193]}
   );
   gpc606_5 gpc1444 (
      {stage0_36[440], stage0_36[441], stage0_36[442], stage0_36[443], stage0_36[444], stage0_36[445]},
      {stage0_38[318], stage0_38[319], stage0_38[320], stage0_38[321], stage0_38[322], stage0_38[323]},
      {stage1_40[53],stage1_39[78],stage1_38[130],stage1_37[142],stage1_36[194]}
   );
   gpc606_5 gpc1445 (
      {stage0_36[446], stage0_36[447], stage0_36[448], stage0_36[449], stage0_36[450], stage0_36[451]},
      {stage0_38[324], stage0_38[325], stage0_38[326], stage0_38[327], stage0_38[328], stage0_38[329]},
      {stage1_40[54],stage1_39[79],stage1_38[131],stage1_37[143],stage1_36[195]}
   );
   gpc606_5 gpc1446 (
      {stage0_36[452], stage0_36[453], stage0_36[454], stage0_36[455], stage0_36[456], stage0_36[457]},
      {stage0_38[330], stage0_38[331], stage0_38[332], stage0_38[333], stage0_38[334], stage0_38[335]},
      {stage1_40[55],stage1_39[80],stage1_38[132],stage1_37[144],stage1_36[196]}
   );
   gpc606_5 gpc1447 (
      {stage0_36[458], stage0_36[459], stage0_36[460], stage0_36[461], stage0_36[462], stage0_36[463]},
      {stage0_38[336], stage0_38[337], stage0_38[338], stage0_38[339], stage0_38[340], stage0_38[341]},
      {stage1_40[56],stage1_39[81],stage1_38[133],stage1_37[145],stage1_36[197]}
   );
   gpc606_5 gpc1448 (
      {stage0_36[464], stage0_36[465], stage0_36[466], stage0_36[467], stage0_36[468], stage0_36[469]},
      {stage0_38[342], stage0_38[343], stage0_38[344], stage0_38[345], stage0_38[346], stage0_38[347]},
      {stage1_40[57],stage1_39[82],stage1_38[134],stage1_37[146],stage1_36[198]}
   );
   gpc606_5 gpc1449 (
      {stage0_36[470], stage0_36[471], stage0_36[472], stage0_36[473], stage0_36[474], stage0_36[475]},
      {stage0_38[348], stage0_38[349], stage0_38[350], stage0_38[351], stage0_38[352], stage0_38[353]},
      {stage1_40[58],stage1_39[83],stage1_38[135],stage1_37[147],stage1_36[199]}
   );
   gpc606_5 gpc1450 (
      {stage0_36[476], stage0_36[477], stage0_36[478], stage0_36[479], stage0_36[480], stage0_36[481]},
      {stage0_38[354], stage0_38[355], stage0_38[356], stage0_38[357], stage0_38[358], stage0_38[359]},
      {stage1_40[59],stage1_39[84],stage1_38[136],stage1_37[148],stage1_36[200]}
   );
   gpc606_5 gpc1451 (
      {stage0_36[482], stage0_36[483], stage0_36[484], stage0_36[485], 1'b0, 1'b0},
      {stage0_38[360], stage0_38[361], stage0_38[362], stage0_38[363], stage0_38[364], stage0_38[365]},
      {stage1_40[60],stage1_39[85],stage1_38[137],stage1_37[149],stage1_36[201]}
   );
   gpc606_5 gpc1452 (
      {stage0_37[193], stage0_37[194], stage0_37[195], stage0_37[196], stage0_37[197], stage0_37[198]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[61],stage1_39[86],stage1_38[138],stage1_37[150]}
   );
   gpc606_5 gpc1453 (
      {stage0_37[199], stage0_37[200], stage0_37[201], stage0_37[202], stage0_37[203], stage0_37[204]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[62],stage1_39[87],stage1_38[139],stage1_37[151]}
   );
   gpc606_5 gpc1454 (
      {stage0_37[205], stage0_37[206], stage0_37[207], stage0_37[208], stage0_37[209], stage0_37[210]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[63],stage1_39[88],stage1_38[140],stage1_37[152]}
   );
   gpc606_5 gpc1455 (
      {stage0_37[211], stage0_37[212], stage0_37[213], stage0_37[214], stage0_37[215], stage0_37[216]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[64],stage1_39[89],stage1_38[141],stage1_37[153]}
   );
   gpc606_5 gpc1456 (
      {stage0_37[217], stage0_37[218], stage0_37[219], stage0_37[220], stage0_37[221], stage0_37[222]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[65],stage1_39[90],stage1_38[142],stage1_37[154]}
   );
   gpc606_5 gpc1457 (
      {stage0_37[223], stage0_37[224], stage0_37[225], stage0_37[226], stage0_37[227], stage0_37[228]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[66],stage1_39[91],stage1_38[143],stage1_37[155]}
   );
   gpc606_5 gpc1458 (
      {stage0_37[229], stage0_37[230], stage0_37[231], stage0_37[232], stage0_37[233], stage0_37[234]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[67],stage1_39[92],stage1_38[144],stage1_37[156]}
   );
   gpc606_5 gpc1459 (
      {stage0_37[235], stage0_37[236], stage0_37[237], stage0_37[238], stage0_37[239], stage0_37[240]},
      {stage0_39[42], stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage1_41[7],stage1_40[68],stage1_39[93],stage1_38[145],stage1_37[157]}
   );
   gpc606_5 gpc1460 (
      {stage0_37[241], stage0_37[242], stage0_37[243], stage0_37[244], stage0_37[245], stage0_37[246]},
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52], stage0_39[53]},
      {stage1_41[8],stage1_40[69],stage1_39[94],stage1_38[146],stage1_37[158]}
   );
   gpc606_5 gpc1461 (
      {stage0_37[247], stage0_37[248], stage0_37[249], stage0_37[250], stage0_37[251], stage0_37[252]},
      {stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59]},
      {stage1_41[9],stage1_40[70],stage1_39[95],stage1_38[147],stage1_37[159]}
   );
   gpc606_5 gpc1462 (
      {stage0_37[253], stage0_37[254], stage0_37[255], stage0_37[256], stage0_37[257], stage0_37[258]},
      {stage0_39[60], stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage1_41[10],stage1_40[71],stage1_39[96],stage1_38[148],stage1_37[160]}
   );
   gpc606_5 gpc1463 (
      {stage0_37[259], stage0_37[260], stage0_37[261], stage0_37[262], stage0_37[263], stage0_37[264]},
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71]},
      {stage1_41[11],stage1_40[72],stage1_39[97],stage1_38[149],stage1_37[161]}
   );
   gpc606_5 gpc1464 (
      {stage0_37[265], stage0_37[266], stage0_37[267], stage0_37[268], stage0_37[269], stage0_37[270]},
      {stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage1_41[12],stage1_40[73],stage1_39[98],stage1_38[150],stage1_37[162]}
   );
   gpc606_5 gpc1465 (
      {stage0_37[271], stage0_37[272], stage0_37[273], stage0_37[274], stage0_37[275], stage0_37[276]},
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82], stage0_39[83]},
      {stage1_41[13],stage1_40[74],stage1_39[99],stage1_38[151],stage1_37[163]}
   );
   gpc606_5 gpc1466 (
      {stage0_37[277], stage0_37[278], stage0_37[279], stage0_37[280], stage0_37[281], stage0_37[282]},
      {stage0_39[84], stage0_39[85], stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89]},
      {stage1_41[14],stage1_40[75],stage1_39[100],stage1_38[152],stage1_37[164]}
   );
   gpc606_5 gpc1467 (
      {stage0_37[283], stage0_37[284], stage0_37[285], stage0_37[286], stage0_37[287], stage0_37[288]},
      {stage0_39[90], stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage1_41[15],stage1_40[76],stage1_39[101],stage1_38[153],stage1_37[165]}
   );
   gpc606_5 gpc1468 (
      {stage0_37[289], stage0_37[290], stage0_37[291], stage0_37[292], stage0_37[293], stage0_37[294]},
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100], stage0_39[101]},
      {stage1_41[16],stage1_40[77],stage1_39[102],stage1_38[154],stage1_37[166]}
   );
   gpc606_5 gpc1469 (
      {stage0_37[295], stage0_37[296], stage0_37[297], stage0_37[298], stage0_37[299], stage0_37[300]},
      {stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105], stage0_39[106], stage0_39[107]},
      {stage1_41[17],stage1_40[78],stage1_39[103],stage1_38[155],stage1_37[167]}
   );
   gpc606_5 gpc1470 (
      {stage0_37[301], stage0_37[302], stage0_37[303], stage0_37[304], stage0_37[305], stage0_37[306]},
      {stage0_39[108], stage0_39[109], stage0_39[110], stage0_39[111], stage0_39[112], stage0_39[113]},
      {stage1_41[18],stage1_40[79],stage1_39[104],stage1_38[156],stage1_37[168]}
   );
   gpc606_5 gpc1471 (
      {stage0_37[307], stage0_37[308], stage0_37[309], stage0_37[310], stage0_37[311], stage0_37[312]},
      {stage0_39[114], stage0_39[115], stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119]},
      {stage1_41[19],stage1_40[80],stage1_39[105],stage1_38[157],stage1_37[169]}
   );
   gpc606_5 gpc1472 (
      {stage0_37[313], stage0_37[314], stage0_37[315], stage0_37[316], stage0_37[317], stage0_37[318]},
      {stage0_39[120], stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage1_41[20],stage1_40[81],stage1_39[106],stage1_38[158],stage1_37[170]}
   );
   gpc606_5 gpc1473 (
      {stage0_37[319], stage0_37[320], stage0_37[321], stage0_37[322], stage0_37[323], stage0_37[324]},
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130], stage0_39[131]},
      {stage1_41[21],stage1_40[82],stage1_39[107],stage1_38[159],stage1_37[171]}
   );
   gpc606_5 gpc1474 (
      {stage0_37[325], stage0_37[326], stage0_37[327], stage0_37[328], stage0_37[329], stage0_37[330]},
      {stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135], stage0_39[136], stage0_39[137]},
      {stage1_41[22],stage1_40[83],stage1_39[108],stage1_38[160],stage1_37[172]}
   );
   gpc606_5 gpc1475 (
      {stage0_37[331], stage0_37[332], stage0_37[333], stage0_37[334], stage0_37[335], stage0_37[336]},
      {stage0_39[138], stage0_39[139], stage0_39[140], stage0_39[141], stage0_39[142], stage0_39[143]},
      {stage1_41[23],stage1_40[84],stage1_39[109],stage1_38[161],stage1_37[173]}
   );
   gpc606_5 gpc1476 (
      {stage0_37[337], stage0_37[338], stage0_37[339], stage0_37[340], stage0_37[341], stage0_37[342]},
      {stage0_39[144], stage0_39[145], stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149]},
      {stage1_41[24],stage1_40[85],stage1_39[110],stage1_38[162],stage1_37[174]}
   );
   gpc606_5 gpc1477 (
      {stage0_37[343], stage0_37[344], stage0_37[345], stage0_37[346], stage0_37[347], stage0_37[348]},
      {stage0_39[150], stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage1_41[25],stage1_40[86],stage1_39[111],stage1_38[163],stage1_37[175]}
   );
   gpc606_5 gpc1478 (
      {stage0_37[349], stage0_37[350], stage0_37[351], stage0_37[352], stage0_37[353], stage0_37[354]},
      {stage0_39[156], stage0_39[157], stage0_39[158], stage0_39[159], stage0_39[160], stage0_39[161]},
      {stage1_41[26],stage1_40[87],stage1_39[112],stage1_38[164],stage1_37[176]}
   );
   gpc615_5 gpc1479 (
      {stage0_38[366], stage0_38[367], stage0_38[368], stage0_38[369], stage0_38[370]},
      {stage0_39[162]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[27],stage1_40[88],stage1_39[113],stage1_38[165]}
   );
   gpc615_5 gpc1480 (
      {stage0_38[371], stage0_38[372], stage0_38[373], stage0_38[374], stage0_38[375]},
      {stage0_39[163]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[28],stage1_40[89],stage1_39[114],stage1_38[166]}
   );
   gpc615_5 gpc1481 (
      {stage0_38[376], stage0_38[377], stage0_38[378], stage0_38[379], stage0_38[380]},
      {stage0_39[164]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[29],stage1_40[90],stage1_39[115],stage1_38[167]}
   );
   gpc615_5 gpc1482 (
      {stage0_38[381], stage0_38[382], stage0_38[383], stage0_38[384], stage0_38[385]},
      {stage0_39[165]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[30],stage1_40[91],stage1_39[116],stage1_38[168]}
   );
   gpc615_5 gpc1483 (
      {stage0_38[386], stage0_38[387], stage0_38[388], stage0_38[389], stage0_38[390]},
      {stage0_39[166]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[31],stage1_40[92],stage1_39[117],stage1_38[169]}
   );
   gpc615_5 gpc1484 (
      {stage0_39[167], stage0_39[168], stage0_39[169], stage0_39[170], stage0_39[171]},
      {stage0_40[30]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[5],stage1_41[32],stage1_40[93],stage1_39[118]}
   );
   gpc615_5 gpc1485 (
      {stage0_39[172], stage0_39[173], stage0_39[174], stage0_39[175], stage0_39[176]},
      {stage0_40[31]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[6],stage1_41[33],stage1_40[94],stage1_39[119]}
   );
   gpc615_5 gpc1486 (
      {stage0_39[177], stage0_39[178], stage0_39[179], stage0_39[180], stage0_39[181]},
      {stage0_40[32]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[7],stage1_41[34],stage1_40[95],stage1_39[120]}
   );
   gpc615_5 gpc1487 (
      {stage0_39[182], stage0_39[183], stage0_39[184], stage0_39[185], stage0_39[186]},
      {stage0_40[33]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[8],stage1_41[35],stage1_40[96],stage1_39[121]}
   );
   gpc615_5 gpc1488 (
      {stage0_39[187], stage0_39[188], stage0_39[189], stage0_39[190], stage0_39[191]},
      {stage0_40[34]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[9],stage1_41[36],stage1_40[97],stage1_39[122]}
   );
   gpc615_5 gpc1489 (
      {stage0_39[192], stage0_39[193], stage0_39[194], stage0_39[195], stage0_39[196]},
      {stage0_40[35]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[10],stage1_41[37],stage1_40[98],stage1_39[123]}
   );
   gpc615_5 gpc1490 (
      {stage0_39[197], stage0_39[198], stage0_39[199], stage0_39[200], stage0_39[201]},
      {stage0_40[36]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[11],stage1_41[38],stage1_40[99],stage1_39[124]}
   );
   gpc615_5 gpc1491 (
      {stage0_39[202], stage0_39[203], stage0_39[204], stage0_39[205], stage0_39[206]},
      {stage0_40[37]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[12],stage1_41[39],stage1_40[100],stage1_39[125]}
   );
   gpc615_5 gpc1492 (
      {stage0_39[207], stage0_39[208], stage0_39[209], stage0_39[210], stage0_39[211]},
      {stage0_40[38]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[13],stage1_41[40],stage1_40[101],stage1_39[126]}
   );
   gpc615_5 gpc1493 (
      {stage0_39[212], stage0_39[213], stage0_39[214], stage0_39[215], stage0_39[216]},
      {stage0_40[39]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[14],stage1_41[41],stage1_40[102],stage1_39[127]}
   );
   gpc615_5 gpc1494 (
      {stage0_39[217], stage0_39[218], stage0_39[219], stage0_39[220], stage0_39[221]},
      {stage0_40[40]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[15],stage1_41[42],stage1_40[103],stage1_39[128]}
   );
   gpc615_5 gpc1495 (
      {stage0_39[222], stage0_39[223], stage0_39[224], stage0_39[225], stage0_39[226]},
      {stage0_40[41]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[16],stage1_41[43],stage1_40[104],stage1_39[129]}
   );
   gpc615_5 gpc1496 (
      {stage0_39[227], stage0_39[228], stage0_39[229], stage0_39[230], stage0_39[231]},
      {stage0_40[42]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[17],stage1_41[44],stage1_40[105],stage1_39[130]}
   );
   gpc615_5 gpc1497 (
      {stage0_39[232], stage0_39[233], stage0_39[234], stage0_39[235], stage0_39[236]},
      {stage0_40[43]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[18],stage1_41[45],stage1_40[106],stage1_39[131]}
   );
   gpc615_5 gpc1498 (
      {stage0_39[237], stage0_39[238], stage0_39[239], stage0_39[240], stage0_39[241]},
      {stage0_40[44]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[19],stage1_41[46],stage1_40[107],stage1_39[132]}
   );
   gpc615_5 gpc1499 (
      {stage0_39[242], stage0_39[243], stage0_39[244], stage0_39[245], stage0_39[246]},
      {stage0_40[45]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage1_43[15],stage1_42[20],stage1_41[47],stage1_40[108],stage1_39[133]}
   );
   gpc615_5 gpc1500 (
      {stage0_39[247], stage0_39[248], stage0_39[249], stage0_39[250], stage0_39[251]},
      {stage0_40[46]},
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage1_43[16],stage1_42[21],stage1_41[48],stage1_40[109],stage1_39[134]}
   );
   gpc615_5 gpc1501 (
      {stage0_39[252], stage0_39[253], stage0_39[254], stage0_39[255], stage0_39[256]},
      {stage0_40[47]},
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage1_43[17],stage1_42[22],stage1_41[49],stage1_40[110],stage1_39[135]}
   );
   gpc615_5 gpc1502 (
      {stage0_39[257], stage0_39[258], stage0_39[259], stage0_39[260], stage0_39[261]},
      {stage0_40[48]},
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage1_43[18],stage1_42[23],stage1_41[50],stage1_40[111],stage1_39[136]}
   );
   gpc615_5 gpc1503 (
      {stage0_39[262], stage0_39[263], stage0_39[264], stage0_39[265], stage0_39[266]},
      {stage0_40[49]},
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage1_43[19],stage1_42[24],stage1_41[51],stage1_40[112],stage1_39[137]}
   );
   gpc615_5 gpc1504 (
      {stage0_39[267], stage0_39[268], stage0_39[269], stage0_39[270], stage0_39[271]},
      {stage0_40[50]},
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage1_43[20],stage1_42[25],stage1_41[52],stage1_40[113],stage1_39[138]}
   );
   gpc615_5 gpc1505 (
      {stage0_39[272], stage0_39[273], stage0_39[274], stage0_39[275], stage0_39[276]},
      {stage0_40[51]},
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage1_43[21],stage1_42[26],stage1_41[53],stage1_40[114],stage1_39[139]}
   );
   gpc615_5 gpc1506 (
      {stage0_39[277], stage0_39[278], stage0_39[279], stage0_39[280], stage0_39[281]},
      {stage0_40[52]},
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage1_43[22],stage1_42[27],stage1_41[54],stage1_40[115],stage1_39[140]}
   );
   gpc615_5 gpc1507 (
      {stage0_39[282], stage0_39[283], stage0_39[284], stage0_39[285], stage0_39[286]},
      {stage0_40[53]},
      {stage0_41[138], stage0_41[139], stage0_41[140], stage0_41[141], stage0_41[142], stage0_41[143]},
      {stage1_43[23],stage1_42[28],stage1_41[55],stage1_40[116],stage1_39[141]}
   );
   gpc615_5 gpc1508 (
      {stage0_39[287], stage0_39[288], stage0_39[289], stage0_39[290], stage0_39[291]},
      {stage0_40[54]},
      {stage0_41[144], stage0_41[145], stage0_41[146], stage0_41[147], stage0_41[148], stage0_41[149]},
      {stage1_43[24],stage1_42[29],stage1_41[56],stage1_40[117],stage1_39[142]}
   );
   gpc615_5 gpc1509 (
      {stage0_39[292], stage0_39[293], stage0_39[294], stage0_39[295], stage0_39[296]},
      {stage0_40[55]},
      {stage0_41[150], stage0_41[151], stage0_41[152], stage0_41[153], stage0_41[154], stage0_41[155]},
      {stage1_43[25],stage1_42[30],stage1_41[57],stage1_40[118],stage1_39[143]}
   );
   gpc615_5 gpc1510 (
      {stage0_39[297], stage0_39[298], stage0_39[299], stage0_39[300], stage0_39[301]},
      {stage0_40[56]},
      {stage0_41[156], stage0_41[157], stage0_41[158], stage0_41[159], stage0_41[160], stage0_41[161]},
      {stage1_43[26],stage1_42[31],stage1_41[58],stage1_40[119],stage1_39[144]}
   );
   gpc615_5 gpc1511 (
      {stage0_39[302], stage0_39[303], stage0_39[304], stage0_39[305], stage0_39[306]},
      {stage0_40[57]},
      {stage0_41[162], stage0_41[163], stage0_41[164], stage0_41[165], stage0_41[166], stage0_41[167]},
      {stage1_43[27],stage1_42[32],stage1_41[59],stage1_40[120],stage1_39[145]}
   );
   gpc615_5 gpc1512 (
      {stage0_39[307], stage0_39[308], stage0_39[309], stage0_39[310], stage0_39[311]},
      {stage0_40[58]},
      {stage0_41[168], stage0_41[169], stage0_41[170], stage0_41[171], stage0_41[172], stage0_41[173]},
      {stage1_43[28],stage1_42[33],stage1_41[60],stage1_40[121],stage1_39[146]}
   );
   gpc615_5 gpc1513 (
      {stage0_39[312], stage0_39[313], stage0_39[314], stage0_39[315], stage0_39[316]},
      {stage0_40[59]},
      {stage0_41[174], stage0_41[175], stage0_41[176], stage0_41[177], stage0_41[178], stage0_41[179]},
      {stage1_43[29],stage1_42[34],stage1_41[61],stage1_40[122],stage1_39[147]}
   );
   gpc615_5 gpc1514 (
      {stage0_39[317], stage0_39[318], stage0_39[319], stage0_39[320], stage0_39[321]},
      {stage0_40[60]},
      {stage0_41[180], stage0_41[181], stage0_41[182], stage0_41[183], stage0_41[184], stage0_41[185]},
      {stage1_43[30],stage1_42[35],stage1_41[62],stage1_40[123],stage1_39[148]}
   );
   gpc615_5 gpc1515 (
      {stage0_39[322], stage0_39[323], stage0_39[324], stage0_39[325], stage0_39[326]},
      {stage0_40[61]},
      {stage0_41[186], stage0_41[187], stage0_41[188], stage0_41[189], stage0_41[190], stage0_41[191]},
      {stage1_43[31],stage1_42[36],stage1_41[63],stage1_40[124],stage1_39[149]}
   );
   gpc615_5 gpc1516 (
      {stage0_39[327], stage0_39[328], stage0_39[329], stage0_39[330], stage0_39[331]},
      {stage0_40[62]},
      {stage0_41[192], stage0_41[193], stage0_41[194], stage0_41[195], stage0_41[196], stage0_41[197]},
      {stage1_43[32],stage1_42[37],stage1_41[64],stage1_40[125],stage1_39[150]}
   );
   gpc615_5 gpc1517 (
      {stage0_39[332], stage0_39[333], stage0_39[334], stage0_39[335], stage0_39[336]},
      {stage0_40[63]},
      {stage0_41[198], stage0_41[199], stage0_41[200], stage0_41[201], stage0_41[202], stage0_41[203]},
      {stage1_43[33],stage1_42[38],stage1_41[65],stage1_40[126],stage1_39[151]}
   );
   gpc615_5 gpc1518 (
      {stage0_39[337], stage0_39[338], stage0_39[339], stage0_39[340], stage0_39[341]},
      {stage0_40[64]},
      {stage0_41[204], stage0_41[205], stage0_41[206], stage0_41[207], stage0_41[208], stage0_41[209]},
      {stage1_43[34],stage1_42[39],stage1_41[66],stage1_40[127],stage1_39[152]}
   );
   gpc615_5 gpc1519 (
      {stage0_39[342], stage0_39[343], stage0_39[344], stage0_39[345], stage0_39[346]},
      {stage0_40[65]},
      {stage0_41[210], stage0_41[211], stage0_41[212], stage0_41[213], stage0_41[214], stage0_41[215]},
      {stage1_43[35],stage1_42[40],stage1_41[67],stage1_40[128],stage1_39[153]}
   );
   gpc615_5 gpc1520 (
      {stage0_39[347], stage0_39[348], stage0_39[349], stage0_39[350], stage0_39[351]},
      {stage0_40[66]},
      {stage0_41[216], stage0_41[217], stage0_41[218], stage0_41[219], stage0_41[220], stage0_41[221]},
      {stage1_43[36],stage1_42[41],stage1_41[68],stage1_40[129],stage1_39[154]}
   );
   gpc615_5 gpc1521 (
      {stage0_39[352], stage0_39[353], stage0_39[354], stage0_39[355], stage0_39[356]},
      {stage0_40[67]},
      {stage0_41[222], stage0_41[223], stage0_41[224], stage0_41[225], stage0_41[226], stage0_41[227]},
      {stage1_43[37],stage1_42[42],stage1_41[69],stage1_40[130],stage1_39[155]}
   );
   gpc615_5 gpc1522 (
      {stage0_39[357], stage0_39[358], stage0_39[359], stage0_39[360], stage0_39[361]},
      {stage0_40[68]},
      {stage0_41[228], stage0_41[229], stage0_41[230], stage0_41[231], stage0_41[232], stage0_41[233]},
      {stage1_43[38],stage1_42[43],stage1_41[70],stage1_40[131],stage1_39[156]}
   );
   gpc615_5 gpc1523 (
      {stage0_39[362], stage0_39[363], stage0_39[364], stage0_39[365], stage0_39[366]},
      {stage0_40[69]},
      {stage0_41[234], stage0_41[235], stage0_41[236], stage0_41[237], stage0_41[238], stage0_41[239]},
      {stage1_43[39],stage1_42[44],stage1_41[71],stage1_40[132],stage1_39[157]}
   );
   gpc615_5 gpc1524 (
      {stage0_39[367], stage0_39[368], stage0_39[369], stage0_39[370], stage0_39[371]},
      {stage0_40[70]},
      {stage0_41[240], stage0_41[241], stage0_41[242], stage0_41[243], stage0_41[244], stage0_41[245]},
      {stage1_43[40],stage1_42[45],stage1_41[72],stage1_40[133],stage1_39[158]}
   );
   gpc615_5 gpc1525 (
      {stage0_39[372], stage0_39[373], stage0_39[374], stage0_39[375], stage0_39[376]},
      {stage0_40[71]},
      {stage0_41[246], stage0_41[247], stage0_41[248], stage0_41[249], stage0_41[250], stage0_41[251]},
      {stage1_43[41],stage1_42[46],stage1_41[73],stage1_40[134],stage1_39[159]}
   );
   gpc615_5 gpc1526 (
      {stage0_39[377], stage0_39[378], stage0_39[379], stage0_39[380], stage0_39[381]},
      {stage0_40[72]},
      {stage0_41[252], stage0_41[253], stage0_41[254], stage0_41[255], stage0_41[256], stage0_41[257]},
      {stage1_43[42],stage1_42[47],stage1_41[74],stage1_40[135],stage1_39[160]}
   );
   gpc615_5 gpc1527 (
      {stage0_39[382], stage0_39[383], stage0_39[384], stage0_39[385], stage0_39[386]},
      {stage0_40[73]},
      {stage0_41[258], stage0_41[259], stage0_41[260], stage0_41[261], stage0_41[262], stage0_41[263]},
      {stage1_43[43],stage1_42[48],stage1_41[75],stage1_40[136],stage1_39[161]}
   );
   gpc615_5 gpc1528 (
      {stage0_39[387], stage0_39[388], stage0_39[389], stage0_39[390], stage0_39[391]},
      {stage0_40[74]},
      {stage0_41[264], stage0_41[265], stage0_41[266], stage0_41[267], stage0_41[268], stage0_41[269]},
      {stage1_43[44],stage1_42[49],stage1_41[76],stage1_40[137],stage1_39[162]}
   );
   gpc615_5 gpc1529 (
      {stage0_39[392], stage0_39[393], stage0_39[394], stage0_39[395], stage0_39[396]},
      {stage0_40[75]},
      {stage0_41[270], stage0_41[271], stage0_41[272], stage0_41[273], stage0_41[274], stage0_41[275]},
      {stage1_43[45],stage1_42[50],stage1_41[77],stage1_40[138],stage1_39[163]}
   );
   gpc615_5 gpc1530 (
      {stage0_39[397], stage0_39[398], stage0_39[399], stage0_39[400], stage0_39[401]},
      {stage0_40[76]},
      {stage0_41[276], stage0_41[277], stage0_41[278], stage0_41[279], stage0_41[280], stage0_41[281]},
      {stage1_43[46],stage1_42[51],stage1_41[78],stage1_40[139],stage1_39[164]}
   );
   gpc615_5 gpc1531 (
      {stage0_39[402], stage0_39[403], stage0_39[404], stage0_39[405], stage0_39[406]},
      {stage0_40[77]},
      {stage0_41[282], stage0_41[283], stage0_41[284], stage0_41[285], stage0_41[286], stage0_41[287]},
      {stage1_43[47],stage1_42[52],stage1_41[79],stage1_40[140],stage1_39[165]}
   );
   gpc615_5 gpc1532 (
      {stage0_39[407], stage0_39[408], stage0_39[409], stage0_39[410], stage0_39[411]},
      {stage0_40[78]},
      {stage0_41[288], stage0_41[289], stage0_41[290], stage0_41[291], stage0_41[292], stage0_41[293]},
      {stage1_43[48],stage1_42[53],stage1_41[80],stage1_40[141],stage1_39[166]}
   );
   gpc615_5 gpc1533 (
      {stage0_39[412], stage0_39[413], stage0_39[414], stage0_39[415], stage0_39[416]},
      {stage0_40[79]},
      {stage0_41[294], stage0_41[295], stage0_41[296], stage0_41[297], stage0_41[298], stage0_41[299]},
      {stage1_43[49],stage1_42[54],stage1_41[81],stage1_40[142],stage1_39[167]}
   );
   gpc615_5 gpc1534 (
      {stage0_39[417], stage0_39[418], stage0_39[419], stage0_39[420], stage0_39[421]},
      {stage0_40[80]},
      {stage0_41[300], stage0_41[301], stage0_41[302], stage0_41[303], stage0_41[304], stage0_41[305]},
      {stage1_43[50],stage1_42[55],stage1_41[82],stage1_40[143],stage1_39[168]}
   );
   gpc615_5 gpc1535 (
      {stage0_39[422], stage0_39[423], stage0_39[424], stage0_39[425], stage0_39[426]},
      {stage0_40[81]},
      {stage0_41[306], stage0_41[307], stage0_41[308], stage0_41[309], stage0_41[310], stage0_41[311]},
      {stage1_43[51],stage1_42[56],stage1_41[83],stage1_40[144],stage1_39[169]}
   );
   gpc615_5 gpc1536 (
      {stage0_39[427], stage0_39[428], stage0_39[429], stage0_39[430], stage0_39[431]},
      {stage0_40[82]},
      {stage0_41[312], stage0_41[313], stage0_41[314], stage0_41[315], stage0_41[316], stage0_41[317]},
      {stage1_43[52],stage1_42[57],stage1_41[84],stage1_40[145],stage1_39[170]}
   );
   gpc615_5 gpc1537 (
      {stage0_39[432], stage0_39[433], stage0_39[434], stage0_39[435], stage0_39[436]},
      {stage0_40[83]},
      {stage0_41[318], stage0_41[319], stage0_41[320], stage0_41[321], stage0_41[322], stage0_41[323]},
      {stage1_43[53],stage1_42[58],stage1_41[85],stage1_40[146],stage1_39[171]}
   );
   gpc615_5 gpc1538 (
      {stage0_39[437], stage0_39[438], stage0_39[439], stage0_39[440], stage0_39[441]},
      {stage0_40[84]},
      {stage0_41[324], stage0_41[325], stage0_41[326], stage0_41[327], stage0_41[328], stage0_41[329]},
      {stage1_43[54],stage1_42[59],stage1_41[86],stage1_40[147],stage1_39[172]}
   );
   gpc615_5 gpc1539 (
      {stage0_39[442], stage0_39[443], stage0_39[444], stage0_39[445], stage0_39[446]},
      {stage0_40[85]},
      {stage0_41[330], stage0_41[331], stage0_41[332], stage0_41[333], stage0_41[334], stage0_41[335]},
      {stage1_43[55],stage1_42[60],stage1_41[87],stage1_40[148],stage1_39[173]}
   );
   gpc606_5 gpc1540 (
      {stage0_40[86], stage0_40[87], stage0_40[88], stage0_40[89], stage0_40[90], stage0_40[91]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[56],stage1_42[61],stage1_41[88],stage1_40[149]}
   );
   gpc606_5 gpc1541 (
      {stage0_40[92], stage0_40[93], stage0_40[94], stage0_40[95], stage0_40[96], stage0_40[97]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[57],stage1_42[62],stage1_41[89],stage1_40[150]}
   );
   gpc606_5 gpc1542 (
      {stage0_40[98], stage0_40[99], stage0_40[100], stage0_40[101], stage0_40[102], stage0_40[103]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[58],stage1_42[63],stage1_41[90],stage1_40[151]}
   );
   gpc606_5 gpc1543 (
      {stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107], stage0_40[108], stage0_40[109]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[59],stage1_42[64],stage1_41[91],stage1_40[152]}
   );
   gpc606_5 gpc1544 (
      {stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113], stage0_40[114], stage0_40[115]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[60],stage1_42[65],stage1_41[92],stage1_40[153]}
   );
   gpc606_5 gpc1545 (
      {stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119], stage0_40[120], stage0_40[121]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[61],stage1_42[66],stage1_41[93],stage1_40[154]}
   );
   gpc606_5 gpc1546 (
      {stage0_40[122], stage0_40[123], stage0_40[124], stage0_40[125], stage0_40[126], stage0_40[127]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[62],stage1_42[67],stage1_41[94],stage1_40[155]}
   );
   gpc606_5 gpc1547 (
      {stage0_40[128], stage0_40[129], stage0_40[130], stage0_40[131], stage0_40[132], stage0_40[133]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[63],stage1_42[68],stage1_41[95],stage1_40[156]}
   );
   gpc606_5 gpc1548 (
      {stage0_40[134], stage0_40[135], stage0_40[136], stage0_40[137], stage0_40[138], stage0_40[139]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[64],stage1_42[69],stage1_41[96],stage1_40[157]}
   );
   gpc606_5 gpc1549 (
      {stage0_40[140], stage0_40[141], stage0_40[142], stage0_40[143], stage0_40[144], stage0_40[145]},
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage1_44[9],stage1_43[65],stage1_42[70],stage1_41[97],stage1_40[158]}
   );
   gpc606_5 gpc1550 (
      {stage0_40[146], stage0_40[147], stage0_40[148], stage0_40[149], stage0_40[150], stage0_40[151]},
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage1_44[10],stage1_43[66],stage1_42[71],stage1_41[98],stage1_40[159]}
   );
   gpc606_5 gpc1551 (
      {stage0_40[152], stage0_40[153], stage0_40[154], stage0_40[155], stage0_40[156], stage0_40[157]},
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage1_44[11],stage1_43[67],stage1_42[72],stage1_41[99],stage1_40[160]}
   );
   gpc606_5 gpc1552 (
      {stage0_40[158], stage0_40[159], stage0_40[160], stage0_40[161], stage0_40[162], stage0_40[163]},
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76], stage0_42[77]},
      {stage1_44[12],stage1_43[68],stage1_42[73],stage1_41[100],stage1_40[161]}
   );
   gpc606_5 gpc1553 (
      {stage0_40[164], stage0_40[165], stage0_40[166], stage0_40[167], stage0_40[168], stage0_40[169]},
      {stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81], stage0_42[82], stage0_42[83]},
      {stage1_44[13],stage1_43[69],stage1_42[74],stage1_41[101],stage1_40[162]}
   );
   gpc606_5 gpc1554 (
      {stage0_40[170], stage0_40[171], stage0_40[172], stage0_40[173], stage0_40[174], stage0_40[175]},
      {stage0_42[84], stage0_42[85], stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89]},
      {stage1_44[14],stage1_43[70],stage1_42[75],stage1_41[102],stage1_40[163]}
   );
   gpc606_5 gpc1555 (
      {stage0_40[176], stage0_40[177], stage0_40[178], stage0_40[179], stage0_40[180], stage0_40[181]},
      {stage0_42[90], stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage1_44[15],stage1_43[71],stage1_42[76],stage1_41[103],stage1_40[164]}
   );
   gpc606_5 gpc1556 (
      {stage0_40[182], stage0_40[183], stage0_40[184], stage0_40[185], stage0_40[186], stage0_40[187]},
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage1_44[16],stage1_43[72],stage1_42[77],stage1_41[104],stage1_40[165]}
   );
   gpc606_5 gpc1557 (
      {stage0_40[188], stage0_40[189], stage0_40[190], stage0_40[191], stage0_40[192], stage0_40[193]},
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106], stage0_42[107]},
      {stage1_44[17],stage1_43[73],stage1_42[78],stage1_41[105],stage1_40[166]}
   );
   gpc606_5 gpc1558 (
      {stage0_40[194], stage0_40[195], stage0_40[196], stage0_40[197], stage0_40[198], stage0_40[199]},
      {stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111], stage0_42[112], stage0_42[113]},
      {stage1_44[18],stage1_43[74],stage1_42[79],stage1_41[106],stage1_40[167]}
   );
   gpc606_5 gpc1559 (
      {stage0_40[200], stage0_40[201], stage0_40[202], stage0_40[203], stage0_40[204], stage0_40[205]},
      {stage0_42[114], stage0_42[115], stage0_42[116], stage0_42[117], stage0_42[118], stage0_42[119]},
      {stage1_44[19],stage1_43[75],stage1_42[80],stage1_41[107],stage1_40[168]}
   );
   gpc606_5 gpc1560 (
      {stage0_40[206], stage0_40[207], stage0_40[208], stage0_40[209], stage0_40[210], stage0_40[211]},
      {stage0_42[120], stage0_42[121], stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125]},
      {stage1_44[20],stage1_43[76],stage1_42[81],stage1_41[108],stage1_40[169]}
   );
   gpc606_5 gpc1561 (
      {stage0_40[212], stage0_40[213], stage0_40[214], stage0_40[215], stage0_40[216], stage0_40[217]},
      {stage0_42[126], stage0_42[127], stage0_42[128], stage0_42[129], stage0_42[130], stage0_42[131]},
      {stage1_44[21],stage1_43[77],stage1_42[82],stage1_41[109],stage1_40[170]}
   );
   gpc606_5 gpc1562 (
      {stage0_40[218], stage0_40[219], stage0_40[220], stage0_40[221], stage0_40[222], stage0_40[223]},
      {stage0_42[132], stage0_42[133], stage0_42[134], stage0_42[135], stage0_42[136], stage0_42[137]},
      {stage1_44[22],stage1_43[78],stage1_42[83],stage1_41[110],stage1_40[171]}
   );
   gpc606_5 gpc1563 (
      {stage0_40[224], stage0_40[225], stage0_40[226], stage0_40[227], stage0_40[228], stage0_40[229]},
      {stage0_42[138], stage0_42[139], stage0_42[140], stage0_42[141], stage0_42[142], stage0_42[143]},
      {stage1_44[23],stage1_43[79],stage1_42[84],stage1_41[111],stage1_40[172]}
   );
   gpc606_5 gpc1564 (
      {stage0_40[230], stage0_40[231], stage0_40[232], stage0_40[233], stage0_40[234], stage0_40[235]},
      {stage0_42[144], stage0_42[145], stage0_42[146], stage0_42[147], stage0_42[148], stage0_42[149]},
      {stage1_44[24],stage1_43[80],stage1_42[85],stage1_41[112],stage1_40[173]}
   );
   gpc606_5 gpc1565 (
      {stage0_40[236], stage0_40[237], stage0_40[238], stage0_40[239], stage0_40[240], stage0_40[241]},
      {stage0_42[150], stage0_42[151], stage0_42[152], stage0_42[153], stage0_42[154], stage0_42[155]},
      {stage1_44[25],stage1_43[81],stage1_42[86],stage1_41[113],stage1_40[174]}
   );
   gpc606_5 gpc1566 (
      {stage0_40[242], stage0_40[243], stage0_40[244], stage0_40[245], stage0_40[246], stage0_40[247]},
      {stage0_42[156], stage0_42[157], stage0_42[158], stage0_42[159], stage0_42[160], stage0_42[161]},
      {stage1_44[26],stage1_43[82],stage1_42[87],stage1_41[114],stage1_40[175]}
   );
   gpc606_5 gpc1567 (
      {stage0_40[248], stage0_40[249], stage0_40[250], stage0_40[251], stage0_40[252], stage0_40[253]},
      {stage0_42[162], stage0_42[163], stage0_42[164], stage0_42[165], stage0_42[166], stage0_42[167]},
      {stage1_44[27],stage1_43[83],stage1_42[88],stage1_41[115],stage1_40[176]}
   );
   gpc606_5 gpc1568 (
      {stage0_40[254], stage0_40[255], stage0_40[256], stage0_40[257], stage0_40[258], stage0_40[259]},
      {stage0_42[168], stage0_42[169], stage0_42[170], stage0_42[171], stage0_42[172], stage0_42[173]},
      {stage1_44[28],stage1_43[84],stage1_42[89],stage1_41[116],stage1_40[177]}
   );
   gpc606_5 gpc1569 (
      {stage0_40[260], stage0_40[261], stage0_40[262], stage0_40[263], stage0_40[264], stage0_40[265]},
      {stage0_42[174], stage0_42[175], stage0_42[176], stage0_42[177], stage0_42[178], stage0_42[179]},
      {stage1_44[29],stage1_43[85],stage1_42[90],stage1_41[117],stage1_40[178]}
   );
   gpc606_5 gpc1570 (
      {stage0_40[266], stage0_40[267], stage0_40[268], stage0_40[269], stage0_40[270], stage0_40[271]},
      {stage0_42[180], stage0_42[181], stage0_42[182], stage0_42[183], stage0_42[184], stage0_42[185]},
      {stage1_44[30],stage1_43[86],stage1_42[91],stage1_41[118],stage1_40[179]}
   );
   gpc606_5 gpc1571 (
      {stage0_40[272], stage0_40[273], stage0_40[274], stage0_40[275], stage0_40[276], stage0_40[277]},
      {stage0_42[186], stage0_42[187], stage0_42[188], stage0_42[189], stage0_42[190], stage0_42[191]},
      {stage1_44[31],stage1_43[87],stage1_42[92],stage1_41[119],stage1_40[180]}
   );
   gpc606_5 gpc1572 (
      {stage0_40[278], stage0_40[279], stage0_40[280], stage0_40[281], stage0_40[282], stage0_40[283]},
      {stage0_42[192], stage0_42[193], stage0_42[194], stage0_42[195], stage0_42[196], stage0_42[197]},
      {stage1_44[32],stage1_43[88],stage1_42[93],stage1_41[120],stage1_40[181]}
   );
   gpc606_5 gpc1573 (
      {stage0_40[284], stage0_40[285], stage0_40[286], stage0_40[287], stage0_40[288], stage0_40[289]},
      {stage0_42[198], stage0_42[199], stage0_42[200], stage0_42[201], stage0_42[202], stage0_42[203]},
      {stage1_44[33],stage1_43[89],stage1_42[94],stage1_41[121],stage1_40[182]}
   );
   gpc606_5 gpc1574 (
      {stage0_40[290], stage0_40[291], stage0_40[292], stage0_40[293], stage0_40[294], stage0_40[295]},
      {stage0_42[204], stage0_42[205], stage0_42[206], stage0_42[207], stage0_42[208], stage0_42[209]},
      {stage1_44[34],stage1_43[90],stage1_42[95],stage1_41[122],stage1_40[183]}
   );
   gpc606_5 gpc1575 (
      {stage0_40[296], stage0_40[297], stage0_40[298], stage0_40[299], stage0_40[300], stage0_40[301]},
      {stage0_42[210], stage0_42[211], stage0_42[212], stage0_42[213], stage0_42[214], stage0_42[215]},
      {stage1_44[35],stage1_43[91],stage1_42[96],stage1_41[123],stage1_40[184]}
   );
   gpc606_5 gpc1576 (
      {stage0_40[302], stage0_40[303], stage0_40[304], stage0_40[305], stage0_40[306], stage0_40[307]},
      {stage0_42[216], stage0_42[217], stage0_42[218], stage0_42[219], stage0_42[220], stage0_42[221]},
      {stage1_44[36],stage1_43[92],stage1_42[97],stage1_41[124],stage1_40[185]}
   );
   gpc606_5 gpc1577 (
      {stage0_40[308], stage0_40[309], stage0_40[310], stage0_40[311], stage0_40[312], stage0_40[313]},
      {stage0_42[222], stage0_42[223], stage0_42[224], stage0_42[225], stage0_42[226], stage0_42[227]},
      {stage1_44[37],stage1_43[93],stage1_42[98],stage1_41[125],stage1_40[186]}
   );
   gpc606_5 gpc1578 (
      {stage0_40[314], stage0_40[315], stage0_40[316], stage0_40[317], stage0_40[318], stage0_40[319]},
      {stage0_42[228], stage0_42[229], stage0_42[230], stage0_42[231], stage0_42[232], stage0_42[233]},
      {stage1_44[38],stage1_43[94],stage1_42[99],stage1_41[126],stage1_40[187]}
   );
   gpc606_5 gpc1579 (
      {stage0_40[320], stage0_40[321], stage0_40[322], stage0_40[323], stage0_40[324], stage0_40[325]},
      {stage0_42[234], stage0_42[235], stage0_42[236], stage0_42[237], stage0_42[238], stage0_42[239]},
      {stage1_44[39],stage1_43[95],stage1_42[100],stage1_41[127],stage1_40[188]}
   );
   gpc606_5 gpc1580 (
      {stage0_40[326], stage0_40[327], stage0_40[328], stage0_40[329], stage0_40[330], stage0_40[331]},
      {stage0_42[240], stage0_42[241], stage0_42[242], stage0_42[243], stage0_42[244], stage0_42[245]},
      {stage1_44[40],stage1_43[96],stage1_42[101],stage1_41[128],stage1_40[189]}
   );
   gpc606_5 gpc1581 (
      {stage0_40[332], stage0_40[333], stage0_40[334], stage0_40[335], stage0_40[336], stage0_40[337]},
      {stage0_42[246], stage0_42[247], stage0_42[248], stage0_42[249], stage0_42[250], stage0_42[251]},
      {stage1_44[41],stage1_43[97],stage1_42[102],stage1_41[129],stage1_40[190]}
   );
   gpc606_5 gpc1582 (
      {stage0_40[338], stage0_40[339], stage0_40[340], stage0_40[341], stage0_40[342], stage0_40[343]},
      {stage0_42[252], stage0_42[253], stage0_42[254], stage0_42[255], stage0_42[256], stage0_42[257]},
      {stage1_44[42],stage1_43[98],stage1_42[103],stage1_41[130],stage1_40[191]}
   );
   gpc606_5 gpc1583 (
      {stage0_40[344], stage0_40[345], stage0_40[346], stage0_40[347], stage0_40[348], stage0_40[349]},
      {stage0_42[258], stage0_42[259], stage0_42[260], stage0_42[261], stage0_42[262], stage0_42[263]},
      {stage1_44[43],stage1_43[99],stage1_42[104],stage1_41[131],stage1_40[192]}
   );
   gpc606_5 gpc1584 (
      {stage0_40[350], stage0_40[351], stage0_40[352], stage0_40[353], stage0_40[354], stage0_40[355]},
      {stage0_42[264], stage0_42[265], stage0_42[266], stage0_42[267], stage0_42[268], stage0_42[269]},
      {stage1_44[44],stage1_43[100],stage1_42[105],stage1_41[132],stage1_40[193]}
   );
   gpc606_5 gpc1585 (
      {stage0_40[356], stage0_40[357], stage0_40[358], stage0_40[359], stage0_40[360], stage0_40[361]},
      {stage0_42[270], stage0_42[271], stage0_42[272], stage0_42[273], stage0_42[274], stage0_42[275]},
      {stage1_44[45],stage1_43[101],stage1_42[106],stage1_41[133],stage1_40[194]}
   );
   gpc606_5 gpc1586 (
      {stage0_40[362], stage0_40[363], stage0_40[364], stage0_40[365], stage0_40[366], stage0_40[367]},
      {stage0_42[276], stage0_42[277], stage0_42[278], stage0_42[279], stage0_42[280], stage0_42[281]},
      {stage1_44[46],stage1_43[102],stage1_42[107],stage1_41[134],stage1_40[195]}
   );
   gpc606_5 gpc1587 (
      {stage0_40[368], stage0_40[369], stage0_40[370], stage0_40[371], stage0_40[372], stage0_40[373]},
      {stage0_42[282], stage0_42[283], stage0_42[284], stage0_42[285], stage0_42[286], stage0_42[287]},
      {stage1_44[47],stage1_43[103],stage1_42[108],stage1_41[135],stage1_40[196]}
   );
   gpc606_5 gpc1588 (
      {stage0_40[374], stage0_40[375], stage0_40[376], stage0_40[377], stage0_40[378], stage0_40[379]},
      {stage0_42[288], stage0_42[289], stage0_42[290], stage0_42[291], stage0_42[292], stage0_42[293]},
      {stage1_44[48],stage1_43[104],stage1_42[109],stage1_41[136],stage1_40[197]}
   );
   gpc606_5 gpc1589 (
      {stage0_41[336], stage0_41[337], stage0_41[338], stage0_41[339], stage0_41[340], stage0_41[341]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[49],stage1_43[105],stage1_42[110],stage1_41[137]}
   );
   gpc606_5 gpc1590 (
      {stage0_41[342], stage0_41[343], stage0_41[344], stage0_41[345], stage0_41[346], stage0_41[347]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[50],stage1_43[106],stage1_42[111],stage1_41[138]}
   );
   gpc606_5 gpc1591 (
      {stage0_41[348], stage0_41[349], stage0_41[350], stage0_41[351], stage0_41[352], stage0_41[353]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[51],stage1_43[107],stage1_42[112],stage1_41[139]}
   );
   gpc606_5 gpc1592 (
      {stage0_41[354], stage0_41[355], stage0_41[356], stage0_41[357], stage0_41[358], stage0_41[359]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[52],stage1_43[108],stage1_42[113],stage1_41[140]}
   );
   gpc606_5 gpc1593 (
      {stage0_41[360], stage0_41[361], stage0_41[362], stage0_41[363], stage0_41[364], stage0_41[365]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[53],stage1_43[109],stage1_42[114],stage1_41[141]}
   );
   gpc606_5 gpc1594 (
      {stage0_41[366], stage0_41[367], stage0_41[368], stage0_41[369], stage0_41[370], stage0_41[371]},
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage1_45[5],stage1_44[54],stage1_43[110],stage1_42[115],stage1_41[142]}
   );
   gpc606_5 gpc1595 (
      {stage0_41[372], stage0_41[373], stage0_41[374], stage0_41[375], stage0_41[376], stage0_41[377]},
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage1_45[6],stage1_44[55],stage1_43[111],stage1_42[116],stage1_41[143]}
   );
   gpc606_5 gpc1596 (
      {stage0_41[378], stage0_41[379], stage0_41[380], stage0_41[381], stage0_41[382], stage0_41[383]},
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage1_45[7],stage1_44[56],stage1_43[112],stage1_42[117],stage1_41[144]}
   );
   gpc606_5 gpc1597 (
      {stage0_41[384], stage0_41[385], stage0_41[386], stage0_41[387], stage0_41[388], stage0_41[389]},
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage1_45[8],stage1_44[57],stage1_43[113],stage1_42[118],stage1_41[145]}
   );
   gpc606_5 gpc1598 (
      {stage0_41[390], stage0_41[391], stage0_41[392], stage0_41[393], stage0_41[394], stage0_41[395]},
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage1_45[9],stage1_44[58],stage1_43[114],stage1_42[119],stage1_41[146]}
   );
   gpc606_5 gpc1599 (
      {stage0_41[396], stage0_41[397], stage0_41[398], stage0_41[399], stage0_41[400], stage0_41[401]},
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage1_45[10],stage1_44[59],stage1_43[115],stage1_42[120],stage1_41[147]}
   );
   gpc606_5 gpc1600 (
      {stage0_41[402], stage0_41[403], stage0_41[404], stage0_41[405], stage0_41[406], stage0_41[407]},
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage1_45[11],stage1_44[60],stage1_43[116],stage1_42[121],stage1_41[148]}
   );
   gpc606_5 gpc1601 (
      {stage0_41[408], stage0_41[409], stage0_41[410], stage0_41[411], stage0_41[412], stage0_41[413]},
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage1_45[12],stage1_44[61],stage1_43[117],stage1_42[122],stage1_41[149]}
   );
   gpc606_5 gpc1602 (
      {stage0_41[414], stage0_41[415], stage0_41[416], stage0_41[417], stage0_41[418], stage0_41[419]},
      {stage0_43[78], stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage1_45[13],stage1_44[62],stage1_43[118],stage1_42[123],stage1_41[150]}
   );
   gpc606_5 gpc1603 (
      {stage0_41[420], stage0_41[421], stage0_41[422], stage0_41[423], stage0_41[424], stage0_41[425]},
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88], stage0_43[89]},
      {stage1_45[14],stage1_44[63],stage1_43[119],stage1_42[124],stage1_41[151]}
   );
   gpc606_5 gpc1604 (
      {stage0_41[426], stage0_41[427], stage0_41[428], stage0_41[429], stage0_41[430], stage0_41[431]},
      {stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93], stage0_43[94], stage0_43[95]},
      {stage1_45[15],stage1_44[64],stage1_43[120],stage1_42[125],stage1_41[152]}
   );
   gpc615_5 gpc1605 (
      {stage0_41[432], stage0_41[433], stage0_41[434], stage0_41[435], stage0_41[436]},
      {stage0_42[294]},
      {stage0_43[96], stage0_43[97], stage0_43[98], stage0_43[99], stage0_43[100], stage0_43[101]},
      {stage1_45[16],stage1_44[65],stage1_43[121],stage1_42[126],stage1_41[153]}
   );
   gpc615_5 gpc1606 (
      {stage0_41[437], stage0_41[438], stage0_41[439], stage0_41[440], stage0_41[441]},
      {stage0_42[295]},
      {stage0_43[102], stage0_43[103], stage0_43[104], stage0_43[105], stage0_43[106], stage0_43[107]},
      {stage1_45[17],stage1_44[66],stage1_43[122],stage1_42[127],stage1_41[154]}
   );
   gpc615_5 gpc1607 (
      {stage0_41[442], stage0_41[443], stage0_41[444], stage0_41[445], stage0_41[446]},
      {stage0_42[296]},
      {stage0_43[108], stage0_43[109], stage0_43[110], stage0_43[111], stage0_43[112], stage0_43[113]},
      {stage1_45[18],stage1_44[67],stage1_43[123],stage1_42[128],stage1_41[155]}
   );
   gpc615_5 gpc1608 (
      {stage0_41[447], stage0_41[448], stage0_41[449], stage0_41[450], stage0_41[451]},
      {stage0_42[297]},
      {stage0_43[114], stage0_43[115], stage0_43[116], stage0_43[117], stage0_43[118], stage0_43[119]},
      {stage1_45[19],stage1_44[68],stage1_43[124],stage1_42[129],stage1_41[156]}
   );
   gpc615_5 gpc1609 (
      {stage0_41[452], stage0_41[453], stage0_41[454], stage0_41[455], stage0_41[456]},
      {stage0_42[298]},
      {stage0_43[120], stage0_43[121], stage0_43[122], stage0_43[123], stage0_43[124], stage0_43[125]},
      {stage1_45[20],stage1_44[69],stage1_43[125],stage1_42[130],stage1_41[157]}
   );
   gpc615_5 gpc1610 (
      {stage0_41[457], stage0_41[458], stage0_41[459], stage0_41[460], stage0_41[461]},
      {stage0_42[299]},
      {stage0_43[126], stage0_43[127], stage0_43[128], stage0_43[129], stage0_43[130], stage0_43[131]},
      {stage1_45[21],stage1_44[70],stage1_43[126],stage1_42[131],stage1_41[158]}
   );
   gpc615_5 gpc1611 (
      {stage0_41[462], stage0_41[463], stage0_41[464], stage0_41[465], stage0_41[466]},
      {stage0_42[300]},
      {stage0_43[132], stage0_43[133], stage0_43[134], stage0_43[135], stage0_43[136], stage0_43[137]},
      {stage1_45[22],stage1_44[71],stage1_43[127],stage1_42[132],stage1_41[159]}
   );
   gpc615_5 gpc1612 (
      {stage0_41[467], stage0_41[468], stage0_41[469], stage0_41[470], stage0_41[471]},
      {stage0_42[301]},
      {stage0_43[138], stage0_43[139], stage0_43[140], stage0_43[141], stage0_43[142], stage0_43[143]},
      {stage1_45[23],stage1_44[72],stage1_43[128],stage1_42[133],stage1_41[160]}
   );
   gpc615_5 gpc1613 (
      {stage0_41[472], stage0_41[473], stage0_41[474], stage0_41[475], stage0_41[476]},
      {stage0_42[302]},
      {stage0_43[144], stage0_43[145], stage0_43[146], stage0_43[147], stage0_43[148], stage0_43[149]},
      {stage1_45[24],stage1_44[73],stage1_43[129],stage1_42[134],stage1_41[161]}
   );
   gpc615_5 gpc1614 (
      {stage0_42[303], stage0_42[304], stage0_42[305], stage0_42[306], stage0_42[307]},
      {stage0_43[150]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[25],stage1_44[74],stage1_43[130],stage1_42[135]}
   );
   gpc615_5 gpc1615 (
      {stage0_42[308], stage0_42[309], stage0_42[310], stage0_42[311], stage0_42[312]},
      {stage0_43[151]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[26],stage1_44[75],stage1_43[131],stage1_42[136]}
   );
   gpc615_5 gpc1616 (
      {stage0_42[313], stage0_42[314], stage0_42[315], stage0_42[316], stage0_42[317]},
      {stage0_43[152]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[27],stage1_44[76],stage1_43[132],stage1_42[137]}
   );
   gpc615_5 gpc1617 (
      {stage0_42[318], stage0_42[319], stage0_42[320], stage0_42[321], stage0_42[322]},
      {stage0_43[153]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[28],stage1_44[77],stage1_43[133],stage1_42[138]}
   );
   gpc615_5 gpc1618 (
      {stage0_42[323], stage0_42[324], stage0_42[325], stage0_42[326], stage0_42[327]},
      {stage0_43[154]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[29],stage1_44[78],stage1_43[134],stage1_42[139]}
   );
   gpc615_5 gpc1619 (
      {stage0_42[328], stage0_42[329], stage0_42[330], stage0_42[331], stage0_42[332]},
      {stage0_43[155]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[30],stage1_44[79],stage1_43[135],stage1_42[140]}
   );
   gpc615_5 gpc1620 (
      {stage0_42[333], stage0_42[334], stage0_42[335], stage0_42[336], stage0_42[337]},
      {stage0_43[156]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[31],stage1_44[80],stage1_43[136],stage1_42[141]}
   );
   gpc615_5 gpc1621 (
      {stage0_42[338], stage0_42[339], stage0_42[340], stage0_42[341], stage0_42[342]},
      {stage0_43[157]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[32],stage1_44[81],stage1_43[137],stage1_42[142]}
   );
   gpc615_5 gpc1622 (
      {stage0_42[343], stage0_42[344], stage0_42[345], stage0_42[346], stage0_42[347]},
      {stage0_43[158]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[33],stage1_44[82],stage1_43[138],stage1_42[143]}
   );
   gpc615_5 gpc1623 (
      {stage0_42[348], stage0_42[349], stage0_42[350], stage0_42[351], stage0_42[352]},
      {stage0_43[159]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[34],stage1_44[83],stage1_43[139],stage1_42[144]}
   );
   gpc615_5 gpc1624 (
      {stage0_42[353], stage0_42[354], stage0_42[355], stage0_42[356], stage0_42[357]},
      {stage0_43[160]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[35],stage1_44[84],stage1_43[140],stage1_42[145]}
   );
   gpc615_5 gpc1625 (
      {stage0_42[358], stage0_42[359], stage0_42[360], stage0_42[361], stage0_42[362]},
      {stage0_43[161]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[36],stage1_44[85],stage1_43[141],stage1_42[146]}
   );
   gpc615_5 gpc1626 (
      {stage0_42[363], stage0_42[364], stage0_42[365], stage0_42[366], stage0_42[367]},
      {stage0_43[162]},
      {stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76], stage0_44[77]},
      {stage1_46[12],stage1_45[37],stage1_44[86],stage1_43[142],stage1_42[147]}
   );
   gpc615_5 gpc1627 (
      {stage0_42[368], stage0_42[369], stage0_42[370], stage0_42[371], stage0_42[372]},
      {stage0_43[163]},
      {stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82], stage0_44[83]},
      {stage1_46[13],stage1_45[38],stage1_44[87],stage1_43[143],stage1_42[148]}
   );
   gpc615_5 gpc1628 (
      {stage0_42[373], stage0_42[374], stage0_42[375], stage0_42[376], stage0_42[377]},
      {stage0_43[164]},
      {stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88], stage0_44[89]},
      {stage1_46[14],stage1_45[39],stage1_44[88],stage1_43[144],stage1_42[149]}
   );
   gpc615_5 gpc1629 (
      {stage0_42[378], stage0_42[379], stage0_42[380], stage0_42[381], stage0_42[382]},
      {stage0_43[165]},
      {stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94], stage0_44[95]},
      {stage1_46[15],stage1_45[40],stage1_44[89],stage1_43[145],stage1_42[150]}
   );
   gpc615_5 gpc1630 (
      {stage0_42[383], stage0_42[384], stage0_42[385], stage0_42[386], stage0_42[387]},
      {stage0_43[166]},
      {stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100], stage0_44[101]},
      {stage1_46[16],stage1_45[41],stage1_44[90],stage1_43[146],stage1_42[151]}
   );
   gpc615_5 gpc1631 (
      {stage0_42[388], stage0_42[389], stage0_42[390], stage0_42[391], stage0_42[392]},
      {stage0_43[167]},
      {stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106], stage0_44[107]},
      {stage1_46[17],stage1_45[42],stage1_44[91],stage1_43[147],stage1_42[152]}
   );
   gpc615_5 gpc1632 (
      {stage0_42[393], stage0_42[394], stage0_42[395], stage0_42[396], stage0_42[397]},
      {stage0_43[168]},
      {stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112], stage0_44[113]},
      {stage1_46[18],stage1_45[43],stage1_44[92],stage1_43[148],stage1_42[153]}
   );
   gpc615_5 gpc1633 (
      {stage0_42[398], stage0_42[399], stage0_42[400], stage0_42[401], stage0_42[402]},
      {stage0_43[169]},
      {stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118], stage0_44[119]},
      {stage1_46[19],stage1_45[44],stage1_44[93],stage1_43[149],stage1_42[154]}
   );
   gpc615_5 gpc1634 (
      {stage0_42[403], stage0_42[404], stage0_42[405], stage0_42[406], stage0_42[407]},
      {stage0_43[170]},
      {stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124], stage0_44[125]},
      {stage1_46[20],stage1_45[45],stage1_44[94],stage1_43[150],stage1_42[155]}
   );
   gpc615_5 gpc1635 (
      {stage0_42[408], stage0_42[409], stage0_42[410], stage0_42[411], stage0_42[412]},
      {stage0_43[171]},
      {stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130], stage0_44[131]},
      {stage1_46[21],stage1_45[46],stage1_44[95],stage1_43[151],stage1_42[156]}
   );
   gpc615_5 gpc1636 (
      {stage0_42[413], stage0_42[414], stage0_42[415], stage0_42[416], stage0_42[417]},
      {stage0_43[172]},
      {stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136], stage0_44[137]},
      {stage1_46[22],stage1_45[47],stage1_44[96],stage1_43[152],stage1_42[157]}
   );
   gpc615_5 gpc1637 (
      {stage0_42[418], stage0_42[419], stage0_42[420], stage0_42[421], stage0_42[422]},
      {stage0_43[173]},
      {stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142], stage0_44[143]},
      {stage1_46[23],stage1_45[48],stage1_44[97],stage1_43[153],stage1_42[158]}
   );
   gpc615_5 gpc1638 (
      {stage0_42[423], stage0_42[424], stage0_42[425], stage0_42[426], stage0_42[427]},
      {stage0_43[174]},
      {stage0_44[144], stage0_44[145], stage0_44[146], stage0_44[147], stage0_44[148], stage0_44[149]},
      {stage1_46[24],stage1_45[49],stage1_44[98],stage1_43[154],stage1_42[159]}
   );
   gpc615_5 gpc1639 (
      {stage0_42[428], stage0_42[429], stage0_42[430], stage0_42[431], stage0_42[432]},
      {stage0_43[175]},
      {stage0_44[150], stage0_44[151], stage0_44[152], stage0_44[153], stage0_44[154], stage0_44[155]},
      {stage1_46[25],stage1_45[50],stage1_44[99],stage1_43[155],stage1_42[160]}
   );
   gpc615_5 gpc1640 (
      {stage0_42[433], stage0_42[434], stage0_42[435], stage0_42[436], stage0_42[437]},
      {stage0_43[176]},
      {stage0_44[156], stage0_44[157], stage0_44[158], stage0_44[159], stage0_44[160], stage0_44[161]},
      {stage1_46[26],stage1_45[51],stage1_44[100],stage1_43[156],stage1_42[161]}
   );
   gpc615_5 gpc1641 (
      {stage0_42[438], stage0_42[439], stage0_42[440], stage0_42[441], stage0_42[442]},
      {stage0_43[177]},
      {stage0_44[162], stage0_44[163], stage0_44[164], stage0_44[165], stage0_44[166], stage0_44[167]},
      {stage1_46[27],stage1_45[52],stage1_44[101],stage1_43[157],stage1_42[162]}
   );
   gpc615_5 gpc1642 (
      {stage0_42[443], stage0_42[444], stage0_42[445], stage0_42[446], stage0_42[447]},
      {stage0_43[178]},
      {stage0_44[168], stage0_44[169], stage0_44[170], stage0_44[171], stage0_44[172], stage0_44[173]},
      {stage1_46[28],stage1_45[53],stage1_44[102],stage1_43[158],stage1_42[163]}
   );
   gpc615_5 gpc1643 (
      {stage0_42[448], stage0_42[449], stage0_42[450], stage0_42[451], stage0_42[452]},
      {stage0_43[179]},
      {stage0_44[174], stage0_44[175], stage0_44[176], stage0_44[177], stage0_44[178], stage0_44[179]},
      {stage1_46[29],stage1_45[54],stage1_44[103],stage1_43[159],stage1_42[164]}
   );
   gpc615_5 gpc1644 (
      {stage0_42[453], stage0_42[454], stage0_42[455], stage0_42[456], stage0_42[457]},
      {stage0_43[180]},
      {stage0_44[180], stage0_44[181], stage0_44[182], stage0_44[183], stage0_44[184], stage0_44[185]},
      {stage1_46[30],stage1_45[55],stage1_44[104],stage1_43[160],stage1_42[165]}
   );
   gpc615_5 gpc1645 (
      {stage0_42[458], stage0_42[459], stage0_42[460], stage0_42[461], stage0_42[462]},
      {stage0_43[181]},
      {stage0_44[186], stage0_44[187], stage0_44[188], stage0_44[189], stage0_44[190], stage0_44[191]},
      {stage1_46[31],stage1_45[56],stage1_44[105],stage1_43[161],stage1_42[166]}
   );
   gpc615_5 gpc1646 (
      {stage0_42[463], stage0_42[464], stage0_42[465], stage0_42[466], stage0_42[467]},
      {stage0_43[182]},
      {stage0_44[192], stage0_44[193], stage0_44[194], stage0_44[195], stage0_44[196], stage0_44[197]},
      {stage1_46[32],stage1_45[57],stage1_44[106],stage1_43[162],stage1_42[167]}
   );
   gpc615_5 gpc1647 (
      {stage0_42[468], stage0_42[469], stage0_42[470], stage0_42[471], stage0_42[472]},
      {stage0_43[183]},
      {stage0_44[198], stage0_44[199], stage0_44[200], stage0_44[201], stage0_44[202], stage0_44[203]},
      {stage1_46[33],stage1_45[58],stage1_44[107],stage1_43[163],stage1_42[168]}
   );
   gpc615_5 gpc1648 (
      {stage0_42[473], stage0_42[474], stage0_42[475], stage0_42[476], stage0_42[477]},
      {stage0_43[184]},
      {stage0_44[204], stage0_44[205], stage0_44[206], stage0_44[207], stage0_44[208], stage0_44[209]},
      {stage1_46[34],stage1_45[59],stage1_44[108],stage1_43[164],stage1_42[169]}
   );
   gpc615_5 gpc1649 (
      {stage0_42[478], stage0_42[479], stage0_42[480], stage0_42[481], stage0_42[482]},
      {stage0_43[185]},
      {stage0_44[210], stage0_44[211], stage0_44[212], stage0_44[213], stage0_44[214], stage0_44[215]},
      {stage1_46[35],stage1_45[60],stage1_44[109],stage1_43[165],stage1_42[170]}
   );
   gpc615_5 gpc1650 (
      {stage0_43[186], stage0_43[187], stage0_43[188], stage0_43[189], stage0_43[190]},
      {stage0_44[216]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[36],stage1_45[61],stage1_44[110],stage1_43[166]}
   );
   gpc615_5 gpc1651 (
      {stage0_43[191], stage0_43[192], stage0_43[193], stage0_43[194], stage0_43[195]},
      {stage0_44[217]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[37],stage1_45[62],stage1_44[111],stage1_43[167]}
   );
   gpc615_5 gpc1652 (
      {stage0_43[196], stage0_43[197], stage0_43[198], stage0_43[199], stage0_43[200]},
      {stage0_44[218]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[38],stage1_45[63],stage1_44[112],stage1_43[168]}
   );
   gpc615_5 gpc1653 (
      {stage0_43[201], stage0_43[202], stage0_43[203], stage0_43[204], stage0_43[205]},
      {stage0_44[219]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[39],stage1_45[64],stage1_44[113],stage1_43[169]}
   );
   gpc615_5 gpc1654 (
      {stage0_43[206], stage0_43[207], stage0_43[208], stage0_43[209], stage0_43[210]},
      {stage0_44[220]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[40],stage1_45[65],stage1_44[114],stage1_43[170]}
   );
   gpc615_5 gpc1655 (
      {stage0_43[211], stage0_43[212], stage0_43[213], stage0_43[214], stage0_43[215]},
      {stage0_44[221]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[41],stage1_45[66],stage1_44[115],stage1_43[171]}
   );
   gpc615_5 gpc1656 (
      {stage0_43[216], stage0_43[217], stage0_43[218], stage0_43[219], stage0_43[220]},
      {stage0_44[222]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[42],stage1_45[67],stage1_44[116],stage1_43[172]}
   );
   gpc615_5 gpc1657 (
      {stage0_43[221], stage0_43[222], stage0_43[223], stage0_43[224], stage0_43[225]},
      {stage0_44[223]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[43],stage1_45[68],stage1_44[117],stage1_43[173]}
   );
   gpc615_5 gpc1658 (
      {stage0_43[226], stage0_43[227], stage0_43[228], stage0_43[229], stage0_43[230]},
      {stage0_44[224]},
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage1_47[8],stage1_46[44],stage1_45[69],stage1_44[118],stage1_43[174]}
   );
   gpc615_5 gpc1659 (
      {stage0_43[231], stage0_43[232], stage0_43[233], stage0_43[234], stage0_43[235]},
      {stage0_44[225]},
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage1_47[9],stage1_46[45],stage1_45[70],stage1_44[119],stage1_43[175]}
   );
   gpc615_5 gpc1660 (
      {stage0_43[236], stage0_43[237], stage0_43[238], stage0_43[239], stage0_43[240]},
      {stage0_44[226]},
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage1_47[10],stage1_46[46],stage1_45[71],stage1_44[120],stage1_43[176]}
   );
   gpc615_5 gpc1661 (
      {stage0_43[241], stage0_43[242], stage0_43[243], stage0_43[244], stage0_43[245]},
      {stage0_44[227]},
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage1_47[11],stage1_46[47],stage1_45[72],stage1_44[121],stage1_43[177]}
   );
   gpc615_5 gpc1662 (
      {stage0_43[246], stage0_43[247], stage0_43[248], stage0_43[249], stage0_43[250]},
      {stage0_44[228]},
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage1_47[12],stage1_46[48],stage1_45[73],stage1_44[122],stage1_43[178]}
   );
   gpc615_5 gpc1663 (
      {stage0_43[251], stage0_43[252], stage0_43[253], stage0_43[254], stage0_43[255]},
      {stage0_44[229]},
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage1_47[13],stage1_46[49],stage1_45[74],stage1_44[123],stage1_43[179]}
   );
   gpc615_5 gpc1664 (
      {stage0_43[256], stage0_43[257], stage0_43[258], stage0_43[259], stage0_43[260]},
      {stage0_44[230]},
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage1_47[14],stage1_46[50],stage1_45[75],stage1_44[124],stage1_43[180]}
   );
   gpc615_5 gpc1665 (
      {stage0_43[261], stage0_43[262], stage0_43[263], stage0_43[264], stage0_43[265]},
      {stage0_44[231]},
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage1_47[15],stage1_46[51],stage1_45[76],stage1_44[125],stage1_43[181]}
   );
   gpc615_5 gpc1666 (
      {stage0_43[266], stage0_43[267], stage0_43[268], stage0_43[269], stage0_43[270]},
      {stage0_44[232]},
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage1_47[16],stage1_46[52],stage1_45[77],stage1_44[126],stage1_43[182]}
   );
   gpc615_5 gpc1667 (
      {stage0_43[271], stage0_43[272], stage0_43[273], stage0_43[274], stage0_43[275]},
      {stage0_44[233]},
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage1_47[17],stage1_46[53],stage1_45[78],stage1_44[127],stage1_43[183]}
   );
   gpc615_5 gpc1668 (
      {stage0_43[276], stage0_43[277], stage0_43[278], stage0_43[279], stage0_43[280]},
      {stage0_44[234]},
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage1_47[18],stage1_46[54],stage1_45[79],stage1_44[128],stage1_43[184]}
   );
   gpc615_5 gpc1669 (
      {stage0_43[281], stage0_43[282], stage0_43[283], stage0_43[284], stage0_43[285]},
      {stage0_44[235]},
      {stage0_45[114], stage0_45[115], stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119]},
      {stage1_47[19],stage1_46[55],stage1_45[80],stage1_44[129],stage1_43[185]}
   );
   gpc615_5 gpc1670 (
      {stage0_43[286], stage0_43[287], stage0_43[288], stage0_43[289], stage0_43[290]},
      {stage0_44[236]},
      {stage0_45[120], stage0_45[121], stage0_45[122], stage0_45[123], stage0_45[124], stage0_45[125]},
      {stage1_47[20],stage1_46[56],stage1_45[81],stage1_44[130],stage1_43[186]}
   );
   gpc615_5 gpc1671 (
      {stage0_43[291], stage0_43[292], stage0_43[293], stage0_43[294], stage0_43[295]},
      {stage0_44[237]},
      {stage0_45[126], stage0_45[127], stage0_45[128], stage0_45[129], stage0_45[130], stage0_45[131]},
      {stage1_47[21],stage1_46[57],stage1_45[82],stage1_44[131],stage1_43[187]}
   );
   gpc615_5 gpc1672 (
      {stage0_43[296], stage0_43[297], stage0_43[298], stage0_43[299], stage0_43[300]},
      {stage0_44[238]},
      {stage0_45[132], stage0_45[133], stage0_45[134], stage0_45[135], stage0_45[136], stage0_45[137]},
      {stage1_47[22],stage1_46[58],stage1_45[83],stage1_44[132],stage1_43[188]}
   );
   gpc615_5 gpc1673 (
      {stage0_43[301], stage0_43[302], stage0_43[303], stage0_43[304], stage0_43[305]},
      {stage0_44[239]},
      {stage0_45[138], stage0_45[139], stage0_45[140], stage0_45[141], stage0_45[142], stage0_45[143]},
      {stage1_47[23],stage1_46[59],stage1_45[84],stage1_44[133],stage1_43[189]}
   );
   gpc615_5 gpc1674 (
      {stage0_43[306], stage0_43[307], stage0_43[308], stage0_43[309], stage0_43[310]},
      {stage0_44[240]},
      {stage0_45[144], stage0_45[145], stage0_45[146], stage0_45[147], stage0_45[148], stage0_45[149]},
      {stage1_47[24],stage1_46[60],stage1_45[85],stage1_44[134],stage1_43[190]}
   );
   gpc615_5 gpc1675 (
      {stage0_43[311], stage0_43[312], stage0_43[313], stage0_43[314], stage0_43[315]},
      {stage0_44[241]},
      {stage0_45[150], stage0_45[151], stage0_45[152], stage0_45[153], stage0_45[154], stage0_45[155]},
      {stage1_47[25],stage1_46[61],stage1_45[86],stage1_44[135],stage1_43[191]}
   );
   gpc615_5 gpc1676 (
      {stage0_43[316], stage0_43[317], stage0_43[318], stage0_43[319], stage0_43[320]},
      {stage0_44[242]},
      {stage0_45[156], stage0_45[157], stage0_45[158], stage0_45[159], stage0_45[160], stage0_45[161]},
      {stage1_47[26],stage1_46[62],stage1_45[87],stage1_44[136],stage1_43[192]}
   );
   gpc615_5 gpc1677 (
      {stage0_43[321], stage0_43[322], stage0_43[323], stage0_43[324], stage0_43[325]},
      {stage0_44[243]},
      {stage0_45[162], stage0_45[163], stage0_45[164], stage0_45[165], stage0_45[166], stage0_45[167]},
      {stage1_47[27],stage1_46[63],stage1_45[88],stage1_44[137],stage1_43[193]}
   );
   gpc615_5 gpc1678 (
      {stage0_43[326], stage0_43[327], stage0_43[328], stage0_43[329], stage0_43[330]},
      {stage0_44[244]},
      {stage0_45[168], stage0_45[169], stage0_45[170], stage0_45[171], stage0_45[172], stage0_45[173]},
      {stage1_47[28],stage1_46[64],stage1_45[89],stage1_44[138],stage1_43[194]}
   );
   gpc615_5 gpc1679 (
      {stage0_43[331], stage0_43[332], stage0_43[333], stage0_43[334], stage0_43[335]},
      {stage0_44[245]},
      {stage0_45[174], stage0_45[175], stage0_45[176], stage0_45[177], stage0_45[178], stage0_45[179]},
      {stage1_47[29],stage1_46[65],stage1_45[90],stage1_44[139],stage1_43[195]}
   );
   gpc615_5 gpc1680 (
      {stage0_43[336], stage0_43[337], stage0_43[338], stage0_43[339], stage0_43[340]},
      {stage0_44[246]},
      {stage0_45[180], stage0_45[181], stage0_45[182], stage0_45[183], stage0_45[184], stage0_45[185]},
      {stage1_47[30],stage1_46[66],stage1_45[91],stage1_44[140],stage1_43[196]}
   );
   gpc615_5 gpc1681 (
      {stage0_43[341], stage0_43[342], stage0_43[343], stage0_43[344], stage0_43[345]},
      {stage0_44[247]},
      {stage0_45[186], stage0_45[187], stage0_45[188], stage0_45[189], stage0_45[190], stage0_45[191]},
      {stage1_47[31],stage1_46[67],stage1_45[92],stage1_44[141],stage1_43[197]}
   );
   gpc615_5 gpc1682 (
      {stage0_43[346], stage0_43[347], stage0_43[348], stage0_43[349], stage0_43[350]},
      {stage0_44[248]},
      {stage0_45[192], stage0_45[193], stage0_45[194], stage0_45[195], stage0_45[196], stage0_45[197]},
      {stage1_47[32],stage1_46[68],stage1_45[93],stage1_44[142],stage1_43[198]}
   );
   gpc615_5 gpc1683 (
      {stage0_43[351], stage0_43[352], stage0_43[353], stage0_43[354], stage0_43[355]},
      {stage0_44[249]},
      {stage0_45[198], stage0_45[199], stage0_45[200], stage0_45[201], stage0_45[202], stage0_45[203]},
      {stage1_47[33],stage1_46[69],stage1_45[94],stage1_44[143],stage1_43[199]}
   );
   gpc615_5 gpc1684 (
      {stage0_43[356], stage0_43[357], stage0_43[358], stage0_43[359], stage0_43[360]},
      {stage0_44[250]},
      {stage0_45[204], stage0_45[205], stage0_45[206], stage0_45[207], stage0_45[208], stage0_45[209]},
      {stage1_47[34],stage1_46[70],stage1_45[95],stage1_44[144],stage1_43[200]}
   );
   gpc615_5 gpc1685 (
      {stage0_43[361], stage0_43[362], stage0_43[363], stage0_43[364], stage0_43[365]},
      {stage0_44[251]},
      {stage0_45[210], stage0_45[211], stage0_45[212], stage0_45[213], stage0_45[214], stage0_45[215]},
      {stage1_47[35],stage1_46[71],stage1_45[96],stage1_44[145],stage1_43[201]}
   );
   gpc615_5 gpc1686 (
      {stage0_43[366], stage0_43[367], stage0_43[368], stage0_43[369], stage0_43[370]},
      {stage0_44[252]},
      {stage0_45[216], stage0_45[217], stage0_45[218], stage0_45[219], stage0_45[220], stage0_45[221]},
      {stage1_47[36],stage1_46[72],stage1_45[97],stage1_44[146],stage1_43[202]}
   );
   gpc615_5 gpc1687 (
      {stage0_43[371], stage0_43[372], stage0_43[373], stage0_43[374], stage0_43[375]},
      {stage0_44[253]},
      {stage0_45[222], stage0_45[223], stage0_45[224], stage0_45[225], stage0_45[226], stage0_45[227]},
      {stage1_47[37],stage1_46[73],stage1_45[98],stage1_44[147],stage1_43[203]}
   );
   gpc615_5 gpc1688 (
      {stage0_43[376], stage0_43[377], stage0_43[378], stage0_43[379], stage0_43[380]},
      {stage0_44[254]},
      {stage0_45[228], stage0_45[229], stage0_45[230], stage0_45[231], stage0_45[232], stage0_45[233]},
      {stage1_47[38],stage1_46[74],stage1_45[99],stage1_44[148],stage1_43[204]}
   );
   gpc615_5 gpc1689 (
      {stage0_43[381], stage0_43[382], stage0_43[383], stage0_43[384], stage0_43[385]},
      {stage0_44[255]},
      {stage0_45[234], stage0_45[235], stage0_45[236], stage0_45[237], stage0_45[238], stage0_45[239]},
      {stage1_47[39],stage1_46[75],stage1_45[100],stage1_44[149],stage1_43[205]}
   );
   gpc615_5 gpc1690 (
      {stage0_43[386], stage0_43[387], stage0_43[388], stage0_43[389], stage0_43[390]},
      {stage0_44[256]},
      {stage0_45[240], stage0_45[241], stage0_45[242], stage0_45[243], stage0_45[244], stage0_45[245]},
      {stage1_47[40],stage1_46[76],stage1_45[101],stage1_44[150],stage1_43[206]}
   );
   gpc615_5 gpc1691 (
      {stage0_43[391], stage0_43[392], stage0_43[393], stage0_43[394], stage0_43[395]},
      {stage0_44[257]},
      {stage0_45[246], stage0_45[247], stage0_45[248], stage0_45[249], stage0_45[250], stage0_45[251]},
      {stage1_47[41],stage1_46[77],stage1_45[102],stage1_44[151],stage1_43[207]}
   );
   gpc615_5 gpc1692 (
      {stage0_43[396], stage0_43[397], stage0_43[398], stage0_43[399], stage0_43[400]},
      {stage0_44[258]},
      {stage0_45[252], stage0_45[253], stage0_45[254], stage0_45[255], stage0_45[256], stage0_45[257]},
      {stage1_47[42],stage1_46[78],stage1_45[103],stage1_44[152],stage1_43[208]}
   );
   gpc615_5 gpc1693 (
      {stage0_43[401], stage0_43[402], stage0_43[403], stage0_43[404], stage0_43[405]},
      {stage0_44[259]},
      {stage0_45[258], stage0_45[259], stage0_45[260], stage0_45[261], stage0_45[262], stage0_45[263]},
      {stage1_47[43],stage1_46[79],stage1_45[104],stage1_44[153],stage1_43[209]}
   );
   gpc615_5 gpc1694 (
      {stage0_43[406], stage0_43[407], stage0_43[408], stage0_43[409], stage0_43[410]},
      {stage0_44[260]},
      {stage0_45[264], stage0_45[265], stage0_45[266], stage0_45[267], stage0_45[268], stage0_45[269]},
      {stage1_47[44],stage1_46[80],stage1_45[105],stage1_44[154],stage1_43[210]}
   );
   gpc615_5 gpc1695 (
      {stage0_43[411], stage0_43[412], stage0_43[413], stage0_43[414], stage0_43[415]},
      {stage0_44[261]},
      {stage0_45[270], stage0_45[271], stage0_45[272], stage0_45[273], stage0_45[274], stage0_45[275]},
      {stage1_47[45],stage1_46[81],stage1_45[106],stage1_44[155],stage1_43[211]}
   );
   gpc615_5 gpc1696 (
      {stage0_43[416], stage0_43[417], stage0_43[418], stage0_43[419], stage0_43[420]},
      {stage0_44[262]},
      {stage0_45[276], stage0_45[277], stage0_45[278], stage0_45[279], stage0_45[280], stage0_45[281]},
      {stage1_47[46],stage1_46[82],stage1_45[107],stage1_44[156],stage1_43[212]}
   );
   gpc615_5 gpc1697 (
      {stage0_43[421], stage0_43[422], stage0_43[423], stage0_43[424], stage0_43[425]},
      {stage0_44[263]},
      {stage0_45[282], stage0_45[283], stage0_45[284], stage0_45[285], stage0_45[286], stage0_45[287]},
      {stage1_47[47],stage1_46[83],stage1_45[108],stage1_44[157],stage1_43[213]}
   );
   gpc615_5 gpc1698 (
      {stage0_43[426], stage0_43[427], stage0_43[428], stage0_43[429], stage0_43[430]},
      {stage0_44[264]},
      {stage0_45[288], stage0_45[289], stage0_45[290], stage0_45[291], stage0_45[292], stage0_45[293]},
      {stage1_47[48],stage1_46[84],stage1_45[109],stage1_44[158],stage1_43[214]}
   );
   gpc615_5 gpc1699 (
      {stage0_43[431], stage0_43[432], stage0_43[433], stage0_43[434], stage0_43[435]},
      {stage0_44[265]},
      {stage0_45[294], stage0_45[295], stage0_45[296], stage0_45[297], stage0_45[298], stage0_45[299]},
      {stage1_47[49],stage1_46[85],stage1_45[110],stage1_44[159],stage1_43[215]}
   );
   gpc615_5 gpc1700 (
      {stage0_43[436], stage0_43[437], stage0_43[438], stage0_43[439], stage0_43[440]},
      {stage0_44[266]},
      {stage0_45[300], stage0_45[301], stage0_45[302], stage0_45[303], stage0_45[304], stage0_45[305]},
      {stage1_47[50],stage1_46[86],stage1_45[111],stage1_44[160],stage1_43[216]}
   );
   gpc615_5 gpc1701 (
      {stage0_43[441], stage0_43[442], stage0_43[443], stage0_43[444], stage0_43[445]},
      {stage0_44[267]},
      {stage0_45[306], stage0_45[307], stage0_45[308], stage0_45[309], stage0_45[310], stage0_45[311]},
      {stage1_47[51],stage1_46[87],stage1_45[112],stage1_44[161],stage1_43[217]}
   );
   gpc615_5 gpc1702 (
      {stage0_43[446], stage0_43[447], stage0_43[448], stage0_43[449], stage0_43[450]},
      {stage0_44[268]},
      {stage0_45[312], stage0_45[313], stage0_45[314], stage0_45[315], stage0_45[316], stage0_45[317]},
      {stage1_47[52],stage1_46[88],stage1_45[113],stage1_44[162],stage1_43[218]}
   );
   gpc615_5 gpc1703 (
      {stage0_44[269], stage0_44[270], stage0_44[271], stage0_44[272], stage0_44[273]},
      {stage0_45[318]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[53],stage1_46[89],stage1_45[114],stage1_44[163]}
   );
   gpc615_5 gpc1704 (
      {stage0_44[274], stage0_44[275], stage0_44[276], stage0_44[277], stage0_44[278]},
      {stage0_45[319]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[54],stage1_46[90],stage1_45[115],stage1_44[164]}
   );
   gpc615_5 gpc1705 (
      {stage0_44[279], stage0_44[280], stage0_44[281], stage0_44[282], stage0_44[283]},
      {stage0_45[320]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[55],stage1_46[91],stage1_45[116],stage1_44[165]}
   );
   gpc615_5 gpc1706 (
      {stage0_44[284], stage0_44[285], stage0_44[286], stage0_44[287], stage0_44[288]},
      {stage0_45[321]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[56],stage1_46[92],stage1_45[117],stage1_44[166]}
   );
   gpc615_5 gpc1707 (
      {stage0_44[289], stage0_44[290], stage0_44[291], stage0_44[292], stage0_44[293]},
      {stage0_45[322]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[57],stage1_46[93],stage1_45[118],stage1_44[167]}
   );
   gpc615_5 gpc1708 (
      {stage0_44[294], stage0_44[295], stage0_44[296], stage0_44[297], stage0_44[298]},
      {stage0_45[323]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[58],stage1_46[94],stage1_45[119],stage1_44[168]}
   );
   gpc615_5 gpc1709 (
      {stage0_44[299], stage0_44[300], stage0_44[301], stage0_44[302], stage0_44[303]},
      {stage0_45[324]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[59],stage1_46[95],stage1_45[120],stage1_44[169]}
   );
   gpc615_5 gpc1710 (
      {stage0_44[304], stage0_44[305], stage0_44[306], stage0_44[307], stage0_44[308]},
      {stage0_45[325]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[60],stage1_46[96],stage1_45[121],stage1_44[170]}
   );
   gpc615_5 gpc1711 (
      {stage0_44[309], stage0_44[310], stage0_44[311], stage0_44[312], stage0_44[313]},
      {stage0_45[326]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[61],stage1_46[97],stage1_45[122],stage1_44[171]}
   );
   gpc615_5 gpc1712 (
      {stage0_44[314], stage0_44[315], stage0_44[316], stage0_44[317], stage0_44[318]},
      {stage0_45[327]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[62],stage1_46[98],stage1_45[123],stage1_44[172]}
   );
   gpc615_5 gpc1713 (
      {stage0_44[319], stage0_44[320], stage0_44[321], stage0_44[322], stage0_44[323]},
      {stage0_45[328]},
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage1_48[10],stage1_47[63],stage1_46[99],stage1_45[124],stage1_44[173]}
   );
   gpc615_5 gpc1714 (
      {stage0_44[324], stage0_44[325], stage0_44[326], stage0_44[327], stage0_44[328]},
      {stage0_45[329]},
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70], stage0_46[71]},
      {stage1_48[11],stage1_47[64],stage1_46[100],stage1_45[125],stage1_44[174]}
   );
   gpc615_5 gpc1715 (
      {stage0_44[329], stage0_44[330], stage0_44[331], stage0_44[332], stage0_44[333]},
      {stage0_45[330]},
      {stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77]},
      {stage1_48[12],stage1_47[65],stage1_46[101],stage1_45[126],stage1_44[175]}
   );
   gpc615_5 gpc1716 (
      {stage0_44[334], stage0_44[335], stage0_44[336], stage0_44[337], stage0_44[338]},
      {stage0_45[331]},
      {stage0_46[78], stage0_46[79], stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83]},
      {stage1_48[13],stage1_47[66],stage1_46[102],stage1_45[127],stage1_44[176]}
   );
   gpc615_5 gpc1717 (
      {stage0_44[339], stage0_44[340], stage0_44[341], stage0_44[342], stage0_44[343]},
      {stage0_45[332]},
      {stage0_46[84], stage0_46[85], stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89]},
      {stage1_48[14],stage1_47[67],stage1_46[103],stage1_45[128],stage1_44[177]}
   );
   gpc615_5 gpc1718 (
      {stage0_44[344], stage0_44[345], stage0_44[346], stage0_44[347], stage0_44[348]},
      {stage0_45[333]},
      {stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage1_48[15],stage1_47[68],stage1_46[104],stage1_45[129],stage1_44[178]}
   );
   gpc615_5 gpc1719 (
      {stage0_44[349], stage0_44[350], stage0_44[351], stage0_44[352], stage0_44[353]},
      {stage0_45[334]},
      {stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100], stage0_46[101]},
      {stage1_48[16],stage1_47[69],stage1_46[105],stage1_45[130],stage1_44[179]}
   );
   gpc615_5 gpc1720 (
      {stage0_44[354], stage0_44[355], stage0_44[356], stage0_44[357], stage0_44[358]},
      {stage0_45[335]},
      {stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage1_48[17],stage1_47[70],stage1_46[106],stage1_45[131],stage1_44[180]}
   );
   gpc615_5 gpc1721 (
      {stage0_44[359], stage0_44[360], stage0_44[361], stage0_44[362], stage0_44[363]},
      {stage0_45[336]},
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113]},
      {stage1_48[18],stage1_47[71],stage1_46[107],stage1_45[132],stage1_44[181]}
   );
   gpc615_5 gpc1722 (
      {stage0_44[364], stage0_44[365], stage0_44[366], stage0_44[367], stage0_44[368]},
      {stage0_45[337]},
      {stage0_46[114], stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119]},
      {stage1_48[19],stage1_47[72],stage1_46[108],stage1_45[133],stage1_44[182]}
   );
   gpc615_5 gpc1723 (
      {stage0_44[369], stage0_44[370], stage0_44[371], stage0_44[372], stage0_44[373]},
      {stage0_45[338]},
      {stage0_46[120], stage0_46[121], stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125]},
      {stage1_48[20],stage1_47[73],stage1_46[109],stage1_45[134],stage1_44[183]}
   );
   gpc615_5 gpc1724 (
      {stage0_44[374], stage0_44[375], stage0_44[376], stage0_44[377], stage0_44[378]},
      {stage0_45[339]},
      {stage0_46[126], stage0_46[127], stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131]},
      {stage1_48[21],stage1_47[74],stage1_46[110],stage1_45[135],stage1_44[184]}
   );
   gpc615_5 gpc1725 (
      {stage0_44[379], stage0_44[380], stage0_44[381], stage0_44[382], stage0_44[383]},
      {stage0_45[340]},
      {stage0_46[132], stage0_46[133], stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137]},
      {stage1_48[22],stage1_47[75],stage1_46[111],stage1_45[136],stage1_44[185]}
   );
   gpc615_5 gpc1726 (
      {stage0_44[384], stage0_44[385], stage0_44[386], stage0_44[387], stage0_44[388]},
      {stage0_45[341]},
      {stage0_46[138], stage0_46[139], stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143]},
      {stage1_48[23],stage1_47[76],stage1_46[112],stage1_45[137],stage1_44[186]}
   );
   gpc615_5 gpc1727 (
      {stage0_44[389], stage0_44[390], stage0_44[391], stage0_44[392], stage0_44[393]},
      {stage0_45[342]},
      {stage0_46[144], stage0_46[145], stage0_46[146], stage0_46[147], stage0_46[148], stage0_46[149]},
      {stage1_48[24],stage1_47[77],stage1_46[113],stage1_45[138],stage1_44[187]}
   );
   gpc615_5 gpc1728 (
      {stage0_44[394], stage0_44[395], stage0_44[396], stage0_44[397], stage0_44[398]},
      {stage0_45[343]},
      {stage0_46[150], stage0_46[151], stage0_46[152], stage0_46[153], stage0_46[154], stage0_46[155]},
      {stage1_48[25],stage1_47[78],stage1_46[114],stage1_45[139],stage1_44[188]}
   );
   gpc615_5 gpc1729 (
      {stage0_44[399], stage0_44[400], stage0_44[401], stage0_44[402], stage0_44[403]},
      {stage0_45[344]},
      {stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159], stage0_46[160], stage0_46[161]},
      {stage1_48[26],stage1_47[79],stage1_46[115],stage1_45[140],stage1_44[189]}
   );
   gpc615_5 gpc1730 (
      {stage0_44[404], stage0_44[405], stage0_44[406], stage0_44[407], stage0_44[408]},
      {stage0_45[345]},
      {stage0_46[162], stage0_46[163], stage0_46[164], stage0_46[165], stage0_46[166], stage0_46[167]},
      {stage1_48[27],stage1_47[80],stage1_46[116],stage1_45[141],stage1_44[190]}
   );
   gpc615_5 gpc1731 (
      {stage0_44[409], stage0_44[410], stage0_44[411], stage0_44[412], stage0_44[413]},
      {stage0_45[346]},
      {stage0_46[168], stage0_46[169], stage0_46[170], stage0_46[171], stage0_46[172], stage0_46[173]},
      {stage1_48[28],stage1_47[81],stage1_46[117],stage1_45[142],stage1_44[191]}
   );
   gpc615_5 gpc1732 (
      {stage0_44[414], stage0_44[415], stage0_44[416], stage0_44[417], stage0_44[418]},
      {stage0_45[347]},
      {stage0_46[174], stage0_46[175], stage0_46[176], stage0_46[177], stage0_46[178], stage0_46[179]},
      {stage1_48[29],stage1_47[82],stage1_46[118],stage1_45[143],stage1_44[192]}
   );
   gpc615_5 gpc1733 (
      {stage0_44[419], stage0_44[420], stage0_44[421], stage0_44[422], stage0_44[423]},
      {stage0_45[348]},
      {stage0_46[180], stage0_46[181], stage0_46[182], stage0_46[183], stage0_46[184], stage0_46[185]},
      {stage1_48[30],stage1_47[83],stage1_46[119],stage1_45[144],stage1_44[193]}
   );
   gpc606_5 gpc1734 (
      {stage0_45[349], stage0_45[350], stage0_45[351], stage0_45[352], stage0_45[353], stage0_45[354]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[31],stage1_47[84],stage1_46[120],stage1_45[145]}
   );
   gpc606_5 gpc1735 (
      {stage0_45[355], stage0_45[356], stage0_45[357], stage0_45[358], stage0_45[359], stage0_45[360]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[32],stage1_47[85],stage1_46[121],stage1_45[146]}
   );
   gpc606_5 gpc1736 (
      {stage0_45[361], stage0_45[362], stage0_45[363], stage0_45[364], stage0_45[365], stage0_45[366]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[33],stage1_47[86],stage1_46[122],stage1_45[147]}
   );
   gpc606_5 gpc1737 (
      {stage0_45[367], stage0_45[368], stage0_45[369], stage0_45[370], stage0_45[371], stage0_45[372]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[34],stage1_47[87],stage1_46[123],stage1_45[148]}
   );
   gpc606_5 gpc1738 (
      {stage0_45[373], stage0_45[374], stage0_45[375], stage0_45[376], stage0_45[377], stage0_45[378]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[35],stage1_47[88],stage1_46[124],stage1_45[149]}
   );
   gpc606_5 gpc1739 (
      {stage0_45[379], stage0_45[380], stage0_45[381], stage0_45[382], stage0_45[383], stage0_45[384]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[36],stage1_47[89],stage1_46[125],stage1_45[150]}
   );
   gpc606_5 gpc1740 (
      {stage0_45[385], stage0_45[386], stage0_45[387], stage0_45[388], stage0_45[389], stage0_45[390]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[37],stage1_47[90],stage1_46[126],stage1_45[151]}
   );
   gpc606_5 gpc1741 (
      {stage0_45[391], stage0_45[392], stage0_45[393], stage0_45[394], stage0_45[395], stage0_45[396]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[38],stage1_47[91],stage1_46[127],stage1_45[152]}
   );
   gpc606_5 gpc1742 (
      {stage0_45[397], stage0_45[398], stage0_45[399], stage0_45[400], stage0_45[401], stage0_45[402]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[39],stage1_47[92],stage1_46[128],stage1_45[153]}
   );
   gpc606_5 gpc1743 (
      {stage0_45[403], stage0_45[404], stage0_45[405], stage0_45[406], stage0_45[407], stage0_45[408]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[40],stage1_47[93],stage1_46[129],stage1_45[154]}
   );
   gpc606_5 gpc1744 (
      {stage0_45[409], stage0_45[410], stage0_45[411], stage0_45[412], stage0_45[413], stage0_45[414]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[41],stage1_47[94],stage1_46[130],stage1_45[155]}
   );
   gpc606_5 gpc1745 (
      {stage0_45[415], stage0_45[416], stage0_45[417], stage0_45[418], stage0_45[419], stage0_45[420]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[42],stage1_47[95],stage1_46[131],stage1_45[156]}
   );
   gpc606_5 gpc1746 (
      {stage0_45[421], stage0_45[422], stage0_45[423], stage0_45[424], stage0_45[425], stage0_45[426]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[43],stage1_47[96],stage1_46[132],stage1_45[157]}
   );
   gpc606_5 gpc1747 (
      {stage0_45[427], stage0_45[428], stage0_45[429], stage0_45[430], stage0_45[431], stage0_45[432]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[44],stage1_47[97],stage1_46[133],stage1_45[158]}
   );
   gpc135_4 gpc1748 (
      {stage0_46[186], stage0_46[187], stage0_46[188], stage0_46[189], stage0_46[190]},
      {stage0_47[84], stage0_47[85], stage0_47[86]},
      {stage0_48[0]},
      {stage1_49[14],stage1_48[45],stage1_47[98],stage1_46[134]}
   );
   gpc135_4 gpc1749 (
      {stage0_46[191], stage0_46[192], stage0_46[193], stage0_46[194], stage0_46[195]},
      {stage0_47[87], stage0_47[88], stage0_47[89]},
      {stage0_48[1]},
      {stage1_49[15],stage1_48[46],stage1_47[99],stage1_46[135]}
   );
   gpc135_4 gpc1750 (
      {stage0_46[196], stage0_46[197], stage0_46[198], stage0_46[199], stage0_46[200]},
      {stage0_47[90], stage0_47[91], stage0_47[92]},
      {stage0_48[2]},
      {stage1_49[16],stage1_48[47],stage1_47[100],stage1_46[136]}
   );
   gpc135_4 gpc1751 (
      {stage0_46[201], stage0_46[202], stage0_46[203], stage0_46[204], stage0_46[205]},
      {stage0_47[93], stage0_47[94], stage0_47[95]},
      {stage0_48[3]},
      {stage1_49[17],stage1_48[48],stage1_47[101],stage1_46[137]}
   );
   gpc135_4 gpc1752 (
      {stage0_46[206], stage0_46[207], stage0_46[208], stage0_46[209], stage0_46[210]},
      {stage0_47[96], stage0_47[97], stage0_47[98]},
      {stage0_48[4]},
      {stage1_49[18],stage1_48[49],stage1_47[102],stage1_46[138]}
   );
   gpc135_4 gpc1753 (
      {stage0_46[211], stage0_46[212], stage0_46[213], stage0_46[214], stage0_46[215]},
      {stage0_47[99], stage0_47[100], stage0_47[101]},
      {stage0_48[5]},
      {stage1_49[19],stage1_48[50],stage1_47[103],stage1_46[139]}
   );
   gpc135_4 gpc1754 (
      {stage0_46[216], stage0_46[217], stage0_46[218], stage0_46[219], stage0_46[220]},
      {stage0_47[102], stage0_47[103], stage0_47[104]},
      {stage0_48[6]},
      {stage1_49[20],stage1_48[51],stage1_47[104],stage1_46[140]}
   );
   gpc135_4 gpc1755 (
      {stage0_46[221], stage0_46[222], stage0_46[223], stage0_46[224], stage0_46[225]},
      {stage0_47[105], stage0_47[106], stage0_47[107]},
      {stage0_48[7]},
      {stage1_49[21],stage1_48[52],stage1_47[105],stage1_46[141]}
   );
   gpc135_4 gpc1756 (
      {stage0_46[226], stage0_46[227], stage0_46[228], stage0_46[229], stage0_46[230]},
      {stage0_47[108], stage0_47[109], stage0_47[110]},
      {stage0_48[8]},
      {stage1_49[22],stage1_48[53],stage1_47[106],stage1_46[142]}
   );
   gpc135_4 gpc1757 (
      {stage0_46[231], stage0_46[232], stage0_46[233], stage0_46[234], stage0_46[235]},
      {stage0_47[111], stage0_47[112], stage0_47[113]},
      {stage0_48[9]},
      {stage1_49[23],stage1_48[54],stage1_47[107],stage1_46[143]}
   );
   gpc615_5 gpc1758 (
      {stage0_46[236], stage0_46[237], stage0_46[238], stage0_46[239], stage0_46[240]},
      {stage0_47[114]},
      {stage0_48[10], stage0_48[11], stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15]},
      {stage1_50[0],stage1_49[24],stage1_48[55],stage1_47[108],stage1_46[144]}
   );
   gpc615_5 gpc1759 (
      {stage0_46[241], stage0_46[242], stage0_46[243], stage0_46[244], stage0_46[245]},
      {stage0_47[115]},
      {stage0_48[16], stage0_48[17], stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21]},
      {stage1_50[1],stage1_49[25],stage1_48[56],stage1_47[109],stage1_46[145]}
   );
   gpc615_5 gpc1760 (
      {stage0_46[246], stage0_46[247], stage0_46[248], stage0_46[249], stage0_46[250]},
      {stage0_47[116]},
      {stage0_48[22], stage0_48[23], stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27]},
      {stage1_50[2],stage1_49[26],stage1_48[57],stage1_47[110],stage1_46[146]}
   );
   gpc615_5 gpc1761 (
      {stage0_46[251], stage0_46[252], stage0_46[253], stage0_46[254], stage0_46[255]},
      {stage0_47[117]},
      {stage0_48[28], stage0_48[29], stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33]},
      {stage1_50[3],stage1_49[27],stage1_48[58],stage1_47[111],stage1_46[147]}
   );
   gpc615_5 gpc1762 (
      {stage0_46[256], stage0_46[257], stage0_46[258], stage0_46[259], stage0_46[260]},
      {stage0_47[118]},
      {stage0_48[34], stage0_48[35], stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39]},
      {stage1_50[4],stage1_49[28],stage1_48[59],stage1_47[112],stage1_46[148]}
   );
   gpc615_5 gpc1763 (
      {stage0_46[261], stage0_46[262], stage0_46[263], stage0_46[264], stage0_46[265]},
      {stage0_47[119]},
      {stage0_48[40], stage0_48[41], stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45]},
      {stage1_50[5],stage1_49[29],stage1_48[60],stage1_47[113],stage1_46[149]}
   );
   gpc615_5 gpc1764 (
      {stage0_46[266], stage0_46[267], stage0_46[268], stage0_46[269], stage0_46[270]},
      {stage0_47[120]},
      {stage0_48[46], stage0_48[47], stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51]},
      {stage1_50[6],stage1_49[30],stage1_48[61],stage1_47[114],stage1_46[150]}
   );
   gpc615_5 gpc1765 (
      {stage0_46[271], stage0_46[272], stage0_46[273], stage0_46[274], stage0_46[275]},
      {stage0_47[121]},
      {stage0_48[52], stage0_48[53], stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57]},
      {stage1_50[7],stage1_49[31],stage1_48[62],stage1_47[115],stage1_46[151]}
   );
   gpc615_5 gpc1766 (
      {stage0_46[276], stage0_46[277], stage0_46[278], stage0_46[279], stage0_46[280]},
      {stage0_47[122]},
      {stage0_48[58], stage0_48[59], stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63]},
      {stage1_50[8],stage1_49[32],stage1_48[63],stage1_47[116],stage1_46[152]}
   );
   gpc615_5 gpc1767 (
      {stage0_46[281], stage0_46[282], stage0_46[283], stage0_46[284], stage0_46[285]},
      {stage0_47[123]},
      {stage0_48[64], stage0_48[65], stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69]},
      {stage1_50[9],stage1_49[33],stage1_48[64],stage1_47[117],stage1_46[153]}
   );
   gpc615_5 gpc1768 (
      {stage0_46[286], stage0_46[287], stage0_46[288], stage0_46[289], stage0_46[290]},
      {stage0_47[124]},
      {stage0_48[70], stage0_48[71], stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75]},
      {stage1_50[10],stage1_49[34],stage1_48[65],stage1_47[118],stage1_46[154]}
   );
   gpc615_5 gpc1769 (
      {stage0_46[291], stage0_46[292], stage0_46[293], stage0_46[294], stage0_46[295]},
      {stage0_47[125]},
      {stage0_48[76], stage0_48[77], stage0_48[78], stage0_48[79], stage0_48[80], stage0_48[81]},
      {stage1_50[11],stage1_49[35],stage1_48[66],stage1_47[119],stage1_46[155]}
   );
   gpc615_5 gpc1770 (
      {stage0_46[296], stage0_46[297], stage0_46[298], stage0_46[299], stage0_46[300]},
      {stage0_47[126]},
      {stage0_48[82], stage0_48[83], stage0_48[84], stage0_48[85], stage0_48[86], stage0_48[87]},
      {stage1_50[12],stage1_49[36],stage1_48[67],stage1_47[120],stage1_46[156]}
   );
   gpc615_5 gpc1771 (
      {stage0_46[301], stage0_46[302], stage0_46[303], stage0_46[304], stage0_46[305]},
      {stage0_47[127]},
      {stage0_48[88], stage0_48[89], stage0_48[90], stage0_48[91], stage0_48[92], stage0_48[93]},
      {stage1_50[13],stage1_49[37],stage1_48[68],stage1_47[121],stage1_46[157]}
   );
   gpc615_5 gpc1772 (
      {stage0_46[306], stage0_46[307], stage0_46[308], stage0_46[309], stage0_46[310]},
      {stage0_47[128]},
      {stage0_48[94], stage0_48[95], stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99]},
      {stage1_50[14],stage1_49[38],stage1_48[69],stage1_47[122],stage1_46[158]}
   );
   gpc615_5 gpc1773 (
      {stage0_46[311], stage0_46[312], stage0_46[313], stage0_46[314], stage0_46[315]},
      {stage0_47[129]},
      {stage0_48[100], stage0_48[101], stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105]},
      {stage1_50[15],stage1_49[39],stage1_48[70],stage1_47[123],stage1_46[159]}
   );
   gpc615_5 gpc1774 (
      {stage0_46[316], stage0_46[317], stage0_46[318], stage0_46[319], stage0_46[320]},
      {stage0_47[130]},
      {stage0_48[106], stage0_48[107], stage0_48[108], stage0_48[109], stage0_48[110], stage0_48[111]},
      {stage1_50[16],stage1_49[40],stage1_48[71],stage1_47[124],stage1_46[160]}
   );
   gpc615_5 gpc1775 (
      {stage0_46[321], stage0_46[322], stage0_46[323], stage0_46[324], stage0_46[325]},
      {stage0_47[131]},
      {stage0_48[112], stage0_48[113], stage0_48[114], stage0_48[115], stage0_48[116], stage0_48[117]},
      {stage1_50[17],stage1_49[41],stage1_48[72],stage1_47[125],stage1_46[161]}
   );
   gpc615_5 gpc1776 (
      {stage0_46[326], stage0_46[327], stage0_46[328], stage0_46[329], stage0_46[330]},
      {stage0_47[132]},
      {stage0_48[118], stage0_48[119], stage0_48[120], stage0_48[121], stage0_48[122], stage0_48[123]},
      {stage1_50[18],stage1_49[42],stage1_48[73],stage1_47[126],stage1_46[162]}
   );
   gpc615_5 gpc1777 (
      {stage0_46[331], stage0_46[332], stage0_46[333], stage0_46[334], stage0_46[335]},
      {stage0_47[133]},
      {stage0_48[124], stage0_48[125], stage0_48[126], stage0_48[127], stage0_48[128], stage0_48[129]},
      {stage1_50[19],stage1_49[43],stage1_48[74],stage1_47[127],stage1_46[163]}
   );
   gpc615_5 gpc1778 (
      {stage0_46[336], stage0_46[337], stage0_46[338], stage0_46[339], stage0_46[340]},
      {stage0_47[134]},
      {stage0_48[130], stage0_48[131], stage0_48[132], stage0_48[133], stage0_48[134], stage0_48[135]},
      {stage1_50[20],stage1_49[44],stage1_48[75],stage1_47[128],stage1_46[164]}
   );
   gpc615_5 gpc1779 (
      {stage0_46[341], stage0_46[342], stage0_46[343], stage0_46[344], stage0_46[345]},
      {stage0_47[135]},
      {stage0_48[136], stage0_48[137], stage0_48[138], stage0_48[139], stage0_48[140], stage0_48[141]},
      {stage1_50[21],stage1_49[45],stage1_48[76],stage1_47[129],stage1_46[165]}
   );
   gpc615_5 gpc1780 (
      {stage0_46[346], stage0_46[347], stage0_46[348], stage0_46[349], stage0_46[350]},
      {stage0_47[136]},
      {stage0_48[142], stage0_48[143], stage0_48[144], stage0_48[145], stage0_48[146], stage0_48[147]},
      {stage1_50[22],stage1_49[46],stage1_48[77],stage1_47[130],stage1_46[166]}
   );
   gpc615_5 gpc1781 (
      {stage0_46[351], stage0_46[352], stage0_46[353], stage0_46[354], stage0_46[355]},
      {stage0_47[137]},
      {stage0_48[148], stage0_48[149], stage0_48[150], stage0_48[151], stage0_48[152], stage0_48[153]},
      {stage1_50[23],stage1_49[47],stage1_48[78],stage1_47[131],stage1_46[167]}
   );
   gpc615_5 gpc1782 (
      {stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141], stage0_47[142]},
      {stage0_48[154]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[24],stage1_49[48],stage1_48[79],stage1_47[132]}
   );
   gpc615_5 gpc1783 (
      {stage0_47[143], stage0_47[144], stage0_47[145], stage0_47[146], stage0_47[147]},
      {stage0_48[155]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[25],stage1_49[49],stage1_48[80],stage1_47[133]}
   );
   gpc615_5 gpc1784 (
      {stage0_47[148], stage0_47[149], stage0_47[150], stage0_47[151], stage0_47[152]},
      {stage0_48[156]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[26],stage1_49[50],stage1_48[81],stage1_47[134]}
   );
   gpc615_5 gpc1785 (
      {stage0_47[153], stage0_47[154], stage0_47[155], stage0_47[156], stage0_47[157]},
      {stage0_48[157]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[27],stage1_49[51],stage1_48[82],stage1_47[135]}
   );
   gpc615_5 gpc1786 (
      {stage0_47[158], stage0_47[159], stage0_47[160], stage0_47[161], stage0_47[162]},
      {stage0_48[158]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[28],stage1_49[52],stage1_48[83],stage1_47[136]}
   );
   gpc615_5 gpc1787 (
      {stage0_47[163], stage0_47[164], stage0_47[165], stage0_47[166], stage0_47[167]},
      {stage0_48[159]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[29],stage1_49[53],stage1_48[84],stage1_47[137]}
   );
   gpc615_5 gpc1788 (
      {stage0_47[168], stage0_47[169], stage0_47[170], stage0_47[171], stage0_47[172]},
      {stage0_48[160]},
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage1_51[6],stage1_50[30],stage1_49[54],stage1_48[85],stage1_47[138]}
   );
   gpc615_5 gpc1789 (
      {stage0_47[173], stage0_47[174], stage0_47[175], stage0_47[176], stage0_47[177]},
      {stage0_48[161]},
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage1_51[7],stage1_50[31],stage1_49[55],stage1_48[86],stage1_47[139]}
   );
   gpc615_5 gpc1790 (
      {stage0_47[178], stage0_47[179], stage0_47[180], stage0_47[181], stage0_47[182]},
      {stage0_48[162]},
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage1_51[8],stage1_50[32],stage1_49[56],stage1_48[87],stage1_47[140]}
   );
   gpc615_5 gpc1791 (
      {stage0_47[183], stage0_47[184], stage0_47[185], stage0_47[186], stage0_47[187]},
      {stage0_48[163]},
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage1_51[9],stage1_50[33],stage1_49[57],stage1_48[88],stage1_47[141]}
   );
   gpc615_5 gpc1792 (
      {stage0_47[188], stage0_47[189], stage0_47[190], stage0_47[191], stage0_47[192]},
      {stage0_48[164]},
      {stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64], stage0_49[65]},
      {stage1_51[10],stage1_50[34],stage1_49[58],stage1_48[89],stage1_47[142]}
   );
   gpc615_5 gpc1793 (
      {stage0_47[193], stage0_47[194], stage0_47[195], stage0_47[196], stage0_47[197]},
      {stage0_48[165]},
      {stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70], stage0_49[71]},
      {stage1_51[11],stage1_50[35],stage1_49[59],stage1_48[90],stage1_47[143]}
   );
   gpc615_5 gpc1794 (
      {stage0_47[198], stage0_47[199], stage0_47[200], stage0_47[201], stage0_47[202]},
      {stage0_48[166]},
      {stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76], stage0_49[77]},
      {stage1_51[12],stage1_50[36],stage1_49[60],stage1_48[91],stage1_47[144]}
   );
   gpc615_5 gpc1795 (
      {stage0_47[203], stage0_47[204], stage0_47[205], stage0_47[206], stage0_47[207]},
      {stage0_48[167]},
      {stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82], stage0_49[83]},
      {stage1_51[13],stage1_50[37],stage1_49[61],stage1_48[92],stage1_47[145]}
   );
   gpc615_5 gpc1796 (
      {stage0_47[208], stage0_47[209], stage0_47[210], stage0_47[211], stage0_47[212]},
      {stage0_48[168]},
      {stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88], stage0_49[89]},
      {stage1_51[14],stage1_50[38],stage1_49[62],stage1_48[93],stage1_47[146]}
   );
   gpc615_5 gpc1797 (
      {stage0_47[213], stage0_47[214], stage0_47[215], stage0_47[216], stage0_47[217]},
      {stage0_48[169]},
      {stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94], stage0_49[95]},
      {stage1_51[15],stage1_50[39],stage1_49[63],stage1_48[94],stage1_47[147]}
   );
   gpc615_5 gpc1798 (
      {stage0_47[218], stage0_47[219], stage0_47[220], stage0_47[221], stage0_47[222]},
      {stage0_48[170]},
      {stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100], stage0_49[101]},
      {stage1_51[16],stage1_50[40],stage1_49[64],stage1_48[95],stage1_47[148]}
   );
   gpc615_5 gpc1799 (
      {stage0_47[223], stage0_47[224], stage0_47[225], stage0_47[226], stage0_47[227]},
      {stage0_48[171]},
      {stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106], stage0_49[107]},
      {stage1_51[17],stage1_50[41],stage1_49[65],stage1_48[96],stage1_47[149]}
   );
   gpc615_5 gpc1800 (
      {stage0_47[228], stage0_47[229], stage0_47[230], stage0_47[231], stage0_47[232]},
      {stage0_48[172]},
      {stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112], stage0_49[113]},
      {stage1_51[18],stage1_50[42],stage1_49[66],stage1_48[97],stage1_47[150]}
   );
   gpc615_5 gpc1801 (
      {stage0_47[233], stage0_47[234], stage0_47[235], stage0_47[236], stage0_47[237]},
      {stage0_48[173]},
      {stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118], stage0_49[119]},
      {stage1_51[19],stage1_50[43],stage1_49[67],stage1_48[98],stage1_47[151]}
   );
   gpc615_5 gpc1802 (
      {stage0_47[238], stage0_47[239], stage0_47[240], stage0_47[241], stage0_47[242]},
      {stage0_48[174]},
      {stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124], stage0_49[125]},
      {stage1_51[20],stage1_50[44],stage1_49[68],stage1_48[99],stage1_47[152]}
   );
   gpc615_5 gpc1803 (
      {stage0_47[243], stage0_47[244], stage0_47[245], stage0_47[246], stage0_47[247]},
      {stage0_48[175]},
      {stage0_49[126], stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130], stage0_49[131]},
      {stage1_51[21],stage1_50[45],stage1_49[69],stage1_48[100],stage1_47[153]}
   );
   gpc615_5 gpc1804 (
      {stage0_47[248], stage0_47[249], stage0_47[250], stage0_47[251], stage0_47[252]},
      {stage0_48[176]},
      {stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136], stage0_49[137]},
      {stage1_51[22],stage1_50[46],stage1_49[70],stage1_48[101],stage1_47[154]}
   );
   gpc615_5 gpc1805 (
      {stage0_47[253], stage0_47[254], stage0_47[255], stage0_47[256], stage0_47[257]},
      {stage0_48[177]},
      {stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141], stage0_49[142], stage0_49[143]},
      {stage1_51[23],stage1_50[47],stage1_49[71],stage1_48[102],stage1_47[155]}
   );
   gpc615_5 gpc1806 (
      {stage0_47[258], stage0_47[259], stage0_47[260], stage0_47[261], stage0_47[262]},
      {stage0_48[178]},
      {stage0_49[144], stage0_49[145], stage0_49[146], stage0_49[147], stage0_49[148], stage0_49[149]},
      {stage1_51[24],stage1_50[48],stage1_49[72],stage1_48[103],stage1_47[156]}
   );
   gpc615_5 gpc1807 (
      {stage0_47[263], stage0_47[264], stage0_47[265], stage0_47[266], stage0_47[267]},
      {stage0_48[179]},
      {stage0_49[150], stage0_49[151], stage0_49[152], stage0_49[153], stage0_49[154], stage0_49[155]},
      {stage1_51[25],stage1_50[49],stage1_49[73],stage1_48[104],stage1_47[157]}
   );
   gpc615_5 gpc1808 (
      {stage0_47[268], stage0_47[269], stage0_47[270], stage0_47[271], stage0_47[272]},
      {stage0_48[180]},
      {stage0_49[156], stage0_49[157], stage0_49[158], stage0_49[159], stage0_49[160], stage0_49[161]},
      {stage1_51[26],stage1_50[50],stage1_49[74],stage1_48[105],stage1_47[158]}
   );
   gpc615_5 gpc1809 (
      {stage0_47[273], stage0_47[274], stage0_47[275], stage0_47[276], stage0_47[277]},
      {stage0_48[181]},
      {stage0_49[162], stage0_49[163], stage0_49[164], stage0_49[165], stage0_49[166], stage0_49[167]},
      {stage1_51[27],stage1_50[51],stage1_49[75],stage1_48[106],stage1_47[159]}
   );
   gpc615_5 gpc1810 (
      {stage0_47[278], stage0_47[279], stage0_47[280], stage0_47[281], stage0_47[282]},
      {stage0_48[182]},
      {stage0_49[168], stage0_49[169], stage0_49[170], stage0_49[171], stage0_49[172], stage0_49[173]},
      {stage1_51[28],stage1_50[52],stage1_49[76],stage1_48[107],stage1_47[160]}
   );
   gpc615_5 gpc1811 (
      {stage0_47[283], stage0_47[284], stage0_47[285], stage0_47[286], stage0_47[287]},
      {stage0_48[183]},
      {stage0_49[174], stage0_49[175], stage0_49[176], stage0_49[177], stage0_49[178], stage0_49[179]},
      {stage1_51[29],stage1_50[53],stage1_49[77],stage1_48[108],stage1_47[161]}
   );
   gpc615_5 gpc1812 (
      {stage0_47[288], stage0_47[289], stage0_47[290], stage0_47[291], stage0_47[292]},
      {stage0_48[184]},
      {stage0_49[180], stage0_49[181], stage0_49[182], stage0_49[183], stage0_49[184], stage0_49[185]},
      {stage1_51[30],stage1_50[54],stage1_49[78],stage1_48[109],stage1_47[162]}
   );
   gpc615_5 gpc1813 (
      {stage0_47[293], stage0_47[294], stage0_47[295], stage0_47[296], stage0_47[297]},
      {stage0_48[185]},
      {stage0_49[186], stage0_49[187], stage0_49[188], stage0_49[189], stage0_49[190], stage0_49[191]},
      {stage1_51[31],stage1_50[55],stage1_49[79],stage1_48[110],stage1_47[163]}
   );
   gpc615_5 gpc1814 (
      {stage0_47[298], stage0_47[299], stage0_47[300], stage0_47[301], stage0_47[302]},
      {stage0_48[186]},
      {stage0_49[192], stage0_49[193], stage0_49[194], stage0_49[195], stage0_49[196], stage0_49[197]},
      {stage1_51[32],stage1_50[56],stage1_49[80],stage1_48[111],stage1_47[164]}
   );
   gpc615_5 gpc1815 (
      {stage0_47[303], stage0_47[304], stage0_47[305], stage0_47[306], stage0_47[307]},
      {stage0_48[187]},
      {stage0_49[198], stage0_49[199], stage0_49[200], stage0_49[201], stage0_49[202], stage0_49[203]},
      {stage1_51[33],stage1_50[57],stage1_49[81],stage1_48[112],stage1_47[165]}
   );
   gpc615_5 gpc1816 (
      {stage0_47[308], stage0_47[309], stage0_47[310], stage0_47[311], stage0_47[312]},
      {stage0_48[188]},
      {stage0_49[204], stage0_49[205], stage0_49[206], stage0_49[207], stage0_49[208], stage0_49[209]},
      {stage1_51[34],stage1_50[58],stage1_49[82],stage1_48[113],stage1_47[166]}
   );
   gpc615_5 gpc1817 (
      {stage0_47[313], stage0_47[314], stage0_47[315], stage0_47[316], stage0_47[317]},
      {stage0_48[189]},
      {stage0_49[210], stage0_49[211], stage0_49[212], stage0_49[213], stage0_49[214], stage0_49[215]},
      {stage1_51[35],stage1_50[59],stage1_49[83],stage1_48[114],stage1_47[167]}
   );
   gpc615_5 gpc1818 (
      {stage0_47[318], stage0_47[319], stage0_47[320], stage0_47[321], stage0_47[322]},
      {stage0_48[190]},
      {stage0_49[216], stage0_49[217], stage0_49[218], stage0_49[219], stage0_49[220], stage0_49[221]},
      {stage1_51[36],stage1_50[60],stage1_49[84],stage1_48[115],stage1_47[168]}
   );
   gpc615_5 gpc1819 (
      {stage0_47[323], stage0_47[324], stage0_47[325], stage0_47[326], stage0_47[327]},
      {stage0_48[191]},
      {stage0_49[222], stage0_49[223], stage0_49[224], stage0_49[225], stage0_49[226], stage0_49[227]},
      {stage1_51[37],stage1_50[61],stage1_49[85],stage1_48[116],stage1_47[169]}
   );
   gpc615_5 gpc1820 (
      {stage0_47[328], stage0_47[329], stage0_47[330], stage0_47[331], stage0_47[332]},
      {stage0_48[192]},
      {stage0_49[228], stage0_49[229], stage0_49[230], stage0_49[231], stage0_49[232], stage0_49[233]},
      {stage1_51[38],stage1_50[62],stage1_49[86],stage1_48[117],stage1_47[170]}
   );
   gpc615_5 gpc1821 (
      {stage0_47[333], stage0_47[334], stage0_47[335], stage0_47[336], stage0_47[337]},
      {stage0_48[193]},
      {stage0_49[234], stage0_49[235], stage0_49[236], stage0_49[237], stage0_49[238], stage0_49[239]},
      {stage1_51[39],stage1_50[63],stage1_49[87],stage1_48[118],stage1_47[171]}
   );
   gpc615_5 gpc1822 (
      {stage0_47[338], stage0_47[339], stage0_47[340], stage0_47[341], stage0_47[342]},
      {stage0_48[194]},
      {stage0_49[240], stage0_49[241], stage0_49[242], stage0_49[243], stage0_49[244], stage0_49[245]},
      {stage1_51[40],stage1_50[64],stage1_49[88],stage1_48[119],stage1_47[172]}
   );
   gpc615_5 gpc1823 (
      {stage0_47[343], stage0_47[344], stage0_47[345], stage0_47[346], stage0_47[347]},
      {stage0_48[195]},
      {stage0_49[246], stage0_49[247], stage0_49[248], stage0_49[249], stage0_49[250], stage0_49[251]},
      {stage1_51[41],stage1_50[65],stage1_49[89],stage1_48[120],stage1_47[173]}
   );
   gpc615_5 gpc1824 (
      {stage0_47[348], stage0_47[349], stage0_47[350], stage0_47[351], stage0_47[352]},
      {stage0_48[196]},
      {stage0_49[252], stage0_49[253], stage0_49[254], stage0_49[255], stage0_49[256], stage0_49[257]},
      {stage1_51[42],stage1_50[66],stage1_49[90],stage1_48[121],stage1_47[174]}
   );
   gpc615_5 gpc1825 (
      {stage0_47[353], stage0_47[354], stage0_47[355], stage0_47[356], stage0_47[357]},
      {stage0_48[197]},
      {stage0_49[258], stage0_49[259], stage0_49[260], stage0_49[261], stage0_49[262], stage0_49[263]},
      {stage1_51[43],stage1_50[67],stage1_49[91],stage1_48[122],stage1_47[175]}
   );
   gpc615_5 gpc1826 (
      {stage0_47[358], stage0_47[359], stage0_47[360], stage0_47[361], stage0_47[362]},
      {stage0_48[198]},
      {stage0_49[264], stage0_49[265], stage0_49[266], stage0_49[267], stage0_49[268], stage0_49[269]},
      {stage1_51[44],stage1_50[68],stage1_49[92],stage1_48[123],stage1_47[176]}
   );
   gpc615_5 gpc1827 (
      {stage0_47[363], stage0_47[364], stage0_47[365], stage0_47[366], stage0_47[367]},
      {stage0_48[199]},
      {stage0_49[270], stage0_49[271], stage0_49[272], stage0_49[273], stage0_49[274], stage0_49[275]},
      {stage1_51[45],stage1_50[69],stage1_49[93],stage1_48[124],stage1_47[177]}
   );
   gpc615_5 gpc1828 (
      {stage0_47[368], stage0_47[369], stage0_47[370], stage0_47[371], stage0_47[372]},
      {stage0_48[200]},
      {stage0_49[276], stage0_49[277], stage0_49[278], stage0_49[279], stage0_49[280], stage0_49[281]},
      {stage1_51[46],stage1_50[70],stage1_49[94],stage1_48[125],stage1_47[178]}
   );
   gpc615_5 gpc1829 (
      {stage0_47[373], stage0_47[374], stage0_47[375], stage0_47[376], stage0_47[377]},
      {stage0_48[201]},
      {stage0_49[282], stage0_49[283], stage0_49[284], stage0_49[285], stage0_49[286], stage0_49[287]},
      {stage1_51[47],stage1_50[71],stage1_49[95],stage1_48[126],stage1_47[179]}
   );
   gpc615_5 gpc1830 (
      {stage0_47[378], stage0_47[379], stage0_47[380], stage0_47[381], stage0_47[382]},
      {stage0_48[202]},
      {stage0_49[288], stage0_49[289], stage0_49[290], stage0_49[291], stage0_49[292], stage0_49[293]},
      {stage1_51[48],stage1_50[72],stage1_49[96],stage1_48[127],stage1_47[180]}
   );
   gpc615_5 gpc1831 (
      {stage0_47[383], stage0_47[384], stage0_47[385], stage0_47[386], stage0_47[387]},
      {stage0_48[203]},
      {stage0_49[294], stage0_49[295], stage0_49[296], stage0_49[297], stage0_49[298], stage0_49[299]},
      {stage1_51[49],stage1_50[73],stage1_49[97],stage1_48[128],stage1_47[181]}
   );
   gpc615_5 gpc1832 (
      {stage0_47[388], stage0_47[389], stage0_47[390], stage0_47[391], stage0_47[392]},
      {stage0_48[204]},
      {stage0_49[300], stage0_49[301], stage0_49[302], stage0_49[303], stage0_49[304], stage0_49[305]},
      {stage1_51[50],stage1_50[74],stage1_49[98],stage1_48[129],stage1_47[182]}
   );
   gpc615_5 gpc1833 (
      {stage0_47[393], stage0_47[394], stage0_47[395], stage0_47[396], stage0_47[397]},
      {stage0_48[205]},
      {stage0_49[306], stage0_49[307], stage0_49[308], stage0_49[309], stage0_49[310], stage0_49[311]},
      {stage1_51[51],stage1_50[75],stage1_49[99],stage1_48[130],stage1_47[183]}
   );
   gpc615_5 gpc1834 (
      {stage0_47[398], stage0_47[399], stage0_47[400], stage0_47[401], stage0_47[402]},
      {stage0_48[206]},
      {stage0_49[312], stage0_49[313], stage0_49[314], stage0_49[315], stage0_49[316], stage0_49[317]},
      {stage1_51[52],stage1_50[76],stage1_49[100],stage1_48[131],stage1_47[184]}
   );
   gpc615_5 gpc1835 (
      {stage0_47[403], stage0_47[404], stage0_47[405], stage0_47[406], stage0_47[407]},
      {stage0_48[207]},
      {stage0_49[318], stage0_49[319], stage0_49[320], stage0_49[321], stage0_49[322], stage0_49[323]},
      {stage1_51[53],stage1_50[77],stage1_49[101],stage1_48[132],stage1_47[185]}
   );
   gpc615_5 gpc1836 (
      {stage0_47[408], stage0_47[409], stage0_47[410], stage0_47[411], stage0_47[412]},
      {stage0_48[208]},
      {stage0_49[324], stage0_49[325], stage0_49[326], stage0_49[327], stage0_49[328], stage0_49[329]},
      {stage1_51[54],stage1_50[78],stage1_49[102],stage1_48[133],stage1_47[186]}
   );
   gpc615_5 gpc1837 (
      {stage0_47[413], stage0_47[414], stage0_47[415], stage0_47[416], stage0_47[417]},
      {stage0_48[209]},
      {stage0_49[330], stage0_49[331], stage0_49[332], stage0_49[333], stage0_49[334], stage0_49[335]},
      {stage1_51[55],stage1_50[79],stage1_49[103],stage1_48[134],stage1_47[187]}
   );
   gpc615_5 gpc1838 (
      {stage0_47[418], stage0_47[419], stage0_47[420], stage0_47[421], stage0_47[422]},
      {stage0_48[210]},
      {stage0_49[336], stage0_49[337], stage0_49[338], stage0_49[339], stage0_49[340], stage0_49[341]},
      {stage1_51[56],stage1_50[80],stage1_49[104],stage1_48[135],stage1_47[188]}
   );
   gpc615_5 gpc1839 (
      {stage0_47[423], stage0_47[424], stage0_47[425], stage0_47[426], stage0_47[427]},
      {stage0_48[211]},
      {stage0_49[342], stage0_49[343], stage0_49[344], stage0_49[345], stage0_49[346], stage0_49[347]},
      {stage1_51[57],stage1_50[81],stage1_49[105],stage1_48[136],stage1_47[189]}
   );
   gpc615_5 gpc1840 (
      {stage0_47[428], stage0_47[429], stage0_47[430], stage0_47[431], stage0_47[432]},
      {stage0_48[212]},
      {stage0_49[348], stage0_49[349], stage0_49[350], stage0_49[351], stage0_49[352], stage0_49[353]},
      {stage1_51[58],stage1_50[82],stage1_49[106],stage1_48[137],stage1_47[190]}
   );
   gpc615_5 gpc1841 (
      {stage0_47[433], stage0_47[434], stage0_47[435], stage0_47[436], stage0_47[437]},
      {stage0_48[213]},
      {stage0_49[354], stage0_49[355], stage0_49[356], stage0_49[357], stage0_49[358], stage0_49[359]},
      {stage1_51[59],stage1_50[83],stage1_49[107],stage1_48[138],stage1_47[191]}
   );
   gpc615_5 gpc1842 (
      {stage0_47[438], stage0_47[439], stage0_47[440], stage0_47[441], stage0_47[442]},
      {stage0_48[214]},
      {stage0_49[360], stage0_49[361], stage0_49[362], stage0_49[363], stage0_49[364], stage0_49[365]},
      {stage1_51[60],stage1_50[84],stage1_49[108],stage1_48[139],stage1_47[192]}
   );
   gpc606_5 gpc1843 (
      {stage0_48[215], stage0_48[216], stage0_48[217], stage0_48[218], stage0_48[219], stage0_48[220]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[61],stage1_50[85],stage1_49[109],stage1_48[140]}
   );
   gpc606_5 gpc1844 (
      {stage0_48[221], stage0_48[222], stage0_48[223], stage0_48[224], stage0_48[225], stage0_48[226]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[62],stage1_50[86],stage1_49[110],stage1_48[141]}
   );
   gpc606_5 gpc1845 (
      {stage0_48[227], stage0_48[228], stage0_48[229], stage0_48[230], stage0_48[231], stage0_48[232]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[63],stage1_50[87],stage1_49[111],stage1_48[142]}
   );
   gpc606_5 gpc1846 (
      {stage0_48[233], stage0_48[234], stage0_48[235], stage0_48[236], stage0_48[237], stage0_48[238]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[64],stage1_50[88],stage1_49[112],stage1_48[143]}
   );
   gpc606_5 gpc1847 (
      {stage0_48[239], stage0_48[240], stage0_48[241], stage0_48[242], stage0_48[243], stage0_48[244]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[65],stage1_50[89],stage1_49[113],stage1_48[144]}
   );
   gpc606_5 gpc1848 (
      {stage0_48[245], stage0_48[246], stage0_48[247], stage0_48[248], stage0_48[249], stage0_48[250]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[66],stage1_50[90],stage1_49[114],stage1_48[145]}
   );
   gpc606_5 gpc1849 (
      {stage0_48[251], stage0_48[252], stage0_48[253], stage0_48[254], stage0_48[255], stage0_48[256]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[67],stage1_50[91],stage1_49[115],stage1_48[146]}
   );
   gpc606_5 gpc1850 (
      {stage0_48[257], stage0_48[258], stage0_48[259], stage0_48[260], stage0_48[261], stage0_48[262]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[68],stage1_50[92],stage1_49[116],stage1_48[147]}
   );
   gpc606_5 gpc1851 (
      {stage0_48[263], stage0_48[264], stage0_48[265], stage0_48[266], stage0_48[267], stage0_48[268]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[69],stage1_50[93],stage1_49[117],stage1_48[148]}
   );
   gpc606_5 gpc1852 (
      {stage0_48[269], stage0_48[270], stage0_48[271], stage0_48[272], stage0_48[273], stage0_48[274]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[70],stage1_50[94],stage1_49[118],stage1_48[149]}
   );
   gpc606_5 gpc1853 (
      {stage0_48[275], stage0_48[276], stage0_48[277], stage0_48[278], stage0_48[279], stage0_48[280]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[71],stage1_50[95],stage1_49[119],stage1_48[150]}
   );
   gpc606_5 gpc1854 (
      {stage0_48[281], stage0_48[282], stage0_48[283], stage0_48[284], stage0_48[285], stage0_48[286]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[72],stage1_50[96],stage1_49[120],stage1_48[151]}
   );
   gpc606_5 gpc1855 (
      {stage0_48[287], stage0_48[288], stage0_48[289], stage0_48[290], stage0_48[291], stage0_48[292]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[73],stage1_50[97],stage1_49[121],stage1_48[152]}
   );
   gpc615_5 gpc1856 (
      {stage0_48[293], stage0_48[294], stage0_48[295], stage0_48[296], stage0_48[297]},
      {stage0_49[366]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[74],stage1_50[98],stage1_49[122],stage1_48[153]}
   );
   gpc615_5 gpc1857 (
      {stage0_48[298], stage0_48[299], stage0_48[300], stage0_48[301], stage0_48[302]},
      {stage0_49[367]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[75],stage1_50[99],stage1_49[123],stage1_48[154]}
   );
   gpc615_5 gpc1858 (
      {stage0_48[303], stage0_48[304], stage0_48[305], stage0_48[306], stage0_48[307]},
      {stage0_49[368]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[76],stage1_50[100],stage1_49[124],stage1_48[155]}
   );
   gpc615_5 gpc1859 (
      {stage0_48[308], stage0_48[309], stage0_48[310], stage0_48[311], stage0_48[312]},
      {stage0_49[369]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[77],stage1_50[101],stage1_49[125],stage1_48[156]}
   );
   gpc615_5 gpc1860 (
      {stage0_48[313], stage0_48[314], stage0_48[315], stage0_48[316], stage0_48[317]},
      {stage0_49[370]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[78],stage1_50[102],stage1_49[126],stage1_48[157]}
   );
   gpc615_5 gpc1861 (
      {stage0_48[318], stage0_48[319], stage0_48[320], stage0_48[321], stage0_48[322]},
      {stage0_49[371]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[79],stage1_50[103],stage1_49[127],stage1_48[158]}
   );
   gpc615_5 gpc1862 (
      {stage0_48[323], stage0_48[324], stage0_48[325], stage0_48[326], stage0_48[327]},
      {stage0_49[372]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[80],stage1_50[104],stage1_49[128],stage1_48[159]}
   );
   gpc615_5 gpc1863 (
      {stage0_48[328], stage0_48[329], stage0_48[330], stage0_48[331], stage0_48[332]},
      {stage0_49[373]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[81],stage1_50[105],stage1_49[129],stage1_48[160]}
   );
   gpc615_5 gpc1864 (
      {stage0_48[333], stage0_48[334], stage0_48[335], stage0_48[336], stage0_48[337]},
      {stage0_49[374]},
      {stage0_50[126], stage0_50[127], stage0_50[128], stage0_50[129], stage0_50[130], stage0_50[131]},
      {stage1_52[21],stage1_51[82],stage1_50[106],stage1_49[130],stage1_48[161]}
   );
   gpc615_5 gpc1865 (
      {stage0_48[338], stage0_48[339], stage0_48[340], stage0_48[341], stage0_48[342]},
      {stage0_49[375]},
      {stage0_50[132], stage0_50[133], stage0_50[134], stage0_50[135], stage0_50[136], stage0_50[137]},
      {stage1_52[22],stage1_51[83],stage1_50[107],stage1_49[131],stage1_48[162]}
   );
   gpc615_5 gpc1866 (
      {stage0_48[343], stage0_48[344], stage0_48[345], stage0_48[346], stage0_48[347]},
      {stage0_49[376]},
      {stage0_50[138], stage0_50[139], stage0_50[140], stage0_50[141], stage0_50[142], stage0_50[143]},
      {stage1_52[23],stage1_51[84],stage1_50[108],stage1_49[132],stage1_48[163]}
   );
   gpc615_5 gpc1867 (
      {stage0_48[348], stage0_48[349], stage0_48[350], stage0_48[351], stage0_48[352]},
      {stage0_49[377]},
      {stage0_50[144], stage0_50[145], stage0_50[146], stage0_50[147], stage0_50[148], stage0_50[149]},
      {stage1_52[24],stage1_51[85],stage1_50[109],stage1_49[133],stage1_48[164]}
   );
   gpc615_5 gpc1868 (
      {stage0_48[353], stage0_48[354], stage0_48[355], stage0_48[356], stage0_48[357]},
      {stage0_49[378]},
      {stage0_50[150], stage0_50[151], stage0_50[152], stage0_50[153], stage0_50[154], stage0_50[155]},
      {stage1_52[25],stage1_51[86],stage1_50[110],stage1_49[134],stage1_48[165]}
   );
   gpc615_5 gpc1869 (
      {stage0_48[358], stage0_48[359], stage0_48[360], stage0_48[361], stage0_48[362]},
      {stage0_49[379]},
      {stage0_50[156], stage0_50[157], stage0_50[158], stage0_50[159], stage0_50[160], stage0_50[161]},
      {stage1_52[26],stage1_51[87],stage1_50[111],stage1_49[135],stage1_48[166]}
   );
   gpc615_5 gpc1870 (
      {stage0_48[363], stage0_48[364], stage0_48[365], stage0_48[366], stage0_48[367]},
      {stage0_49[380]},
      {stage0_50[162], stage0_50[163], stage0_50[164], stage0_50[165], stage0_50[166], stage0_50[167]},
      {stage1_52[27],stage1_51[88],stage1_50[112],stage1_49[136],stage1_48[167]}
   );
   gpc615_5 gpc1871 (
      {stage0_48[368], stage0_48[369], stage0_48[370], stage0_48[371], stage0_48[372]},
      {stage0_49[381]},
      {stage0_50[168], stage0_50[169], stage0_50[170], stage0_50[171], stage0_50[172], stage0_50[173]},
      {stage1_52[28],stage1_51[89],stage1_50[113],stage1_49[137],stage1_48[168]}
   );
   gpc615_5 gpc1872 (
      {stage0_48[373], stage0_48[374], stage0_48[375], stage0_48[376], stage0_48[377]},
      {stage0_49[382]},
      {stage0_50[174], stage0_50[175], stage0_50[176], stage0_50[177], stage0_50[178], stage0_50[179]},
      {stage1_52[29],stage1_51[90],stage1_50[114],stage1_49[138],stage1_48[169]}
   );
   gpc615_5 gpc1873 (
      {stage0_48[378], stage0_48[379], stage0_48[380], stage0_48[381], stage0_48[382]},
      {stage0_49[383]},
      {stage0_50[180], stage0_50[181], stage0_50[182], stage0_50[183], stage0_50[184], stage0_50[185]},
      {stage1_52[30],stage1_51[91],stage1_50[115],stage1_49[139],stage1_48[170]}
   );
   gpc615_5 gpc1874 (
      {stage0_48[383], stage0_48[384], stage0_48[385], stage0_48[386], stage0_48[387]},
      {stage0_49[384]},
      {stage0_50[186], stage0_50[187], stage0_50[188], stage0_50[189], stage0_50[190], stage0_50[191]},
      {stage1_52[31],stage1_51[92],stage1_50[116],stage1_49[140],stage1_48[171]}
   );
   gpc615_5 gpc1875 (
      {stage0_48[388], stage0_48[389], stage0_48[390], stage0_48[391], stage0_48[392]},
      {stage0_49[385]},
      {stage0_50[192], stage0_50[193], stage0_50[194], stage0_50[195], stage0_50[196], stage0_50[197]},
      {stage1_52[32],stage1_51[93],stage1_50[117],stage1_49[141],stage1_48[172]}
   );
   gpc615_5 gpc1876 (
      {stage0_48[393], stage0_48[394], stage0_48[395], stage0_48[396], stage0_48[397]},
      {stage0_49[386]},
      {stage0_50[198], stage0_50[199], stage0_50[200], stage0_50[201], stage0_50[202], stage0_50[203]},
      {stage1_52[33],stage1_51[94],stage1_50[118],stage1_49[142],stage1_48[173]}
   );
   gpc615_5 gpc1877 (
      {stage0_48[398], stage0_48[399], stage0_48[400], stage0_48[401], stage0_48[402]},
      {stage0_49[387]},
      {stage0_50[204], stage0_50[205], stage0_50[206], stage0_50[207], stage0_50[208], stage0_50[209]},
      {stage1_52[34],stage1_51[95],stage1_50[119],stage1_49[143],stage1_48[174]}
   );
   gpc615_5 gpc1878 (
      {stage0_48[403], stage0_48[404], stage0_48[405], stage0_48[406], stage0_48[407]},
      {stage0_49[388]},
      {stage0_50[210], stage0_50[211], stage0_50[212], stage0_50[213], stage0_50[214], stage0_50[215]},
      {stage1_52[35],stage1_51[96],stage1_50[120],stage1_49[144],stage1_48[175]}
   );
   gpc615_5 gpc1879 (
      {stage0_48[408], stage0_48[409], stage0_48[410], stage0_48[411], stage0_48[412]},
      {stage0_49[389]},
      {stage0_50[216], stage0_50[217], stage0_50[218], stage0_50[219], stage0_50[220], stage0_50[221]},
      {stage1_52[36],stage1_51[97],stage1_50[121],stage1_49[145],stage1_48[176]}
   );
   gpc615_5 gpc1880 (
      {stage0_48[413], stage0_48[414], stage0_48[415], stage0_48[416], stage0_48[417]},
      {stage0_49[390]},
      {stage0_50[222], stage0_50[223], stage0_50[224], stage0_50[225], stage0_50[226], stage0_50[227]},
      {stage1_52[37],stage1_51[98],stage1_50[122],stage1_49[146],stage1_48[177]}
   );
   gpc615_5 gpc1881 (
      {stage0_48[418], stage0_48[419], stage0_48[420], stage0_48[421], stage0_48[422]},
      {stage0_49[391]},
      {stage0_50[228], stage0_50[229], stage0_50[230], stage0_50[231], stage0_50[232], stage0_50[233]},
      {stage1_52[38],stage1_51[99],stage1_50[123],stage1_49[147],stage1_48[178]}
   );
   gpc615_5 gpc1882 (
      {stage0_48[423], stage0_48[424], stage0_48[425], stage0_48[426], stage0_48[427]},
      {stage0_49[392]},
      {stage0_50[234], stage0_50[235], stage0_50[236], stage0_50[237], stage0_50[238], stage0_50[239]},
      {stage1_52[39],stage1_51[100],stage1_50[124],stage1_49[148],stage1_48[179]}
   );
   gpc615_5 gpc1883 (
      {stage0_48[428], stage0_48[429], stage0_48[430], stage0_48[431], stage0_48[432]},
      {stage0_49[393]},
      {stage0_50[240], stage0_50[241], stage0_50[242], stage0_50[243], stage0_50[244], stage0_50[245]},
      {stage1_52[40],stage1_51[101],stage1_50[125],stage1_49[149],stage1_48[180]}
   );
   gpc615_5 gpc1884 (
      {stage0_48[433], stage0_48[434], stage0_48[435], stage0_48[436], stage0_48[437]},
      {stage0_49[394]},
      {stage0_50[246], stage0_50[247], stage0_50[248], stage0_50[249], stage0_50[250], stage0_50[251]},
      {stage1_52[41],stage1_51[102],stage1_50[126],stage1_49[150],stage1_48[181]}
   );
   gpc615_5 gpc1885 (
      {stage0_48[438], stage0_48[439], stage0_48[440], stage0_48[441], stage0_48[442]},
      {stage0_49[395]},
      {stage0_50[252], stage0_50[253], stage0_50[254], stage0_50[255], stage0_50[256], stage0_50[257]},
      {stage1_52[42],stage1_51[103],stage1_50[127],stage1_49[151],stage1_48[182]}
   );
   gpc615_5 gpc1886 (
      {stage0_48[443], stage0_48[444], stage0_48[445], stage0_48[446], stage0_48[447]},
      {stage0_49[396]},
      {stage0_50[258], stage0_50[259], stage0_50[260], stage0_50[261], stage0_50[262], stage0_50[263]},
      {stage1_52[43],stage1_51[104],stage1_50[128],stage1_49[152],stage1_48[183]}
   );
   gpc615_5 gpc1887 (
      {stage0_48[448], stage0_48[449], stage0_48[450], stage0_48[451], stage0_48[452]},
      {stage0_49[397]},
      {stage0_50[264], stage0_50[265], stage0_50[266], stage0_50[267], stage0_50[268], stage0_50[269]},
      {stage1_52[44],stage1_51[105],stage1_50[129],stage1_49[153],stage1_48[184]}
   );
   gpc615_5 gpc1888 (
      {stage0_48[453], stage0_48[454], stage0_48[455], stage0_48[456], stage0_48[457]},
      {stage0_49[398]},
      {stage0_50[270], stage0_50[271], stage0_50[272], stage0_50[273], stage0_50[274], stage0_50[275]},
      {stage1_52[45],stage1_51[106],stage1_50[130],stage1_49[154],stage1_48[185]}
   );
   gpc615_5 gpc1889 (
      {stage0_48[458], stage0_48[459], stage0_48[460], stage0_48[461], stage0_48[462]},
      {stage0_49[399]},
      {stage0_50[276], stage0_50[277], stage0_50[278], stage0_50[279], stage0_50[280], stage0_50[281]},
      {stage1_52[46],stage1_51[107],stage1_50[131],stage1_49[155],stage1_48[186]}
   );
   gpc615_5 gpc1890 (
      {stage0_48[463], stage0_48[464], stage0_48[465], stage0_48[466], stage0_48[467]},
      {stage0_49[400]},
      {stage0_50[282], stage0_50[283], stage0_50[284], stage0_50[285], stage0_50[286], stage0_50[287]},
      {stage1_52[47],stage1_51[108],stage1_50[132],stage1_49[156],stage1_48[187]}
   );
   gpc615_5 gpc1891 (
      {stage0_48[468], stage0_48[469], stage0_48[470], stage0_48[471], stage0_48[472]},
      {stage0_49[401]},
      {stage0_50[288], stage0_50[289], stage0_50[290], stage0_50[291], stage0_50[292], stage0_50[293]},
      {stage1_52[48],stage1_51[109],stage1_50[133],stage1_49[157],stage1_48[188]}
   );
   gpc615_5 gpc1892 (
      {stage0_48[473], stage0_48[474], stage0_48[475], stage0_48[476], stage0_48[477]},
      {stage0_49[402]},
      {stage0_50[294], stage0_50[295], stage0_50[296], stage0_50[297], stage0_50[298], stage0_50[299]},
      {stage1_52[49],stage1_51[110],stage1_50[134],stage1_49[158],stage1_48[189]}
   );
   gpc606_5 gpc1893 (
      {stage0_49[403], stage0_49[404], stage0_49[405], stage0_49[406], stage0_49[407], stage0_49[408]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[50],stage1_51[111],stage1_50[135],stage1_49[159]}
   );
   gpc606_5 gpc1894 (
      {stage0_49[409], stage0_49[410], stage0_49[411], stage0_49[412], stage0_49[413], stage0_49[414]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[51],stage1_51[112],stage1_50[136],stage1_49[160]}
   );
   gpc606_5 gpc1895 (
      {stage0_49[415], stage0_49[416], stage0_49[417], stage0_49[418], stage0_49[419], stage0_49[420]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[52],stage1_51[113],stage1_50[137],stage1_49[161]}
   );
   gpc606_5 gpc1896 (
      {stage0_49[421], stage0_49[422], stage0_49[423], stage0_49[424], stage0_49[425], stage0_49[426]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[53],stage1_51[114],stage1_50[138],stage1_49[162]}
   );
   gpc606_5 gpc1897 (
      {stage0_49[427], stage0_49[428], stage0_49[429], stage0_49[430], stage0_49[431], stage0_49[432]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[54],stage1_51[115],stage1_50[139],stage1_49[163]}
   );
   gpc606_5 gpc1898 (
      {stage0_49[433], stage0_49[434], stage0_49[435], stage0_49[436], stage0_49[437], stage0_49[438]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[55],stage1_51[116],stage1_50[140],stage1_49[164]}
   );
   gpc606_5 gpc1899 (
      {stage0_49[439], stage0_49[440], stage0_49[441], stage0_49[442], stage0_49[443], stage0_49[444]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[56],stage1_51[117],stage1_50[141],stage1_49[165]}
   );
   gpc606_5 gpc1900 (
      {stage0_49[445], stage0_49[446], stage0_49[447], stage0_49[448], stage0_49[449], stage0_49[450]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[57],stage1_51[118],stage1_50[142],stage1_49[166]}
   );
   gpc606_5 gpc1901 (
      {stage0_49[451], stage0_49[452], stage0_49[453], stage0_49[454], stage0_49[455], stage0_49[456]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[58],stage1_51[119],stage1_50[143],stage1_49[167]}
   );
   gpc606_5 gpc1902 (
      {stage0_49[457], stage0_49[458], stage0_49[459], stage0_49[460], stage0_49[461], stage0_49[462]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[59],stage1_51[120],stage1_50[144],stage1_49[168]}
   );
   gpc606_5 gpc1903 (
      {stage0_49[463], stage0_49[464], stage0_49[465], stage0_49[466], stage0_49[467], stage0_49[468]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[60],stage1_51[121],stage1_50[145],stage1_49[169]}
   );
   gpc606_5 gpc1904 (
      {stage0_49[469], stage0_49[470], stage0_49[471], stage0_49[472], stage0_49[473], stage0_49[474]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[61],stage1_51[122],stage1_50[146],stage1_49[170]}
   );
   gpc606_5 gpc1905 (
      {stage0_49[475], stage0_49[476], stage0_49[477], stage0_49[478], stage0_49[479], stage0_49[480]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[62],stage1_51[123],stage1_50[147],stage1_49[171]}
   );
   gpc615_5 gpc1906 (
      {stage0_49[481], stage0_49[482], stage0_49[483], stage0_49[484], stage0_49[485]},
      {stage0_50[300]},
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage1_53[13],stage1_52[63],stage1_51[124],stage1_50[148],stage1_49[172]}
   );
   gpc615_5 gpc1907 (
      {stage0_50[301], stage0_50[302], stage0_50[303], stage0_50[304], stage0_50[305]},
      {stage0_51[84]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[14],stage1_52[64],stage1_51[125],stage1_50[149]}
   );
   gpc615_5 gpc1908 (
      {stage0_50[306], stage0_50[307], stage0_50[308], stage0_50[309], stage0_50[310]},
      {stage0_51[85]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[15],stage1_52[65],stage1_51[126],stage1_50[150]}
   );
   gpc615_5 gpc1909 (
      {stage0_50[311], stage0_50[312], stage0_50[313], stage0_50[314], stage0_50[315]},
      {stage0_51[86]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[16],stage1_52[66],stage1_51[127],stage1_50[151]}
   );
   gpc615_5 gpc1910 (
      {stage0_50[316], stage0_50[317], stage0_50[318], stage0_50[319], stage0_50[320]},
      {stage0_51[87]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[17],stage1_52[67],stage1_51[128],stage1_50[152]}
   );
   gpc615_5 gpc1911 (
      {stage0_50[321], stage0_50[322], stage0_50[323], stage0_50[324], stage0_50[325]},
      {stage0_51[88]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[18],stage1_52[68],stage1_51[129],stage1_50[153]}
   );
   gpc615_5 gpc1912 (
      {stage0_50[326], stage0_50[327], stage0_50[328], stage0_50[329], stage0_50[330]},
      {stage0_51[89]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[19],stage1_52[69],stage1_51[130],stage1_50[154]}
   );
   gpc615_5 gpc1913 (
      {stage0_50[331], stage0_50[332], stage0_50[333], stage0_50[334], stage0_50[335]},
      {stage0_51[90]},
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage1_54[6],stage1_53[20],stage1_52[70],stage1_51[131],stage1_50[155]}
   );
   gpc615_5 gpc1914 (
      {stage0_50[336], stage0_50[337], stage0_50[338], stage0_50[339], stage0_50[340]},
      {stage0_51[91]},
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage1_54[7],stage1_53[21],stage1_52[71],stage1_51[132],stage1_50[156]}
   );
   gpc615_5 gpc1915 (
      {stage0_50[341], stage0_50[342], stage0_50[343], stage0_50[344], stage0_50[345]},
      {stage0_51[92]},
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage1_54[8],stage1_53[22],stage1_52[72],stage1_51[133],stage1_50[157]}
   );
   gpc615_5 gpc1916 (
      {stage0_50[346], stage0_50[347], stage0_50[348], stage0_50[349], stage0_50[350]},
      {stage0_51[93]},
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage1_54[9],stage1_53[23],stage1_52[73],stage1_51[134],stage1_50[158]}
   );
   gpc615_5 gpc1917 (
      {stage0_50[351], stage0_50[352], stage0_50[353], stage0_50[354], stage0_50[355]},
      {stage0_51[94]},
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage1_54[10],stage1_53[24],stage1_52[74],stage1_51[135],stage1_50[159]}
   );
   gpc615_5 gpc1918 (
      {stage0_50[356], stage0_50[357], stage0_50[358], stage0_50[359], stage0_50[360]},
      {stage0_51[95]},
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage1_54[11],stage1_53[25],stage1_52[75],stage1_51[136],stage1_50[160]}
   );
   gpc615_5 gpc1919 (
      {stage0_50[361], stage0_50[362], stage0_50[363], stage0_50[364], stage0_50[365]},
      {stage0_51[96]},
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage1_54[12],stage1_53[26],stage1_52[76],stage1_51[137],stage1_50[161]}
   );
   gpc615_5 gpc1920 (
      {stage0_50[366], stage0_50[367], stage0_50[368], stage0_50[369], stage0_50[370]},
      {stage0_51[97]},
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage1_54[13],stage1_53[27],stage1_52[77],stage1_51[138],stage1_50[162]}
   );
   gpc615_5 gpc1921 (
      {stage0_50[371], stage0_50[372], stage0_50[373], stage0_50[374], stage0_50[375]},
      {stage0_51[98]},
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage1_54[14],stage1_53[28],stage1_52[78],stage1_51[139],stage1_50[163]}
   );
   gpc615_5 gpc1922 (
      {stage0_50[376], stage0_50[377], stage0_50[378], stage0_50[379], stage0_50[380]},
      {stage0_51[99]},
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage1_54[15],stage1_53[29],stage1_52[79],stage1_51[140],stage1_50[164]}
   );
   gpc615_5 gpc1923 (
      {stage0_50[381], stage0_50[382], stage0_50[383], stage0_50[384], stage0_50[385]},
      {stage0_51[100]},
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage1_54[16],stage1_53[30],stage1_52[80],stage1_51[141],stage1_50[165]}
   );
   gpc615_5 gpc1924 (
      {stage0_50[386], stage0_50[387], stage0_50[388], stage0_50[389], stage0_50[390]},
      {stage0_51[101]},
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage1_54[17],stage1_53[31],stage1_52[81],stage1_51[142],stage1_50[166]}
   );
   gpc615_5 gpc1925 (
      {stage0_50[391], stage0_50[392], stage0_50[393], stage0_50[394], stage0_50[395]},
      {stage0_51[102]},
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage1_54[18],stage1_53[32],stage1_52[82],stage1_51[143],stage1_50[167]}
   );
   gpc615_5 gpc1926 (
      {stage0_50[396], stage0_50[397], stage0_50[398], stage0_50[399], stage0_50[400]},
      {stage0_51[103]},
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage1_54[19],stage1_53[33],stage1_52[83],stage1_51[144],stage1_50[168]}
   );
   gpc615_5 gpc1927 (
      {stage0_50[401], stage0_50[402], stage0_50[403], stage0_50[404], stage0_50[405]},
      {stage0_51[104]},
      {stage0_52[120], stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125]},
      {stage1_54[20],stage1_53[34],stage1_52[84],stage1_51[145],stage1_50[169]}
   );
   gpc615_5 gpc1928 (
      {stage0_50[406], stage0_50[407], stage0_50[408], stage0_50[409], stage0_50[410]},
      {stage0_51[105]},
      {stage0_52[126], stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131]},
      {stage1_54[21],stage1_53[35],stage1_52[85],stage1_51[146],stage1_50[170]}
   );
   gpc615_5 gpc1929 (
      {stage0_50[411], stage0_50[412], stage0_50[413], stage0_50[414], stage0_50[415]},
      {stage0_51[106]},
      {stage0_52[132], stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137]},
      {stage1_54[22],stage1_53[36],stage1_52[86],stage1_51[147],stage1_50[171]}
   );
   gpc615_5 gpc1930 (
      {stage0_50[416], stage0_50[417], stage0_50[418], stage0_50[419], stage0_50[420]},
      {stage0_51[107]},
      {stage0_52[138], stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142], stage0_52[143]},
      {stage1_54[23],stage1_53[37],stage1_52[87],stage1_51[148],stage1_50[172]}
   );
   gpc615_5 gpc1931 (
      {stage0_50[421], stage0_50[422], stage0_50[423], stage0_50[424], stage0_50[425]},
      {stage0_51[108]},
      {stage0_52[144], stage0_52[145], stage0_52[146], stage0_52[147], stage0_52[148], stage0_52[149]},
      {stage1_54[24],stage1_53[38],stage1_52[88],stage1_51[149],stage1_50[173]}
   );
   gpc615_5 gpc1932 (
      {stage0_50[426], stage0_50[427], stage0_50[428], stage0_50[429], stage0_50[430]},
      {stage0_51[109]},
      {stage0_52[150], stage0_52[151], stage0_52[152], stage0_52[153], stage0_52[154], stage0_52[155]},
      {stage1_54[25],stage1_53[39],stage1_52[89],stage1_51[150],stage1_50[174]}
   );
   gpc615_5 gpc1933 (
      {stage0_50[431], stage0_50[432], stage0_50[433], stage0_50[434], stage0_50[435]},
      {stage0_51[110]},
      {stage0_52[156], stage0_52[157], stage0_52[158], stage0_52[159], stage0_52[160], stage0_52[161]},
      {stage1_54[26],stage1_53[40],stage1_52[90],stage1_51[151],stage1_50[175]}
   );
   gpc615_5 gpc1934 (
      {stage0_50[436], stage0_50[437], stage0_50[438], stage0_50[439], stage0_50[440]},
      {stage0_51[111]},
      {stage0_52[162], stage0_52[163], stage0_52[164], stage0_52[165], stage0_52[166], stage0_52[167]},
      {stage1_54[27],stage1_53[41],stage1_52[91],stage1_51[152],stage1_50[176]}
   );
   gpc615_5 gpc1935 (
      {stage0_50[441], stage0_50[442], stage0_50[443], stage0_50[444], stage0_50[445]},
      {stage0_51[112]},
      {stage0_52[168], stage0_52[169], stage0_52[170], stage0_52[171], stage0_52[172], stage0_52[173]},
      {stage1_54[28],stage1_53[42],stage1_52[92],stage1_51[153],stage1_50[177]}
   );
   gpc615_5 gpc1936 (
      {stage0_50[446], stage0_50[447], stage0_50[448], stage0_50[449], stage0_50[450]},
      {stage0_51[113]},
      {stage0_52[174], stage0_52[175], stage0_52[176], stage0_52[177], stage0_52[178], stage0_52[179]},
      {stage1_54[29],stage1_53[43],stage1_52[93],stage1_51[154],stage1_50[178]}
   );
   gpc615_5 gpc1937 (
      {stage0_50[451], stage0_50[452], stage0_50[453], stage0_50[454], stage0_50[455]},
      {stage0_51[114]},
      {stage0_52[180], stage0_52[181], stage0_52[182], stage0_52[183], stage0_52[184], stage0_52[185]},
      {stage1_54[30],stage1_53[44],stage1_52[94],stage1_51[155],stage1_50[179]}
   );
   gpc615_5 gpc1938 (
      {stage0_50[456], stage0_50[457], stage0_50[458], stage0_50[459], stage0_50[460]},
      {stage0_51[115]},
      {stage0_52[186], stage0_52[187], stage0_52[188], stage0_52[189], stage0_52[190], stage0_52[191]},
      {stage1_54[31],stage1_53[45],stage1_52[95],stage1_51[156],stage1_50[180]}
   );
   gpc615_5 gpc1939 (
      {stage0_50[461], stage0_50[462], stage0_50[463], stage0_50[464], stage0_50[465]},
      {stage0_51[116]},
      {stage0_52[192], stage0_52[193], stage0_52[194], stage0_52[195], stage0_52[196], stage0_52[197]},
      {stage1_54[32],stage1_53[46],stage1_52[96],stage1_51[157],stage1_50[181]}
   );
   gpc615_5 gpc1940 (
      {stage0_50[466], stage0_50[467], stage0_50[468], stage0_50[469], stage0_50[470]},
      {stage0_51[117]},
      {stage0_52[198], stage0_52[199], stage0_52[200], stage0_52[201], stage0_52[202], stage0_52[203]},
      {stage1_54[33],stage1_53[47],stage1_52[97],stage1_51[158],stage1_50[182]}
   );
   gpc615_5 gpc1941 (
      {stage0_50[471], stage0_50[472], stage0_50[473], stage0_50[474], stage0_50[475]},
      {stage0_51[118]},
      {stage0_52[204], stage0_52[205], stage0_52[206], stage0_52[207], stage0_52[208], stage0_52[209]},
      {stage1_54[34],stage1_53[48],stage1_52[98],stage1_51[159],stage1_50[183]}
   );
   gpc615_5 gpc1942 (
      {stage0_50[476], stage0_50[477], stage0_50[478], stage0_50[479], stage0_50[480]},
      {stage0_51[119]},
      {stage0_52[210], stage0_52[211], stage0_52[212], stage0_52[213], stage0_52[214], stage0_52[215]},
      {stage1_54[35],stage1_53[49],stage1_52[99],stage1_51[160],stage1_50[184]}
   );
   gpc615_5 gpc1943 (
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124]},
      {stage0_52[216]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[36],stage1_53[50],stage1_52[100],stage1_51[161]}
   );
   gpc615_5 gpc1944 (
      {stage0_51[125], stage0_51[126], stage0_51[127], stage0_51[128], stage0_51[129]},
      {stage0_52[217]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[37],stage1_53[51],stage1_52[101],stage1_51[162]}
   );
   gpc615_5 gpc1945 (
      {stage0_51[130], stage0_51[131], stage0_51[132], stage0_51[133], stage0_51[134]},
      {stage0_52[218]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[38],stage1_53[52],stage1_52[102],stage1_51[163]}
   );
   gpc615_5 gpc1946 (
      {stage0_51[135], stage0_51[136], stage0_51[137], stage0_51[138], stage0_51[139]},
      {stage0_52[219]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[39],stage1_53[53],stage1_52[103],stage1_51[164]}
   );
   gpc615_5 gpc1947 (
      {stage0_51[140], stage0_51[141], stage0_51[142], stage0_51[143], stage0_51[144]},
      {stage0_52[220]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[40],stage1_53[54],stage1_52[104],stage1_51[165]}
   );
   gpc615_5 gpc1948 (
      {stage0_51[145], stage0_51[146], stage0_51[147], stage0_51[148], stage0_51[149]},
      {stage0_52[221]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[41],stage1_53[55],stage1_52[105],stage1_51[166]}
   );
   gpc615_5 gpc1949 (
      {stage0_51[150], stage0_51[151], stage0_51[152], stage0_51[153], stage0_51[154]},
      {stage0_52[222]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[42],stage1_53[56],stage1_52[106],stage1_51[167]}
   );
   gpc615_5 gpc1950 (
      {stage0_51[155], stage0_51[156], stage0_51[157], stage0_51[158], stage0_51[159]},
      {stage0_52[223]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[43],stage1_53[57],stage1_52[107],stage1_51[168]}
   );
   gpc615_5 gpc1951 (
      {stage0_51[160], stage0_51[161], stage0_51[162], stage0_51[163], stage0_51[164]},
      {stage0_52[224]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[44],stage1_53[58],stage1_52[108],stage1_51[169]}
   );
   gpc615_5 gpc1952 (
      {stage0_51[165], stage0_51[166], stage0_51[167], stage0_51[168], stage0_51[169]},
      {stage0_52[225]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[45],stage1_53[59],stage1_52[109],stage1_51[170]}
   );
   gpc615_5 gpc1953 (
      {stage0_51[170], stage0_51[171], stage0_51[172], stage0_51[173], stage0_51[174]},
      {stage0_52[226]},
      {stage0_53[60], stage0_53[61], stage0_53[62], stage0_53[63], stage0_53[64], stage0_53[65]},
      {stage1_55[10],stage1_54[46],stage1_53[60],stage1_52[110],stage1_51[171]}
   );
   gpc615_5 gpc1954 (
      {stage0_51[175], stage0_51[176], stage0_51[177], stage0_51[178], stage0_51[179]},
      {stage0_52[227]},
      {stage0_53[66], stage0_53[67], stage0_53[68], stage0_53[69], stage0_53[70], stage0_53[71]},
      {stage1_55[11],stage1_54[47],stage1_53[61],stage1_52[111],stage1_51[172]}
   );
   gpc615_5 gpc1955 (
      {stage0_51[180], stage0_51[181], stage0_51[182], stage0_51[183], stage0_51[184]},
      {stage0_52[228]},
      {stage0_53[72], stage0_53[73], stage0_53[74], stage0_53[75], stage0_53[76], stage0_53[77]},
      {stage1_55[12],stage1_54[48],stage1_53[62],stage1_52[112],stage1_51[173]}
   );
   gpc615_5 gpc1956 (
      {stage0_51[185], stage0_51[186], stage0_51[187], stage0_51[188], stage0_51[189]},
      {stage0_52[229]},
      {stage0_53[78], stage0_53[79], stage0_53[80], stage0_53[81], stage0_53[82], stage0_53[83]},
      {stage1_55[13],stage1_54[49],stage1_53[63],stage1_52[113],stage1_51[174]}
   );
   gpc615_5 gpc1957 (
      {stage0_51[190], stage0_51[191], stage0_51[192], stage0_51[193], stage0_51[194]},
      {stage0_52[230]},
      {stage0_53[84], stage0_53[85], stage0_53[86], stage0_53[87], stage0_53[88], stage0_53[89]},
      {stage1_55[14],stage1_54[50],stage1_53[64],stage1_52[114],stage1_51[175]}
   );
   gpc615_5 gpc1958 (
      {stage0_51[195], stage0_51[196], stage0_51[197], stage0_51[198], stage0_51[199]},
      {stage0_52[231]},
      {stage0_53[90], stage0_53[91], stage0_53[92], stage0_53[93], stage0_53[94], stage0_53[95]},
      {stage1_55[15],stage1_54[51],stage1_53[65],stage1_52[115],stage1_51[176]}
   );
   gpc615_5 gpc1959 (
      {stage0_51[200], stage0_51[201], stage0_51[202], stage0_51[203], stage0_51[204]},
      {stage0_52[232]},
      {stage0_53[96], stage0_53[97], stage0_53[98], stage0_53[99], stage0_53[100], stage0_53[101]},
      {stage1_55[16],stage1_54[52],stage1_53[66],stage1_52[116],stage1_51[177]}
   );
   gpc615_5 gpc1960 (
      {stage0_51[205], stage0_51[206], stage0_51[207], stage0_51[208], stage0_51[209]},
      {stage0_52[233]},
      {stage0_53[102], stage0_53[103], stage0_53[104], stage0_53[105], stage0_53[106], stage0_53[107]},
      {stage1_55[17],stage1_54[53],stage1_53[67],stage1_52[117],stage1_51[178]}
   );
   gpc615_5 gpc1961 (
      {stage0_51[210], stage0_51[211], stage0_51[212], stage0_51[213], stage0_51[214]},
      {stage0_52[234]},
      {stage0_53[108], stage0_53[109], stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113]},
      {stage1_55[18],stage1_54[54],stage1_53[68],stage1_52[118],stage1_51[179]}
   );
   gpc615_5 gpc1962 (
      {stage0_51[215], stage0_51[216], stage0_51[217], stage0_51[218], stage0_51[219]},
      {stage0_52[235]},
      {stage0_53[114], stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage1_55[19],stage1_54[55],stage1_53[69],stage1_52[119],stage1_51[180]}
   );
   gpc615_5 gpc1963 (
      {stage0_51[220], stage0_51[221], stage0_51[222], stage0_51[223], stage0_51[224]},
      {stage0_52[236]},
      {stage0_53[120], stage0_53[121], stage0_53[122], stage0_53[123], stage0_53[124], stage0_53[125]},
      {stage1_55[20],stage1_54[56],stage1_53[70],stage1_52[120],stage1_51[181]}
   );
   gpc615_5 gpc1964 (
      {stage0_51[225], stage0_51[226], stage0_51[227], stage0_51[228], stage0_51[229]},
      {stage0_52[237]},
      {stage0_53[126], stage0_53[127], stage0_53[128], stage0_53[129], stage0_53[130], stage0_53[131]},
      {stage1_55[21],stage1_54[57],stage1_53[71],stage1_52[121],stage1_51[182]}
   );
   gpc615_5 gpc1965 (
      {stage0_51[230], stage0_51[231], stage0_51[232], stage0_51[233], stage0_51[234]},
      {stage0_52[238]},
      {stage0_53[132], stage0_53[133], stage0_53[134], stage0_53[135], stage0_53[136], stage0_53[137]},
      {stage1_55[22],stage1_54[58],stage1_53[72],stage1_52[122],stage1_51[183]}
   );
   gpc615_5 gpc1966 (
      {stage0_51[235], stage0_51[236], stage0_51[237], stage0_51[238], stage0_51[239]},
      {stage0_52[239]},
      {stage0_53[138], stage0_53[139], stage0_53[140], stage0_53[141], stage0_53[142], stage0_53[143]},
      {stage1_55[23],stage1_54[59],stage1_53[73],stage1_52[123],stage1_51[184]}
   );
   gpc615_5 gpc1967 (
      {stage0_51[240], stage0_51[241], stage0_51[242], stage0_51[243], stage0_51[244]},
      {stage0_52[240]},
      {stage0_53[144], stage0_53[145], stage0_53[146], stage0_53[147], stage0_53[148], stage0_53[149]},
      {stage1_55[24],stage1_54[60],stage1_53[74],stage1_52[124],stage1_51[185]}
   );
   gpc615_5 gpc1968 (
      {stage0_51[245], stage0_51[246], stage0_51[247], stage0_51[248], stage0_51[249]},
      {stage0_52[241]},
      {stage0_53[150], stage0_53[151], stage0_53[152], stage0_53[153], stage0_53[154], stage0_53[155]},
      {stage1_55[25],stage1_54[61],stage1_53[75],stage1_52[125],stage1_51[186]}
   );
   gpc615_5 gpc1969 (
      {stage0_51[250], stage0_51[251], stage0_51[252], stage0_51[253], stage0_51[254]},
      {stage0_52[242]},
      {stage0_53[156], stage0_53[157], stage0_53[158], stage0_53[159], stage0_53[160], stage0_53[161]},
      {stage1_55[26],stage1_54[62],stage1_53[76],stage1_52[126],stage1_51[187]}
   );
   gpc615_5 gpc1970 (
      {stage0_51[255], stage0_51[256], stage0_51[257], stage0_51[258], stage0_51[259]},
      {stage0_52[243]},
      {stage0_53[162], stage0_53[163], stage0_53[164], stage0_53[165], stage0_53[166], stage0_53[167]},
      {stage1_55[27],stage1_54[63],stage1_53[77],stage1_52[127],stage1_51[188]}
   );
   gpc615_5 gpc1971 (
      {stage0_51[260], stage0_51[261], stage0_51[262], stage0_51[263], stage0_51[264]},
      {stage0_52[244]},
      {stage0_53[168], stage0_53[169], stage0_53[170], stage0_53[171], stage0_53[172], stage0_53[173]},
      {stage1_55[28],stage1_54[64],stage1_53[78],stage1_52[128],stage1_51[189]}
   );
   gpc615_5 gpc1972 (
      {stage0_51[265], stage0_51[266], stage0_51[267], stage0_51[268], stage0_51[269]},
      {stage0_52[245]},
      {stage0_53[174], stage0_53[175], stage0_53[176], stage0_53[177], stage0_53[178], stage0_53[179]},
      {stage1_55[29],stage1_54[65],stage1_53[79],stage1_52[129],stage1_51[190]}
   );
   gpc615_5 gpc1973 (
      {stage0_51[270], stage0_51[271], stage0_51[272], stage0_51[273], stage0_51[274]},
      {stage0_52[246]},
      {stage0_53[180], stage0_53[181], stage0_53[182], stage0_53[183], stage0_53[184], stage0_53[185]},
      {stage1_55[30],stage1_54[66],stage1_53[80],stage1_52[130],stage1_51[191]}
   );
   gpc615_5 gpc1974 (
      {stage0_51[275], stage0_51[276], stage0_51[277], stage0_51[278], stage0_51[279]},
      {stage0_52[247]},
      {stage0_53[186], stage0_53[187], stage0_53[188], stage0_53[189], stage0_53[190], stage0_53[191]},
      {stage1_55[31],stage1_54[67],stage1_53[81],stage1_52[131],stage1_51[192]}
   );
   gpc615_5 gpc1975 (
      {stage0_51[280], stage0_51[281], stage0_51[282], stage0_51[283], stage0_51[284]},
      {stage0_52[248]},
      {stage0_53[192], stage0_53[193], stage0_53[194], stage0_53[195], stage0_53[196], stage0_53[197]},
      {stage1_55[32],stage1_54[68],stage1_53[82],stage1_52[132],stage1_51[193]}
   );
   gpc615_5 gpc1976 (
      {stage0_51[285], stage0_51[286], stage0_51[287], stage0_51[288], stage0_51[289]},
      {stage0_52[249]},
      {stage0_53[198], stage0_53[199], stage0_53[200], stage0_53[201], stage0_53[202], stage0_53[203]},
      {stage1_55[33],stage1_54[69],stage1_53[83],stage1_52[133],stage1_51[194]}
   );
   gpc615_5 gpc1977 (
      {stage0_51[290], stage0_51[291], stage0_51[292], stage0_51[293], stage0_51[294]},
      {stage0_52[250]},
      {stage0_53[204], stage0_53[205], stage0_53[206], stage0_53[207], stage0_53[208], stage0_53[209]},
      {stage1_55[34],stage1_54[70],stage1_53[84],stage1_52[134],stage1_51[195]}
   );
   gpc615_5 gpc1978 (
      {stage0_51[295], stage0_51[296], stage0_51[297], stage0_51[298], stage0_51[299]},
      {stage0_52[251]},
      {stage0_53[210], stage0_53[211], stage0_53[212], stage0_53[213], stage0_53[214], stage0_53[215]},
      {stage1_55[35],stage1_54[71],stage1_53[85],stage1_52[135],stage1_51[196]}
   );
   gpc615_5 gpc1979 (
      {stage0_51[300], stage0_51[301], stage0_51[302], stage0_51[303], stage0_51[304]},
      {stage0_52[252]},
      {stage0_53[216], stage0_53[217], stage0_53[218], stage0_53[219], stage0_53[220], stage0_53[221]},
      {stage1_55[36],stage1_54[72],stage1_53[86],stage1_52[136],stage1_51[197]}
   );
   gpc615_5 gpc1980 (
      {stage0_51[305], stage0_51[306], stage0_51[307], stage0_51[308], stage0_51[309]},
      {stage0_52[253]},
      {stage0_53[222], stage0_53[223], stage0_53[224], stage0_53[225], stage0_53[226], stage0_53[227]},
      {stage1_55[37],stage1_54[73],stage1_53[87],stage1_52[137],stage1_51[198]}
   );
   gpc615_5 gpc1981 (
      {stage0_51[310], stage0_51[311], stage0_51[312], stage0_51[313], stage0_51[314]},
      {stage0_52[254]},
      {stage0_53[228], stage0_53[229], stage0_53[230], stage0_53[231], stage0_53[232], stage0_53[233]},
      {stage1_55[38],stage1_54[74],stage1_53[88],stage1_52[138],stage1_51[199]}
   );
   gpc615_5 gpc1982 (
      {stage0_51[315], stage0_51[316], stage0_51[317], stage0_51[318], stage0_51[319]},
      {stage0_52[255]},
      {stage0_53[234], stage0_53[235], stage0_53[236], stage0_53[237], stage0_53[238], stage0_53[239]},
      {stage1_55[39],stage1_54[75],stage1_53[89],stage1_52[139],stage1_51[200]}
   );
   gpc615_5 gpc1983 (
      {stage0_51[320], stage0_51[321], stage0_51[322], stage0_51[323], stage0_51[324]},
      {stage0_52[256]},
      {stage0_53[240], stage0_53[241], stage0_53[242], stage0_53[243], stage0_53[244], stage0_53[245]},
      {stage1_55[40],stage1_54[76],stage1_53[90],stage1_52[140],stage1_51[201]}
   );
   gpc615_5 gpc1984 (
      {stage0_51[325], stage0_51[326], stage0_51[327], stage0_51[328], stage0_51[329]},
      {stage0_52[257]},
      {stage0_53[246], stage0_53[247], stage0_53[248], stage0_53[249], stage0_53[250], stage0_53[251]},
      {stage1_55[41],stage1_54[77],stage1_53[91],stage1_52[141],stage1_51[202]}
   );
   gpc615_5 gpc1985 (
      {stage0_51[330], stage0_51[331], stage0_51[332], stage0_51[333], stage0_51[334]},
      {stage0_52[258]},
      {stage0_53[252], stage0_53[253], stage0_53[254], stage0_53[255], stage0_53[256], stage0_53[257]},
      {stage1_55[42],stage1_54[78],stage1_53[92],stage1_52[142],stage1_51[203]}
   );
   gpc615_5 gpc1986 (
      {stage0_51[335], stage0_51[336], stage0_51[337], stage0_51[338], stage0_51[339]},
      {stage0_52[259]},
      {stage0_53[258], stage0_53[259], stage0_53[260], stage0_53[261], stage0_53[262], stage0_53[263]},
      {stage1_55[43],stage1_54[79],stage1_53[93],stage1_52[143],stage1_51[204]}
   );
   gpc615_5 gpc1987 (
      {stage0_51[340], stage0_51[341], stage0_51[342], stage0_51[343], stage0_51[344]},
      {stage0_52[260]},
      {stage0_53[264], stage0_53[265], stage0_53[266], stage0_53[267], stage0_53[268], stage0_53[269]},
      {stage1_55[44],stage1_54[80],stage1_53[94],stage1_52[144],stage1_51[205]}
   );
   gpc615_5 gpc1988 (
      {stage0_51[345], stage0_51[346], stage0_51[347], stage0_51[348], stage0_51[349]},
      {stage0_52[261]},
      {stage0_53[270], stage0_53[271], stage0_53[272], stage0_53[273], stage0_53[274], stage0_53[275]},
      {stage1_55[45],stage1_54[81],stage1_53[95],stage1_52[145],stage1_51[206]}
   );
   gpc615_5 gpc1989 (
      {stage0_51[350], stage0_51[351], stage0_51[352], stage0_51[353], stage0_51[354]},
      {stage0_52[262]},
      {stage0_53[276], stage0_53[277], stage0_53[278], stage0_53[279], stage0_53[280], stage0_53[281]},
      {stage1_55[46],stage1_54[82],stage1_53[96],stage1_52[146],stage1_51[207]}
   );
   gpc615_5 gpc1990 (
      {stage0_51[355], stage0_51[356], stage0_51[357], stage0_51[358], stage0_51[359]},
      {stage0_52[263]},
      {stage0_53[282], stage0_53[283], stage0_53[284], stage0_53[285], stage0_53[286], stage0_53[287]},
      {stage1_55[47],stage1_54[83],stage1_53[97],stage1_52[147],stage1_51[208]}
   );
   gpc615_5 gpc1991 (
      {stage0_51[360], stage0_51[361], stage0_51[362], stage0_51[363], stage0_51[364]},
      {stage0_52[264]},
      {stage0_53[288], stage0_53[289], stage0_53[290], stage0_53[291], stage0_53[292], stage0_53[293]},
      {stage1_55[48],stage1_54[84],stage1_53[98],stage1_52[148],stage1_51[209]}
   );
   gpc615_5 gpc1992 (
      {stage0_51[365], stage0_51[366], stage0_51[367], stage0_51[368], stage0_51[369]},
      {stage0_52[265]},
      {stage0_53[294], stage0_53[295], stage0_53[296], stage0_53[297], stage0_53[298], stage0_53[299]},
      {stage1_55[49],stage1_54[85],stage1_53[99],stage1_52[149],stage1_51[210]}
   );
   gpc615_5 gpc1993 (
      {stage0_51[370], stage0_51[371], stage0_51[372], stage0_51[373], stage0_51[374]},
      {stage0_52[266]},
      {stage0_53[300], stage0_53[301], stage0_53[302], stage0_53[303], stage0_53[304], stage0_53[305]},
      {stage1_55[50],stage1_54[86],stage1_53[100],stage1_52[150],stage1_51[211]}
   );
   gpc615_5 gpc1994 (
      {stage0_51[375], stage0_51[376], stage0_51[377], stage0_51[378], stage0_51[379]},
      {stage0_52[267]},
      {stage0_53[306], stage0_53[307], stage0_53[308], stage0_53[309], stage0_53[310], stage0_53[311]},
      {stage1_55[51],stage1_54[87],stage1_53[101],stage1_52[151],stage1_51[212]}
   );
   gpc615_5 gpc1995 (
      {stage0_51[380], stage0_51[381], stage0_51[382], stage0_51[383], stage0_51[384]},
      {stage0_52[268]},
      {stage0_53[312], stage0_53[313], stage0_53[314], stage0_53[315], stage0_53[316], stage0_53[317]},
      {stage1_55[52],stage1_54[88],stage1_53[102],stage1_52[152],stage1_51[213]}
   );
   gpc615_5 gpc1996 (
      {stage0_51[385], stage0_51[386], stage0_51[387], stage0_51[388], stage0_51[389]},
      {stage0_52[269]},
      {stage0_53[318], stage0_53[319], stage0_53[320], stage0_53[321], stage0_53[322], stage0_53[323]},
      {stage1_55[53],stage1_54[89],stage1_53[103],stage1_52[153],stage1_51[214]}
   );
   gpc615_5 gpc1997 (
      {stage0_51[390], stage0_51[391], stage0_51[392], stage0_51[393], stage0_51[394]},
      {stage0_52[270]},
      {stage0_53[324], stage0_53[325], stage0_53[326], stage0_53[327], stage0_53[328], stage0_53[329]},
      {stage1_55[54],stage1_54[90],stage1_53[104],stage1_52[154],stage1_51[215]}
   );
   gpc615_5 gpc1998 (
      {stage0_51[395], stage0_51[396], stage0_51[397], stage0_51[398], stage0_51[399]},
      {stage0_52[271]},
      {stage0_53[330], stage0_53[331], stage0_53[332], stage0_53[333], stage0_53[334], stage0_53[335]},
      {stage1_55[55],stage1_54[91],stage1_53[105],stage1_52[155],stage1_51[216]}
   );
   gpc615_5 gpc1999 (
      {stage0_51[400], stage0_51[401], stage0_51[402], stage0_51[403], stage0_51[404]},
      {stage0_52[272]},
      {stage0_53[336], stage0_53[337], stage0_53[338], stage0_53[339], stage0_53[340], stage0_53[341]},
      {stage1_55[56],stage1_54[92],stage1_53[106],stage1_52[156],stage1_51[217]}
   );
   gpc615_5 gpc2000 (
      {stage0_51[405], stage0_51[406], stage0_51[407], stage0_51[408], stage0_51[409]},
      {stage0_52[273]},
      {stage0_53[342], stage0_53[343], stage0_53[344], stage0_53[345], stage0_53[346], stage0_53[347]},
      {stage1_55[57],stage1_54[93],stage1_53[107],stage1_52[157],stage1_51[218]}
   );
   gpc615_5 gpc2001 (
      {stage0_51[410], stage0_51[411], stage0_51[412], stage0_51[413], stage0_51[414]},
      {stage0_52[274]},
      {stage0_53[348], stage0_53[349], stage0_53[350], stage0_53[351], stage0_53[352], stage0_53[353]},
      {stage1_55[58],stage1_54[94],stage1_53[108],stage1_52[158],stage1_51[219]}
   );
   gpc615_5 gpc2002 (
      {stage0_51[415], stage0_51[416], stage0_51[417], stage0_51[418], stage0_51[419]},
      {stage0_52[275]},
      {stage0_53[354], stage0_53[355], stage0_53[356], stage0_53[357], stage0_53[358], stage0_53[359]},
      {stage1_55[59],stage1_54[95],stage1_53[109],stage1_52[159],stage1_51[220]}
   );
   gpc615_5 gpc2003 (
      {stage0_51[420], stage0_51[421], stage0_51[422], stage0_51[423], stage0_51[424]},
      {stage0_52[276]},
      {stage0_53[360], stage0_53[361], stage0_53[362], stage0_53[363], stage0_53[364], stage0_53[365]},
      {stage1_55[60],stage1_54[96],stage1_53[110],stage1_52[160],stage1_51[221]}
   );
   gpc615_5 gpc2004 (
      {stage0_51[425], stage0_51[426], stage0_51[427], stage0_51[428], stage0_51[429]},
      {stage0_52[277]},
      {stage0_53[366], stage0_53[367], stage0_53[368], stage0_53[369], stage0_53[370], stage0_53[371]},
      {stage1_55[61],stage1_54[97],stage1_53[111],stage1_52[161],stage1_51[222]}
   );
   gpc615_5 gpc2005 (
      {stage0_51[430], stage0_51[431], stage0_51[432], stage0_51[433], stage0_51[434]},
      {stage0_52[278]},
      {stage0_53[372], stage0_53[373], stage0_53[374], stage0_53[375], stage0_53[376], stage0_53[377]},
      {stage1_55[62],stage1_54[98],stage1_53[112],stage1_52[162],stage1_51[223]}
   );
   gpc606_5 gpc2006 (
      {stage0_52[279], stage0_52[280], stage0_52[281], stage0_52[282], stage0_52[283], stage0_52[284]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[63],stage1_54[99],stage1_53[113],stage1_52[163]}
   );
   gpc606_5 gpc2007 (
      {stage0_52[285], stage0_52[286], stage0_52[287], stage0_52[288], stage0_52[289], stage0_52[290]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[64],stage1_54[100],stage1_53[114],stage1_52[164]}
   );
   gpc606_5 gpc2008 (
      {stage0_52[291], stage0_52[292], stage0_52[293], stage0_52[294], stage0_52[295], stage0_52[296]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[65],stage1_54[101],stage1_53[115],stage1_52[165]}
   );
   gpc606_5 gpc2009 (
      {stage0_52[297], stage0_52[298], stage0_52[299], stage0_52[300], stage0_52[301], stage0_52[302]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[66],stage1_54[102],stage1_53[116],stage1_52[166]}
   );
   gpc606_5 gpc2010 (
      {stage0_52[303], stage0_52[304], stage0_52[305], stage0_52[306], stage0_52[307], stage0_52[308]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[67],stage1_54[103],stage1_53[117],stage1_52[167]}
   );
   gpc606_5 gpc2011 (
      {stage0_52[309], stage0_52[310], stage0_52[311], stage0_52[312], stage0_52[313], stage0_52[314]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[68],stage1_54[104],stage1_53[118],stage1_52[168]}
   );
   gpc606_5 gpc2012 (
      {stage0_52[315], stage0_52[316], stage0_52[317], stage0_52[318], stage0_52[319], stage0_52[320]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[69],stage1_54[105],stage1_53[119],stage1_52[169]}
   );
   gpc606_5 gpc2013 (
      {stage0_52[321], stage0_52[322], stage0_52[323], stage0_52[324], stage0_52[325], stage0_52[326]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[70],stage1_54[106],stage1_53[120],stage1_52[170]}
   );
   gpc606_5 gpc2014 (
      {stage0_52[327], stage0_52[328], stage0_52[329], stage0_52[330], stage0_52[331], stage0_52[332]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[71],stage1_54[107],stage1_53[121],stage1_52[171]}
   );
   gpc606_5 gpc2015 (
      {stage0_52[333], stage0_52[334], stage0_52[335], stage0_52[336], stage0_52[337], stage0_52[338]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[72],stage1_54[108],stage1_53[122],stage1_52[172]}
   );
   gpc606_5 gpc2016 (
      {stage0_52[339], stage0_52[340], stage0_52[341], stage0_52[342], stage0_52[343], stage0_52[344]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[73],stage1_54[109],stage1_53[123],stage1_52[173]}
   );
   gpc606_5 gpc2017 (
      {stage0_52[345], stage0_52[346], stage0_52[347], stage0_52[348], stage0_52[349], stage0_52[350]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[74],stage1_54[110],stage1_53[124],stage1_52[174]}
   );
   gpc606_5 gpc2018 (
      {stage0_52[351], stage0_52[352], stage0_52[353], stage0_52[354], stage0_52[355], stage0_52[356]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[75],stage1_54[111],stage1_53[125],stage1_52[175]}
   );
   gpc606_5 gpc2019 (
      {stage0_52[357], stage0_52[358], stage0_52[359], stage0_52[360], stage0_52[361], stage0_52[362]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[76],stage1_54[112],stage1_53[126],stage1_52[176]}
   );
   gpc606_5 gpc2020 (
      {stage0_52[363], stage0_52[364], stage0_52[365], stage0_52[366], stage0_52[367], stage0_52[368]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[77],stage1_54[113],stage1_53[127],stage1_52[177]}
   );
   gpc606_5 gpc2021 (
      {stage0_52[369], stage0_52[370], stage0_52[371], stage0_52[372], stage0_52[373], stage0_52[374]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[78],stage1_54[114],stage1_53[128],stage1_52[178]}
   );
   gpc606_5 gpc2022 (
      {stage0_52[375], stage0_52[376], stage0_52[377], stage0_52[378], stage0_52[379], stage0_52[380]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[79],stage1_54[115],stage1_53[129],stage1_52[179]}
   );
   gpc606_5 gpc2023 (
      {stage0_52[381], stage0_52[382], stage0_52[383], stage0_52[384], stage0_52[385], stage0_52[386]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[80],stage1_54[116],stage1_53[130],stage1_52[180]}
   );
   gpc606_5 gpc2024 (
      {stage0_52[387], stage0_52[388], stage0_52[389], stage0_52[390], stage0_52[391], stage0_52[392]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[81],stage1_54[117],stage1_53[131],stage1_52[181]}
   );
   gpc606_5 gpc2025 (
      {stage0_52[393], stage0_52[394], stage0_52[395], stage0_52[396], stage0_52[397], stage0_52[398]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[82],stage1_54[118],stage1_53[132],stage1_52[182]}
   );
   gpc606_5 gpc2026 (
      {stage0_52[399], stage0_52[400], stage0_52[401], stage0_52[402], stage0_52[403], stage0_52[404]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[83],stage1_54[119],stage1_53[133],stage1_52[183]}
   );
   gpc606_5 gpc2027 (
      {stage0_52[405], stage0_52[406], stage0_52[407], stage0_52[408], stage0_52[409], stage0_52[410]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[84],stage1_54[120],stage1_53[134],stage1_52[184]}
   );
   gpc606_5 gpc2028 (
      {stage0_52[411], stage0_52[412], stage0_52[413], stage0_52[414], stage0_52[415], stage0_52[416]},
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136], stage0_54[137]},
      {stage1_56[22],stage1_55[85],stage1_54[121],stage1_53[135],stage1_52[185]}
   );
   gpc606_5 gpc2029 (
      {stage0_52[417], stage0_52[418], stage0_52[419], stage0_52[420], stage0_52[421], stage0_52[422]},
      {stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141], stage0_54[142], stage0_54[143]},
      {stage1_56[23],stage1_55[86],stage1_54[122],stage1_53[136],stage1_52[186]}
   );
   gpc606_5 gpc2030 (
      {stage0_52[423], stage0_52[424], stage0_52[425], stage0_52[426], stage0_52[427], stage0_52[428]},
      {stage0_54[144], stage0_54[145], stage0_54[146], stage0_54[147], stage0_54[148], stage0_54[149]},
      {stage1_56[24],stage1_55[87],stage1_54[123],stage1_53[137],stage1_52[187]}
   );
   gpc606_5 gpc2031 (
      {stage0_52[429], stage0_52[430], stage0_52[431], stage0_52[432], stage0_52[433], stage0_52[434]},
      {stage0_54[150], stage0_54[151], stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155]},
      {stage1_56[25],stage1_55[88],stage1_54[124],stage1_53[138],stage1_52[188]}
   );
   gpc606_5 gpc2032 (
      {stage0_52[435], stage0_52[436], stage0_52[437], stage0_52[438], stage0_52[439], stage0_52[440]},
      {stage0_54[156], stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage1_56[26],stage1_55[89],stage1_54[125],stage1_53[139],stage1_52[189]}
   );
   gpc606_5 gpc2033 (
      {stage0_52[441], stage0_52[442], stage0_52[443], stage0_52[444], stage0_52[445], stage0_52[446]},
      {stage0_54[162], stage0_54[163], stage0_54[164], stage0_54[165], stage0_54[166], stage0_54[167]},
      {stage1_56[27],stage1_55[90],stage1_54[126],stage1_53[140],stage1_52[190]}
   );
   gpc615_5 gpc2034 (
      {stage0_52[447], stage0_52[448], stage0_52[449], stage0_52[450], stage0_52[451]},
      {stage0_53[378]},
      {stage0_54[168], stage0_54[169], stage0_54[170], stage0_54[171], stage0_54[172], stage0_54[173]},
      {stage1_56[28],stage1_55[91],stage1_54[127],stage1_53[141],stage1_52[191]}
   );
   gpc615_5 gpc2035 (
      {stage0_52[452], stage0_52[453], stage0_52[454], stage0_52[455], stage0_52[456]},
      {stage0_53[379]},
      {stage0_54[174], stage0_54[175], stage0_54[176], stage0_54[177], stage0_54[178], stage0_54[179]},
      {stage1_56[29],stage1_55[92],stage1_54[128],stage1_53[142],stage1_52[192]}
   );
   gpc615_5 gpc2036 (
      {stage0_52[457], stage0_52[458], stage0_52[459], stage0_52[460], stage0_52[461]},
      {stage0_53[380]},
      {stage0_54[180], stage0_54[181], stage0_54[182], stage0_54[183], stage0_54[184], stage0_54[185]},
      {stage1_56[30],stage1_55[93],stage1_54[129],stage1_53[143],stage1_52[193]}
   );
   gpc615_5 gpc2037 (
      {stage0_52[462], stage0_52[463], stage0_52[464], stage0_52[465], stage0_52[466]},
      {stage0_53[381]},
      {stage0_54[186], stage0_54[187], stage0_54[188], stage0_54[189], stage0_54[190], stage0_54[191]},
      {stage1_56[31],stage1_55[94],stage1_54[130],stage1_53[144],stage1_52[194]}
   );
   gpc615_5 gpc2038 (
      {stage0_52[467], stage0_52[468], stage0_52[469], stage0_52[470], stage0_52[471]},
      {stage0_53[382]},
      {stage0_54[192], stage0_54[193], stage0_54[194], stage0_54[195], stage0_54[196], stage0_54[197]},
      {stage1_56[32],stage1_55[95],stage1_54[131],stage1_53[145],stage1_52[195]}
   );
   gpc615_5 gpc2039 (
      {stage0_52[472], stage0_52[473], stage0_52[474], stage0_52[475], stage0_52[476]},
      {stage0_53[383]},
      {stage0_54[198], stage0_54[199], stage0_54[200], stage0_54[201], stage0_54[202], stage0_54[203]},
      {stage1_56[33],stage1_55[96],stage1_54[132],stage1_53[146],stage1_52[196]}
   );
   gpc615_5 gpc2040 (
      {stage0_52[477], stage0_52[478], stage0_52[479], stage0_52[480], stage0_52[481]},
      {stage0_53[384]},
      {stage0_54[204], stage0_54[205], stage0_54[206], stage0_54[207], stage0_54[208], stage0_54[209]},
      {stage1_56[34],stage1_55[97],stage1_54[133],stage1_53[147],stage1_52[197]}
   );
   gpc615_5 gpc2041 (
      {stage0_52[482], stage0_52[483], stage0_52[484], stage0_52[485], 1'b0},
      {stage0_53[385]},
      {stage0_54[210], stage0_54[211], stage0_54[212], stage0_54[213], stage0_54[214], stage0_54[215]},
      {stage1_56[35],stage1_55[98],stage1_54[134],stage1_53[148],stage1_52[198]}
   );
   gpc615_5 gpc2042 (
      {stage0_53[386], stage0_53[387], stage0_53[388], stage0_53[389], stage0_53[390]},
      {stage0_54[216]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[36],stage1_55[99],stage1_54[135],stage1_53[149]}
   );
   gpc615_5 gpc2043 (
      {stage0_53[391], stage0_53[392], stage0_53[393], stage0_53[394], stage0_53[395]},
      {stage0_54[217]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[37],stage1_55[100],stage1_54[136],stage1_53[150]}
   );
   gpc615_5 gpc2044 (
      {stage0_53[396], stage0_53[397], stage0_53[398], stage0_53[399], stage0_53[400]},
      {stage0_54[218]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[38],stage1_55[101],stage1_54[137],stage1_53[151]}
   );
   gpc615_5 gpc2045 (
      {stage0_53[401], stage0_53[402], stage0_53[403], stage0_53[404], stage0_53[405]},
      {stage0_54[219]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[39],stage1_55[102],stage1_54[138],stage1_53[152]}
   );
   gpc615_5 gpc2046 (
      {stage0_53[406], stage0_53[407], stage0_53[408], stage0_53[409], stage0_53[410]},
      {stage0_54[220]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[40],stage1_55[103],stage1_54[139],stage1_53[153]}
   );
   gpc615_5 gpc2047 (
      {stage0_53[411], stage0_53[412], stage0_53[413], stage0_53[414], stage0_53[415]},
      {stage0_54[221]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[41],stage1_55[104],stage1_54[140],stage1_53[154]}
   );
   gpc615_5 gpc2048 (
      {stage0_53[416], stage0_53[417], stage0_53[418], stage0_53[419], stage0_53[420]},
      {stage0_54[222]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[42],stage1_55[105],stage1_54[141],stage1_53[155]}
   );
   gpc615_5 gpc2049 (
      {stage0_53[421], stage0_53[422], stage0_53[423], stage0_53[424], stage0_53[425]},
      {stage0_54[223]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[43],stage1_55[106],stage1_54[142],stage1_53[156]}
   );
   gpc615_5 gpc2050 (
      {stage0_53[426], stage0_53[427], stage0_53[428], stage0_53[429], stage0_53[430]},
      {stage0_54[224]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[44],stage1_55[107],stage1_54[143],stage1_53[157]}
   );
   gpc615_5 gpc2051 (
      {stage0_53[431], stage0_53[432], stage0_53[433], stage0_53[434], stage0_53[435]},
      {stage0_54[225]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[45],stage1_55[108],stage1_54[144],stage1_53[158]}
   );
   gpc615_5 gpc2052 (
      {stage0_53[436], stage0_53[437], stage0_53[438], stage0_53[439], stage0_53[440]},
      {stage0_54[226]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[46],stage1_55[109],stage1_54[145],stage1_53[159]}
   );
   gpc615_5 gpc2053 (
      {stage0_53[441], stage0_53[442], stage0_53[443], stage0_53[444], stage0_53[445]},
      {stage0_54[227]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[47],stage1_55[110],stage1_54[146],stage1_53[160]}
   );
   gpc615_5 gpc2054 (
      {stage0_53[446], stage0_53[447], stage0_53[448], stage0_53[449], stage0_53[450]},
      {stage0_54[228]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[48],stage1_55[111],stage1_54[147],stage1_53[161]}
   );
   gpc615_5 gpc2055 (
      {stage0_53[451], stage0_53[452], stage0_53[453], stage0_53[454], stage0_53[455]},
      {stage0_54[229]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[49],stage1_55[112],stage1_54[148],stage1_53[162]}
   );
   gpc615_5 gpc2056 (
      {stage0_53[456], stage0_53[457], stage0_53[458], stage0_53[459], stage0_53[460]},
      {stage0_54[230]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[50],stage1_55[113],stage1_54[149],stage1_53[163]}
   );
   gpc615_5 gpc2057 (
      {stage0_53[461], stage0_53[462], stage0_53[463], stage0_53[464], stage0_53[465]},
      {stage0_54[231]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[51],stage1_55[114],stage1_54[150],stage1_53[164]}
   );
   gpc615_5 gpc2058 (
      {stage0_53[466], stage0_53[467], stage0_53[468], stage0_53[469], stage0_53[470]},
      {stage0_54[232]},
      {stage0_55[96], stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101]},
      {stage1_57[16],stage1_56[52],stage1_55[115],stage1_54[151],stage1_53[165]}
   );
   gpc615_5 gpc2059 (
      {stage0_53[471], stage0_53[472], stage0_53[473], stage0_53[474], stage0_53[475]},
      {stage0_54[233]},
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage1_57[17],stage1_56[53],stage1_55[116],stage1_54[152],stage1_53[166]}
   );
   gpc615_5 gpc2060 (
      {stage0_53[476], stage0_53[477], stage0_53[478], stage0_53[479], stage0_53[480]},
      {stage0_54[234]},
      {stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111], stage0_55[112], stage0_55[113]},
      {stage1_57[18],stage1_56[54],stage1_55[117],stage1_54[153],stage1_53[167]}
   );
   gpc615_5 gpc2061 (
      {stage0_53[481], stage0_53[482], stage0_53[483], stage0_53[484], stage0_53[485]},
      {stage0_54[235]},
      {stage0_55[114], stage0_55[115], stage0_55[116], stage0_55[117], stage0_55[118], stage0_55[119]},
      {stage1_57[19],stage1_56[55],stage1_55[118],stage1_54[154],stage1_53[168]}
   );
   gpc117_4 gpc2062 (
      {stage0_54[236], stage0_54[237], stage0_54[238], stage0_54[239], stage0_54[240], stage0_54[241], stage0_54[242]},
      {stage0_55[120]},
      {stage0_56[0]},
      {stage1_57[20],stage1_56[56],stage1_55[119],stage1_54[155]}
   );
   gpc615_5 gpc2063 (
      {stage0_54[243], stage0_54[244], stage0_54[245], stage0_54[246], stage0_54[247]},
      {stage0_55[121]},
      {stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5], stage0_56[6]},
      {stage1_58[0],stage1_57[21],stage1_56[57],stage1_55[120],stage1_54[156]}
   );
   gpc615_5 gpc2064 (
      {stage0_54[248], stage0_54[249], stage0_54[250], stage0_54[251], stage0_54[252]},
      {stage0_55[122]},
      {stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11], stage0_56[12]},
      {stage1_58[1],stage1_57[22],stage1_56[58],stage1_55[121],stage1_54[157]}
   );
   gpc615_5 gpc2065 (
      {stage0_54[253], stage0_54[254], stage0_54[255], stage0_54[256], stage0_54[257]},
      {stage0_55[123]},
      {stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17], stage0_56[18]},
      {stage1_58[2],stage1_57[23],stage1_56[59],stage1_55[122],stage1_54[158]}
   );
   gpc615_5 gpc2066 (
      {stage0_54[258], stage0_54[259], stage0_54[260], stage0_54[261], stage0_54[262]},
      {stage0_55[124]},
      {stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23], stage0_56[24]},
      {stage1_58[3],stage1_57[24],stage1_56[60],stage1_55[123],stage1_54[159]}
   );
   gpc615_5 gpc2067 (
      {stage0_54[263], stage0_54[264], stage0_54[265], stage0_54[266], stage0_54[267]},
      {stage0_55[125]},
      {stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29], stage0_56[30]},
      {stage1_58[4],stage1_57[25],stage1_56[61],stage1_55[124],stage1_54[160]}
   );
   gpc615_5 gpc2068 (
      {stage0_54[268], stage0_54[269], stage0_54[270], stage0_54[271], stage0_54[272]},
      {stage0_55[126]},
      {stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35], stage0_56[36]},
      {stage1_58[5],stage1_57[26],stage1_56[62],stage1_55[125],stage1_54[161]}
   );
   gpc615_5 gpc2069 (
      {stage0_54[273], stage0_54[274], stage0_54[275], stage0_54[276], stage0_54[277]},
      {stage0_55[127]},
      {stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41], stage0_56[42]},
      {stage1_58[6],stage1_57[27],stage1_56[63],stage1_55[126],stage1_54[162]}
   );
   gpc615_5 gpc2070 (
      {stage0_54[278], stage0_54[279], stage0_54[280], stage0_54[281], stage0_54[282]},
      {stage0_55[128]},
      {stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47], stage0_56[48]},
      {stage1_58[7],stage1_57[28],stage1_56[64],stage1_55[127],stage1_54[163]}
   );
   gpc615_5 gpc2071 (
      {stage0_54[283], stage0_54[284], stage0_54[285], stage0_54[286], stage0_54[287]},
      {stage0_55[129]},
      {stage0_56[49], stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53], stage0_56[54]},
      {stage1_58[8],stage1_57[29],stage1_56[65],stage1_55[128],stage1_54[164]}
   );
   gpc615_5 gpc2072 (
      {stage0_54[288], stage0_54[289], stage0_54[290], stage0_54[291], stage0_54[292]},
      {stage0_55[130]},
      {stage0_56[55], stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60]},
      {stage1_58[9],stage1_57[30],stage1_56[66],stage1_55[129],stage1_54[165]}
   );
   gpc615_5 gpc2073 (
      {stage0_54[293], stage0_54[294], stage0_54[295], stage0_54[296], stage0_54[297]},
      {stage0_55[131]},
      {stage0_56[61], stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65], stage0_56[66]},
      {stage1_58[10],stage1_57[31],stage1_56[67],stage1_55[130],stage1_54[166]}
   );
   gpc615_5 gpc2074 (
      {stage0_54[298], stage0_54[299], stage0_54[300], stage0_54[301], stage0_54[302]},
      {stage0_55[132]},
      {stage0_56[67], stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71], stage0_56[72]},
      {stage1_58[11],stage1_57[32],stage1_56[68],stage1_55[131],stage1_54[167]}
   );
   gpc615_5 gpc2075 (
      {stage0_54[303], stage0_54[304], stage0_54[305], stage0_54[306], stage0_54[307]},
      {stage0_55[133]},
      {stage0_56[73], stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77], stage0_56[78]},
      {stage1_58[12],stage1_57[33],stage1_56[69],stage1_55[132],stage1_54[168]}
   );
   gpc615_5 gpc2076 (
      {stage0_54[308], stage0_54[309], stage0_54[310], stage0_54[311], stage0_54[312]},
      {stage0_55[134]},
      {stage0_56[79], stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83], stage0_56[84]},
      {stage1_58[13],stage1_57[34],stage1_56[70],stage1_55[133],stage1_54[169]}
   );
   gpc615_5 gpc2077 (
      {stage0_54[313], stage0_54[314], stage0_54[315], stage0_54[316], stage0_54[317]},
      {stage0_55[135]},
      {stage0_56[85], stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89], stage0_56[90]},
      {stage1_58[14],stage1_57[35],stage1_56[71],stage1_55[134],stage1_54[170]}
   );
   gpc615_5 gpc2078 (
      {stage0_54[318], stage0_54[319], stage0_54[320], stage0_54[321], stage0_54[322]},
      {stage0_55[136]},
      {stage0_56[91], stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95], stage0_56[96]},
      {stage1_58[15],stage1_57[36],stage1_56[72],stage1_55[135],stage1_54[171]}
   );
   gpc615_5 gpc2079 (
      {stage0_54[323], stage0_54[324], stage0_54[325], stage0_54[326], stage0_54[327]},
      {stage0_55[137]},
      {stage0_56[97], stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101], stage0_56[102]},
      {stage1_58[16],stage1_57[37],stage1_56[73],stage1_55[136],stage1_54[172]}
   );
   gpc615_5 gpc2080 (
      {stage0_54[328], stage0_54[329], stage0_54[330], stage0_54[331], stage0_54[332]},
      {stage0_55[138]},
      {stage0_56[103], stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107], stage0_56[108]},
      {stage1_58[17],stage1_57[38],stage1_56[74],stage1_55[137],stage1_54[173]}
   );
   gpc615_5 gpc2081 (
      {stage0_54[333], stage0_54[334], stage0_54[335], stage0_54[336], stage0_54[337]},
      {stage0_55[139]},
      {stage0_56[109], stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113], stage0_56[114]},
      {stage1_58[18],stage1_57[39],stage1_56[75],stage1_55[138],stage1_54[174]}
   );
   gpc615_5 gpc2082 (
      {stage0_54[338], stage0_54[339], stage0_54[340], stage0_54[341], stage0_54[342]},
      {stage0_55[140]},
      {stage0_56[115], stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119], stage0_56[120]},
      {stage1_58[19],stage1_57[40],stage1_56[76],stage1_55[139],stage1_54[175]}
   );
   gpc615_5 gpc2083 (
      {stage0_54[343], stage0_54[344], stage0_54[345], stage0_54[346], stage0_54[347]},
      {stage0_55[141]},
      {stage0_56[121], stage0_56[122], stage0_56[123], stage0_56[124], stage0_56[125], stage0_56[126]},
      {stage1_58[20],stage1_57[41],stage1_56[77],stage1_55[140],stage1_54[176]}
   );
   gpc615_5 gpc2084 (
      {stage0_54[348], stage0_54[349], stage0_54[350], stage0_54[351], stage0_54[352]},
      {stage0_55[142]},
      {stage0_56[127], stage0_56[128], stage0_56[129], stage0_56[130], stage0_56[131], stage0_56[132]},
      {stage1_58[21],stage1_57[42],stage1_56[78],stage1_55[141],stage1_54[177]}
   );
   gpc615_5 gpc2085 (
      {stage0_54[353], stage0_54[354], stage0_54[355], stage0_54[356], stage0_54[357]},
      {stage0_55[143]},
      {stage0_56[133], stage0_56[134], stage0_56[135], stage0_56[136], stage0_56[137], stage0_56[138]},
      {stage1_58[22],stage1_57[43],stage1_56[79],stage1_55[142],stage1_54[178]}
   );
   gpc615_5 gpc2086 (
      {stage0_54[358], stage0_54[359], stage0_54[360], stage0_54[361], stage0_54[362]},
      {stage0_55[144]},
      {stage0_56[139], stage0_56[140], stage0_56[141], stage0_56[142], stage0_56[143], stage0_56[144]},
      {stage1_58[23],stage1_57[44],stage1_56[80],stage1_55[143],stage1_54[179]}
   );
   gpc615_5 gpc2087 (
      {stage0_54[363], stage0_54[364], stage0_54[365], stage0_54[366], stage0_54[367]},
      {stage0_55[145]},
      {stage0_56[145], stage0_56[146], stage0_56[147], stage0_56[148], stage0_56[149], stage0_56[150]},
      {stage1_58[24],stage1_57[45],stage1_56[81],stage1_55[144],stage1_54[180]}
   );
   gpc615_5 gpc2088 (
      {stage0_54[368], stage0_54[369], stage0_54[370], stage0_54[371], stage0_54[372]},
      {stage0_55[146]},
      {stage0_56[151], stage0_56[152], stage0_56[153], stage0_56[154], stage0_56[155], stage0_56[156]},
      {stage1_58[25],stage1_57[46],stage1_56[82],stage1_55[145],stage1_54[181]}
   );
   gpc615_5 gpc2089 (
      {stage0_54[373], stage0_54[374], stage0_54[375], stage0_54[376], stage0_54[377]},
      {stage0_55[147]},
      {stage0_56[157], stage0_56[158], stage0_56[159], stage0_56[160], stage0_56[161], stage0_56[162]},
      {stage1_58[26],stage1_57[47],stage1_56[83],stage1_55[146],stage1_54[182]}
   );
   gpc615_5 gpc2090 (
      {stage0_54[378], stage0_54[379], stage0_54[380], stage0_54[381], stage0_54[382]},
      {stage0_55[148]},
      {stage0_56[163], stage0_56[164], stage0_56[165], stage0_56[166], stage0_56[167], stage0_56[168]},
      {stage1_58[27],stage1_57[48],stage1_56[84],stage1_55[147],stage1_54[183]}
   );
   gpc615_5 gpc2091 (
      {stage0_54[383], stage0_54[384], stage0_54[385], stage0_54[386], stage0_54[387]},
      {stage0_55[149]},
      {stage0_56[169], stage0_56[170], stage0_56[171], stage0_56[172], stage0_56[173], stage0_56[174]},
      {stage1_58[28],stage1_57[49],stage1_56[85],stage1_55[148],stage1_54[184]}
   );
   gpc615_5 gpc2092 (
      {stage0_54[388], stage0_54[389], stage0_54[390], stage0_54[391], stage0_54[392]},
      {stage0_55[150]},
      {stage0_56[175], stage0_56[176], stage0_56[177], stage0_56[178], stage0_56[179], stage0_56[180]},
      {stage1_58[29],stage1_57[50],stage1_56[86],stage1_55[149],stage1_54[185]}
   );
   gpc615_5 gpc2093 (
      {stage0_54[393], stage0_54[394], stage0_54[395], stage0_54[396], stage0_54[397]},
      {stage0_55[151]},
      {stage0_56[181], stage0_56[182], stage0_56[183], stage0_56[184], stage0_56[185], stage0_56[186]},
      {stage1_58[30],stage1_57[51],stage1_56[87],stage1_55[150],stage1_54[186]}
   );
   gpc615_5 gpc2094 (
      {stage0_54[398], stage0_54[399], stage0_54[400], stage0_54[401], stage0_54[402]},
      {stage0_55[152]},
      {stage0_56[187], stage0_56[188], stage0_56[189], stage0_56[190], stage0_56[191], stage0_56[192]},
      {stage1_58[31],stage1_57[52],stage1_56[88],stage1_55[151],stage1_54[187]}
   );
   gpc615_5 gpc2095 (
      {stage0_54[403], stage0_54[404], stage0_54[405], stage0_54[406], stage0_54[407]},
      {stage0_55[153]},
      {stage0_56[193], stage0_56[194], stage0_56[195], stage0_56[196], stage0_56[197], stage0_56[198]},
      {stage1_58[32],stage1_57[53],stage1_56[89],stage1_55[152],stage1_54[188]}
   );
   gpc615_5 gpc2096 (
      {stage0_54[408], stage0_54[409], stage0_54[410], stage0_54[411], stage0_54[412]},
      {stage0_55[154]},
      {stage0_56[199], stage0_56[200], stage0_56[201], stage0_56[202], stage0_56[203], stage0_56[204]},
      {stage1_58[33],stage1_57[54],stage1_56[90],stage1_55[153],stage1_54[189]}
   );
   gpc615_5 gpc2097 (
      {stage0_54[413], stage0_54[414], stage0_54[415], stage0_54[416], stage0_54[417]},
      {stage0_55[155]},
      {stage0_56[205], stage0_56[206], stage0_56[207], stage0_56[208], stage0_56[209], stage0_56[210]},
      {stage1_58[34],stage1_57[55],stage1_56[91],stage1_55[154],stage1_54[190]}
   );
   gpc615_5 gpc2098 (
      {stage0_54[418], stage0_54[419], stage0_54[420], stage0_54[421], stage0_54[422]},
      {stage0_55[156]},
      {stage0_56[211], stage0_56[212], stage0_56[213], stage0_56[214], stage0_56[215], stage0_56[216]},
      {stage1_58[35],stage1_57[56],stage1_56[92],stage1_55[155],stage1_54[191]}
   );
   gpc615_5 gpc2099 (
      {stage0_54[423], stage0_54[424], stage0_54[425], stage0_54[426], stage0_54[427]},
      {stage0_55[157]},
      {stage0_56[217], stage0_56[218], stage0_56[219], stage0_56[220], stage0_56[221], stage0_56[222]},
      {stage1_58[36],stage1_57[57],stage1_56[93],stage1_55[156],stage1_54[192]}
   );
   gpc615_5 gpc2100 (
      {stage0_54[428], stage0_54[429], stage0_54[430], stage0_54[431], stage0_54[432]},
      {stage0_55[158]},
      {stage0_56[223], stage0_56[224], stage0_56[225], stage0_56[226], stage0_56[227], stage0_56[228]},
      {stage1_58[37],stage1_57[58],stage1_56[94],stage1_55[157],stage1_54[193]}
   );
   gpc615_5 gpc2101 (
      {stage0_54[433], stage0_54[434], stage0_54[435], stage0_54[436], stage0_54[437]},
      {stage0_55[159]},
      {stage0_56[229], stage0_56[230], stage0_56[231], stage0_56[232], stage0_56[233], stage0_56[234]},
      {stage1_58[38],stage1_57[59],stage1_56[95],stage1_55[158],stage1_54[194]}
   );
   gpc615_5 gpc2102 (
      {stage0_54[438], stage0_54[439], stage0_54[440], stage0_54[441], stage0_54[442]},
      {stage0_55[160]},
      {stage0_56[235], stage0_56[236], stage0_56[237], stage0_56[238], stage0_56[239], stage0_56[240]},
      {stage1_58[39],stage1_57[60],stage1_56[96],stage1_55[159],stage1_54[195]}
   );
   gpc615_5 gpc2103 (
      {stage0_54[443], stage0_54[444], stage0_54[445], stage0_54[446], stage0_54[447]},
      {stage0_55[161]},
      {stage0_56[241], stage0_56[242], stage0_56[243], stage0_56[244], stage0_56[245], stage0_56[246]},
      {stage1_58[40],stage1_57[61],stage1_56[97],stage1_55[160],stage1_54[196]}
   );
   gpc615_5 gpc2104 (
      {stage0_54[448], stage0_54[449], stage0_54[450], stage0_54[451], stage0_54[452]},
      {stage0_55[162]},
      {stage0_56[247], stage0_56[248], stage0_56[249], stage0_56[250], stage0_56[251], stage0_56[252]},
      {stage1_58[41],stage1_57[62],stage1_56[98],stage1_55[161],stage1_54[197]}
   );
   gpc606_5 gpc2105 (
      {stage0_55[163], stage0_55[164], stage0_55[165], stage0_55[166], stage0_55[167], stage0_55[168]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[42],stage1_57[63],stage1_56[99],stage1_55[162]}
   );
   gpc606_5 gpc2106 (
      {stage0_55[169], stage0_55[170], stage0_55[171], stage0_55[172], stage0_55[173], stage0_55[174]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[43],stage1_57[64],stage1_56[100],stage1_55[163]}
   );
   gpc606_5 gpc2107 (
      {stage0_55[175], stage0_55[176], stage0_55[177], stage0_55[178], stage0_55[179], stage0_55[180]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[44],stage1_57[65],stage1_56[101],stage1_55[164]}
   );
   gpc606_5 gpc2108 (
      {stage0_55[181], stage0_55[182], stage0_55[183], stage0_55[184], stage0_55[185], stage0_55[186]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[45],stage1_57[66],stage1_56[102],stage1_55[165]}
   );
   gpc606_5 gpc2109 (
      {stage0_55[187], stage0_55[188], stage0_55[189], stage0_55[190], stage0_55[191], stage0_55[192]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[46],stage1_57[67],stage1_56[103],stage1_55[166]}
   );
   gpc606_5 gpc2110 (
      {stage0_55[193], stage0_55[194], stage0_55[195], stage0_55[196], stage0_55[197], stage0_55[198]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[47],stage1_57[68],stage1_56[104],stage1_55[167]}
   );
   gpc606_5 gpc2111 (
      {stage0_55[199], stage0_55[200], stage0_55[201], stage0_55[202], stage0_55[203], stage0_55[204]},
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage1_59[6],stage1_58[48],stage1_57[69],stage1_56[105],stage1_55[168]}
   );
   gpc606_5 gpc2112 (
      {stage0_55[205], stage0_55[206], stage0_55[207], stage0_55[208], stage0_55[209], stage0_55[210]},
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage1_59[7],stage1_58[49],stage1_57[70],stage1_56[106],stage1_55[169]}
   );
   gpc606_5 gpc2113 (
      {stage0_55[211], stage0_55[212], stage0_55[213], stage0_55[214], stage0_55[215], stage0_55[216]},
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage1_59[8],stage1_58[50],stage1_57[71],stage1_56[107],stage1_55[170]}
   );
   gpc606_5 gpc2114 (
      {stage0_55[217], stage0_55[218], stage0_55[219], stage0_55[220], stage0_55[221], stage0_55[222]},
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage1_59[9],stage1_58[51],stage1_57[72],stage1_56[108],stage1_55[171]}
   );
   gpc606_5 gpc2115 (
      {stage0_55[223], stage0_55[224], stage0_55[225], stage0_55[226], stage0_55[227], stage0_55[228]},
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage1_59[10],stage1_58[52],stage1_57[73],stage1_56[109],stage1_55[172]}
   );
   gpc606_5 gpc2116 (
      {stage0_55[229], stage0_55[230], stage0_55[231], stage0_55[232], stage0_55[233], stage0_55[234]},
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage1_59[11],stage1_58[53],stage1_57[74],stage1_56[110],stage1_55[173]}
   );
   gpc606_5 gpc2117 (
      {stage0_55[235], stage0_55[236], stage0_55[237], stage0_55[238], stage0_55[239], stage0_55[240]},
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage1_59[12],stage1_58[54],stage1_57[75],stage1_56[111],stage1_55[174]}
   );
   gpc606_5 gpc2118 (
      {stage0_55[241], stage0_55[242], stage0_55[243], stage0_55[244], stage0_55[245], stage0_55[246]},
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage1_59[13],stage1_58[55],stage1_57[76],stage1_56[112],stage1_55[175]}
   );
   gpc606_5 gpc2119 (
      {stage0_55[247], stage0_55[248], stage0_55[249], stage0_55[250], stage0_55[251], stage0_55[252]},
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage1_59[14],stage1_58[56],stage1_57[77],stage1_56[113],stage1_55[176]}
   );
   gpc606_5 gpc2120 (
      {stage0_55[253], stage0_55[254], stage0_55[255], stage0_55[256], stage0_55[257], stage0_55[258]},
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage1_59[15],stage1_58[57],stage1_57[78],stage1_56[114],stage1_55[177]}
   );
   gpc606_5 gpc2121 (
      {stage0_55[259], stage0_55[260], stage0_55[261], stage0_55[262], stage0_55[263], stage0_55[264]},
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage1_59[16],stage1_58[58],stage1_57[79],stage1_56[115],stage1_55[178]}
   );
   gpc606_5 gpc2122 (
      {stage0_55[265], stage0_55[266], stage0_55[267], stage0_55[268], stage0_55[269], stage0_55[270]},
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage1_59[17],stage1_58[59],stage1_57[80],stage1_56[116],stage1_55[179]}
   );
   gpc606_5 gpc2123 (
      {stage0_55[271], stage0_55[272], stage0_55[273], stage0_55[274], stage0_55[275], stage0_55[276]},
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage1_59[18],stage1_58[60],stage1_57[81],stage1_56[117],stage1_55[180]}
   );
   gpc606_5 gpc2124 (
      {stage0_55[277], stage0_55[278], stage0_55[279], stage0_55[280], stage0_55[281], stage0_55[282]},
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage1_59[19],stage1_58[61],stage1_57[82],stage1_56[118],stage1_55[181]}
   );
   gpc606_5 gpc2125 (
      {stage0_55[283], stage0_55[284], stage0_55[285], stage0_55[286], stage0_55[287], stage0_55[288]},
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage1_59[20],stage1_58[62],stage1_57[83],stage1_56[119],stage1_55[182]}
   );
   gpc606_5 gpc2126 (
      {stage0_55[289], stage0_55[290], stage0_55[291], stage0_55[292], stage0_55[293], stage0_55[294]},
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage1_59[21],stage1_58[63],stage1_57[84],stage1_56[120],stage1_55[183]}
   );
   gpc606_5 gpc2127 (
      {stage0_55[295], stage0_55[296], stage0_55[297], stage0_55[298], stage0_55[299], stage0_55[300]},
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage1_59[22],stage1_58[64],stage1_57[85],stage1_56[121],stage1_55[184]}
   );
   gpc606_5 gpc2128 (
      {stage0_55[301], stage0_55[302], stage0_55[303], stage0_55[304], stage0_55[305], stage0_55[306]},
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage1_59[23],stage1_58[65],stage1_57[86],stage1_56[122],stage1_55[185]}
   );
   gpc606_5 gpc2129 (
      {stage0_55[307], stage0_55[308], stage0_55[309], stage0_55[310], stage0_55[311], stage0_55[312]},
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage1_59[24],stage1_58[66],stage1_57[87],stage1_56[123],stage1_55[186]}
   );
   gpc606_5 gpc2130 (
      {stage0_55[313], stage0_55[314], stage0_55[315], stage0_55[316], stage0_55[317], stage0_55[318]},
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage1_59[25],stage1_58[67],stage1_57[88],stage1_56[124],stage1_55[187]}
   );
   gpc606_5 gpc2131 (
      {stage0_55[319], stage0_55[320], stage0_55[321], stage0_55[322], stage0_55[323], stage0_55[324]},
      {stage0_57[156], stage0_57[157], stage0_57[158], stage0_57[159], stage0_57[160], stage0_57[161]},
      {stage1_59[26],stage1_58[68],stage1_57[89],stage1_56[125],stage1_55[188]}
   );
   gpc606_5 gpc2132 (
      {stage0_55[325], stage0_55[326], stage0_55[327], stage0_55[328], stage0_55[329], stage0_55[330]},
      {stage0_57[162], stage0_57[163], stage0_57[164], stage0_57[165], stage0_57[166], stage0_57[167]},
      {stage1_59[27],stage1_58[69],stage1_57[90],stage1_56[126],stage1_55[189]}
   );
   gpc606_5 gpc2133 (
      {stage0_55[331], stage0_55[332], stage0_55[333], stage0_55[334], stage0_55[335], stage0_55[336]},
      {stage0_57[168], stage0_57[169], stage0_57[170], stage0_57[171], stage0_57[172], stage0_57[173]},
      {stage1_59[28],stage1_58[70],stage1_57[91],stage1_56[127],stage1_55[190]}
   );
   gpc606_5 gpc2134 (
      {stage0_55[337], stage0_55[338], stage0_55[339], stage0_55[340], stage0_55[341], stage0_55[342]},
      {stage0_57[174], stage0_57[175], stage0_57[176], stage0_57[177], stage0_57[178], stage0_57[179]},
      {stage1_59[29],stage1_58[71],stage1_57[92],stage1_56[128],stage1_55[191]}
   );
   gpc606_5 gpc2135 (
      {stage0_55[343], stage0_55[344], stage0_55[345], stage0_55[346], stage0_55[347], stage0_55[348]},
      {stage0_57[180], stage0_57[181], stage0_57[182], stage0_57[183], stage0_57[184], stage0_57[185]},
      {stage1_59[30],stage1_58[72],stage1_57[93],stage1_56[129],stage1_55[192]}
   );
   gpc606_5 gpc2136 (
      {stage0_55[349], stage0_55[350], stage0_55[351], stage0_55[352], stage0_55[353], stage0_55[354]},
      {stage0_57[186], stage0_57[187], stage0_57[188], stage0_57[189], stage0_57[190], stage0_57[191]},
      {stage1_59[31],stage1_58[73],stage1_57[94],stage1_56[130],stage1_55[193]}
   );
   gpc606_5 gpc2137 (
      {stage0_55[355], stage0_55[356], stage0_55[357], stage0_55[358], stage0_55[359], stage0_55[360]},
      {stage0_57[192], stage0_57[193], stage0_57[194], stage0_57[195], stage0_57[196], stage0_57[197]},
      {stage1_59[32],stage1_58[74],stage1_57[95],stage1_56[131],stage1_55[194]}
   );
   gpc606_5 gpc2138 (
      {stage0_55[361], stage0_55[362], stage0_55[363], stage0_55[364], stage0_55[365], stage0_55[366]},
      {stage0_57[198], stage0_57[199], stage0_57[200], stage0_57[201], stage0_57[202], stage0_57[203]},
      {stage1_59[33],stage1_58[75],stage1_57[96],stage1_56[132],stage1_55[195]}
   );
   gpc606_5 gpc2139 (
      {stage0_55[367], stage0_55[368], stage0_55[369], stage0_55[370], stage0_55[371], stage0_55[372]},
      {stage0_57[204], stage0_57[205], stage0_57[206], stage0_57[207], stage0_57[208], stage0_57[209]},
      {stage1_59[34],stage1_58[76],stage1_57[97],stage1_56[133],stage1_55[196]}
   );
   gpc606_5 gpc2140 (
      {stage0_55[373], stage0_55[374], stage0_55[375], stage0_55[376], stage0_55[377], stage0_55[378]},
      {stage0_57[210], stage0_57[211], stage0_57[212], stage0_57[213], stage0_57[214], stage0_57[215]},
      {stage1_59[35],stage1_58[77],stage1_57[98],stage1_56[134],stage1_55[197]}
   );
   gpc606_5 gpc2141 (
      {stage0_55[379], stage0_55[380], stage0_55[381], stage0_55[382], stage0_55[383], stage0_55[384]},
      {stage0_57[216], stage0_57[217], stage0_57[218], stage0_57[219], stage0_57[220], stage0_57[221]},
      {stage1_59[36],stage1_58[78],stage1_57[99],stage1_56[135],stage1_55[198]}
   );
   gpc606_5 gpc2142 (
      {stage0_55[385], stage0_55[386], stage0_55[387], stage0_55[388], stage0_55[389], stage0_55[390]},
      {stage0_57[222], stage0_57[223], stage0_57[224], stage0_57[225], stage0_57[226], stage0_57[227]},
      {stage1_59[37],stage1_58[79],stage1_57[100],stage1_56[136],stage1_55[199]}
   );
   gpc606_5 gpc2143 (
      {stage0_55[391], stage0_55[392], stage0_55[393], stage0_55[394], stage0_55[395], stage0_55[396]},
      {stage0_57[228], stage0_57[229], stage0_57[230], stage0_57[231], stage0_57[232], stage0_57[233]},
      {stage1_59[38],stage1_58[80],stage1_57[101],stage1_56[137],stage1_55[200]}
   );
   gpc606_5 gpc2144 (
      {stage0_55[397], stage0_55[398], stage0_55[399], stage0_55[400], stage0_55[401], stage0_55[402]},
      {stage0_57[234], stage0_57[235], stage0_57[236], stage0_57[237], stage0_57[238], stage0_57[239]},
      {stage1_59[39],stage1_58[81],stage1_57[102],stage1_56[138],stage1_55[201]}
   );
   gpc606_5 gpc2145 (
      {stage0_55[403], stage0_55[404], stage0_55[405], stage0_55[406], stage0_55[407], stage0_55[408]},
      {stage0_57[240], stage0_57[241], stage0_57[242], stage0_57[243], stage0_57[244], stage0_57[245]},
      {stage1_59[40],stage1_58[82],stage1_57[103],stage1_56[139],stage1_55[202]}
   );
   gpc606_5 gpc2146 (
      {stage0_55[409], stage0_55[410], stage0_55[411], stage0_55[412], stage0_55[413], stage0_55[414]},
      {stage0_57[246], stage0_57[247], stage0_57[248], stage0_57[249], stage0_57[250], stage0_57[251]},
      {stage1_59[41],stage1_58[83],stage1_57[104],stage1_56[140],stage1_55[203]}
   );
   gpc615_5 gpc2147 (
      {stage0_55[415], stage0_55[416], stage0_55[417], stage0_55[418], stage0_55[419]},
      {stage0_56[253]},
      {stage0_57[252], stage0_57[253], stage0_57[254], stage0_57[255], stage0_57[256], stage0_57[257]},
      {stage1_59[42],stage1_58[84],stage1_57[105],stage1_56[141],stage1_55[204]}
   );
   gpc615_5 gpc2148 (
      {stage0_55[420], stage0_55[421], stage0_55[422], stage0_55[423], stage0_55[424]},
      {stage0_56[254]},
      {stage0_57[258], stage0_57[259], stage0_57[260], stage0_57[261], stage0_57[262], stage0_57[263]},
      {stage1_59[43],stage1_58[85],stage1_57[106],stage1_56[142],stage1_55[205]}
   );
   gpc606_5 gpc2149 (
      {stage0_56[255], stage0_56[256], stage0_56[257], stage0_56[258], stage0_56[259], stage0_56[260]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[44],stage1_58[86],stage1_57[107],stage1_56[143]}
   );
   gpc606_5 gpc2150 (
      {stage0_56[261], stage0_56[262], stage0_56[263], stage0_56[264], stage0_56[265], stage0_56[266]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[45],stage1_58[87],stage1_57[108],stage1_56[144]}
   );
   gpc606_5 gpc2151 (
      {stage0_56[267], stage0_56[268], stage0_56[269], stage0_56[270], stage0_56[271], stage0_56[272]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[46],stage1_58[88],stage1_57[109],stage1_56[145]}
   );
   gpc606_5 gpc2152 (
      {stage0_56[273], stage0_56[274], stage0_56[275], stage0_56[276], stage0_56[277], stage0_56[278]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[47],stage1_58[89],stage1_57[110],stage1_56[146]}
   );
   gpc606_5 gpc2153 (
      {stage0_56[279], stage0_56[280], stage0_56[281], stage0_56[282], stage0_56[283], stage0_56[284]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[48],stage1_58[90],stage1_57[111],stage1_56[147]}
   );
   gpc606_5 gpc2154 (
      {stage0_56[285], stage0_56[286], stage0_56[287], stage0_56[288], stage0_56[289], stage0_56[290]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[49],stage1_58[91],stage1_57[112],stage1_56[148]}
   );
   gpc606_5 gpc2155 (
      {stage0_56[291], stage0_56[292], stage0_56[293], stage0_56[294], stage0_56[295], stage0_56[296]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[50],stage1_58[92],stage1_57[113],stage1_56[149]}
   );
   gpc606_5 gpc2156 (
      {stage0_56[297], stage0_56[298], stage0_56[299], stage0_56[300], stage0_56[301], stage0_56[302]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[51],stage1_58[93],stage1_57[114],stage1_56[150]}
   );
   gpc606_5 gpc2157 (
      {stage0_56[303], stage0_56[304], stage0_56[305], stage0_56[306], stage0_56[307], stage0_56[308]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[52],stage1_58[94],stage1_57[115],stage1_56[151]}
   );
   gpc606_5 gpc2158 (
      {stage0_56[309], stage0_56[310], stage0_56[311], stage0_56[312], stage0_56[313], stage0_56[314]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[53],stage1_58[95],stage1_57[116],stage1_56[152]}
   );
   gpc606_5 gpc2159 (
      {stage0_56[315], stage0_56[316], stage0_56[317], stage0_56[318], stage0_56[319], stage0_56[320]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[54],stage1_58[96],stage1_57[117],stage1_56[153]}
   );
   gpc615_5 gpc2160 (
      {stage0_56[321], stage0_56[322], stage0_56[323], stage0_56[324], stage0_56[325]},
      {stage0_57[264]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[55],stage1_58[97],stage1_57[118],stage1_56[154]}
   );
   gpc615_5 gpc2161 (
      {stage0_56[326], stage0_56[327], stage0_56[328], stage0_56[329], stage0_56[330]},
      {stage0_57[265]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[56],stage1_58[98],stage1_57[119],stage1_56[155]}
   );
   gpc615_5 gpc2162 (
      {stage0_56[331], stage0_56[332], stage0_56[333], stage0_56[334], stage0_56[335]},
      {stage0_57[266]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[57],stage1_58[99],stage1_57[120],stage1_56[156]}
   );
   gpc615_5 gpc2163 (
      {stage0_56[336], stage0_56[337], stage0_56[338], stage0_56[339], stage0_56[340]},
      {stage0_57[267]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[58],stage1_58[100],stage1_57[121],stage1_56[157]}
   );
   gpc615_5 gpc2164 (
      {stage0_56[341], stage0_56[342], stage0_56[343], stage0_56[344], stage0_56[345]},
      {stage0_57[268]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[59],stage1_58[101],stage1_57[122],stage1_56[158]}
   );
   gpc615_5 gpc2165 (
      {stage0_56[346], stage0_56[347], stage0_56[348], stage0_56[349], stage0_56[350]},
      {stage0_57[269]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[60],stage1_58[102],stage1_57[123],stage1_56[159]}
   );
   gpc615_5 gpc2166 (
      {stage0_56[351], stage0_56[352], stage0_56[353], stage0_56[354], stage0_56[355]},
      {stage0_57[270]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[61],stage1_58[103],stage1_57[124],stage1_56[160]}
   );
   gpc615_5 gpc2167 (
      {stage0_56[356], stage0_56[357], stage0_56[358], stage0_56[359], stage0_56[360]},
      {stage0_57[271]},
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage1_60[18],stage1_59[62],stage1_58[104],stage1_57[125],stage1_56[161]}
   );
   gpc615_5 gpc2168 (
      {stage0_56[361], stage0_56[362], stage0_56[363], stage0_56[364], stage0_56[365]},
      {stage0_57[272]},
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage1_60[19],stage1_59[63],stage1_58[105],stage1_57[126],stage1_56[162]}
   );
   gpc615_5 gpc2169 (
      {stage0_56[366], stage0_56[367], stage0_56[368], stage0_56[369], stage0_56[370]},
      {stage0_57[273]},
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage1_60[20],stage1_59[64],stage1_58[106],stage1_57[127],stage1_56[163]}
   );
   gpc615_5 gpc2170 (
      {stage0_56[371], stage0_56[372], stage0_56[373], stage0_56[374], stage0_56[375]},
      {stage0_57[274]},
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage1_60[21],stage1_59[65],stage1_58[107],stage1_57[128],stage1_56[164]}
   );
   gpc615_5 gpc2171 (
      {stage0_56[376], stage0_56[377], stage0_56[378], stage0_56[379], stage0_56[380]},
      {stage0_57[275]},
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage1_60[22],stage1_59[66],stage1_58[108],stage1_57[129],stage1_56[165]}
   );
   gpc615_5 gpc2172 (
      {stage0_56[381], stage0_56[382], stage0_56[383], stage0_56[384], stage0_56[385]},
      {stage0_57[276]},
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage1_60[23],stage1_59[67],stage1_58[109],stage1_57[130],stage1_56[166]}
   );
   gpc615_5 gpc2173 (
      {stage0_56[386], stage0_56[387], stage0_56[388], stage0_56[389], stage0_56[390]},
      {stage0_57[277]},
      {stage0_58[144], stage0_58[145], stage0_58[146], stage0_58[147], stage0_58[148], stage0_58[149]},
      {stage1_60[24],stage1_59[68],stage1_58[110],stage1_57[131],stage1_56[167]}
   );
   gpc615_5 gpc2174 (
      {stage0_56[391], stage0_56[392], stage0_56[393], stage0_56[394], stage0_56[395]},
      {stage0_57[278]},
      {stage0_58[150], stage0_58[151], stage0_58[152], stage0_58[153], stage0_58[154], stage0_58[155]},
      {stage1_60[25],stage1_59[69],stage1_58[111],stage1_57[132],stage1_56[168]}
   );
   gpc615_5 gpc2175 (
      {stage0_56[396], stage0_56[397], stage0_56[398], stage0_56[399], stage0_56[400]},
      {stage0_57[279]},
      {stage0_58[156], stage0_58[157], stage0_58[158], stage0_58[159], stage0_58[160], stage0_58[161]},
      {stage1_60[26],stage1_59[70],stage1_58[112],stage1_57[133],stage1_56[169]}
   );
   gpc615_5 gpc2176 (
      {stage0_56[401], stage0_56[402], stage0_56[403], stage0_56[404], stage0_56[405]},
      {stage0_57[280]},
      {stage0_58[162], stage0_58[163], stage0_58[164], stage0_58[165], stage0_58[166], stage0_58[167]},
      {stage1_60[27],stage1_59[71],stage1_58[113],stage1_57[134],stage1_56[170]}
   );
   gpc615_5 gpc2177 (
      {stage0_56[406], stage0_56[407], stage0_56[408], stage0_56[409], stage0_56[410]},
      {stage0_57[281]},
      {stage0_58[168], stage0_58[169], stage0_58[170], stage0_58[171], stage0_58[172], stage0_58[173]},
      {stage1_60[28],stage1_59[72],stage1_58[114],stage1_57[135],stage1_56[171]}
   );
   gpc615_5 gpc2178 (
      {stage0_56[411], stage0_56[412], stage0_56[413], stage0_56[414], stage0_56[415]},
      {stage0_57[282]},
      {stage0_58[174], stage0_58[175], stage0_58[176], stage0_58[177], stage0_58[178], stage0_58[179]},
      {stage1_60[29],stage1_59[73],stage1_58[115],stage1_57[136],stage1_56[172]}
   );
   gpc615_5 gpc2179 (
      {stage0_56[416], stage0_56[417], stage0_56[418], stage0_56[419], stage0_56[420]},
      {stage0_57[283]},
      {stage0_58[180], stage0_58[181], stage0_58[182], stage0_58[183], stage0_58[184], stage0_58[185]},
      {stage1_60[30],stage1_59[74],stage1_58[116],stage1_57[137],stage1_56[173]}
   );
   gpc615_5 gpc2180 (
      {stage0_56[421], stage0_56[422], stage0_56[423], stage0_56[424], stage0_56[425]},
      {stage0_57[284]},
      {stage0_58[186], stage0_58[187], stage0_58[188], stage0_58[189], stage0_58[190], stage0_58[191]},
      {stage1_60[31],stage1_59[75],stage1_58[117],stage1_57[138],stage1_56[174]}
   );
   gpc615_5 gpc2181 (
      {stage0_56[426], stage0_56[427], stage0_56[428], stage0_56[429], stage0_56[430]},
      {stage0_57[285]},
      {stage0_58[192], stage0_58[193], stage0_58[194], stage0_58[195], stage0_58[196], stage0_58[197]},
      {stage1_60[32],stage1_59[76],stage1_58[118],stage1_57[139],stage1_56[175]}
   );
   gpc615_5 gpc2182 (
      {stage0_56[431], stage0_56[432], stage0_56[433], stage0_56[434], stage0_56[435]},
      {stage0_57[286]},
      {stage0_58[198], stage0_58[199], stage0_58[200], stage0_58[201], stage0_58[202], stage0_58[203]},
      {stage1_60[33],stage1_59[77],stage1_58[119],stage1_57[140],stage1_56[176]}
   );
   gpc615_5 gpc2183 (
      {stage0_56[436], stage0_56[437], stage0_56[438], stage0_56[439], stage0_56[440]},
      {stage0_57[287]},
      {stage0_58[204], stage0_58[205], stage0_58[206], stage0_58[207], stage0_58[208], stage0_58[209]},
      {stage1_60[34],stage1_59[78],stage1_58[120],stage1_57[141],stage1_56[177]}
   );
   gpc615_5 gpc2184 (
      {stage0_56[441], stage0_56[442], stage0_56[443], stage0_56[444], stage0_56[445]},
      {stage0_57[288]},
      {stage0_58[210], stage0_58[211], stage0_58[212], stage0_58[213], stage0_58[214], stage0_58[215]},
      {stage1_60[35],stage1_59[79],stage1_58[121],stage1_57[142],stage1_56[178]}
   );
   gpc615_5 gpc2185 (
      {stage0_56[446], stage0_56[447], stage0_56[448], stage0_56[449], stage0_56[450]},
      {stage0_57[289]},
      {stage0_58[216], stage0_58[217], stage0_58[218], stage0_58[219], stage0_58[220], stage0_58[221]},
      {stage1_60[36],stage1_59[80],stage1_58[122],stage1_57[143],stage1_56[179]}
   );
   gpc615_5 gpc2186 (
      {stage0_56[451], stage0_56[452], stage0_56[453], stage0_56[454], stage0_56[455]},
      {stage0_57[290]},
      {stage0_58[222], stage0_58[223], stage0_58[224], stage0_58[225], stage0_58[226], stage0_58[227]},
      {stage1_60[37],stage1_59[81],stage1_58[123],stage1_57[144],stage1_56[180]}
   );
   gpc615_5 gpc2187 (
      {stage0_56[456], stage0_56[457], stage0_56[458], stage0_56[459], stage0_56[460]},
      {stage0_57[291]},
      {stage0_58[228], stage0_58[229], stage0_58[230], stage0_58[231], stage0_58[232], stage0_58[233]},
      {stage1_60[38],stage1_59[82],stage1_58[124],stage1_57[145],stage1_56[181]}
   );
   gpc615_5 gpc2188 (
      {stage0_56[461], stage0_56[462], stage0_56[463], stage0_56[464], stage0_56[465]},
      {stage0_57[292]},
      {stage0_58[234], stage0_58[235], stage0_58[236], stage0_58[237], stage0_58[238], stage0_58[239]},
      {stage1_60[39],stage1_59[83],stage1_58[125],stage1_57[146],stage1_56[182]}
   );
   gpc615_5 gpc2189 (
      {stage0_56[466], stage0_56[467], stage0_56[468], stage0_56[469], stage0_56[470]},
      {stage0_57[293]},
      {stage0_58[240], stage0_58[241], stage0_58[242], stage0_58[243], stage0_58[244], stage0_58[245]},
      {stage1_60[40],stage1_59[84],stage1_58[126],stage1_57[147],stage1_56[183]}
   );
   gpc615_5 gpc2190 (
      {stage0_56[471], stage0_56[472], stage0_56[473], stage0_56[474], stage0_56[475]},
      {stage0_57[294]},
      {stage0_58[246], stage0_58[247], stage0_58[248], stage0_58[249], stage0_58[250], stage0_58[251]},
      {stage1_60[41],stage1_59[85],stage1_58[127],stage1_57[148],stage1_56[184]}
   );
   gpc615_5 gpc2191 (
      {stage0_56[476], stage0_56[477], stage0_56[478], stage0_56[479], stage0_56[480]},
      {stage0_57[295]},
      {stage0_58[252], stage0_58[253], stage0_58[254], stage0_58[255], stage0_58[256], stage0_58[257]},
      {stage1_60[42],stage1_59[86],stage1_58[128],stage1_57[149],stage1_56[185]}
   );
   gpc615_5 gpc2192 (
      {stage0_56[481], stage0_56[482], stage0_56[483], stage0_56[484], stage0_56[485]},
      {stage0_57[296]},
      {stage0_58[258], stage0_58[259], stage0_58[260], stage0_58[261], stage0_58[262], stage0_58[263]},
      {stage1_60[43],stage1_59[87],stage1_58[129],stage1_57[150],stage1_56[186]}
   );
   gpc615_5 gpc2193 (
      {stage0_57[297], stage0_57[298], stage0_57[299], stage0_57[300], stage0_57[301]},
      {stage0_58[264]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[44],stage1_59[88],stage1_58[130],stage1_57[151]}
   );
   gpc615_5 gpc2194 (
      {stage0_57[302], stage0_57[303], stage0_57[304], stage0_57[305], stage0_57[306]},
      {stage0_58[265]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[45],stage1_59[89],stage1_58[131],stage1_57[152]}
   );
   gpc615_5 gpc2195 (
      {stage0_57[307], stage0_57[308], stage0_57[309], stage0_57[310], stage0_57[311]},
      {stage0_58[266]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[46],stage1_59[90],stage1_58[132],stage1_57[153]}
   );
   gpc615_5 gpc2196 (
      {stage0_57[312], stage0_57[313], stage0_57[314], stage0_57[315], stage0_57[316]},
      {stage0_58[267]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[47],stage1_59[91],stage1_58[133],stage1_57[154]}
   );
   gpc615_5 gpc2197 (
      {stage0_57[317], stage0_57[318], stage0_57[319], stage0_57[320], stage0_57[321]},
      {stage0_58[268]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[48],stage1_59[92],stage1_58[134],stage1_57[155]}
   );
   gpc615_5 gpc2198 (
      {stage0_57[322], stage0_57[323], stage0_57[324], stage0_57[325], stage0_57[326]},
      {stage0_58[269]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[49],stage1_59[93],stage1_58[135],stage1_57[156]}
   );
   gpc615_5 gpc2199 (
      {stage0_57[327], stage0_57[328], stage0_57[329], stage0_57[330], stage0_57[331]},
      {stage0_58[270]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[50],stage1_59[94],stage1_58[136],stage1_57[157]}
   );
   gpc615_5 gpc2200 (
      {stage0_57[332], stage0_57[333], stage0_57[334], stage0_57[335], stage0_57[336]},
      {stage0_58[271]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[51],stage1_59[95],stage1_58[137],stage1_57[158]}
   );
   gpc615_5 gpc2201 (
      {stage0_57[337], stage0_57[338], stage0_57[339], stage0_57[340], stage0_57[341]},
      {stage0_58[272]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[52],stage1_59[96],stage1_58[138],stage1_57[159]}
   );
   gpc615_5 gpc2202 (
      {stage0_57[342], stage0_57[343], stage0_57[344], stage0_57[345], stage0_57[346]},
      {stage0_58[273]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[53],stage1_59[97],stage1_58[139],stage1_57[160]}
   );
   gpc615_5 gpc2203 (
      {stage0_57[347], stage0_57[348], stage0_57[349], stage0_57[350], stage0_57[351]},
      {stage0_58[274]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[54],stage1_59[98],stage1_58[140],stage1_57[161]}
   );
   gpc615_5 gpc2204 (
      {stage0_57[352], stage0_57[353], stage0_57[354], stage0_57[355], stage0_57[356]},
      {stage0_58[275]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[55],stage1_59[99],stage1_58[141],stage1_57[162]}
   );
   gpc615_5 gpc2205 (
      {stage0_57[357], stage0_57[358], stage0_57[359], stage0_57[360], stage0_57[361]},
      {stage0_58[276]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[56],stage1_59[100],stage1_58[142],stage1_57[163]}
   );
   gpc615_5 gpc2206 (
      {stage0_57[362], stage0_57[363], stage0_57[364], stage0_57[365], stage0_57[366]},
      {stage0_58[277]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[57],stage1_59[101],stage1_58[143],stage1_57[164]}
   );
   gpc615_5 gpc2207 (
      {stage0_57[367], stage0_57[368], stage0_57[369], stage0_57[370], stage0_57[371]},
      {stage0_58[278]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[58],stage1_59[102],stage1_58[144],stage1_57[165]}
   );
   gpc615_5 gpc2208 (
      {stage0_57[372], stage0_57[373], stage0_57[374], stage0_57[375], stage0_57[376]},
      {stage0_58[279]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[59],stage1_59[103],stage1_58[145],stage1_57[166]}
   );
   gpc615_5 gpc2209 (
      {stage0_57[377], stage0_57[378], stage0_57[379], stage0_57[380], stage0_57[381]},
      {stage0_58[280]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[60],stage1_59[104],stage1_58[146],stage1_57[167]}
   );
   gpc615_5 gpc2210 (
      {stage0_57[382], stage0_57[383], stage0_57[384], stage0_57[385], stage0_57[386]},
      {stage0_58[281]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[61],stage1_59[105],stage1_58[147],stage1_57[168]}
   );
   gpc615_5 gpc2211 (
      {stage0_57[387], stage0_57[388], stage0_57[389], stage0_57[390], stage0_57[391]},
      {stage0_58[282]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[62],stage1_59[106],stage1_58[148],stage1_57[169]}
   );
   gpc615_5 gpc2212 (
      {stage0_57[392], stage0_57[393], stage0_57[394], stage0_57[395], stage0_57[396]},
      {stage0_58[283]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[63],stage1_59[107],stage1_58[149],stage1_57[170]}
   );
   gpc615_5 gpc2213 (
      {stage0_57[397], stage0_57[398], stage0_57[399], stage0_57[400], stage0_57[401]},
      {stage0_58[284]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[64],stage1_59[108],stage1_58[150],stage1_57[171]}
   );
   gpc615_5 gpc2214 (
      {stage0_57[402], stage0_57[403], stage0_57[404], stage0_57[405], stage0_57[406]},
      {stage0_58[285]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[65],stage1_59[109],stage1_58[151],stage1_57[172]}
   );
   gpc615_5 gpc2215 (
      {stage0_57[407], stage0_57[408], stage0_57[409], stage0_57[410], stage0_57[411]},
      {stage0_58[286]},
      {stage0_59[132], stage0_59[133], stage0_59[134], stage0_59[135], stage0_59[136], stage0_59[137]},
      {stage1_61[22],stage1_60[66],stage1_59[110],stage1_58[152],stage1_57[173]}
   );
   gpc615_5 gpc2216 (
      {stage0_57[412], stage0_57[413], stage0_57[414], stage0_57[415], stage0_57[416]},
      {stage0_58[287]},
      {stage0_59[138], stage0_59[139], stage0_59[140], stage0_59[141], stage0_59[142], stage0_59[143]},
      {stage1_61[23],stage1_60[67],stage1_59[111],stage1_58[153],stage1_57[174]}
   );
   gpc615_5 gpc2217 (
      {stage0_57[417], stage0_57[418], stage0_57[419], stage0_57[420], stage0_57[421]},
      {stage0_58[288]},
      {stage0_59[144], stage0_59[145], stage0_59[146], stage0_59[147], stage0_59[148], stage0_59[149]},
      {stage1_61[24],stage1_60[68],stage1_59[112],stage1_58[154],stage1_57[175]}
   );
   gpc615_5 gpc2218 (
      {stage0_57[422], stage0_57[423], stage0_57[424], stage0_57[425], stage0_57[426]},
      {stage0_58[289]},
      {stage0_59[150], stage0_59[151], stage0_59[152], stage0_59[153], stage0_59[154], stage0_59[155]},
      {stage1_61[25],stage1_60[69],stage1_59[113],stage1_58[155],stage1_57[176]}
   );
   gpc615_5 gpc2219 (
      {stage0_57[427], stage0_57[428], stage0_57[429], stage0_57[430], stage0_57[431]},
      {stage0_58[290]},
      {stage0_59[156], stage0_59[157], stage0_59[158], stage0_59[159], stage0_59[160], stage0_59[161]},
      {stage1_61[26],stage1_60[70],stage1_59[114],stage1_58[156],stage1_57[177]}
   );
   gpc615_5 gpc2220 (
      {stage0_57[432], stage0_57[433], stage0_57[434], stage0_57[435], stage0_57[436]},
      {stage0_58[291]},
      {stage0_59[162], stage0_59[163], stage0_59[164], stage0_59[165], stage0_59[166], stage0_59[167]},
      {stage1_61[27],stage1_60[71],stage1_59[115],stage1_58[157],stage1_57[178]}
   );
   gpc615_5 gpc2221 (
      {stage0_57[437], stage0_57[438], stage0_57[439], stage0_57[440], stage0_57[441]},
      {stage0_58[292]},
      {stage0_59[168], stage0_59[169], stage0_59[170], stage0_59[171], stage0_59[172], stage0_59[173]},
      {stage1_61[28],stage1_60[72],stage1_59[116],stage1_58[158],stage1_57[179]}
   );
   gpc615_5 gpc2222 (
      {stage0_57[442], stage0_57[443], stage0_57[444], stage0_57[445], stage0_57[446]},
      {stage0_58[293]},
      {stage0_59[174], stage0_59[175], stage0_59[176], stage0_59[177], stage0_59[178], stage0_59[179]},
      {stage1_61[29],stage1_60[73],stage1_59[117],stage1_58[159],stage1_57[180]}
   );
   gpc615_5 gpc2223 (
      {stage0_57[447], stage0_57[448], stage0_57[449], stage0_57[450], stage0_57[451]},
      {stage0_58[294]},
      {stage0_59[180], stage0_59[181], stage0_59[182], stage0_59[183], stage0_59[184], stage0_59[185]},
      {stage1_61[30],stage1_60[74],stage1_59[118],stage1_58[160],stage1_57[181]}
   );
   gpc615_5 gpc2224 (
      {stage0_57[452], stage0_57[453], stage0_57[454], stage0_57[455], stage0_57[456]},
      {stage0_58[295]},
      {stage0_59[186], stage0_59[187], stage0_59[188], stage0_59[189], stage0_59[190], stage0_59[191]},
      {stage1_61[31],stage1_60[75],stage1_59[119],stage1_58[161],stage1_57[182]}
   );
   gpc615_5 gpc2225 (
      {stage0_57[457], stage0_57[458], stage0_57[459], stage0_57[460], stage0_57[461]},
      {stage0_58[296]},
      {stage0_59[192], stage0_59[193], stage0_59[194], stage0_59[195], stage0_59[196], stage0_59[197]},
      {stage1_61[32],stage1_60[76],stage1_59[120],stage1_58[162],stage1_57[183]}
   );
   gpc615_5 gpc2226 (
      {stage0_57[462], stage0_57[463], stage0_57[464], stage0_57[465], stage0_57[466]},
      {stage0_58[297]},
      {stage0_59[198], stage0_59[199], stage0_59[200], stage0_59[201], stage0_59[202], stage0_59[203]},
      {stage1_61[33],stage1_60[77],stage1_59[121],stage1_58[163],stage1_57[184]}
   );
   gpc615_5 gpc2227 (
      {stage0_57[467], stage0_57[468], stage0_57[469], stage0_57[470], stage0_57[471]},
      {stage0_58[298]},
      {stage0_59[204], stage0_59[205], stage0_59[206], stage0_59[207], stage0_59[208], stage0_59[209]},
      {stage1_61[34],stage1_60[78],stage1_59[122],stage1_58[164],stage1_57[185]}
   );
   gpc615_5 gpc2228 (
      {stage0_57[472], stage0_57[473], stage0_57[474], stage0_57[475], stage0_57[476]},
      {stage0_58[299]},
      {stage0_59[210], stage0_59[211], stage0_59[212], stage0_59[213], stage0_59[214], stage0_59[215]},
      {stage1_61[35],stage1_60[79],stage1_59[123],stage1_58[165],stage1_57[186]}
   );
   gpc615_5 gpc2229 (
      {stage0_57[477], stage0_57[478], stage0_57[479], stage0_57[480], stage0_57[481]},
      {stage0_58[300]},
      {stage0_59[216], stage0_59[217], stage0_59[218], stage0_59[219], stage0_59[220], stage0_59[221]},
      {stage1_61[36],stage1_60[80],stage1_59[124],stage1_58[166],stage1_57[187]}
   );
   gpc615_5 gpc2230 (
      {stage0_57[482], stage0_57[483], stage0_57[484], stage0_57[485], 1'b0},
      {stage0_58[301]},
      {stage0_59[222], stage0_59[223], stage0_59[224], stage0_59[225], stage0_59[226], stage0_59[227]},
      {stage1_61[37],stage1_60[81],stage1_59[125],stage1_58[167],stage1_57[188]}
   );
   gpc7_3 gpc2231 (
      {stage0_58[302], stage0_58[303], stage0_58[304], stage0_58[305], stage0_58[306], stage0_58[307], stage0_58[308]},
      {stage1_60[82],stage1_59[126],stage1_58[168]}
   );
   gpc7_3 gpc2232 (
      {stage0_58[309], stage0_58[310], stage0_58[311], stage0_58[312], stage0_58[313], stage0_58[314], stage0_58[315]},
      {stage1_60[83],stage1_59[127],stage1_58[169]}
   );
   gpc7_3 gpc2233 (
      {stage0_58[316], stage0_58[317], stage0_58[318], stage0_58[319], stage0_58[320], stage0_58[321], stage0_58[322]},
      {stage1_60[84],stage1_59[128],stage1_58[170]}
   );
   gpc7_3 gpc2234 (
      {stage0_58[323], stage0_58[324], stage0_58[325], stage0_58[326], stage0_58[327], stage0_58[328], stage0_58[329]},
      {stage1_60[85],stage1_59[129],stage1_58[171]}
   );
   gpc7_3 gpc2235 (
      {stage0_58[330], stage0_58[331], stage0_58[332], stage0_58[333], stage0_58[334], stage0_58[335], stage0_58[336]},
      {stage1_60[86],stage1_59[130],stage1_58[172]}
   );
   gpc7_3 gpc2236 (
      {stage0_58[337], stage0_58[338], stage0_58[339], stage0_58[340], stage0_58[341], stage0_58[342], stage0_58[343]},
      {stage1_60[87],stage1_59[131],stage1_58[173]}
   );
   gpc606_5 gpc2237 (
      {stage0_58[344], stage0_58[345], stage0_58[346], stage0_58[347], stage0_58[348], stage0_58[349]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[38],stage1_60[88],stage1_59[132],stage1_58[174]}
   );
   gpc606_5 gpc2238 (
      {stage0_58[350], stage0_58[351], stage0_58[352], stage0_58[353], stage0_58[354], stage0_58[355]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[39],stage1_60[89],stage1_59[133],stage1_58[175]}
   );
   gpc606_5 gpc2239 (
      {stage0_58[356], stage0_58[357], stage0_58[358], stage0_58[359], stage0_58[360], stage0_58[361]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[40],stage1_60[90],stage1_59[134],stage1_58[176]}
   );
   gpc606_5 gpc2240 (
      {stage0_58[362], stage0_58[363], stage0_58[364], stage0_58[365], stage0_58[366], stage0_58[367]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[41],stage1_60[91],stage1_59[135],stage1_58[177]}
   );
   gpc606_5 gpc2241 (
      {stage0_58[368], stage0_58[369], stage0_58[370], stage0_58[371], stage0_58[372], stage0_58[373]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[42],stage1_60[92],stage1_59[136],stage1_58[178]}
   );
   gpc606_5 gpc2242 (
      {stage0_58[374], stage0_58[375], stage0_58[376], stage0_58[377], stage0_58[378], stage0_58[379]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[43],stage1_60[93],stage1_59[137],stage1_58[179]}
   );
   gpc606_5 gpc2243 (
      {stage0_58[380], stage0_58[381], stage0_58[382], stage0_58[383], stage0_58[384], stage0_58[385]},
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage1_62[6],stage1_61[44],stage1_60[94],stage1_59[138],stage1_58[180]}
   );
   gpc606_5 gpc2244 (
      {stage0_58[386], stage0_58[387], stage0_58[388], stage0_58[389], stage0_58[390], stage0_58[391]},
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage1_62[7],stage1_61[45],stage1_60[95],stage1_59[139],stage1_58[181]}
   );
   gpc606_5 gpc2245 (
      {stage0_58[392], stage0_58[393], stage0_58[394], stage0_58[395], stage0_58[396], stage0_58[397]},
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage1_62[8],stage1_61[46],stage1_60[96],stage1_59[140],stage1_58[182]}
   );
   gpc606_5 gpc2246 (
      {stage0_58[398], stage0_58[399], stage0_58[400], stage0_58[401], stage0_58[402], stage0_58[403]},
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage1_62[9],stage1_61[47],stage1_60[97],stage1_59[141],stage1_58[183]}
   );
   gpc606_5 gpc2247 (
      {stage0_58[404], stage0_58[405], stage0_58[406], stage0_58[407], stage0_58[408], stage0_58[409]},
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage1_62[10],stage1_61[48],stage1_60[98],stage1_59[142],stage1_58[184]}
   );
   gpc606_5 gpc2248 (
      {stage0_58[410], stage0_58[411], stage0_58[412], stage0_58[413], stage0_58[414], stage0_58[415]},
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage1_62[11],stage1_61[49],stage1_60[99],stage1_59[143],stage1_58[185]}
   );
   gpc606_5 gpc2249 (
      {stage0_58[416], stage0_58[417], stage0_58[418], stage0_58[419], stage0_58[420], stage0_58[421]},
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage1_62[12],stage1_61[50],stage1_60[100],stage1_59[144],stage1_58[186]}
   );
   gpc606_5 gpc2250 (
      {stage0_58[422], stage0_58[423], stage0_58[424], stage0_58[425], stage0_58[426], stage0_58[427]},
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage1_62[13],stage1_61[51],stage1_60[101],stage1_59[145],stage1_58[187]}
   );
   gpc606_5 gpc2251 (
      {stage0_58[428], stage0_58[429], stage0_58[430], stage0_58[431], stage0_58[432], stage0_58[433]},
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage1_62[14],stage1_61[52],stage1_60[102],stage1_59[146],stage1_58[188]}
   );
   gpc606_5 gpc2252 (
      {stage0_58[434], stage0_58[435], stage0_58[436], stage0_58[437], stage0_58[438], stage0_58[439]},
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage1_62[15],stage1_61[53],stage1_60[103],stage1_59[147],stage1_58[189]}
   );
   gpc615_5 gpc2253 (
      {stage0_58[440], stage0_58[441], stage0_58[442], stage0_58[443], stage0_58[444]},
      {stage0_59[228]},
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage1_62[16],stage1_61[54],stage1_60[104],stage1_59[148],stage1_58[190]}
   );
   gpc615_5 gpc2254 (
      {stage0_58[445], stage0_58[446], stage0_58[447], stage0_58[448], stage0_58[449]},
      {stage0_59[229]},
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage1_62[17],stage1_61[55],stage1_60[105],stage1_59[149],stage1_58[191]}
   );
   gpc615_5 gpc2255 (
      {stage0_58[450], stage0_58[451], stage0_58[452], stage0_58[453], stage0_58[454]},
      {stage0_59[230]},
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage1_62[18],stage1_61[56],stage1_60[106],stage1_59[150],stage1_58[192]}
   );
   gpc615_5 gpc2256 (
      {stage0_58[455], stage0_58[456], stage0_58[457], stage0_58[458], stage0_58[459]},
      {stage0_59[231]},
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage1_62[19],stage1_61[57],stage1_60[107],stage1_59[151],stage1_58[193]}
   );
   gpc117_4 gpc2257 (
      {stage0_59[232], stage0_59[233], stage0_59[234], stage0_59[235], stage0_59[236], stage0_59[237], stage0_59[238]},
      {stage0_60[120]},
      {stage0_61[0]},
      {stage1_62[20],stage1_61[58],stage1_60[108],stage1_59[152]}
   );
   gpc117_4 gpc2258 (
      {stage0_59[239], stage0_59[240], stage0_59[241], stage0_59[242], stage0_59[243], stage0_59[244], stage0_59[245]},
      {stage0_60[121]},
      {stage0_61[1]},
      {stage1_62[21],stage1_61[59],stage1_60[109],stage1_59[153]}
   );
   gpc117_4 gpc2259 (
      {stage0_59[246], stage0_59[247], stage0_59[248], stage0_59[249], stage0_59[250], stage0_59[251], stage0_59[252]},
      {stage0_60[122]},
      {stage0_61[2]},
      {stage1_62[22],stage1_61[60],stage1_60[110],stage1_59[154]}
   );
   gpc117_4 gpc2260 (
      {stage0_59[253], stage0_59[254], stage0_59[255], stage0_59[256], stage0_59[257], stage0_59[258], stage0_59[259]},
      {stage0_60[123]},
      {stage0_61[3]},
      {stage1_62[23],stage1_61[61],stage1_60[111],stage1_59[155]}
   );
   gpc117_4 gpc2261 (
      {stage0_59[260], stage0_59[261], stage0_59[262], stage0_59[263], stage0_59[264], stage0_59[265], stage0_59[266]},
      {stage0_60[124]},
      {stage0_61[4]},
      {stage1_62[24],stage1_61[62],stage1_60[112],stage1_59[156]}
   );
   gpc117_4 gpc2262 (
      {stage0_59[267], stage0_59[268], stage0_59[269], stage0_59[270], stage0_59[271], stage0_59[272], stage0_59[273]},
      {stage0_60[125]},
      {stage0_61[5]},
      {stage1_62[25],stage1_61[63],stage1_60[113],stage1_59[157]}
   );
   gpc117_4 gpc2263 (
      {stage0_59[274], stage0_59[275], stage0_59[276], stage0_59[277], stage0_59[278], stage0_59[279], stage0_59[280]},
      {stage0_60[126]},
      {stage0_61[6]},
      {stage1_62[26],stage1_61[64],stage1_60[114],stage1_59[158]}
   );
   gpc117_4 gpc2264 (
      {stage0_59[281], stage0_59[282], stage0_59[283], stage0_59[284], stage0_59[285], stage0_59[286], stage0_59[287]},
      {stage0_60[127]},
      {stage0_61[7]},
      {stage1_62[27],stage1_61[65],stage1_60[115],stage1_59[159]}
   );
   gpc117_4 gpc2265 (
      {stage0_59[288], stage0_59[289], stage0_59[290], stage0_59[291], stage0_59[292], stage0_59[293], stage0_59[294]},
      {stage0_60[128]},
      {stage0_61[8]},
      {stage1_62[28],stage1_61[66],stage1_60[116],stage1_59[160]}
   );
   gpc117_4 gpc2266 (
      {stage0_59[295], stage0_59[296], stage0_59[297], stage0_59[298], stage0_59[299], stage0_59[300], stage0_59[301]},
      {stage0_60[129]},
      {stage0_61[9]},
      {stage1_62[29],stage1_61[67],stage1_60[117],stage1_59[161]}
   );
   gpc117_4 gpc2267 (
      {stage0_59[302], stage0_59[303], stage0_59[304], stage0_59[305], stage0_59[306], stage0_59[307], stage0_59[308]},
      {stage0_60[130]},
      {stage0_61[10]},
      {stage1_62[30],stage1_61[68],stage1_60[118],stage1_59[162]}
   );
   gpc117_4 gpc2268 (
      {stage0_59[309], stage0_59[310], stage0_59[311], stage0_59[312], stage0_59[313], stage0_59[314], stage0_59[315]},
      {stage0_60[131]},
      {stage0_61[11]},
      {stage1_62[31],stage1_61[69],stage1_60[119],stage1_59[163]}
   );
   gpc117_4 gpc2269 (
      {stage0_59[316], stage0_59[317], stage0_59[318], stage0_59[319], stage0_59[320], stage0_59[321], stage0_59[322]},
      {stage0_60[132]},
      {stage0_61[12]},
      {stage1_62[32],stage1_61[70],stage1_60[120],stage1_59[164]}
   );
   gpc117_4 gpc2270 (
      {stage0_59[323], stage0_59[324], stage0_59[325], stage0_59[326], stage0_59[327], stage0_59[328], stage0_59[329]},
      {stage0_60[133]},
      {stage0_61[13]},
      {stage1_62[33],stage1_61[71],stage1_60[121],stage1_59[165]}
   );
   gpc117_4 gpc2271 (
      {stage0_59[330], stage0_59[331], stage0_59[332], stage0_59[333], stage0_59[334], stage0_59[335], stage0_59[336]},
      {stage0_60[134]},
      {stage0_61[14]},
      {stage1_62[34],stage1_61[72],stage1_60[122],stage1_59[166]}
   );
   gpc606_5 gpc2272 (
      {stage0_59[337], stage0_59[338], stage0_59[339], stage0_59[340], stage0_59[341], stage0_59[342]},
      {stage0_61[15], stage0_61[16], stage0_61[17], stage0_61[18], stage0_61[19], stage0_61[20]},
      {stage1_63[0],stage1_62[35],stage1_61[73],stage1_60[123],stage1_59[167]}
   );
   gpc606_5 gpc2273 (
      {stage0_59[343], stage0_59[344], stage0_59[345], stage0_59[346], stage0_59[347], stage0_59[348]},
      {stage0_61[21], stage0_61[22], stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26]},
      {stage1_63[1],stage1_62[36],stage1_61[74],stage1_60[124],stage1_59[168]}
   );
   gpc606_5 gpc2274 (
      {stage0_59[349], stage0_59[350], stage0_59[351], stage0_59[352], stage0_59[353], stage0_59[354]},
      {stage0_61[27], stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31], stage0_61[32]},
      {stage1_63[2],stage1_62[37],stage1_61[75],stage1_60[125],stage1_59[169]}
   );
   gpc606_5 gpc2275 (
      {stage0_59[355], stage0_59[356], stage0_59[357], stage0_59[358], stage0_59[359], stage0_59[360]},
      {stage0_61[33], stage0_61[34], stage0_61[35], stage0_61[36], stage0_61[37], stage0_61[38]},
      {stage1_63[3],stage1_62[38],stage1_61[76],stage1_60[126],stage1_59[170]}
   );
   gpc606_5 gpc2276 (
      {stage0_59[361], stage0_59[362], stage0_59[363], stage0_59[364], stage0_59[365], stage0_59[366]},
      {stage0_61[39], stage0_61[40], stage0_61[41], stage0_61[42], stage0_61[43], stage0_61[44]},
      {stage1_63[4],stage1_62[39],stage1_61[77],stage1_60[127],stage1_59[171]}
   );
   gpc606_5 gpc2277 (
      {stage0_59[367], stage0_59[368], stage0_59[369], stage0_59[370], stage0_59[371], stage0_59[372]},
      {stage0_61[45], stage0_61[46], stage0_61[47], stage0_61[48], stage0_61[49], stage0_61[50]},
      {stage1_63[5],stage1_62[40],stage1_61[78],stage1_60[128],stage1_59[172]}
   );
   gpc606_5 gpc2278 (
      {stage0_59[373], stage0_59[374], stage0_59[375], stage0_59[376], stage0_59[377], stage0_59[378]},
      {stage0_61[51], stage0_61[52], stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56]},
      {stage1_63[6],stage1_62[41],stage1_61[79],stage1_60[129],stage1_59[173]}
   );
   gpc606_5 gpc2279 (
      {stage0_59[379], stage0_59[380], stage0_59[381], stage0_59[382], stage0_59[383], stage0_59[384]},
      {stage0_61[57], stage0_61[58], stage0_61[59], stage0_61[60], stage0_61[61], stage0_61[62]},
      {stage1_63[7],stage1_62[42],stage1_61[80],stage1_60[130],stage1_59[174]}
   );
   gpc606_5 gpc2280 (
      {stage0_59[385], stage0_59[386], stage0_59[387], stage0_59[388], stage0_59[389], stage0_59[390]},
      {stage0_61[63], stage0_61[64], stage0_61[65], stage0_61[66], stage0_61[67], stage0_61[68]},
      {stage1_63[8],stage1_62[43],stage1_61[81],stage1_60[131],stage1_59[175]}
   );
   gpc606_5 gpc2281 (
      {stage0_59[391], stage0_59[392], stage0_59[393], stage0_59[394], stage0_59[395], stage0_59[396]},
      {stage0_61[69], stage0_61[70], stage0_61[71], stage0_61[72], stage0_61[73], stage0_61[74]},
      {stage1_63[9],stage1_62[44],stage1_61[82],stage1_60[132],stage1_59[176]}
   );
   gpc606_5 gpc2282 (
      {stage0_59[397], stage0_59[398], stage0_59[399], stage0_59[400], stage0_59[401], stage0_59[402]},
      {stage0_61[75], stage0_61[76], stage0_61[77], stage0_61[78], stage0_61[79], stage0_61[80]},
      {stage1_63[10],stage1_62[45],stage1_61[83],stage1_60[133],stage1_59[177]}
   );
   gpc606_5 gpc2283 (
      {stage0_59[403], stage0_59[404], stage0_59[405], stage0_59[406], stage0_59[407], stage0_59[408]},
      {stage0_61[81], stage0_61[82], stage0_61[83], stage0_61[84], stage0_61[85], stage0_61[86]},
      {stage1_63[11],stage1_62[46],stage1_61[84],stage1_60[134],stage1_59[178]}
   );
   gpc606_5 gpc2284 (
      {stage0_59[409], stage0_59[410], stage0_59[411], stage0_59[412], stage0_59[413], stage0_59[414]},
      {stage0_61[87], stage0_61[88], stage0_61[89], stage0_61[90], stage0_61[91], stage0_61[92]},
      {stage1_63[12],stage1_62[47],stage1_61[85],stage1_60[135],stage1_59[179]}
   );
   gpc606_5 gpc2285 (
      {stage0_59[415], stage0_59[416], stage0_59[417], stage0_59[418], stage0_59[419], stage0_59[420]},
      {stage0_61[93], stage0_61[94], stage0_61[95], stage0_61[96], stage0_61[97], stage0_61[98]},
      {stage1_63[13],stage1_62[48],stage1_61[86],stage1_60[136],stage1_59[180]}
   );
   gpc606_5 gpc2286 (
      {stage0_59[421], stage0_59[422], stage0_59[423], stage0_59[424], stage0_59[425], stage0_59[426]},
      {stage0_61[99], stage0_61[100], stage0_61[101], stage0_61[102], stage0_61[103], stage0_61[104]},
      {stage1_63[14],stage1_62[49],stage1_61[87],stage1_60[137],stage1_59[181]}
   );
   gpc606_5 gpc2287 (
      {stage0_59[427], stage0_59[428], stage0_59[429], stage0_59[430], stage0_59[431], stage0_59[432]},
      {stage0_61[105], stage0_61[106], stage0_61[107], stage0_61[108], stage0_61[109], stage0_61[110]},
      {stage1_63[15],stage1_62[50],stage1_61[88],stage1_60[138],stage1_59[182]}
   );
   gpc606_5 gpc2288 (
      {stage0_59[433], stage0_59[434], stage0_59[435], stage0_59[436], stage0_59[437], stage0_59[438]},
      {stage0_61[111], stage0_61[112], stage0_61[113], stage0_61[114], stage0_61[115], stage0_61[116]},
      {stage1_63[16],stage1_62[51],stage1_61[89],stage1_60[139],stage1_59[183]}
   );
   gpc606_5 gpc2289 (
      {stage0_59[439], stage0_59[440], stage0_59[441], stage0_59[442], stage0_59[443], stage0_59[444]},
      {stage0_61[117], stage0_61[118], stage0_61[119], stage0_61[120], stage0_61[121], stage0_61[122]},
      {stage1_63[17],stage1_62[52],stage1_61[90],stage1_60[140],stage1_59[184]}
   );
   gpc606_5 gpc2290 (
      {stage0_59[445], stage0_59[446], stage0_59[447], stage0_59[448], stage0_59[449], stage0_59[450]},
      {stage0_61[123], stage0_61[124], stage0_61[125], stage0_61[126], stage0_61[127], stage0_61[128]},
      {stage1_63[18],stage1_62[53],stage1_61[91],stage1_60[141],stage1_59[185]}
   );
   gpc606_5 gpc2291 (
      {stage0_59[451], stage0_59[452], stage0_59[453], stage0_59[454], stage0_59[455], stage0_59[456]},
      {stage0_61[129], stage0_61[130], stage0_61[131], stage0_61[132], stage0_61[133], stage0_61[134]},
      {stage1_63[19],stage1_62[54],stage1_61[92],stage1_60[142],stage1_59[186]}
   );
   gpc606_5 gpc2292 (
      {stage0_59[457], stage0_59[458], stage0_59[459], stage0_59[460], stage0_59[461], stage0_59[462]},
      {stage0_61[135], stage0_61[136], stage0_61[137], stage0_61[138], stage0_61[139], stage0_61[140]},
      {stage1_63[20],stage1_62[55],stage1_61[93],stage1_60[143],stage1_59[187]}
   );
   gpc606_5 gpc2293 (
      {stage0_59[463], stage0_59[464], stage0_59[465], stage0_59[466], stage0_59[467], stage0_59[468]},
      {stage0_61[141], stage0_61[142], stage0_61[143], stage0_61[144], stage0_61[145], stage0_61[146]},
      {stage1_63[21],stage1_62[56],stage1_61[94],stage1_60[144],stage1_59[188]}
   );
   gpc606_5 gpc2294 (
      {stage0_60[135], stage0_60[136], stage0_60[137], stage0_60[138], stage0_60[139], stage0_60[140]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[22],stage1_62[57],stage1_61[95],stage1_60[145]}
   );
   gpc615_5 gpc2295 (
      {stage0_60[141], stage0_60[142], stage0_60[143], stage0_60[144], stage0_60[145]},
      {stage0_61[147]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[23],stage1_62[58],stage1_61[96],stage1_60[146]}
   );
   gpc615_5 gpc2296 (
      {stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149], stage0_60[150]},
      {stage0_61[148]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[24],stage1_62[59],stage1_61[97],stage1_60[147]}
   );
   gpc615_5 gpc2297 (
      {stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155]},
      {stage0_61[149]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[25],stage1_62[60],stage1_61[98],stage1_60[148]}
   );
   gpc615_5 gpc2298 (
      {stage0_60[156], stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160]},
      {stage0_61[150]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[26],stage1_62[61],stage1_61[99],stage1_60[149]}
   );
   gpc615_5 gpc2299 (
      {stage0_60[161], stage0_60[162], stage0_60[163], stage0_60[164], stage0_60[165]},
      {stage0_61[151]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[27],stage1_62[62],stage1_61[100],stage1_60[150]}
   );
   gpc615_5 gpc2300 (
      {stage0_60[166], stage0_60[167], stage0_60[168], stage0_60[169], stage0_60[170]},
      {stage0_61[152]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[28],stage1_62[63],stage1_61[101],stage1_60[151]}
   );
   gpc615_5 gpc2301 (
      {stage0_60[171], stage0_60[172], stage0_60[173], stage0_60[174], stage0_60[175]},
      {stage0_61[153]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[29],stage1_62[64],stage1_61[102],stage1_60[152]}
   );
   gpc615_5 gpc2302 (
      {stage0_60[176], stage0_60[177], stage0_60[178], stage0_60[179], stage0_60[180]},
      {stage0_61[154]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[30],stage1_62[65],stage1_61[103],stage1_60[153]}
   );
   gpc615_5 gpc2303 (
      {stage0_60[181], stage0_60[182], stage0_60[183], stage0_60[184], stage0_60[185]},
      {stage0_61[155]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[31],stage1_62[66],stage1_61[104],stage1_60[154]}
   );
   gpc615_5 gpc2304 (
      {stage0_60[186], stage0_60[187], stage0_60[188], stage0_60[189], stage0_60[190]},
      {stage0_61[156]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[32],stage1_62[67],stage1_61[105],stage1_60[155]}
   );
   gpc615_5 gpc2305 (
      {stage0_60[191], stage0_60[192], stage0_60[193], stage0_60[194], stage0_60[195]},
      {stage0_61[157]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[33],stage1_62[68],stage1_61[106],stage1_60[156]}
   );
   gpc615_5 gpc2306 (
      {stage0_60[196], stage0_60[197], stage0_60[198], stage0_60[199], stage0_60[200]},
      {stage0_61[158]},
      {stage0_62[72], stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77]},
      {stage1_64[12],stage1_63[34],stage1_62[69],stage1_61[107],stage1_60[157]}
   );
   gpc615_5 gpc2307 (
      {stage0_60[201], stage0_60[202], stage0_60[203], stage0_60[204], stage0_60[205]},
      {stage0_61[159]},
      {stage0_62[78], stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83]},
      {stage1_64[13],stage1_63[35],stage1_62[70],stage1_61[108],stage1_60[158]}
   );
   gpc615_5 gpc2308 (
      {stage0_60[206], stage0_60[207], stage0_60[208], stage0_60[209], stage0_60[210]},
      {stage0_61[160]},
      {stage0_62[84], stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89]},
      {stage1_64[14],stage1_63[36],stage1_62[71],stage1_61[109],stage1_60[159]}
   );
   gpc615_5 gpc2309 (
      {stage0_60[211], stage0_60[212], stage0_60[213], stage0_60[214], stage0_60[215]},
      {stage0_61[161]},
      {stage0_62[90], stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95]},
      {stage1_64[15],stage1_63[37],stage1_62[72],stage1_61[110],stage1_60[160]}
   );
   gpc615_5 gpc2310 (
      {stage0_60[216], stage0_60[217], stage0_60[218], stage0_60[219], stage0_60[220]},
      {stage0_61[162]},
      {stage0_62[96], stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101]},
      {stage1_64[16],stage1_63[38],stage1_62[73],stage1_61[111],stage1_60[161]}
   );
   gpc615_5 gpc2311 (
      {stage0_60[221], stage0_60[222], stage0_60[223], stage0_60[224], stage0_60[225]},
      {stage0_61[163]},
      {stage0_62[102], stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107]},
      {stage1_64[17],stage1_63[39],stage1_62[74],stage1_61[112],stage1_60[162]}
   );
   gpc615_5 gpc2312 (
      {stage0_60[226], stage0_60[227], stage0_60[228], stage0_60[229], stage0_60[230]},
      {stage0_61[164]},
      {stage0_62[108], stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113]},
      {stage1_64[18],stage1_63[40],stage1_62[75],stage1_61[113],stage1_60[163]}
   );
   gpc615_5 gpc2313 (
      {stage0_60[231], stage0_60[232], stage0_60[233], stage0_60[234], stage0_60[235]},
      {stage0_61[165]},
      {stage0_62[114], stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119]},
      {stage1_64[19],stage1_63[41],stage1_62[76],stage1_61[114],stage1_60[164]}
   );
   gpc615_5 gpc2314 (
      {stage0_60[236], stage0_60[237], stage0_60[238], stage0_60[239], stage0_60[240]},
      {stage0_61[166]},
      {stage0_62[120], stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125]},
      {stage1_64[20],stage1_63[42],stage1_62[77],stage1_61[115],stage1_60[165]}
   );
   gpc615_5 gpc2315 (
      {stage0_60[241], stage0_60[242], stage0_60[243], stage0_60[244], stage0_60[245]},
      {stage0_61[167]},
      {stage0_62[126], stage0_62[127], stage0_62[128], stage0_62[129], stage0_62[130], stage0_62[131]},
      {stage1_64[21],stage1_63[43],stage1_62[78],stage1_61[116],stage1_60[166]}
   );
   gpc615_5 gpc2316 (
      {stage0_60[246], stage0_60[247], stage0_60[248], stage0_60[249], stage0_60[250]},
      {stage0_61[168]},
      {stage0_62[132], stage0_62[133], stage0_62[134], stage0_62[135], stage0_62[136], stage0_62[137]},
      {stage1_64[22],stage1_63[44],stage1_62[79],stage1_61[117],stage1_60[167]}
   );
   gpc615_5 gpc2317 (
      {stage0_60[251], stage0_60[252], stage0_60[253], stage0_60[254], stage0_60[255]},
      {stage0_61[169]},
      {stage0_62[138], stage0_62[139], stage0_62[140], stage0_62[141], stage0_62[142], stage0_62[143]},
      {stage1_64[23],stage1_63[45],stage1_62[80],stage1_61[118],stage1_60[168]}
   );
   gpc615_5 gpc2318 (
      {stage0_60[256], stage0_60[257], stage0_60[258], stage0_60[259], stage0_60[260]},
      {stage0_61[170]},
      {stage0_62[144], stage0_62[145], stage0_62[146], stage0_62[147], stage0_62[148], stage0_62[149]},
      {stage1_64[24],stage1_63[46],stage1_62[81],stage1_61[119],stage1_60[169]}
   );
   gpc615_5 gpc2319 (
      {stage0_60[261], stage0_60[262], stage0_60[263], stage0_60[264], stage0_60[265]},
      {stage0_61[171]},
      {stage0_62[150], stage0_62[151], stage0_62[152], stage0_62[153], stage0_62[154], stage0_62[155]},
      {stage1_64[25],stage1_63[47],stage1_62[82],stage1_61[120],stage1_60[170]}
   );
   gpc615_5 gpc2320 (
      {stage0_60[266], stage0_60[267], stage0_60[268], stage0_60[269], stage0_60[270]},
      {stage0_61[172]},
      {stage0_62[156], stage0_62[157], stage0_62[158], stage0_62[159], stage0_62[160], stage0_62[161]},
      {stage1_64[26],stage1_63[48],stage1_62[83],stage1_61[121],stage1_60[171]}
   );
   gpc615_5 gpc2321 (
      {stage0_60[271], stage0_60[272], stage0_60[273], stage0_60[274], stage0_60[275]},
      {stage0_61[173]},
      {stage0_62[162], stage0_62[163], stage0_62[164], stage0_62[165], stage0_62[166], stage0_62[167]},
      {stage1_64[27],stage1_63[49],stage1_62[84],stage1_61[122],stage1_60[172]}
   );
   gpc615_5 gpc2322 (
      {stage0_60[276], stage0_60[277], stage0_60[278], stage0_60[279], stage0_60[280]},
      {stage0_61[174]},
      {stage0_62[168], stage0_62[169], stage0_62[170], stage0_62[171], stage0_62[172], stage0_62[173]},
      {stage1_64[28],stage1_63[50],stage1_62[85],stage1_61[123],stage1_60[173]}
   );
   gpc615_5 gpc2323 (
      {stage0_60[281], stage0_60[282], stage0_60[283], stage0_60[284], stage0_60[285]},
      {stage0_61[175]},
      {stage0_62[174], stage0_62[175], stage0_62[176], stage0_62[177], stage0_62[178], stage0_62[179]},
      {stage1_64[29],stage1_63[51],stage1_62[86],stage1_61[124],stage1_60[174]}
   );
   gpc615_5 gpc2324 (
      {stage0_60[286], stage0_60[287], stage0_60[288], stage0_60[289], stage0_60[290]},
      {stage0_61[176]},
      {stage0_62[180], stage0_62[181], stage0_62[182], stage0_62[183], stage0_62[184], stage0_62[185]},
      {stage1_64[30],stage1_63[52],stage1_62[87],stage1_61[125],stage1_60[175]}
   );
   gpc615_5 gpc2325 (
      {stage0_60[291], stage0_60[292], stage0_60[293], stage0_60[294], stage0_60[295]},
      {stage0_61[177]},
      {stage0_62[186], stage0_62[187], stage0_62[188], stage0_62[189], stage0_62[190], stage0_62[191]},
      {stage1_64[31],stage1_63[53],stage1_62[88],stage1_61[126],stage1_60[176]}
   );
   gpc615_5 gpc2326 (
      {stage0_60[296], stage0_60[297], stage0_60[298], stage0_60[299], stage0_60[300]},
      {stage0_61[178]},
      {stage0_62[192], stage0_62[193], stage0_62[194], stage0_62[195], stage0_62[196], stage0_62[197]},
      {stage1_64[32],stage1_63[54],stage1_62[89],stage1_61[127],stage1_60[177]}
   );
   gpc615_5 gpc2327 (
      {stage0_60[301], stage0_60[302], stage0_60[303], stage0_60[304], stage0_60[305]},
      {stage0_61[179]},
      {stage0_62[198], stage0_62[199], stage0_62[200], stage0_62[201], stage0_62[202], stage0_62[203]},
      {stage1_64[33],stage1_63[55],stage1_62[90],stage1_61[128],stage1_60[178]}
   );
   gpc615_5 gpc2328 (
      {stage0_60[306], stage0_60[307], stage0_60[308], stage0_60[309], stage0_60[310]},
      {stage0_61[180]},
      {stage0_62[204], stage0_62[205], stage0_62[206], stage0_62[207], stage0_62[208], stage0_62[209]},
      {stage1_64[34],stage1_63[56],stage1_62[91],stage1_61[129],stage1_60[179]}
   );
   gpc615_5 gpc2329 (
      {stage0_60[311], stage0_60[312], stage0_60[313], stage0_60[314], stage0_60[315]},
      {stage0_61[181]},
      {stage0_62[210], stage0_62[211], stage0_62[212], stage0_62[213], stage0_62[214], stage0_62[215]},
      {stage1_64[35],stage1_63[57],stage1_62[92],stage1_61[130],stage1_60[180]}
   );
   gpc615_5 gpc2330 (
      {stage0_60[316], stage0_60[317], stage0_60[318], stage0_60[319], stage0_60[320]},
      {stage0_61[182]},
      {stage0_62[216], stage0_62[217], stage0_62[218], stage0_62[219], stage0_62[220], stage0_62[221]},
      {stage1_64[36],stage1_63[58],stage1_62[93],stage1_61[131],stage1_60[181]}
   );
   gpc615_5 gpc2331 (
      {stage0_60[321], stage0_60[322], stage0_60[323], stage0_60[324], stage0_60[325]},
      {stage0_61[183]},
      {stage0_62[222], stage0_62[223], stage0_62[224], stage0_62[225], stage0_62[226], stage0_62[227]},
      {stage1_64[37],stage1_63[59],stage1_62[94],stage1_61[132],stage1_60[182]}
   );
   gpc615_5 gpc2332 (
      {stage0_60[326], stage0_60[327], stage0_60[328], stage0_60[329], stage0_60[330]},
      {stage0_61[184]},
      {stage0_62[228], stage0_62[229], stage0_62[230], stage0_62[231], stage0_62[232], stage0_62[233]},
      {stage1_64[38],stage1_63[60],stage1_62[95],stage1_61[133],stage1_60[183]}
   );
   gpc615_5 gpc2333 (
      {stage0_60[331], stage0_60[332], stage0_60[333], stage0_60[334], stage0_60[335]},
      {stage0_61[185]},
      {stage0_62[234], stage0_62[235], stage0_62[236], stage0_62[237], stage0_62[238], stage0_62[239]},
      {stage1_64[39],stage1_63[61],stage1_62[96],stage1_61[134],stage1_60[184]}
   );
   gpc615_5 gpc2334 (
      {stage0_60[336], stage0_60[337], stage0_60[338], stage0_60[339], stage0_60[340]},
      {stage0_61[186]},
      {stage0_62[240], stage0_62[241], stage0_62[242], stage0_62[243], stage0_62[244], stage0_62[245]},
      {stage1_64[40],stage1_63[62],stage1_62[97],stage1_61[135],stage1_60[185]}
   );
   gpc615_5 gpc2335 (
      {stage0_60[341], stage0_60[342], stage0_60[343], stage0_60[344], stage0_60[345]},
      {stage0_61[187]},
      {stage0_62[246], stage0_62[247], stage0_62[248], stage0_62[249], stage0_62[250], stage0_62[251]},
      {stage1_64[41],stage1_63[63],stage1_62[98],stage1_61[136],stage1_60[186]}
   );
   gpc615_5 gpc2336 (
      {stage0_60[346], stage0_60[347], stage0_60[348], stage0_60[349], stage0_60[350]},
      {stage0_61[188]},
      {stage0_62[252], stage0_62[253], stage0_62[254], stage0_62[255], stage0_62[256], stage0_62[257]},
      {stage1_64[42],stage1_63[64],stage1_62[99],stage1_61[137],stage1_60[187]}
   );
   gpc615_5 gpc2337 (
      {stage0_60[351], stage0_60[352], stage0_60[353], stage0_60[354], stage0_60[355]},
      {stage0_61[189]},
      {stage0_62[258], stage0_62[259], stage0_62[260], stage0_62[261], stage0_62[262], stage0_62[263]},
      {stage1_64[43],stage1_63[65],stage1_62[100],stage1_61[138],stage1_60[188]}
   );
   gpc615_5 gpc2338 (
      {stage0_60[356], stage0_60[357], stage0_60[358], stage0_60[359], stage0_60[360]},
      {stage0_61[190]},
      {stage0_62[264], stage0_62[265], stage0_62[266], stage0_62[267], stage0_62[268], stage0_62[269]},
      {stage1_64[44],stage1_63[66],stage1_62[101],stage1_61[139],stage1_60[189]}
   );
   gpc615_5 gpc2339 (
      {stage0_60[361], stage0_60[362], stage0_60[363], stage0_60[364], stage0_60[365]},
      {stage0_61[191]},
      {stage0_62[270], stage0_62[271], stage0_62[272], stage0_62[273], stage0_62[274], stage0_62[275]},
      {stage1_64[45],stage1_63[67],stage1_62[102],stage1_61[140],stage1_60[190]}
   );
   gpc615_5 gpc2340 (
      {stage0_60[366], stage0_60[367], stage0_60[368], stage0_60[369], stage0_60[370]},
      {stage0_61[192]},
      {stage0_62[276], stage0_62[277], stage0_62[278], stage0_62[279], stage0_62[280], stage0_62[281]},
      {stage1_64[46],stage1_63[68],stage1_62[103],stage1_61[141],stage1_60[191]}
   );
   gpc615_5 gpc2341 (
      {stage0_60[371], stage0_60[372], stage0_60[373], stage0_60[374], stage0_60[375]},
      {stage0_61[193]},
      {stage0_62[282], stage0_62[283], stage0_62[284], stage0_62[285], stage0_62[286], stage0_62[287]},
      {stage1_64[47],stage1_63[69],stage1_62[104],stage1_61[142],stage1_60[192]}
   );
   gpc615_5 gpc2342 (
      {stage0_60[376], stage0_60[377], stage0_60[378], stage0_60[379], stage0_60[380]},
      {stage0_61[194]},
      {stage0_62[288], stage0_62[289], stage0_62[290], stage0_62[291], stage0_62[292], stage0_62[293]},
      {stage1_64[48],stage1_63[70],stage1_62[105],stage1_61[143],stage1_60[193]}
   );
   gpc615_5 gpc2343 (
      {stage0_60[381], stage0_60[382], stage0_60[383], stage0_60[384], stage0_60[385]},
      {stage0_61[195]},
      {stage0_62[294], stage0_62[295], stage0_62[296], stage0_62[297], stage0_62[298], stage0_62[299]},
      {stage1_64[49],stage1_63[71],stage1_62[106],stage1_61[144],stage1_60[194]}
   );
   gpc615_5 gpc2344 (
      {stage0_60[386], stage0_60[387], stage0_60[388], stage0_60[389], stage0_60[390]},
      {stage0_61[196]},
      {stage0_62[300], stage0_62[301], stage0_62[302], stage0_62[303], stage0_62[304], stage0_62[305]},
      {stage1_64[50],stage1_63[72],stage1_62[107],stage1_61[145],stage1_60[195]}
   );
   gpc615_5 gpc2345 (
      {stage0_60[391], stage0_60[392], stage0_60[393], stage0_60[394], stage0_60[395]},
      {stage0_61[197]},
      {stage0_62[306], stage0_62[307], stage0_62[308], stage0_62[309], stage0_62[310], stage0_62[311]},
      {stage1_64[51],stage1_63[73],stage1_62[108],stage1_61[146],stage1_60[196]}
   );
   gpc615_5 gpc2346 (
      {stage0_60[396], stage0_60[397], stage0_60[398], stage0_60[399], stage0_60[400]},
      {stage0_61[198]},
      {stage0_62[312], stage0_62[313], stage0_62[314], stage0_62[315], stage0_62[316], stage0_62[317]},
      {stage1_64[52],stage1_63[74],stage1_62[109],stage1_61[147],stage1_60[197]}
   );
   gpc615_5 gpc2347 (
      {stage0_60[401], stage0_60[402], stage0_60[403], stage0_60[404], stage0_60[405]},
      {stage0_61[199]},
      {stage0_62[318], stage0_62[319], stage0_62[320], stage0_62[321], stage0_62[322], stage0_62[323]},
      {stage1_64[53],stage1_63[75],stage1_62[110],stage1_61[148],stage1_60[198]}
   );
   gpc615_5 gpc2348 (
      {stage0_60[406], stage0_60[407], stage0_60[408], stage0_60[409], stage0_60[410]},
      {stage0_61[200]},
      {stage0_62[324], stage0_62[325], stage0_62[326], stage0_62[327], stage0_62[328], stage0_62[329]},
      {stage1_64[54],stage1_63[76],stage1_62[111],stage1_61[149],stage1_60[199]}
   );
   gpc615_5 gpc2349 (
      {stage0_60[411], stage0_60[412], stage0_60[413], stage0_60[414], stage0_60[415]},
      {stage0_61[201]},
      {stage0_62[330], stage0_62[331], stage0_62[332], stage0_62[333], stage0_62[334], stage0_62[335]},
      {stage1_64[55],stage1_63[77],stage1_62[112],stage1_61[150],stage1_60[200]}
   );
   gpc615_5 gpc2350 (
      {stage0_60[416], stage0_60[417], stage0_60[418], stage0_60[419], stage0_60[420]},
      {stage0_61[202]},
      {stage0_62[336], stage0_62[337], stage0_62[338], stage0_62[339], stage0_62[340], stage0_62[341]},
      {stage1_64[56],stage1_63[78],stage1_62[113],stage1_61[151],stage1_60[201]}
   );
   gpc615_5 gpc2351 (
      {stage0_60[421], stage0_60[422], stage0_60[423], stage0_60[424], stage0_60[425]},
      {stage0_61[203]},
      {stage0_62[342], stage0_62[343], stage0_62[344], stage0_62[345], stage0_62[346], stage0_62[347]},
      {stage1_64[57],stage1_63[79],stage1_62[114],stage1_61[152],stage1_60[202]}
   );
   gpc615_5 gpc2352 (
      {stage0_60[426], stage0_60[427], stage0_60[428], stage0_60[429], stage0_60[430]},
      {stage0_61[204]},
      {stage0_62[348], stage0_62[349], stage0_62[350], stage0_62[351], stage0_62[352], stage0_62[353]},
      {stage1_64[58],stage1_63[80],stage1_62[115],stage1_61[153],stage1_60[203]}
   );
   gpc615_5 gpc2353 (
      {stage0_60[431], stage0_60[432], stage0_60[433], stage0_60[434], stage0_60[435]},
      {stage0_61[205]},
      {stage0_62[354], stage0_62[355], stage0_62[356], stage0_62[357], stage0_62[358], stage0_62[359]},
      {stage1_64[59],stage1_63[81],stage1_62[116],stage1_61[154],stage1_60[204]}
   );
   gpc615_5 gpc2354 (
      {stage0_60[436], stage0_60[437], stage0_60[438], stage0_60[439], stage0_60[440]},
      {stage0_61[206]},
      {stage0_62[360], stage0_62[361], stage0_62[362], stage0_62[363], stage0_62[364], stage0_62[365]},
      {stage1_64[60],stage1_63[82],stage1_62[117],stage1_61[155],stage1_60[205]}
   );
   gpc615_5 gpc2355 (
      {stage0_60[441], stage0_60[442], stage0_60[443], stage0_60[444], stage0_60[445]},
      {stage0_61[207]},
      {stage0_62[366], stage0_62[367], stage0_62[368], stage0_62[369], stage0_62[370], stage0_62[371]},
      {stage1_64[61],stage1_63[83],stage1_62[118],stage1_61[156],stage1_60[206]}
   );
   gpc615_5 gpc2356 (
      {stage0_60[446], stage0_60[447], stage0_60[448], stage0_60[449], stage0_60[450]},
      {stage0_61[208]},
      {stage0_62[372], stage0_62[373], stage0_62[374], stage0_62[375], stage0_62[376], stage0_62[377]},
      {stage1_64[62],stage1_63[84],stage1_62[119],stage1_61[157],stage1_60[207]}
   );
   gpc615_5 gpc2357 (
      {stage0_60[451], stage0_60[452], stage0_60[453], stage0_60[454], stage0_60[455]},
      {stage0_61[209]},
      {stage0_62[378], stage0_62[379], stage0_62[380], stage0_62[381], stage0_62[382], stage0_62[383]},
      {stage1_64[63],stage1_63[85],stage1_62[120],stage1_61[158],stage1_60[208]}
   );
   gpc615_5 gpc2358 (
      {stage0_60[456], stage0_60[457], stage0_60[458], stage0_60[459], stage0_60[460]},
      {stage0_61[210]},
      {stage0_62[384], stage0_62[385], stage0_62[386], stage0_62[387], stage0_62[388], stage0_62[389]},
      {stage1_64[64],stage1_63[86],stage1_62[121],stage1_61[159],stage1_60[209]}
   );
   gpc615_5 gpc2359 (
      {stage0_60[461], stage0_60[462], stage0_60[463], stage0_60[464], stage0_60[465]},
      {stage0_61[211]},
      {stage0_62[390], stage0_62[391], stage0_62[392], stage0_62[393], stage0_62[394], stage0_62[395]},
      {stage1_64[65],stage1_63[87],stage1_62[122],stage1_61[160],stage1_60[210]}
   );
   gpc615_5 gpc2360 (
      {stage0_60[466], stage0_60[467], stage0_60[468], stage0_60[469], stage0_60[470]},
      {stage0_61[212]},
      {stage0_62[396], stage0_62[397], stage0_62[398], stage0_62[399], stage0_62[400], stage0_62[401]},
      {stage1_64[66],stage1_63[88],stage1_62[123],stage1_61[161],stage1_60[211]}
   );
   gpc615_5 gpc2361 (
      {stage0_60[471], stage0_60[472], stage0_60[473], stage0_60[474], stage0_60[475]},
      {stage0_61[213]},
      {stage0_62[402], stage0_62[403], stage0_62[404], stage0_62[405], stage0_62[406], stage0_62[407]},
      {stage1_64[67],stage1_63[89],stage1_62[124],stage1_61[162],stage1_60[212]}
   );
   gpc615_5 gpc2362 (
      {stage0_60[476], stage0_60[477], stage0_60[478], stage0_60[479], stage0_60[480]},
      {stage0_61[214]},
      {stage0_62[408], stage0_62[409], stage0_62[410], stage0_62[411], stage0_62[412], stage0_62[413]},
      {stage1_64[68],stage1_63[90],stage1_62[125],stage1_61[163],stage1_60[213]}
   );
   gpc615_5 gpc2363 (
      {stage0_60[481], stage0_60[482], stage0_60[483], stage0_60[484], stage0_60[485]},
      {stage0_61[215]},
      {stage0_62[414], stage0_62[415], stage0_62[416], stage0_62[417], stage0_62[418], stage0_62[419]},
      {stage1_64[69],stage1_63[91],stage1_62[126],stage1_61[164],stage1_60[214]}
   );
   gpc615_5 gpc2364 (
      {stage0_61[216], stage0_61[217], stage0_61[218], stage0_61[219], stage0_61[220]},
      {stage0_62[420]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[70],stage1_63[92],stage1_62[127],stage1_61[165]}
   );
   gpc615_5 gpc2365 (
      {stage0_61[221], stage0_61[222], stage0_61[223], stage0_61[224], stage0_61[225]},
      {stage0_62[421]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[71],stage1_63[93],stage1_62[128],stage1_61[166]}
   );
   gpc615_5 gpc2366 (
      {stage0_61[226], stage0_61[227], stage0_61[228], stage0_61[229], stage0_61[230]},
      {stage0_62[422]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[72],stage1_63[94],stage1_62[129],stage1_61[167]}
   );
   gpc615_5 gpc2367 (
      {stage0_61[231], stage0_61[232], stage0_61[233], stage0_61[234], stage0_61[235]},
      {stage0_62[423]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[73],stage1_63[95],stage1_62[130],stage1_61[168]}
   );
   gpc615_5 gpc2368 (
      {stage0_61[236], stage0_61[237], stage0_61[238], stage0_61[239], stage0_61[240]},
      {stage0_62[424]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[74],stage1_63[96],stage1_62[131],stage1_61[169]}
   );
   gpc615_5 gpc2369 (
      {stage0_61[241], stage0_61[242], stage0_61[243], stage0_61[244], stage0_61[245]},
      {stage0_62[425]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[75],stage1_63[97],stage1_62[132],stage1_61[170]}
   );
   gpc615_5 gpc2370 (
      {stage0_61[246], stage0_61[247], stage0_61[248], stage0_61[249], stage0_61[250]},
      {stage0_62[426]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[76],stage1_63[98],stage1_62[133],stage1_61[171]}
   );
   gpc615_5 gpc2371 (
      {stage0_61[251], stage0_61[252], stage0_61[253], stage0_61[254], stage0_61[255]},
      {stage0_62[427]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[77],stage1_63[99],stage1_62[134],stage1_61[172]}
   );
   gpc615_5 gpc2372 (
      {stage0_61[256], stage0_61[257], stage0_61[258], stage0_61[259], stage0_61[260]},
      {stage0_62[428]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[78],stage1_63[100],stage1_62[135],stage1_61[173]}
   );
   gpc615_5 gpc2373 (
      {stage0_61[261], stage0_61[262], stage0_61[263], stage0_61[264], stage0_61[265]},
      {stage0_62[429]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[79],stage1_63[101],stage1_62[136],stage1_61[174]}
   );
   gpc615_5 gpc2374 (
      {stage0_61[266], stage0_61[267], stage0_61[268], stage0_61[269], stage0_61[270]},
      {stage0_62[430]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[80],stage1_63[102],stage1_62[137],stage1_61[175]}
   );
   gpc615_5 gpc2375 (
      {stage0_61[271], stage0_61[272], stage0_61[273], stage0_61[274], stage0_61[275]},
      {stage0_62[431]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[81],stage1_63[103],stage1_62[138],stage1_61[176]}
   );
   gpc615_5 gpc2376 (
      {stage0_61[276], stage0_61[277], stage0_61[278], stage0_61[279], stage0_61[280]},
      {stage0_62[432]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[82],stage1_63[104],stage1_62[139],stage1_61[177]}
   );
   gpc615_5 gpc2377 (
      {stage0_61[281], stage0_61[282], stage0_61[283], stage0_61[284], stage0_61[285]},
      {stage0_62[433]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[83],stage1_63[105],stage1_62[140],stage1_61[178]}
   );
   gpc615_5 gpc2378 (
      {stage0_61[286], stage0_61[287], stage0_61[288], stage0_61[289], stage0_61[290]},
      {stage0_62[434]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[84],stage1_63[106],stage1_62[141],stage1_61[179]}
   );
   gpc615_5 gpc2379 (
      {stage0_61[291], stage0_61[292], stage0_61[293], stage0_61[294], stage0_61[295]},
      {stage0_62[435]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[85],stage1_63[107],stage1_62[142],stage1_61[180]}
   );
   gpc615_5 gpc2380 (
      {stage0_61[296], stage0_61[297], stage0_61[298], stage0_61[299], stage0_61[300]},
      {stage0_62[436]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[86],stage1_63[108],stage1_62[143],stage1_61[181]}
   );
   gpc615_5 gpc2381 (
      {stage0_61[301], stage0_61[302], stage0_61[303], stage0_61[304], stage0_61[305]},
      {stage0_62[437]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[87],stage1_63[109],stage1_62[144],stage1_61[182]}
   );
   gpc615_5 gpc2382 (
      {stage0_61[306], stage0_61[307], stage0_61[308], stage0_61[309], stage0_61[310]},
      {stage0_62[438]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[88],stage1_63[110],stage1_62[145],stage1_61[183]}
   );
   gpc615_5 gpc2383 (
      {stage0_61[311], stage0_61[312], stage0_61[313], stage0_61[314], stage0_61[315]},
      {stage0_62[439]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[89],stage1_63[111],stage1_62[146],stage1_61[184]}
   );
   gpc615_5 gpc2384 (
      {stage0_61[316], stage0_61[317], stage0_61[318], stage0_61[319], stage0_61[320]},
      {stage0_62[440]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[90],stage1_63[112],stage1_62[147],stage1_61[185]}
   );
   gpc615_5 gpc2385 (
      {stage0_61[321], stage0_61[322], stage0_61[323], stage0_61[324], stage0_61[325]},
      {stage0_62[441]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[91],stage1_63[113],stage1_62[148],stage1_61[186]}
   );
   gpc615_5 gpc2386 (
      {stage0_61[326], stage0_61[327], stage0_61[328], stage0_61[329], stage0_61[330]},
      {stage0_62[442]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[92],stage1_63[114],stage1_62[149],stage1_61[187]}
   );
   gpc615_5 gpc2387 (
      {stage0_61[331], stage0_61[332], stage0_61[333], stage0_61[334], stage0_61[335]},
      {stage0_62[443]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[93],stage1_63[115],stage1_62[150],stage1_61[188]}
   );
   gpc615_5 gpc2388 (
      {stage0_61[336], stage0_61[337], stage0_61[338], stage0_61[339], stage0_61[340]},
      {stage0_62[444]},
      {stage0_63[144], stage0_63[145], stage0_63[146], stage0_63[147], stage0_63[148], stage0_63[149]},
      {stage1_65[24],stage1_64[94],stage1_63[116],stage1_62[151],stage1_61[189]}
   );
   gpc615_5 gpc2389 (
      {stage0_61[341], stage0_61[342], stage0_61[343], stage0_61[344], stage0_61[345]},
      {stage0_62[445]},
      {stage0_63[150], stage0_63[151], stage0_63[152], stage0_63[153], stage0_63[154], stage0_63[155]},
      {stage1_65[25],stage1_64[95],stage1_63[117],stage1_62[152],stage1_61[190]}
   );
   gpc615_5 gpc2390 (
      {stage0_61[346], stage0_61[347], stage0_61[348], stage0_61[349], stage0_61[350]},
      {stage0_62[446]},
      {stage0_63[156], stage0_63[157], stage0_63[158], stage0_63[159], stage0_63[160], stage0_63[161]},
      {stage1_65[26],stage1_64[96],stage1_63[118],stage1_62[153],stage1_61[191]}
   );
   gpc615_5 gpc2391 (
      {stage0_61[351], stage0_61[352], stage0_61[353], stage0_61[354], stage0_61[355]},
      {stage0_62[447]},
      {stage0_63[162], stage0_63[163], stage0_63[164], stage0_63[165], stage0_63[166], stage0_63[167]},
      {stage1_65[27],stage1_64[97],stage1_63[119],stage1_62[154],stage1_61[192]}
   );
   gpc615_5 gpc2392 (
      {stage0_61[356], stage0_61[357], stage0_61[358], stage0_61[359], stage0_61[360]},
      {stage0_62[448]},
      {stage0_63[168], stage0_63[169], stage0_63[170], stage0_63[171], stage0_63[172], stage0_63[173]},
      {stage1_65[28],stage1_64[98],stage1_63[120],stage1_62[155],stage1_61[193]}
   );
   gpc615_5 gpc2393 (
      {stage0_61[361], stage0_61[362], stage0_61[363], stage0_61[364], stage0_61[365]},
      {stage0_62[449]},
      {stage0_63[174], stage0_63[175], stage0_63[176], stage0_63[177], stage0_63[178], stage0_63[179]},
      {stage1_65[29],stage1_64[99],stage1_63[121],stage1_62[156],stage1_61[194]}
   );
   gpc615_5 gpc2394 (
      {stage0_61[366], stage0_61[367], stage0_61[368], stage0_61[369], stage0_61[370]},
      {stage0_62[450]},
      {stage0_63[180], stage0_63[181], stage0_63[182], stage0_63[183], stage0_63[184], stage0_63[185]},
      {stage1_65[30],stage1_64[100],stage1_63[122],stage1_62[157],stage1_61[195]}
   );
   gpc615_5 gpc2395 (
      {stage0_61[371], stage0_61[372], stage0_61[373], stage0_61[374], stage0_61[375]},
      {stage0_62[451]},
      {stage0_63[186], stage0_63[187], stage0_63[188], stage0_63[189], stage0_63[190], stage0_63[191]},
      {stage1_65[31],stage1_64[101],stage1_63[123],stage1_62[158],stage1_61[196]}
   );
   gpc615_5 gpc2396 (
      {stage0_61[376], stage0_61[377], stage0_61[378], stage0_61[379], stage0_61[380]},
      {stage0_62[452]},
      {stage0_63[192], stage0_63[193], stage0_63[194], stage0_63[195], stage0_63[196], stage0_63[197]},
      {stage1_65[32],stage1_64[102],stage1_63[124],stage1_62[159],stage1_61[197]}
   );
   gpc615_5 gpc2397 (
      {stage0_61[381], stage0_61[382], stage0_61[383], stage0_61[384], stage0_61[385]},
      {stage0_62[453]},
      {stage0_63[198], stage0_63[199], stage0_63[200], stage0_63[201], stage0_63[202], stage0_63[203]},
      {stage1_65[33],stage1_64[103],stage1_63[125],stage1_62[160],stage1_61[198]}
   );
   gpc615_5 gpc2398 (
      {stage0_61[386], stage0_61[387], stage0_61[388], stage0_61[389], stage0_61[390]},
      {stage0_62[454]},
      {stage0_63[204], stage0_63[205], stage0_63[206], stage0_63[207], stage0_63[208], stage0_63[209]},
      {stage1_65[34],stage1_64[104],stage1_63[126],stage1_62[161],stage1_61[199]}
   );
   gpc615_5 gpc2399 (
      {stage0_61[391], stage0_61[392], stage0_61[393], stage0_61[394], stage0_61[395]},
      {stage0_62[455]},
      {stage0_63[210], stage0_63[211], stage0_63[212], stage0_63[213], stage0_63[214], stage0_63[215]},
      {stage1_65[35],stage1_64[105],stage1_63[127],stage1_62[162],stage1_61[200]}
   );
   gpc615_5 gpc2400 (
      {stage0_61[396], stage0_61[397], stage0_61[398], stage0_61[399], stage0_61[400]},
      {stage0_62[456]},
      {stage0_63[216], stage0_63[217], stage0_63[218], stage0_63[219], stage0_63[220], stage0_63[221]},
      {stage1_65[36],stage1_64[106],stage1_63[128],stage1_62[163],stage1_61[201]}
   );
   gpc615_5 gpc2401 (
      {stage0_61[401], stage0_61[402], stage0_61[403], stage0_61[404], stage0_61[405]},
      {stage0_62[457]},
      {stage0_63[222], stage0_63[223], stage0_63[224], stage0_63[225], stage0_63[226], stage0_63[227]},
      {stage1_65[37],stage1_64[107],stage1_63[129],stage1_62[164],stage1_61[202]}
   );
   gpc615_5 gpc2402 (
      {stage0_61[406], stage0_61[407], stage0_61[408], stage0_61[409], stage0_61[410]},
      {stage0_62[458]},
      {stage0_63[228], stage0_63[229], stage0_63[230], stage0_63[231], stage0_63[232], stage0_63[233]},
      {stage1_65[38],stage1_64[108],stage1_63[130],stage1_62[165],stage1_61[203]}
   );
   gpc615_5 gpc2403 (
      {stage0_61[411], stage0_61[412], stage0_61[413], stage0_61[414], stage0_61[415]},
      {stage0_62[459]},
      {stage0_63[234], stage0_63[235], stage0_63[236], stage0_63[237], stage0_63[238], stage0_63[239]},
      {stage1_65[39],stage1_64[109],stage1_63[131],stage1_62[166],stage1_61[204]}
   );
   gpc615_5 gpc2404 (
      {stage0_61[416], stage0_61[417], stage0_61[418], stage0_61[419], stage0_61[420]},
      {stage0_62[460]},
      {stage0_63[240], stage0_63[241], stage0_63[242], stage0_63[243], stage0_63[244], stage0_63[245]},
      {stage1_65[40],stage1_64[110],stage1_63[132],stage1_62[167],stage1_61[205]}
   );
   gpc615_5 gpc2405 (
      {stage0_61[421], stage0_61[422], stage0_61[423], stage0_61[424], stage0_61[425]},
      {stage0_62[461]},
      {stage0_63[246], stage0_63[247], stage0_63[248], stage0_63[249], stage0_63[250], stage0_63[251]},
      {stage1_65[41],stage1_64[111],stage1_63[133],stage1_62[168],stage1_61[206]}
   );
   gpc615_5 gpc2406 (
      {stage0_61[426], stage0_61[427], stage0_61[428], stage0_61[429], stage0_61[430]},
      {stage0_62[462]},
      {stage0_63[252], stage0_63[253], stage0_63[254], stage0_63[255], stage0_63[256], stage0_63[257]},
      {stage1_65[42],stage1_64[112],stage1_63[134],stage1_62[169],stage1_61[207]}
   );
   gpc615_5 gpc2407 (
      {stage0_61[431], stage0_61[432], stage0_61[433], stage0_61[434], stage0_61[435]},
      {stage0_62[463]},
      {stage0_63[258], stage0_63[259], stage0_63[260], stage0_63[261], stage0_63[262], stage0_63[263]},
      {stage1_65[43],stage1_64[113],stage1_63[135],stage1_62[170],stage1_61[208]}
   );
   gpc615_5 gpc2408 (
      {stage0_61[436], stage0_61[437], stage0_61[438], stage0_61[439], stage0_61[440]},
      {stage0_62[464]},
      {stage0_63[264], stage0_63[265], stage0_63[266], stage0_63[267], stage0_63[268], stage0_63[269]},
      {stage1_65[44],stage1_64[114],stage1_63[136],stage1_62[171],stage1_61[209]}
   );
   gpc615_5 gpc2409 (
      {stage0_61[441], stage0_61[442], stage0_61[443], stage0_61[444], stage0_61[445]},
      {stage0_62[465]},
      {stage0_63[270], stage0_63[271], stage0_63[272], stage0_63[273], stage0_63[274], stage0_63[275]},
      {stage1_65[45],stage1_64[115],stage1_63[137],stage1_62[172],stage1_61[210]}
   );
   gpc615_5 gpc2410 (
      {stage0_61[446], stage0_61[447], stage0_61[448], stage0_61[449], stage0_61[450]},
      {stage0_62[466]},
      {stage0_63[276], stage0_63[277], stage0_63[278], stage0_63[279], stage0_63[280], stage0_63[281]},
      {stage1_65[46],stage1_64[116],stage1_63[138],stage1_62[173],stage1_61[211]}
   );
   gpc615_5 gpc2411 (
      {stage0_61[451], stage0_61[452], stage0_61[453], stage0_61[454], stage0_61[455]},
      {stage0_62[467]},
      {stage0_63[282], stage0_63[283], stage0_63[284], stage0_63[285], stage0_63[286], stage0_63[287]},
      {stage1_65[47],stage1_64[117],stage1_63[139],stage1_62[174],stage1_61[212]}
   );
   gpc615_5 gpc2412 (
      {stage0_61[456], stage0_61[457], stage0_61[458], stage0_61[459], stage0_61[460]},
      {stage0_62[468]},
      {stage0_63[288], stage0_63[289], stage0_63[290], stage0_63[291], stage0_63[292], stage0_63[293]},
      {stage1_65[48],stage1_64[118],stage1_63[140],stage1_62[175],stage1_61[213]}
   );
   gpc615_5 gpc2413 (
      {stage0_61[461], stage0_61[462], stage0_61[463], stage0_61[464], stage0_61[465]},
      {stage0_62[469]},
      {stage0_63[294], stage0_63[295], stage0_63[296], stage0_63[297], stage0_63[298], stage0_63[299]},
      {stage1_65[49],stage1_64[119],stage1_63[141],stage1_62[176],stage1_61[214]}
   );
   gpc615_5 gpc2414 (
      {stage0_61[466], stage0_61[467], stage0_61[468], stage0_61[469], stage0_61[470]},
      {stage0_62[470]},
      {stage0_63[300], stage0_63[301], stage0_63[302], stage0_63[303], stage0_63[304], stage0_63[305]},
      {stage1_65[50],stage1_64[120],stage1_63[142],stage1_62[177],stage1_61[215]}
   );
   gpc615_5 gpc2415 (
      {stage0_61[471], stage0_61[472], stage0_61[473], stage0_61[474], stage0_61[475]},
      {stage0_62[471]},
      {stage0_63[306], stage0_63[307], stage0_63[308], stage0_63[309], stage0_63[310], stage0_63[311]},
      {stage1_65[51],stage1_64[121],stage1_63[143],stage1_62[178],stage1_61[216]}
   );
   gpc615_5 gpc2416 (
      {stage0_61[476], stage0_61[477], stage0_61[478], stage0_61[479], stage0_61[480]},
      {stage0_62[472]},
      {stage0_63[312], stage0_63[313], stage0_63[314], stage0_63[315], stage0_63[316], stage0_63[317]},
      {stage1_65[52],stage1_64[122],stage1_63[144],stage1_62[179],stage1_61[217]}
   );
   gpc615_5 gpc2417 (
      {stage0_61[481], stage0_61[482], stage0_61[483], stage0_61[484], stage0_61[485]},
      {stage0_62[473]},
      {stage0_63[318], stage0_63[319], stage0_63[320], stage0_63[321], stage0_63[322], stage0_63[323]},
      {stage1_65[53],stage1_64[123],stage1_63[145],stage1_62[180],stage1_61[218]}
   );
   gpc1_1 gpc2418 (
      {stage0_0[448]},
      {stage1_0[87]}
   );
   gpc1_1 gpc2419 (
      {stage0_0[449]},
      {stage1_0[88]}
   );
   gpc1_1 gpc2420 (
      {stage0_0[450]},
      {stage1_0[89]}
   );
   gpc1_1 gpc2421 (
      {stage0_0[451]},
      {stage1_0[90]}
   );
   gpc1_1 gpc2422 (
      {stage0_0[452]},
      {stage1_0[91]}
   );
   gpc1_1 gpc2423 (
      {stage0_0[453]},
      {stage1_0[92]}
   );
   gpc1_1 gpc2424 (
      {stage0_0[454]},
      {stage1_0[93]}
   );
   gpc1_1 gpc2425 (
      {stage0_0[455]},
      {stage1_0[94]}
   );
   gpc1_1 gpc2426 (
      {stage0_0[456]},
      {stage1_0[95]}
   );
   gpc1_1 gpc2427 (
      {stage0_0[457]},
      {stage1_0[96]}
   );
   gpc1_1 gpc2428 (
      {stage0_0[458]},
      {stage1_0[97]}
   );
   gpc1_1 gpc2429 (
      {stage0_0[459]},
      {stage1_0[98]}
   );
   gpc1_1 gpc2430 (
      {stage0_0[460]},
      {stage1_0[99]}
   );
   gpc1_1 gpc2431 (
      {stage0_0[461]},
      {stage1_0[100]}
   );
   gpc1_1 gpc2432 (
      {stage0_0[462]},
      {stage1_0[101]}
   );
   gpc1_1 gpc2433 (
      {stage0_0[463]},
      {stage1_0[102]}
   );
   gpc1_1 gpc2434 (
      {stage0_0[464]},
      {stage1_0[103]}
   );
   gpc1_1 gpc2435 (
      {stage0_0[465]},
      {stage1_0[104]}
   );
   gpc1_1 gpc2436 (
      {stage0_0[466]},
      {stage1_0[105]}
   );
   gpc1_1 gpc2437 (
      {stage0_0[467]},
      {stage1_0[106]}
   );
   gpc1_1 gpc2438 (
      {stage0_0[468]},
      {stage1_0[107]}
   );
   gpc1_1 gpc2439 (
      {stage0_0[469]},
      {stage1_0[108]}
   );
   gpc1_1 gpc2440 (
      {stage0_0[470]},
      {stage1_0[109]}
   );
   gpc1_1 gpc2441 (
      {stage0_0[471]},
      {stage1_0[110]}
   );
   gpc1_1 gpc2442 (
      {stage0_0[472]},
      {stage1_0[111]}
   );
   gpc1_1 gpc2443 (
      {stage0_0[473]},
      {stage1_0[112]}
   );
   gpc1_1 gpc2444 (
      {stage0_0[474]},
      {stage1_0[113]}
   );
   gpc1_1 gpc2445 (
      {stage0_0[475]},
      {stage1_0[114]}
   );
   gpc1_1 gpc2446 (
      {stage0_0[476]},
      {stage1_0[115]}
   );
   gpc1_1 gpc2447 (
      {stage0_0[477]},
      {stage1_0[116]}
   );
   gpc1_1 gpc2448 (
      {stage0_0[478]},
      {stage1_0[117]}
   );
   gpc1_1 gpc2449 (
      {stage0_0[479]},
      {stage1_0[118]}
   );
   gpc1_1 gpc2450 (
      {stage0_0[480]},
      {stage1_0[119]}
   );
   gpc1_1 gpc2451 (
      {stage0_0[481]},
      {stage1_0[120]}
   );
   gpc1_1 gpc2452 (
      {stage0_0[482]},
      {stage1_0[121]}
   );
   gpc1_1 gpc2453 (
      {stage0_0[483]},
      {stage1_0[122]}
   );
   gpc1_1 gpc2454 (
      {stage0_0[484]},
      {stage1_0[123]}
   );
   gpc1_1 gpc2455 (
      {stage0_0[485]},
      {stage1_0[124]}
   );
   gpc1_1 gpc2456 (
      {stage0_1[439]},
      {stage1_1[129]}
   );
   gpc1_1 gpc2457 (
      {stage0_1[440]},
      {stage1_1[130]}
   );
   gpc1_1 gpc2458 (
      {stage0_1[441]},
      {stage1_1[131]}
   );
   gpc1_1 gpc2459 (
      {stage0_1[442]},
      {stage1_1[132]}
   );
   gpc1_1 gpc2460 (
      {stage0_1[443]},
      {stage1_1[133]}
   );
   gpc1_1 gpc2461 (
      {stage0_1[444]},
      {stage1_1[134]}
   );
   gpc1_1 gpc2462 (
      {stage0_1[445]},
      {stage1_1[135]}
   );
   gpc1_1 gpc2463 (
      {stage0_1[446]},
      {stage1_1[136]}
   );
   gpc1_1 gpc2464 (
      {stage0_1[447]},
      {stage1_1[137]}
   );
   gpc1_1 gpc2465 (
      {stage0_1[448]},
      {stage1_1[138]}
   );
   gpc1_1 gpc2466 (
      {stage0_1[449]},
      {stage1_1[139]}
   );
   gpc1_1 gpc2467 (
      {stage0_1[450]},
      {stage1_1[140]}
   );
   gpc1_1 gpc2468 (
      {stage0_1[451]},
      {stage1_1[141]}
   );
   gpc1_1 gpc2469 (
      {stage0_1[452]},
      {stage1_1[142]}
   );
   gpc1_1 gpc2470 (
      {stage0_1[453]},
      {stage1_1[143]}
   );
   gpc1_1 gpc2471 (
      {stage0_1[454]},
      {stage1_1[144]}
   );
   gpc1_1 gpc2472 (
      {stage0_1[455]},
      {stage1_1[145]}
   );
   gpc1_1 gpc2473 (
      {stage0_1[456]},
      {stage1_1[146]}
   );
   gpc1_1 gpc2474 (
      {stage0_1[457]},
      {stage1_1[147]}
   );
   gpc1_1 gpc2475 (
      {stage0_1[458]},
      {stage1_1[148]}
   );
   gpc1_1 gpc2476 (
      {stage0_1[459]},
      {stage1_1[149]}
   );
   gpc1_1 gpc2477 (
      {stage0_1[460]},
      {stage1_1[150]}
   );
   gpc1_1 gpc2478 (
      {stage0_1[461]},
      {stage1_1[151]}
   );
   gpc1_1 gpc2479 (
      {stage0_1[462]},
      {stage1_1[152]}
   );
   gpc1_1 gpc2480 (
      {stage0_1[463]},
      {stage1_1[153]}
   );
   gpc1_1 gpc2481 (
      {stage0_1[464]},
      {stage1_1[154]}
   );
   gpc1_1 gpc2482 (
      {stage0_1[465]},
      {stage1_1[155]}
   );
   gpc1_1 gpc2483 (
      {stage0_1[466]},
      {stage1_1[156]}
   );
   gpc1_1 gpc2484 (
      {stage0_1[467]},
      {stage1_1[157]}
   );
   gpc1_1 gpc2485 (
      {stage0_1[468]},
      {stage1_1[158]}
   );
   gpc1_1 gpc2486 (
      {stage0_1[469]},
      {stage1_1[159]}
   );
   gpc1_1 gpc2487 (
      {stage0_1[470]},
      {stage1_1[160]}
   );
   gpc1_1 gpc2488 (
      {stage0_1[471]},
      {stage1_1[161]}
   );
   gpc1_1 gpc2489 (
      {stage0_1[472]},
      {stage1_1[162]}
   );
   gpc1_1 gpc2490 (
      {stage0_1[473]},
      {stage1_1[163]}
   );
   gpc1_1 gpc2491 (
      {stage0_1[474]},
      {stage1_1[164]}
   );
   gpc1_1 gpc2492 (
      {stage0_1[475]},
      {stage1_1[165]}
   );
   gpc1_1 gpc2493 (
      {stage0_1[476]},
      {stage1_1[166]}
   );
   gpc1_1 gpc2494 (
      {stage0_1[477]},
      {stage1_1[167]}
   );
   gpc1_1 gpc2495 (
      {stage0_1[478]},
      {stage1_1[168]}
   );
   gpc1_1 gpc2496 (
      {stage0_1[479]},
      {stage1_1[169]}
   );
   gpc1_1 gpc2497 (
      {stage0_1[480]},
      {stage1_1[170]}
   );
   gpc1_1 gpc2498 (
      {stage0_1[481]},
      {stage1_1[171]}
   );
   gpc1_1 gpc2499 (
      {stage0_1[482]},
      {stage1_1[172]}
   );
   gpc1_1 gpc2500 (
      {stage0_1[483]},
      {stage1_1[173]}
   );
   gpc1_1 gpc2501 (
      {stage0_1[484]},
      {stage1_1[174]}
   );
   gpc1_1 gpc2502 (
      {stage0_1[485]},
      {stage1_1[175]}
   );
   gpc1_1 gpc2503 (
      {stage0_3[466]},
      {stage1_3[195]}
   );
   gpc1_1 gpc2504 (
      {stage0_3[467]},
      {stage1_3[196]}
   );
   gpc1_1 gpc2505 (
      {stage0_3[468]},
      {stage1_3[197]}
   );
   gpc1_1 gpc2506 (
      {stage0_3[469]},
      {stage1_3[198]}
   );
   gpc1_1 gpc2507 (
      {stage0_3[470]},
      {stage1_3[199]}
   );
   gpc1_1 gpc2508 (
      {stage0_3[471]},
      {stage1_3[200]}
   );
   gpc1_1 gpc2509 (
      {stage0_3[472]},
      {stage1_3[201]}
   );
   gpc1_1 gpc2510 (
      {stage0_3[473]},
      {stage1_3[202]}
   );
   gpc1_1 gpc2511 (
      {stage0_3[474]},
      {stage1_3[203]}
   );
   gpc1_1 gpc2512 (
      {stage0_3[475]},
      {stage1_3[204]}
   );
   gpc1_1 gpc2513 (
      {stage0_3[476]},
      {stage1_3[205]}
   );
   gpc1_1 gpc2514 (
      {stage0_3[477]},
      {stage1_3[206]}
   );
   gpc1_1 gpc2515 (
      {stage0_3[478]},
      {stage1_3[207]}
   );
   gpc1_1 gpc2516 (
      {stage0_3[479]},
      {stage1_3[208]}
   );
   gpc1_1 gpc2517 (
      {stage0_3[480]},
      {stage1_3[209]}
   );
   gpc1_1 gpc2518 (
      {stage0_3[481]},
      {stage1_3[210]}
   );
   gpc1_1 gpc2519 (
      {stage0_3[482]},
      {stage1_3[211]}
   );
   gpc1_1 gpc2520 (
      {stage0_3[483]},
      {stage1_3[212]}
   );
   gpc1_1 gpc2521 (
      {stage0_3[484]},
      {stage1_3[213]}
   );
   gpc1_1 gpc2522 (
      {stage0_3[485]},
      {stage1_3[214]}
   );
   gpc1_1 gpc2523 (
      {stage0_6[466]},
      {stage1_6[194]}
   );
   gpc1_1 gpc2524 (
      {stage0_6[467]},
      {stage1_6[195]}
   );
   gpc1_1 gpc2525 (
      {stage0_6[468]},
      {stage1_6[196]}
   );
   gpc1_1 gpc2526 (
      {stage0_6[469]},
      {stage1_6[197]}
   );
   gpc1_1 gpc2527 (
      {stage0_6[470]},
      {stage1_6[198]}
   );
   gpc1_1 gpc2528 (
      {stage0_6[471]},
      {stage1_6[199]}
   );
   gpc1_1 gpc2529 (
      {stage0_6[472]},
      {stage1_6[200]}
   );
   gpc1_1 gpc2530 (
      {stage0_6[473]},
      {stage1_6[201]}
   );
   gpc1_1 gpc2531 (
      {stage0_6[474]},
      {stage1_6[202]}
   );
   gpc1_1 gpc2532 (
      {stage0_6[475]},
      {stage1_6[203]}
   );
   gpc1_1 gpc2533 (
      {stage0_6[476]},
      {stage1_6[204]}
   );
   gpc1_1 gpc2534 (
      {stage0_6[477]},
      {stage1_6[205]}
   );
   gpc1_1 gpc2535 (
      {stage0_6[478]},
      {stage1_6[206]}
   );
   gpc1_1 gpc2536 (
      {stage0_6[479]},
      {stage1_6[207]}
   );
   gpc1_1 gpc2537 (
      {stage0_6[480]},
      {stage1_6[208]}
   );
   gpc1_1 gpc2538 (
      {stage0_6[481]},
      {stage1_6[209]}
   );
   gpc1_1 gpc2539 (
      {stage0_6[482]},
      {stage1_6[210]}
   );
   gpc1_1 gpc2540 (
      {stage0_6[483]},
      {stage1_6[211]}
   );
   gpc1_1 gpc2541 (
      {stage0_6[484]},
      {stage1_6[212]}
   );
   gpc1_1 gpc2542 (
      {stage0_6[485]},
      {stage1_6[213]}
   );
   gpc1_1 gpc2543 (
      {stage0_7[462]},
      {stage1_7[197]}
   );
   gpc1_1 gpc2544 (
      {stage0_7[463]},
      {stage1_7[198]}
   );
   gpc1_1 gpc2545 (
      {stage0_7[464]},
      {stage1_7[199]}
   );
   gpc1_1 gpc2546 (
      {stage0_7[465]},
      {stage1_7[200]}
   );
   gpc1_1 gpc2547 (
      {stage0_7[466]},
      {stage1_7[201]}
   );
   gpc1_1 gpc2548 (
      {stage0_7[467]},
      {stage1_7[202]}
   );
   gpc1_1 gpc2549 (
      {stage0_7[468]},
      {stage1_7[203]}
   );
   gpc1_1 gpc2550 (
      {stage0_7[469]},
      {stage1_7[204]}
   );
   gpc1_1 gpc2551 (
      {stage0_7[470]},
      {stage1_7[205]}
   );
   gpc1_1 gpc2552 (
      {stage0_7[471]},
      {stage1_7[206]}
   );
   gpc1_1 gpc2553 (
      {stage0_7[472]},
      {stage1_7[207]}
   );
   gpc1_1 gpc2554 (
      {stage0_7[473]},
      {stage1_7[208]}
   );
   gpc1_1 gpc2555 (
      {stage0_7[474]},
      {stage1_7[209]}
   );
   gpc1_1 gpc2556 (
      {stage0_7[475]},
      {stage1_7[210]}
   );
   gpc1_1 gpc2557 (
      {stage0_7[476]},
      {stage1_7[211]}
   );
   gpc1_1 gpc2558 (
      {stage0_7[477]},
      {stage1_7[212]}
   );
   gpc1_1 gpc2559 (
      {stage0_7[478]},
      {stage1_7[213]}
   );
   gpc1_1 gpc2560 (
      {stage0_7[479]},
      {stage1_7[214]}
   );
   gpc1_1 gpc2561 (
      {stage0_7[480]},
      {stage1_7[215]}
   );
   gpc1_1 gpc2562 (
      {stage0_7[481]},
      {stage1_7[216]}
   );
   gpc1_1 gpc2563 (
      {stage0_7[482]},
      {stage1_7[217]}
   );
   gpc1_1 gpc2564 (
      {stage0_7[483]},
      {stage1_7[218]}
   );
   gpc1_1 gpc2565 (
      {stage0_7[484]},
      {stage1_7[219]}
   );
   gpc1_1 gpc2566 (
      {stage0_7[485]},
      {stage1_7[220]}
   );
   gpc1_1 gpc2567 (
      {stage0_8[476]},
      {stage1_8[196]}
   );
   gpc1_1 gpc2568 (
      {stage0_8[477]},
      {stage1_8[197]}
   );
   gpc1_1 gpc2569 (
      {stage0_8[478]},
      {stage1_8[198]}
   );
   gpc1_1 gpc2570 (
      {stage0_8[479]},
      {stage1_8[199]}
   );
   gpc1_1 gpc2571 (
      {stage0_8[480]},
      {stage1_8[200]}
   );
   gpc1_1 gpc2572 (
      {stage0_8[481]},
      {stage1_8[201]}
   );
   gpc1_1 gpc2573 (
      {stage0_8[482]},
      {stage1_8[202]}
   );
   gpc1_1 gpc2574 (
      {stage0_8[483]},
      {stage1_8[203]}
   );
   gpc1_1 gpc2575 (
      {stage0_8[484]},
      {stage1_8[204]}
   );
   gpc1_1 gpc2576 (
      {stage0_8[485]},
      {stage1_8[205]}
   );
   gpc1_1 gpc2577 (
      {stage0_9[468]},
      {stage1_9[196]}
   );
   gpc1_1 gpc2578 (
      {stage0_9[469]},
      {stage1_9[197]}
   );
   gpc1_1 gpc2579 (
      {stage0_9[470]},
      {stage1_9[198]}
   );
   gpc1_1 gpc2580 (
      {stage0_9[471]},
      {stage1_9[199]}
   );
   gpc1_1 gpc2581 (
      {stage0_9[472]},
      {stage1_9[200]}
   );
   gpc1_1 gpc2582 (
      {stage0_9[473]},
      {stage1_9[201]}
   );
   gpc1_1 gpc2583 (
      {stage0_9[474]},
      {stage1_9[202]}
   );
   gpc1_1 gpc2584 (
      {stage0_9[475]},
      {stage1_9[203]}
   );
   gpc1_1 gpc2585 (
      {stage0_9[476]},
      {stage1_9[204]}
   );
   gpc1_1 gpc2586 (
      {stage0_9[477]},
      {stage1_9[205]}
   );
   gpc1_1 gpc2587 (
      {stage0_9[478]},
      {stage1_9[206]}
   );
   gpc1_1 gpc2588 (
      {stage0_9[479]},
      {stage1_9[207]}
   );
   gpc1_1 gpc2589 (
      {stage0_9[480]},
      {stage1_9[208]}
   );
   gpc1_1 gpc2590 (
      {stage0_9[481]},
      {stage1_9[209]}
   );
   gpc1_1 gpc2591 (
      {stage0_9[482]},
      {stage1_9[210]}
   );
   gpc1_1 gpc2592 (
      {stage0_9[483]},
      {stage1_9[211]}
   );
   gpc1_1 gpc2593 (
      {stage0_9[484]},
      {stage1_9[212]}
   );
   gpc1_1 gpc2594 (
      {stage0_9[485]},
      {stage1_9[213]}
   );
   gpc1_1 gpc2595 (
      {stage0_10[384]},
      {stage1_10[183]}
   );
   gpc1_1 gpc2596 (
      {stage0_10[385]},
      {stage1_10[184]}
   );
   gpc1_1 gpc2597 (
      {stage0_10[386]},
      {stage1_10[185]}
   );
   gpc1_1 gpc2598 (
      {stage0_10[387]},
      {stage1_10[186]}
   );
   gpc1_1 gpc2599 (
      {stage0_10[388]},
      {stage1_10[187]}
   );
   gpc1_1 gpc2600 (
      {stage0_10[389]},
      {stage1_10[188]}
   );
   gpc1_1 gpc2601 (
      {stage0_10[390]},
      {stage1_10[189]}
   );
   gpc1_1 gpc2602 (
      {stage0_10[391]},
      {stage1_10[190]}
   );
   gpc1_1 gpc2603 (
      {stage0_10[392]},
      {stage1_10[191]}
   );
   gpc1_1 gpc2604 (
      {stage0_10[393]},
      {stage1_10[192]}
   );
   gpc1_1 gpc2605 (
      {stage0_10[394]},
      {stage1_10[193]}
   );
   gpc1_1 gpc2606 (
      {stage0_10[395]},
      {stage1_10[194]}
   );
   gpc1_1 gpc2607 (
      {stage0_10[396]},
      {stage1_10[195]}
   );
   gpc1_1 gpc2608 (
      {stage0_10[397]},
      {stage1_10[196]}
   );
   gpc1_1 gpc2609 (
      {stage0_10[398]},
      {stage1_10[197]}
   );
   gpc1_1 gpc2610 (
      {stage0_10[399]},
      {stage1_10[198]}
   );
   gpc1_1 gpc2611 (
      {stage0_10[400]},
      {stage1_10[199]}
   );
   gpc1_1 gpc2612 (
      {stage0_10[401]},
      {stage1_10[200]}
   );
   gpc1_1 gpc2613 (
      {stage0_10[402]},
      {stage1_10[201]}
   );
   gpc1_1 gpc2614 (
      {stage0_10[403]},
      {stage1_10[202]}
   );
   gpc1_1 gpc2615 (
      {stage0_10[404]},
      {stage1_10[203]}
   );
   gpc1_1 gpc2616 (
      {stage0_10[405]},
      {stage1_10[204]}
   );
   gpc1_1 gpc2617 (
      {stage0_10[406]},
      {stage1_10[205]}
   );
   gpc1_1 gpc2618 (
      {stage0_10[407]},
      {stage1_10[206]}
   );
   gpc1_1 gpc2619 (
      {stage0_10[408]},
      {stage1_10[207]}
   );
   gpc1_1 gpc2620 (
      {stage0_10[409]},
      {stage1_10[208]}
   );
   gpc1_1 gpc2621 (
      {stage0_10[410]},
      {stage1_10[209]}
   );
   gpc1_1 gpc2622 (
      {stage0_10[411]},
      {stage1_10[210]}
   );
   gpc1_1 gpc2623 (
      {stage0_10[412]},
      {stage1_10[211]}
   );
   gpc1_1 gpc2624 (
      {stage0_10[413]},
      {stage1_10[212]}
   );
   gpc1_1 gpc2625 (
      {stage0_10[414]},
      {stage1_10[213]}
   );
   gpc1_1 gpc2626 (
      {stage0_10[415]},
      {stage1_10[214]}
   );
   gpc1_1 gpc2627 (
      {stage0_10[416]},
      {stage1_10[215]}
   );
   gpc1_1 gpc2628 (
      {stage0_10[417]},
      {stage1_10[216]}
   );
   gpc1_1 gpc2629 (
      {stage0_10[418]},
      {stage1_10[217]}
   );
   gpc1_1 gpc2630 (
      {stage0_10[419]},
      {stage1_10[218]}
   );
   gpc1_1 gpc2631 (
      {stage0_10[420]},
      {stage1_10[219]}
   );
   gpc1_1 gpc2632 (
      {stage0_10[421]},
      {stage1_10[220]}
   );
   gpc1_1 gpc2633 (
      {stage0_10[422]},
      {stage1_10[221]}
   );
   gpc1_1 gpc2634 (
      {stage0_10[423]},
      {stage1_10[222]}
   );
   gpc1_1 gpc2635 (
      {stage0_10[424]},
      {stage1_10[223]}
   );
   gpc1_1 gpc2636 (
      {stage0_10[425]},
      {stage1_10[224]}
   );
   gpc1_1 gpc2637 (
      {stage0_10[426]},
      {stage1_10[225]}
   );
   gpc1_1 gpc2638 (
      {stage0_10[427]},
      {stage1_10[226]}
   );
   gpc1_1 gpc2639 (
      {stage0_10[428]},
      {stage1_10[227]}
   );
   gpc1_1 gpc2640 (
      {stage0_10[429]},
      {stage1_10[228]}
   );
   gpc1_1 gpc2641 (
      {stage0_10[430]},
      {stage1_10[229]}
   );
   gpc1_1 gpc2642 (
      {stage0_10[431]},
      {stage1_10[230]}
   );
   gpc1_1 gpc2643 (
      {stage0_10[432]},
      {stage1_10[231]}
   );
   gpc1_1 gpc2644 (
      {stage0_10[433]},
      {stage1_10[232]}
   );
   gpc1_1 gpc2645 (
      {stage0_10[434]},
      {stage1_10[233]}
   );
   gpc1_1 gpc2646 (
      {stage0_10[435]},
      {stage1_10[234]}
   );
   gpc1_1 gpc2647 (
      {stage0_10[436]},
      {stage1_10[235]}
   );
   gpc1_1 gpc2648 (
      {stage0_10[437]},
      {stage1_10[236]}
   );
   gpc1_1 gpc2649 (
      {stage0_10[438]},
      {stage1_10[237]}
   );
   gpc1_1 gpc2650 (
      {stage0_10[439]},
      {stage1_10[238]}
   );
   gpc1_1 gpc2651 (
      {stage0_10[440]},
      {stage1_10[239]}
   );
   gpc1_1 gpc2652 (
      {stage0_10[441]},
      {stage1_10[240]}
   );
   gpc1_1 gpc2653 (
      {stage0_10[442]},
      {stage1_10[241]}
   );
   gpc1_1 gpc2654 (
      {stage0_10[443]},
      {stage1_10[242]}
   );
   gpc1_1 gpc2655 (
      {stage0_10[444]},
      {stage1_10[243]}
   );
   gpc1_1 gpc2656 (
      {stage0_10[445]},
      {stage1_10[244]}
   );
   gpc1_1 gpc2657 (
      {stage0_10[446]},
      {stage1_10[245]}
   );
   gpc1_1 gpc2658 (
      {stage0_10[447]},
      {stage1_10[246]}
   );
   gpc1_1 gpc2659 (
      {stage0_10[448]},
      {stage1_10[247]}
   );
   gpc1_1 gpc2660 (
      {stage0_10[449]},
      {stage1_10[248]}
   );
   gpc1_1 gpc2661 (
      {stage0_10[450]},
      {stage1_10[249]}
   );
   gpc1_1 gpc2662 (
      {stage0_10[451]},
      {stage1_10[250]}
   );
   gpc1_1 gpc2663 (
      {stage0_10[452]},
      {stage1_10[251]}
   );
   gpc1_1 gpc2664 (
      {stage0_10[453]},
      {stage1_10[252]}
   );
   gpc1_1 gpc2665 (
      {stage0_10[454]},
      {stage1_10[253]}
   );
   gpc1_1 gpc2666 (
      {stage0_10[455]},
      {stage1_10[254]}
   );
   gpc1_1 gpc2667 (
      {stage0_10[456]},
      {stage1_10[255]}
   );
   gpc1_1 gpc2668 (
      {stage0_10[457]},
      {stage1_10[256]}
   );
   gpc1_1 gpc2669 (
      {stage0_10[458]},
      {stage1_10[257]}
   );
   gpc1_1 gpc2670 (
      {stage0_10[459]},
      {stage1_10[258]}
   );
   gpc1_1 gpc2671 (
      {stage0_10[460]},
      {stage1_10[259]}
   );
   gpc1_1 gpc2672 (
      {stage0_10[461]},
      {stage1_10[260]}
   );
   gpc1_1 gpc2673 (
      {stage0_10[462]},
      {stage1_10[261]}
   );
   gpc1_1 gpc2674 (
      {stage0_10[463]},
      {stage1_10[262]}
   );
   gpc1_1 gpc2675 (
      {stage0_10[464]},
      {stage1_10[263]}
   );
   gpc1_1 gpc2676 (
      {stage0_10[465]},
      {stage1_10[264]}
   );
   gpc1_1 gpc2677 (
      {stage0_10[466]},
      {stage1_10[265]}
   );
   gpc1_1 gpc2678 (
      {stage0_10[467]},
      {stage1_10[266]}
   );
   gpc1_1 gpc2679 (
      {stage0_10[468]},
      {stage1_10[267]}
   );
   gpc1_1 gpc2680 (
      {stage0_10[469]},
      {stage1_10[268]}
   );
   gpc1_1 gpc2681 (
      {stage0_10[470]},
      {stage1_10[269]}
   );
   gpc1_1 gpc2682 (
      {stage0_10[471]},
      {stage1_10[270]}
   );
   gpc1_1 gpc2683 (
      {stage0_10[472]},
      {stage1_10[271]}
   );
   gpc1_1 gpc2684 (
      {stage0_10[473]},
      {stage1_10[272]}
   );
   gpc1_1 gpc2685 (
      {stage0_10[474]},
      {stage1_10[273]}
   );
   gpc1_1 gpc2686 (
      {stage0_10[475]},
      {stage1_10[274]}
   );
   gpc1_1 gpc2687 (
      {stage0_10[476]},
      {stage1_10[275]}
   );
   gpc1_1 gpc2688 (
      {stage0_10[477]},
      {stage1_10[276]}
   );
   gpc1_1 gpc2689 (
      {stage0_10[478]},
      {stage1_10[277]}
   );
   gpc1_1 gpc2690 (
      {stage0_10[479]},
      {stage1_10[278]}
   );
   gpc1_1 gpc2691 (
      {stage0_10[480]},
      {stage1_10[279]}
   );
   gpc1_1 gpc2692 (
      {stage0_10[481]},
      {stage1_10[280]}
   );
   gpc1_1 gpc2693 (
      {stage0_10[482]},
      {stage1_10[281]}
   );
   gpc1_1 gpc2694 (
      {stage0_10[483]},
      {stage1_10[282]}
   );
   gpc1_1 gpc2695 (
      {stage0_10[484]},
      {stage1_10[283]}
   );
   gpc1_1 gpc2696 (
      {stage0_10[485]},
      {stage1_10[284]}
   );
   gpc1_1 gpc2697 (
      {stage0_11[367]},
      {stage1_11[158]}
   );
   gpc1_1 gpc2698 (
      {stage0_11[368]},
      {stage1_11[159]}
   );
   gpc1_1 gpc2699 (
      {stage0_11[369]},
      {stage1_11[160]}
   );
   gpc1_1 gpc2700 (
      {stage0_11[370]},
      {stage1_11[161]}
   );
   gpc1_1 gpc2701 (
      {stage0_11[371]},
      {stage1_11[162]}
   );
   gpc1_1 gpc2702 (
      {stage0_11[372]},
      {stage1_11[163]}
   );
   gpc1_1 gpc2703 (
      {stage0_11[373]},
      {stage1_11[164]}
   );
   gpc1_1 gpc2704 (
      {stage0_11[374]},
      {stage1_11[165]}
   );
   gpc1_1 gpc2705 (
      {stage0_11[375]},
      {stage1_11[166]}
   );
   gpc1_1 gpc2706 (
      {stage0_11[376]},
      {stage1_11[167]}
   );
   gpc1_1 gpc2707 (
      {stage0_11[377]},
      {stage1_11[168]}
   );
   gpc1_1 gpc2708 (
      {stage0_11[378]},
      {stage1_11[169]}
   );
   gpc1_1 gpc2709 (
      {stage0_11[379]},
      {stage1_11[170]}
   );
   gpc1_1 gpc2710 (
      {stage0_11[380]},
      {stage1_11[171]}
   );
   gpc1_1 gpc2711 (
      {stage0_11[381]},
      {stage1_11[172]}
   );
   gpc1_1 gpc2712 (
      {stage0_11[382]},
      {stage1_11[173]}
   );
   gpc1_1 gpc2713 (
      {stage0_11[383]},
      {stage1_11[174]}
   );
   gpc1_1 gpc2714 (
      {stage0_11[384]},
      {stage1_11[175]}
   );
   gpc1_1 gpc2715 (
      {stage0_11[385]},
      {stage1_11[176]}
   );
   gpc1_1 gpc2716 (
      {stage0_11[386]},
      {stage1_11[177]}
   );
   gpc1_1 gpc2717 (
      {stage0_11[387]},
      {stage1_11[178]}
   );
   gpc1_1 gpc2718 (
      {stage0_11[388]},
      {stage1_11[179]}
   );
   gpc1_1 gpc2719 (
      {stage0_11[389]},
      {stage1_11[180]}
   );
   gpc1_1 gpc2720 (
      {stage0_11[390]},
      {stage1_11[181]}
   );
   gpc1_1 gpc2721 (
      {stage0_11[391]},
      {stage1_11[182]}
   );
   gpc1_1 gpc2722 (
      {stage0_11[392]},
      {stage1_11[183]}
   );
   gpc1_1 gpc2723 (
      {stage0_11[393]},
      {stage1_11[184]}
   );
   gpc1_1 gpc2724 (
      {stage0_11[394]},
      {stage1_11[185]}
   );
   gpc1_1 gpc2725 (
      {stage0_11[395]},
      {stage1_11[186]}
   );
   gpc1_1 gpc2726 (
      {stage0_11[396]},
      {stage1_11[187]}
   );
   gpc1_1 gpc2727 (
      {stage0_11[397]},
      {stage1_11[188]}
   );
   gpc1_1 gpc2728 (
      {stage0_11[398]},
      {stage1_11[189]}
   );
   gpc1_1 gpc2729 (
      {stage0_11[399]},
      {stage1_11[190]}
   );
   gpc1_1 gpc2730 (
      {stage0_11[400]},
      {stage1_11[191]}
   );
   gpc1_1 gpc2731 (
      {stage0_11[401]},
      {stage1_11[192]}
   );
   gpc1_1 gpc2732 (
      {stage0_11[402]},
      {stage1_11[193]}
   );
   gpc1_1 gpc2733 (
      {stage0_11[403]},
      {stage1_11[194]}
   );
   gpc1_1 gpc2734 (
      {stage0_11[404]},
      {stage1_11[195]}
   );
   gpc1_1 gpc2735 (
      {stage0_11[405]},
      {stage1_11[196]}
   );
   gpc1_1 gpc2736 (
      {stage0_11[406]},
      {stage1_11[197]}
   );
   gpc1_1 gpc2737 (
      {stage0_11[407]},
      {stage1_11[198]}
   );
   gpc1_1 gpc2738 (
      {stage0_11[408]},
      {stage1_11[199]}
   );
   gpc1_1 gpc2739 (
      {stage0_11[409]},
      {stage1_11[200]}
   );
   gpc1_1 gpc2740 (
      {stage0_11[410]},
      {stage1_11[201]}
   );
   gpc1_1 gpc2741 (
      {stage0_11[411]},
      {stage1_11[202]}
   );
   gpc1_1 gpc2742 (
      {stage0_11[412]},
      {stage1_11[203]}
   );
   gpc1_1 gpc2743 (
      {stage0_11[413]},
      {stage1_11[204]}
   );
   gpc1_1 gpc2744 (
      {stage0_11[414]},
      {stage1_11[205]}
   );
   gpc1_1 gpc2745 (
      {stage0_11[415]},
      {stage1_11[206]}
   );
   gpc1_1 gpc2746 (
      {stage0_11[416]},
      {stage1_11[207]}
   );
   gpc1_1 gpc2747 (
      {stage0_11[417]},
      {stage1_11[208]}
   );
   gpc1_1 gpc2748 (
      {stage0_11[418]},
      {stage1_11[209]}
   );
   gpc1_1 gpc2749 (
      {stage0_11[419]},
      {stage1_11[210]}
   );
   gpc1_1 gpc2750 (
      {stage0_11[420]},
      {stage1_11[211]}
   );
   gpc1_1 gpc2751 (
      {stage0_11[421]},
      {stage1_11[212]}
   );
   gpc1_1 gpc2752 (
      {stage0_11[422]},
      {stage1_11[213]}
   );
   gpc1_1 gpc2753 (
      {stage0_11[423]},
      {stage1_11[214]}
   );
   gpc1_1 gpc2754 (
      {stage0_11[424]},
      {stage1_11[215]}
   );
   gpc1_1 gpc2755 (
      {stage0_11[425]},
      {stage1_11[216]}
   );
   gpc1_1 gpc2756 (
      {stage0_11[426]},
      {stage1_11[217]}
   );
   gpc1_1 gpc2757 (
      {stage0_11[427]},
      {stage1_11[218]}
   );
   gpc1_1 gpc2758 (
      {stage0_11[428]},
      {stage1_11[219]}
   );
   gpc1_1 gpc2759 (
      {stage0_11[429]},
      {stage1_11[220]}
   );
   gpc1_1 gpc2760 (
      {stage0_11[430]},
      {stage1_11[221]}
   );
   gpc1_1 gpc2761 (
      {stage0_11[431]},
      {stage1_11[222]}
   );
   gpc1_1 gpc2762 (
      {stage0_11[432]},
      {stage1_11[223]}
   );
   gpc1_1 gpc2763 (
      {stage0_11[433]},
      {stage1_11[224]}
   );
   gpc1_1 gpc2764 (
      {stage0_11[434]},
      {stage1_11[225]}
   );
   gpc1_1 gpc2765 (
      {stage0_11[435]},
      {stage1_11[226]}
   );
   gpc1_1 gpc2766 (
      {stage0_11[436]},
      {stage1_11[227]}
   );
   gpc1_1 gpc2767 (
      {stage0_11[437]},
      {stage1_11[228]}
   );
   gpc1_1 gpc2768 (
      {stage0_11[438]},
      {stage1_11[229]}
   );
   gpc1_1 gpc2769 (
      {stage0_11[439]},
      {stage1_11[230]}
   );
   gpc1_1 gpc2770 (
      {stage0_11[440]},
      {stage1_11[231]}
   );
   gpc1_1 gpc2771 (
      {stage0_11[441]},
      {stage1_11[232]}
   );
   gpc1_1 gpc2772 (
      {stage0_11[442]},
      {stage1_11[233]}
   );
   gpc1_1 gpc2773 (
      {stage0_11[443]},
      {stage1_11[234]}
   );
   gpc1_1 gpc2774 (
      {stage0_11[444]},
      {stage1_11[235]}
   );
   gpc1_1 gpc2775 (
      {stage0_11[445]},
      {stage1_11[236]}
   );
   gpc1_1 gpc2776 (
      {stage0_11[446]},
      {stage1_11[237]}
   );
   gpc1_1 gpc2777 (
      {stage0_11[447]},
      {stage1_11[238]}
   );
   gpc1_1 gpc2778 (
      {stage0_11[448]},
      {stage1_11[239]}
   );
   gpc1_1 gpc2779 (
      {stage0_11[449]},
      {stage1_11[240]}
   );
   gpc1_1 gpc2780 (
      {stage0_11[450]},
      {stage1_11[241]}
   );
   gpc1_1 gpc2781 (
      {stage0_11[451]},
      {stage1_11[242]}
   );
   gpc1_1 gpc2782 (
      {stage0_11[452]},
      {stage1_11[243]}
   );
   gpc1_1 gpc2783 (
      {stage0_11[453]},
      {stage1_11[244]}
   );
   gpc1_1 gpc2784 (
      {stage0_11[454]},
      {stage1_11[245]}
   );
   gpc1_1 gpc2785 (
      {stage0_11[455]},
      {stage1_11[246]}
   );
   gpc1_1 gpc2786 (
      {stage0_11[456]},
      {stage1_11[247]}
   );
   gpc1_1 gpc2787 (
      {stage0_11[457]},
      {stage1_11[248]}
   );
   gpc1_1 gpc2788 (
      {stage0_11[458]},
      {stage1_11[249]}
   );
   gpc1_1 gpc2789 (
      {stage0_11[459]},
      {stage1_11[250]}
   );
   gpc1_1 gpc2790 (
      {stage0_11[460]},
      {stage1_11[251]}
   );
   gpc1_1 gpc2791 (
      {stage0_11[461]},
      {stage1_11[252]}
   );
   gpc1_1 gpc2792 (
      {stage0_11[462]},
      {stage1_11[253]}
   );
   gpc1_1 gpc2793 (
      {stage0_11[463]},
      {stage1_11[254]}
   );
   gpc1_1 gpc2794 (
      {stage0_11[464]},
      {stage1_11[255]}
   );
   gpc1_1 gpc2795 (
      {stage0_11[465]},
      {stage1_11[256]}
   );
   gpc1_1 gpc2796 (
      {stage0_11[466]},
      {stage1_11[257]}
   );
   gpc1_1 gpc2797 (
      {stage0_11[467]},
      {stage1_11[258]}
   );
   gpc1_1 gpc2798 (
      {stage0_11[468]},
      {stage1_11[259]}
   );
   gpc1_1 gpc2799 (
      {stage0_11[469]},
      {stage1_11[260]}
   );
   gpc1_1 gpc2800 (
      {stage0_11[470]},
      {stage1_11[261]}
   );
   gpc1_1 gpc2801 (
      {stage0_11[471]},
      {stage1_11[262]}
   );
   gpc1_1 gpc2802 (
      {stage0_11[472]},
      {stage1_11[263]}
   );
   gpc1_1 gpc2803 (
      {stage0_11[473]},
      {stage1_11[264]}
   );
   gpc1_1 gpc2804 (
      {stage0_11[474]},
      {stage1_11[265]}
   );
   gpc1_1 gpc2805 (
      {stage0_11[475]},
      {stage1_11[266]}
   );
   gpc1_1 gpc2806 (
      {stage0_11[476]},
      {stage1_11[267]}
   );
   gpc1_1 gpc2807 (
      {stage0_11[477]},
      {stage1_11[268]}
   );
   gpc1_1 gpc2808 (
      {stage0_11[478]},
      {stage1_11[269]}
   );
   gpc1_1 gpc2809 (
      {stage0_11[479]},
      {stage1_11[270]}
   );
   gpc1_1 gpc2810 (
      {stage0_11[480]},
      {stage1_11[271]}
   );
   gpc1_1 gpc2811 (
      {stage0_11[481]},
      {stage1_11[272]}
   );
   gpc1_1 gpc2812 (
      {stage0_11[482]},
      {stage1_11[273]}
   );
   gpc1_1 gpc2813 (
      {stage0_11[483]},
      {stage1_11[274]}
   );
   gpc1_1 gpc2814 (
      {stage0_11[484]},
      {stage1_11[275]}
   );
   gpc1_1 gpc2815 (
      {stage0_11[485]},
      {stage1_11[276]}
   );
   gpc1_1 gpc2816 (
      {stage0_12[484]},
      {stage1_12[187]}
   );
   gpc1_1 gpc2817 (
      {stage0_12[485]},
      {stage1_12[188]}
   );
   gpc1_1 gpc2818 (
      {stage0_13[376]},
      {stage1_13[195]}
   );
   gpc1_1 gpc2819 (
      {stage0_13[377]},
      {stage1_13[196]}
   );
   gpc1_1 gpc2820 (
      {stage0_13[378]},
      {stage1_13[197]}
   );
   gpc1_1 gpc2821 (
      {stage0_13[379]},
      {stage1_13[198]}
   );
   gpc1_1 gpc2822 (
      {stage0_13[380]},
      {stage1_13[199]}
   );
   gpc1_1 gpc2823 (
      {stage0_13[381]},
      {stage1_13[200]}
   );
   gpc1_1 gpc2824 (
      {stage0_13[382]},
      {stage1_13[201]}
   );
   gpc1_1 gpc2825 (
      {stage0_13[383]},
      {stage1_13[202]}
   );
   gpc1_1 gpc2826 (
      {stage0_13[384]},
      {stage1_13[203]}
   );
   gpc1_1 gpc2827 (
      {stage0_13[385]},
      {stage1_13[204]}
   );
   gpc1_1 gpc2828 (
      {stage0_13[386]},
      {stage1_13[205]}
   );
   gpc1_1 gpc2829 (
      {stage0_13[387]},
      {stage1_13[206]}
   );
   gpc1_1 gpc2830 (
      {stage0_13[388]},
      {stage1_13[207]}
   );
   gpc1_1 gpc2831 (
      {stage0_13[389]},
      {stage1_13[208]}
   );
   gpc1_1 gpc2832 (
      {stage0_13[390]},
      {stage1_13[209]}
   );
   gpc1_1 gpc2833 (
      {stage0_13[391]},
      {stage1_13[210]}
   );
   gpc1_1 gpc2834 (
      {stage0_13[392]},
      {stage1_13[211]}
   );
   gpc1_1 gpc2835 (
      {stage0_13[393]},
      {stage1_13[212]}
   );
   gpc1_1 gpc2836 (
      {stage0_13[394]},
      {stage1_13[213]}
   );
   gpc1_1 gpc2837 (
      {stage0_13[395]},
      {stage1_13[214]}
   );
   gpc1_1 gpc2838 (
      {stage0_13[396]},
      {stage1_13[215]}
   );
   gpc1_1 gpc2839 (
      {stage0_13[397]},
      {stage1_13[216]}
   );
   gpc1_1 gpc2840 (
      {stage0_13[398]},
      {stage1_13[217]}
   );
   gpc1_1 gpc2841 (
      {stage0_13[399]},
      {stage1_13[218]}
   );
   gpc1_1 gpc2842 (
      {stage0_13[400]},
      {stage1_13[219]}
   );
   gpc1_1 gpc2843 (
      {stage0_13[401]},
      {stage1_13[220]}
   );
   gpc1_1 gpc2844 (
      {stage0_13[402]},
      {stage1_13[221]}
   );
   gpc1_1 gpc2845 (
      {stage0_13[403]},
      {stage1_13[222]}
   );
   gpc1_1 gpc2846 (
      {stage0_13[404]},
      {stage1_13[223]}
   );
   gpc1_1 gpc2847 (
      {stage0_13[405]},
      {stage1_13[224]}
   );
   gpc1_1 gpc2848 (
      {stage0_13[406]},
      {stage1_13[225]}
   );
   gpc1_1 gpc2849 (
      {stage0_13[407]},
      {stage1_13[226]}
   );
   gpc1_1 gpc2850 (
      {stage0_13[408]},
      {stage1_13[227]}
   );
   gpc1_1 gpc2851 (
      {stage0_13[409]},
      {stage1_13[228]}
   );
   gpc1_1 gpc2852 (
      {stage0_13[410]},
      {stage1_13[229]}
   );
   gpc1_1 gpc2853 (
      {stage0_13[411]},
      {stage1_13[230]}
   );
   gpc1_1 gpc2854 (
      {stage0_13[412]},
      {stage1_13[231]}
   );
   gpc1_1 gpc2855 (
      {stage0_13[413]},
      {stage1_13[232]}
   );
   gpc1_1 gpc2856 (
      {stage0_13[414]},
      {stage1_13[233]}
   );
   gpc1_1 gpc2857 (
      {stage0_13[415]},
      {stage1_13[234]}
   );
   gpc1_1 gpc2858 (
      {stage0_13[416]},
      {stage1_13[235]}
   );
   gpc1_1 gpc2859 (
      {stage0_13[417]},
      {stage1_13[236]}
   );
   gpc1_1 gpc2860 (
      {stage0_13[418]},
      {stage1_13[237]}
   );
   gpc1_1 gpc2861 (
      {stage0_13[419]},
      {stage1_13[238]}
   );
   gpc1_1 gpc2862 (
      {stage0_13[420]},
      {stage1_13[239]}
   );
   gpc1_1 gpc2863 (
      {stage0_13[421]},
      {stage1_13[240]}
   );
   gpc1_1 gpc2864 (
      {stage0_13[422]},
      {stage1_13[241]}
   );
   gpc1_1 gpc2865 (
      {stage0_13[423]},
      {stage1_13[242]}
   );
   gpc1_1 gpc2866 (
      {stage0_13[424]},
      {stage1_13[243]}
   );
   gpc1_1 gpc2867 (
      {stage0_13[425]},
      {stage1_13[244]}
   );
   gpc1_1 gpc2868 (
      {stage0_13[426]},
      {stage1_13[245]}
   );
   gpc1_1 gpc2869 (
      {stage0_13[427]},
      {stage1_13[246]}
   );
   gpc1_1 gpc2870 (
      {stage0_13[428]},
      {stage1_13[247]}
   );
   gpc1_1 gpc2871 (
      {stage0_13[429]},
      {stage1_13[248]}
   );
   gpc1_1 gpc2872 (
      {stage0_13[430]},
      {stage1_13[249]}
   );
   gpc1_1 gpc2873 (
      {stage0_13[431]},
      {stage1_13[250]}
   );
   gpc1_1 gpc2874 (
      {stage0_13[432]},
      {stage1_13[251]}
   );
   gpc1_1 gpc2875 (
      {stage0_13[433]},
      {stage1_13[252]}
   );
   gpc1_1 gpc2876 (
      {stage0_13[434]},
      {stage1_13[253]}
   );
   gpc1_1 gpc2877 (
      {stage0_13[435]},
      {stage1_13[254]}
   );
   gpc1_1 gpc2878 (
      {stage0_13[436]},
      {stage1_13[255]}
   );
   gpc1_1 gpc2879 (
      {stage0_13[437]},
      {stage1_13[256]}
   );
   gpc1_1 gpc2880 (
      {stage0_13[438]},
      {stage1_13[257]}
   );
   gpc1_1 gpc2881 (
      {stage0_13[439]},
      {stage1_13[258]}
   );
   gpc1_1 gpc2882 (
      {stage0_13[440]},
      {stage1_13[259]}
   );
   gpc1_1 gpc2883 (
      {stage0_13[441]},
      {stage1_13[260]}
   );
   gpc1_1 gpc2884 (
      {stage0_13[442]},
      {stage1_13[261]}
   );
   gpc1_1 gpc2885 (
      {stage0_13[443]},
      {stage1_13[262]}
   );
   gpc1_1 gpc2886 (
      {stage0_13[444]},
      {stage1_13[263]}
   );
   gpc1_1 gpc2887 (
      {stage0_13[445]},
      {stage1_13[264]}
   );
   gpc1_1 gpc2888 (
      {stage0_13[446]},
      {stage1_13[265]}
   );
   gpc1_1 gpc2889 (
      {stage0_13[447]},
      {stage1_13[266]}
   );
   gpc1_1 gpc2890 (
      {stage0_13[448]},
      {stage1_13[267]}
   );
   gpc1_1 gpc2891 (
      {stage0_13[449]},
      {stage1_13[268]}
   );
   gpc1_1 gpc2892 (
      {stage0_13[450]},
      {stage1_13[269]}
   );
   gpc1_1 gpc2893 (
      {stage0_13[451]},
      {stage1_13[270]}
   );
   gpc1_1 gpc2894 (
      {stage0_13[452]},
      {stage1_13[271]}
   );
   gpc1_1 gpc2895 (
      {stage0_13[453]},
      {stage1_13[272]}
   );
   gpc1_1 gpc2896 (
      {stage0_13[454]},
      {stage1_13[273]}
   );
   gpc1_1 gpc2897 (
      {stage0_13[455]},
      {stage1_13[274]}
   );
   gpc1_1 gpc2898 (
      {stage0_13[456]},
      {stage1_13[275]}
   );
   gpc1_1 gpc2899 (
      {stage0_13[457]},
      {stage1_13[276]}
   );
   gpc1_1 gpc2900 (
      {stage0_13[458]},
      {stage1_13[277]}
   );
   gpc1_1 gpc2901 (
      {stage0_13[459]},
      {stage1_13[278]}
   );
   gpc1_1 gpc2902 (
      {stage0_13[460]},
      {stage1_13[279]}
   );
   gpc1_1 gpc2903 (
      {stage0_13[461]},
      {stage1_13[280]}
   );
   gpc1_1 gpc2904 (
      {stage0_13[462]},
      {stage1_13[281]}
   );
   gpc1_1 gpc2905 (
      {stage0_13[463]},
      {stage1_13[282]}
   );
   gpc1_1 gpc2906 (
      {stage0_13[464]},
      {stage1_13[283]}
   );
   gpc1_1 gpc2907 (
      {stage0_13[465]},
      {stage1_13[284]}
   );
   gpc1_1 gpc2908 (
      {stage0_13[466]},
      {stage1_13[285]}
   );
   gpc1_1 gpc2909 (
      {stage0_13[467]},
      {stage1_13[286]}
   );
   gpc1_1 gpc2910 (
      {stage0_13[468]},
      {stage1_13[287]}
   );
   gpc1_1 gpc2911 (
      {stage0_13[469]},
      {stage1_13[288]}
   );
   gpc1_1 gpc2912 (
      {stage0_13[470]},
      {stage1_13[289]}
   );
   gpc1_1 gpc2913 (
      {stage0_13[471]},
      {stage1_13[290]}
   );
   gpc1_1 gpc2914 (
      {stage0_13[472]},
      {stage1_13[291]}
   );
   gpc1_1 gpc2915 (
      {stage0_13[473]},
      {stage1_13[292]}
   );
   gpc1_1 gpc2916 (
      {stage0_13[474]},
      {stage1_13[293]}
   );
   gpc1_1 gpc2917 (
      {stage0_13[475]},
      {stage1_13[294]}
   );
   gpc1_1 gpc2918 (
      {stage0_13[476]},
      {stage1_13[295]}
   );
   gpc1_1 gpc2919 (
      {stage0_13[477]},
      {stage1_13[296]}
   );
   gpc1_1 gpc2920 (
      {stage0_13[478]},
      {stage1_13[297]}
   );
   gpc1_1 gpc2921 (
      {stage0_13[479]},
      {stage1_13[298]}
   );
   gpc1_1 gpc2922 (
      {stage0_13[480]},
      {stage1_13[299]}
   );
   gpc1_1 gpc2923 (
      {stage0_13[481]},
      {stage1_13[300]}
   );
   gpc1_1 gpc2924 (
      {stage0_13[482]},
      {stage1_13[301]}
   );
   gpc1_1 gpc2925 (
      {stage0_13[483]},
      {stage1_13[302]}
   );
   gpc1_1 gpc2926 (
      {stage0_13[484]},
      {stage1_13[303]}
   );
   gpc1_1 gpc2927 (
      {stage0_13[485]},
      {stage1_13[304]}
   );
   gpc1_1 gpc2928 (
      {stage0_14[419]},
      {stage1_14[152]}
   );
   gpc1_1 gpc2929 (
      {stage0_14[420]},
      {stage1_14[153]}
   );
   gpc1_1 gpc2930 (
      {stage0_14[421]},
      {stage1_14[154]}
   );
   gpc1_1 gpc2931 (
      {stage0_14[422]},
      {stage1_14[155]}
   );
   gpc1_1 gpc2932 (
      {stage0_14[423]},
      {stage1_14[156]}
   );
   gpc1_1 gpc2933 (
      {stage0_14[424]},
      {stage1_14[157]}
   );
   gpc1_1 gpc2934 (
      {stage0_14[425]},
      {stage1_14[158]}
   );
   gpc1_1 gpc2935 (
      {stage0_14[426]},
      {stage1_14[159]}
   );
   gpc1_1 gpc2936 (
      {stage0_14[427]},
      {stage1_14[160]}
   );
   gpc1_1 gpc2937 (
      {stage0_14[428]},
      {stage1_14[161]}
   );
   gpc1_1 gpc2938 (
      {stage0_14[429]},
      {stage1_14[162]}
   );
   gpc1_1 gpc2939 (
      {stage0_14[430]},
      {stage1_14[163]}
   );
   gpc1_1 gpc2940 (
      {stage0_14[431]},
      {stage1_14[164]}
   );
   gpc1_1 gpc2941 (
      {stage0_14[432]},
      {stage1_14[165]}
   );
   gpc1_1 gpc2942 (
      {stage0_14[433]},
      {stage1_14[166]}
   );
   gpc1_1 gpc2943 (
      {stage0_14[434]},
      {stage1_14[167]}
   );
   gpc1_1 gpc2944 (
      {stage0_14[435]},
      {stage1_14[168]}
   );
   gpc1_1 gpc2945 (
      {stage0_14[436]},
      {stage1_14[169]}
   );
   gpc1_1 gpc2946 (
      {stage0_14[437]},
      {stage1_14[170]}
   );
   gpc1_1 gpc2947 (
      {stage0_14[438]},
      {stage1_14[171]}
   );
   gpc1_1 gpc2948 (
      {stage0_14[439]},
      {stage1_14[172]}
   );
   gpc1_1 gpc2949 (
      {stage0_14[440]},
      {stage1_14[173]}
   );
   gpc1_1 gpc2950 (
      {stage0_14[441]},
      {stage1_14[174]}
   );
   gpc1_1 gpc2951 (
      {stage0_14[442]},
      {stage1_14[175]}
   );
   gpc1_1 gpc2952 (
      {stage0_14[443]},
      {stage1_14[176]}
   );
   gpc1_1 gpc2953 (
      {stage0_14[444]},
      {stage1_14[177]}
   );
   gpc1_1 gpc2954 (
      {stage0_14[445]},
      {stage1_14[178]}
   );
   gpc1_1 gpc2955 (
      {stage0_14[446]},
      {stage1_14[179]}
   );
   gpc1_1 gpc2956 (
      {stage0_14[447]},
      {stage1_14[180]}
   );
   gpc1_1 gpc2957 (
      {stage0_14[448]},
      {stage1_14[181]}
   );
   gpc1_1 gpc2958 (
      {stage0_14[449]},
      {stage1_14[182]}
   );
   gpc1_1 gpc2959 (
      {stage0_14[450]},
      {stage1_14[183]}
   );
   gpc1_1 gpc2960 (
      {stage0_14[451]},
      {stage1_14[184]}
   );
   gpc1_1 gpc2961 (
      {stage0_14[452]},
      {stage1_14[185]}
   );
   gpc1_1 gpc2962 (
      {stage0_14[453]},
      {stage1_14[186]}
   );
   gpc1_1 gpc2963 (
      {stage0_14[454]},
      {stage1_14[187]}
   );
   gpc1_1 gpc2964 (
      {stage0_14[455]},
      {stage1_14[188]}
   );
   gpc1_1 gpc2965 (
      {stage0_14[456]},
      {stage1_14[189]}
   );
   gpc1_1 gpc2966 (
      {stage0_14[457]},
      {stage1_14[190]}
   );
   gpc1_1 gpc2967 (
      {stage0_14[458]},
      {stage1_14[191]}
   );
   gpc1_1 gpc2968 (
      {stage0_14[459]},
      {stage1_14[192]}
   );
   gpc1_1 gpc2969 (
      {stage0_14[460]},
      {stage1_14[193]}
   );
   gpc1_1 gpc2970 (
      {stage0_14[461]},
      {stage1_14[194]}
   );
   gpc1_1 gpc2971 (
      {stage0_14[462]},
      {stage1_14[195]}
   );
   gpc1_1 gpc2972 (
      {stage0_14[463]},
      {stage1_14[196]}
   );
   gpc1_1 gpc2973 (
      {stage0_14[464]},
      {stage1_14[197]}
   );
   gpc1_1 gpc2974 (
      {stage0_14[465]},
      {stage1_14[198]}
   );
   gpc1_1 gpc2975 (
      {stage0_14[466]},
      {stage1_14[199]}
   );
   gpc1_1 gpc2976 (
      {stage0_14[467]},
      {stage1_14[200]}
   );
   gpc1_1 gpc2977 (
      {stage0_14[468]},
      {stage1_14[201]}
   );
   gpc1_1 gpc2978 (
      {stage0_14[469]},
      {stage1_14[202]}
   );
   gpc1_1 gpc2979 (
      {stage0_14[470]},
      {stage1_14[203]}
   );
   gpc1_1 gpc2980 (
      {stage0_14[471]},
      {stage1_14[204]}
   );
   gpc1_1 gpc2981 (
      {stage0_14[472]},
      {stage1_14[205]}
   );
   gpc1_1 gpc2982 (
      {stage0_14[473]},
      {stage1_14[206]}
   );
   gpc1_1 gpc2983 (
      {stage0_14[474]},
      {stage1_14[207]}
   );
   gpc1_1 gpc2984 (
      {stage0_14[475]},
      {stage1_14[208]}
   );
   gpc1_1 gpc2985 (
      {stage0_14[476]},
      {stage1_14[209]}
   );
   gpc1_1 gpc2986 (
      {stage0_14[477]},
      {stage1_14[210]}
   );
   gpc1_1 gpc2987 (
      {stage0_14[478]},
      {stage1_14[211]}
   );
   gpc1_1 gpc2988 (
      {stage0_14[479]},
      {stage1_14[212]}
   );
   gpc1_1 gpc2989 (
      {stage0_14[480]},
      {stage1_14[213]}
   );
   gpc1_1 gpc2990 (
      {stage0_14[481]},
      {stage1_14[214]}
   );
   gpc1_1 gpc2991 (
      {stage0_14[482]},
      {stage1_14[215]}
   );
   gpc1_1 gpc2992 (
      {stage0_14[483]},
      {stage1_14[216]}
   );
   gpc1_1 gpc2993 (
      {stage0_14[484]},
      {stage1_14[217]}
   );
   gpc1_1 gpc2994 (
      {stage0_14[485]},
      {stage1_14[218]}
   );
   gpc1_1 gpc2995 (
      {stage0_15[479]},
      {stage1_15[164]}
   );
   gpc1_1 gpc2996 (
      {stage0_15[480]},
      {stage1_15[165]}
   );
   gpc1_1 gpc2997 (
      {stage0_15[481]},
      {stage1_15[166]}
   );
   gpc1_1 gpc2998 (
      {stage0_15[482]},
      {stage1_15[167]}
   );
   gpc1_1 gpc2999 (
      {stage0_15[483]},
      {stage1_15[168]}
   );
   gpc1_1 gpc3000 (
      {stage0_15[484]},
      {stage1_15[169]}
   );
   gpc1_1 gpc3001 (
      {stage0_15[485]},
      {stage1_15[170]}
   );
   gpc1_1 gpc3002 (
      {stage0_17[450]},
      {stage1_17[193]}
   );
   gpc1_1 gpc3003 (
      {stage0_17[451]},
      {stage1_17[194]}
   );
   gpc1_1 gpc3004 (
      {stage0_17[452]},
      {stage1_17[195]}
   );
   gpc1_1 gpc3005 (
      {stage0_17[453]},
      {stage1_17[196]}
   );
   gpc1_1 gpc3006 (
      {stage0_17[454]},
      {stage1_17[197]}
   );
   gpc1_1 gpc3007 (
      {stage0_17[455]},
      {stage1_17[198]}
   );
   gpc1_1 gpc3008 (
      {stage0_17[456]},
      {stage1_17[199]}
   );
   gpc1_1 gpc3009 (
      {stage0_17[457]},
      {stage1_17[200]}
   );
   gpc1_1 gpc3010 (
      {stage0_17[458]},
      {stage1_17[201]}
   );
   gpc1_1 gpc3011 (
      {stage0_17[459]},
      {stage1_17[202]}
   );
   gpc1_1 gpc3012 (
      {stage0_17[460]},
      {stage1_17[203]}
   );
   gpc1_1 gpc3013 (
      {stage0_17[461]},
      {stage1_17[204]}
   );
   gpc1_1 gpc3014 (
      {stage0_17[462]},
      {stage1_17[205]}
   );
   gpc1_1 gpc3015 (
      {stage0_17[463]},
      {stage1_17[206]}
   );
   gpc1_1 gpc3016 (
      {stage0_17[464]},
      {stage1_17[207]}
   );
   gpc1_1 gpc3017 (
      {stage0_17[465]},
      {stage1_17[208]}
   );
   gpc1_1 gpc3018 (
      {stage0_17[466]},
      {stage1_17[209]}
   );
   gpc1_1 gpc3019 (
      {stage0_17[467]},
      {stage1_17[210]}
   );
   gpc1_1 gpc3020 (
      {stage0_17[468]},
      {stage1_17[211]}
   );
   gpc1_1 gpc3021 (
      {stage0_17[469]},
      {stage1_17[212]}
   );
   gpc1_1 gpc3022 (
      {stage0_17[470]},
      {stage1_17[213]}
   );
   gpc1_1 gpc3023 (
      {stage0_17[471]},
      {stage1_17[214]}
   );
   gpc1_1 gpc3024 (
      {stage0_17[472]},
      {stage1_17[215]}
   );
   gpc1_1 gpc3025 (
      {stage0_17[473]},
      {stage1_17[216]}
   );
   gpc1_1 gpc3026 (
      {stage0_17[474]},
      {stage1_17[217]}
   );
   gpc1_1 gpc3027 (
      {stage0_17[475]},
      {stage1_17[218]}
   );
   gpc1_1 gpc3028 (
      {stage0_17[476]},
      {stage1_17[219]}
   );
   gpc1_1 gpc3029 (
      {stage0_17[477]},
      {stage1_17[220]}
   );
   gpc1_1 gpc3030 (
      {stage0_17[478]},
      {stage1_17[221]}
   );
   gpc1_1 gpc3031 (
      {stage0_17[479]},
      {stage1_17[222]}
   );
   gpc1_1 gpc3032 (
      {stage0_17[480]},
      {stage1_17[223]}
   );
   gpc1_1 gpc3033 (
      {stage0_17[481]},
      {stage1_17[224]}
   );
   gpc1_1 gpc3034 (
      {stage0_17[482]},
      {stage1_17[225]}
   );
   gpc1_1 gpc3035 (
      {stage0_17[483]},
      {stage1_17[226]}
   );
   gpc1_1 gpc3036 (
      {stage0_17[484]},
      {stage1_17[227]}
   );
   gpc1_1 gpc3037 (
      {stage0_17[485]},
      {stage1_17[228]}
   );
   gpc1_1 gpc3038 (
      {stage0_18[426]},
      {stage1_18[149]}
   );
   gpc1_1 gpc3039 (
      {stage0_18[427]},
      {stage1_18[150]}
   );
   gpc1_1 gpc3040 (
      {stage0_18[428]},
      {stage1_18[151]}
   );
   gpc1_1 gpc3041 (
      {stage0_18[429]},
      {stage1_18[152]}
   );
   gpc1_1 gpc3042 (
      {stage0_18[430]},
      {stage1_18[153]}
   );
   gpc1_1 gpc3043 (
      {stage0_18[431]},
      {stage1_18[154]}
   );
   gpc1_1 gpc3044 (
      {stage0_18[432]},
      {stage1_18[155]}
   );
   gpc1_1 gpc3045 (
      {stage0_18[433]},
      {stage1_18[156]}
   );
   gpc1_1 gpc3046 (
      {stage0_18[434]},
      {stage1_18[157]}
   );
   gpc1_1 gpc3047 (
      {stage0_18[435]},
      {stage1_18[158]}
   );
   gpc1_1 gpc3048 (
      {stage0_18[436]},
      {stage1_18[159]}
   );
   gpc1_1 gpc3049 (
      {stage0_18[437]},
      {stage1_18[160]}
   );
   gpc1_1 gpc3050 (
      {stage0_18[438]},
      {stage1_18[161]}
   );
   gpc1_1 gpc3051 (
      {stage0_18[439]},
      {stage1_18[162]}
   );
   gpc1_1 gpc3052 (
      {stage0_18[440]},
      {stage1_18[163]}
   );
   gpc1_1 gpc3053 (
      {stage0_18[441]},
      {stage1_18[164]}
   );
   gpc1_1 gpc3054 (
      {stage0_18[442]},
      {stage1_18[165]}
   );
   gpc1_1 gpc3055 (
      {stage0_18[443]},
      {stage1_18[166]}
   );
   gpc1_1 gpc3056 (
      {stage0_18[444]},
      {stage1_18[167]}
   );
   gpc1_1 gpc3057 (
      {stage0_18[445]},
      {stage1_18[168]}
   );
   gpc1_1 gpc3058 (
      {stage0_18[446]},
      {stage1_18[169]}
   );
   gpc1_1 gpc3059 (
      {stage0_18[447]},
      {stage1_18[170]}
   );
   gpc1_1 gpc3060 (
      {stage0_18[448]},
      {stage1_18[171]}
   );
   gpc1_1 gpc3061 (
      {stage0_18[449]},
      {stage1_18[172]}
   );
   gpc1_1 gpc3062 (
      {stage0_18[450]},
      {stage1_18[173]}
   );
   gpc1_1 gpc3063 (
      {stage0_18[451]},
      {stage1_18[174]}
   );
   gpc1_1 gpc3064 (
      {stage0_18[452]},
      {stage1_18[175]}
   );
   gpc1_1 gpc3065 (
      {stage0_18[453]},
      {stage1_18[176]}
   );
   gpc1_1 gpc3066 (
      {stage0_18[454]},
      {stage1_18[177]}
   );
   gpc1_1 gpc3067 (
      {stage0_18[455]},
      {stage1_18[178]}
   );
   gpc1_1 gpc3068 (
      {stage0_18[456]},
      {stage1_18[179]}
   );
   gpc1_1 gpc3069 (
      {stage0_18[457]},
      {stage1_18[180]}
   );
   gpc1_1 gpc3070 (
      {stage0_18[458]},
      {stage1_18[181]}
   );
   gpc1_1 gpc3071 (
      {stage0_18[459]},
      {stage1_18[182]}
   );
   gpc1_1 gpc3072 (
      {stage0_18[460]},
      {stage1_18[183]}
   );
   gpc1_1 gpc3073 (
      {stage0_18[461]},
      {stage1_18[184]}
   );
   gpc1_1 gpc3074 (
      {stage0_18[462]},
      {stage1_18[185]}
   );
   gpc1_1 gpc3075 (
      {stage0_18[463]},
      {stage1_18[186]}
   );
   gpc1_1 gpc3076 (
      {stage0_18[464]},
      {stage1_18[187]}
   );
   gpc1_1 gpc3077 (
      {stage0_18[465]},
      {stage1_18[188]}
   );
   gpc1_1 gpc3078 (
      {stage0_18[466]},
      {stage1_18[189]}
   );
   gpc1_1 gpc3079 (
      {stage0_18[467]},
      {stage1_18[190]}
   );
   gpc1_1 gpc3080 (
      {stage0_18[468]},
      {stage1_18[191]}
   );
   gpc1_1 gpc3081 (
      {stage0_18[469]},
      {stage1_18[192]}
   );
   gpc1_1 gpc3082 (
      {stage0_18[470]},
      {stage1_18[193]}
   );
   gpc1_1 gpc3083 (
      {stage0_18[471]},
      {stage1_18[194]}
   );
   gpc1_1 gpc3084 (
      {stage0_18[472]},
      {stage1_18[195]}
   );
   gpc1_1 gpc3085 (
      {stage0_18[473]},
      {stage1_18[196]}
   );
   gpc1_1 gpc3086 (
      {stage0_18[474]},
      {stage1_18[197]}
   );
   gpc1_1 gpc3087 (
      {stage0_18[475]},
      {stage1_18[198]}
   );
   gpc1_1 gpc3088 (
      {stage0_18[476]},
      {stage1_18[199]}
   );
   gpc1_1 gpc3089 (
      {stage0_18[477]},
      {stage1_18[200]}
   );
   gpc1_1 gpc3090 (
      {stage0_18[478]},
      {stage1_18[201]}
   );
   gpc1_1 gpc3091 (
      {stage0_18[479]},
      {stage1_18[202]}
   );
   gpc1_1 gpc3092 (
      {stage0_18[480]},
      {stage1_18[203]}
   );
   gpc1_1 gpc3093 (
      {stage0_18[481]},
      {stage1_18[204]}
   );
   gpc1_1 gpc3094 (
      {stage0_18[482]},
      {stage1_18[205]}
   );
   gpc1_1 gpc3095 (
      {stage0_18[483]},
      {stage1_18[206]}
   );
   gpc1_1 gpc3096 (
      {stage0_18[484]},
      {stage1_18[207]}
   );
   gpc1_1 gpc3097 (
      {stage0_18[485]},
      {stage1_18[208]}
   );
   gpc1_1 gpc3098 (
      {stage0_19[397]},
      {stage1_19[187]}
   );
   gpc1_1 gpc3099 (
      {stage0_19[398]},
      {stage1_19[188]}
   );
   gpc1_1 gpc3100 (
      {stage0_19[399]},
      {stage1_19[189]}
   );
   gpc1_1 gpc3101 (
      {stage0_19[400]},
      {stage1_19[190]}
   );
   gpc1_1 gpc3102 (
      {stage0_19[401]},
      {stage1_19[191]}
   );
   gpc1_1 gpc3103 (
      {stage0_19[402]},
      {stage1_19[192]}
   );
   gpc1_1 gpc3104 (
      {stage0_19[403]},
      {stage1_19[193]}
   );
   gpc1_1 gpc3105 (
      {stage0_19[404]},
      {stage1_19[194]}
   );
   gpc1_1 gpc3106 (
      {stage0_19[405]},
      {stage1_19[195]}
   );
   gpc1_1 gpc3107 (
      {stage0_19[406]},
      {stage1_19[196]}
   );
   gpc1_1 gpc3108 (
      {stage0_19[407]},
      {stage1_19[197]}
   );
   gpc1_1 gpc3109 (
      {stage0_19[408]},
      {stage1_19[198]}
   );
   gpc1_1 gpc3110 (
      {stage0_19[409]},
      {stage1_19[199]}
   );
   gpc1_1 gpc3111 (
      {stage0_19[410]},
      {stage1_19[200]}
   );
   gpc1_1 gpc3112 (
      {stage0_19[411]},
      {stage1_19[201]}
   );
   gpc1_1 gpc3113 (
      {stage0_19[412]},
      {stage1_19[202]}
   );
   gpc1_1 gpc3114 (
      {stage0_19[413]},
      {stage1_19[203]}
   );
   gpc1_1 gpc3115 (
      {stage0_19[414]},
      {stage1_19[204]}
   );
   gpc1_1 gpc3116 (
      {stage0_19[415]},
      {stage1_19[205]}
   );
   gpc1_1 gpc3117 (
      {stage0_19[416]},
      {stage1_19[206]}
   );
   gpc1_1 gpc3118 (
      {stage0_19[417]},
      {stage1_19[207]}
   );
   gpc1_1 gpc3119 (
      {stage0_19[418]},
      {stage1_19[208]}
   );
   gpc1_1 gpc3120 (
      {stage0_19[419]},
      {stage1_19[209]}
   );
   gpc1_1 gpc3121 (
      {stage0_19[420]},
      {stage1_19[210]}
   );
   gpc1_1 gpc3122 (
      {stage0_19[421]},
      {stage1_19[211]}
   );
   gpc1_1 gpc3123 (
      {stage0_19[422]},
      {stage1_19[212]}
   );
   gpc1_1 gpc3124 (
      {stage0_19[423]},
      {stage1_19[213]}
   );
   gpc1_1 gpc3125 (
      {stage0_19[424]},
      {stage1_19[214]}
   );
   gpc1_1 gpc3126 (
      {stage0_19[425]},
      {stage1_19[215]}
   );
   gpc1_1 gpc3127 (
      {stage0_19[426]},
      {stage1_19[216]}
   );
   gpc1_1 gpc3128 (
      {stage0_19[427]},
      {stage1_19[217]}
   );
   gpc1_1 gpc3129 (
      {stage0_19[428]},
      {stage1_19[218]}
   );
   gpc1_1 gpc3130 (
      {stage0_19[429]},
      {stage1_19[219]}
   );
   gpc1_1 gpc3131 (
      {stage0_19[430]},
      {stage1_19[220]}
   );
   gpc1_1 gpc3132 (
      {stage0_19[431]},
      {stage1_19[221]}
   );
   gpc1_1 gpc3133 (
      {stage0_19[432]},
      {stage1_19[222]}
   );
   gpc1_1 gpc3134 (
      {stage0_19[433]},
      {stage1_19[223]}
   );
   gpc1_1 gpc3135 (
      {stage0_19[434]},
      {stage1_19[224]}
   );
   gpc1_1 gpc3136 (
      {stage0_19[435]},
      {stage1_19[225]}
   );
   gpc1_1 gpc3137 (
      {stage0_19[436]},
      {stage1_19[226]}
   );
   gpc1_1 gpc3138 (
      {stage0_19[437]},
      {stage1_19[227]}
   );
   gpc1_1 gpc3139 (
      {stage0_19[438]},
      {stage1_19[228]}
   );
   gpc1_1 gpc3140 (
      {stage0_19[439]},
      {stage1_19[229]}
   );
   gpc1_1 gpc3141 (
      {stage0_19[440]},
      {stage1_19[230]}
   );
   gpc1_1 gpc3142 (
      {stage0_19[441]},
      {stage1_19[231]}
   );
   gpc1_1 gpc3143 (
      {stage0_19[442]},
      {stage1_19[232]}
   );
   gpc1_1 gpc3144 (
      {stage0_19[443]},
      {stage1_19[233]}
   );
   gpc1_1 gpc3145 (
      {stage0_19[444]},
      {stage1_19[234]}
   );
   gpc1_1 gpc3146 (
      {stage0_19[445]},
      {stage1_19[235]}
   );
   gpc1_1 gpc3147 (
      {stage0_19[446]},
      {stage1_19[236]}
   );
   gpc1_1 gpc3148 (
      {stage0_19[447]},
      {stage1_19[237]}
   );
   gpc1_1 gpc3149 (
      {stage0_19[448]},
      {stage1_19[238]}
   );
   gpc1_1 gpc3150 (
      {stage0_19[449]},
      {stage1_19[239]}
   );
   gpc1_1 gpc3151 (
      {stage0_19[450]},
      {stage1_19[240]}
   );
   gpc1_1 gpc3152 (
      {stage0_19[451]},
      {stage1_19[241]}
   );
   gpc1_1 gpc3153 (
      {stage0_19[452]},
      {stage1_19[242]}
   );
   gpc1_1 gpc3154 (
      {stage0_19[453]},
      {stage1_19[243]}
   );
   gpc1_1 gpc3155 (
      {stage0_19[454]},
      {stage1_19[244]}
   );
   gpc1_1 gpc3156 (
      {stage0_19[455]},
      {stage1_19[245]}
   );
   gpc1_1 gpc3157 (
      {stage0_19[456]},
      {stage1_19[246]}
   );
   gpc1_1 gpc3158 (
      {stage0_19[457]},
      {stage1_19[247]}
   );
   gpc1_1 gpc3159 (
      {stage0_19[458]},
      {stage1_19[248]}
   );
   gpc1_1 gpc3160 (
      {stage0_19[459]},
      {stage1_19[249]}
   );
   gpc1_1 gpc3161 (
      {stage0_19[460]},
      {stage1_19[250]}
   );
   gpc1_1 gpc3162 (
      {stage0_19[461]},
      {stage1_19[251]}
   );
   gpc1_1 gpc3163 (
      {stage0_19[462]},
      {stage1_19[252]}
   );
   gpc1_1 gpc3164 (
      {stage0_19[463]},
      {stage1_19[253]}
   );
   gpc1_1 gpc3165 (
      {stage0_19[464]},
      {stage1_19[254]}
   );
   gpc1_1 gpc3166 (
      {stage0_19[465]},
      {stage1_19[255]}
   );
   gpc1_1 gpc3167 (
      {stage0_19[466]},
      {stage1_19[256]}
   );
   gpc1_1 gpc3168 (
      {stage0_19[467]},
      {stage1_19[257]}
   );
   gpc1_1 gpc3169 (
      {stage0_19[468]},
      {stage1_19[258]}
   );
   gpc1_1 gpc3170 (
      {stage0_19[469]},
      {stage1_19[259]}
   );
   gpc1_1 gpc3171 (
      {stage0_19[470]},
      {stage1_19[260]}
   );
   gpc1_1 gpc3172 (
      {stage0_19[471]},
      {stage1_19[261]}
   );
   gpc1_1 gpc3173 (
      {stage0_19[472]},
      {stage1_19[262]}
   );
   gpc1_1 gpc3174 (
      {stage0_19[473]},
      {stage1_19[263]}
   );
   gpc1_1 gpc3175 (
      {stage0_19[474]},
      {stage1_19[264]}
   );
   gpc1_1 gpc3176 (
      {stage0_19[475]},
      {stage1_19[265]}
   );
   gpc1_1 gpc3177 (
      {stage0_19[476]},
      {stage1_19[266]}
   );
   gpc1_1 gpc3178 (
      {stage0_19[477]},
      {stage1_19[267]}
   );
   gpc1_1 gpc3179 (
      {stage0_19[478]},
      {stage1_19[268]}
   );
   gpc1_1 gpc3180 (
      {stage0_19[479]},
      {stage1_19[269]}
   );
   gpc1_1 gpc3181 (
      {stage0_19[480]},
      {stage1_19[270]}
   );
   gpc1_1 gpc3182 (
      {stage0_19[481]},
      {stage1_19[271]}
   );
   gpc1_1 gpc3183 (
      {stage0_19[482]},
      {stage1_19[272]}
   );
   gpc1_1 gpc3184 (
      {stage0_19[483]},
      {stage1_19[273]}
   );
   gpc1_1 gpc3185 (
      {stage0_19[484]},
      {stage1_19[274]}
   );
   gpc1_1 gpc3186 (
      {stage0_19[485]},
      {stage1_19[275]}
   );
   gpc1_1 gpc3187 (
      {stage0_20[432]},
      {stage1_20[214]}
   );
   gpc1_1 gpc3188 (
      {stage0_20[433]},
      {stage1_20[215]}
   );
   gpc1_1 gpc3189 (
      {stage0_20[434]},
      {stage1_20[216]}
   );
   gpc1_1 gpc3190 (
      {stage0_20[435]},
      {stage1_20[217]}
   );
   gpc1_1 gpc3191 (
      {stage0_20[436]},
      {stage1_20[218]}
   );
   gpc1_1 gpc3192 (
      {stage0_20[437]},
      {stage1_20[219]}
   );
   gpc1_1 gpc3193 (
      {stage0_20[438]},
      {stage1_20[220]}
   );
   gpc1_1 gpc3194 (
      {stage0_20[439]},
      {stage1_20[221]}
   );
   gpc1_1 gpc3195 (
      {stage0_20[440]},
      {stage1_20[222]}
   );
   gpc1_1 gpc3196 (
      {stage0_20[441]},
      {stage1_20[223]}
   );
   gpc1_1 gpc3197 (
      {stage0_20[442]},
      {stage1_20[224]}
   );
   gpc1_1 gpc3198 (
      {stage0_20[443]},
      {stage1_20[225]}
   );
   gpc1_1 gpc3199 (
      {stage0_20[444]},
      {stage1_20[226]}
   );
   gpc1_1 gpc3200 (
      {stage0_20[445]},
      {stage1_20[227]}
   );
   gpc1_1 gpc3201 (
      {stage0_20[446]},
      {stage1_20[228]}
   );
   gpc1_1 gpc3202 (
      {stage0_20[447]},
      {stage1_20[229]}
   );
   gpc1_1 gpc3203 (
      {stage0_20[448]},
      {stage1_20[230]}
   );
   gpc1_1 gpc3204 (
      {stage0_20[449]},
      {stage1_20[231]}
   );
   gpc1_1 gpc3205 (
      {stage0_20[450]},
      {stage1_20[232]}
   );
   gpc1_1 gpc3206 (
      {stage0_20[451]},
      {stage1_20[233]}
   );
   gpc1_1 gpc3207 (
      {stage0_20[452]},
      {stage1_20[234]}
   );
   gpc1_1 gpc3208 (
      {stage0_20[453]},
      {stage1_20[235]}
   );
   gpc1_1 gpc3209 (
      {stage0_20[454]},
      {stage1_20[236]}
   );
   gpc1_1 gpc3210 (
      {stage0_20[455]},
      {stage1_20[237]}
   );
   gpc1_1 gpc3211 (
      {stage0_20[456]},
      {stage1_20[238]}
   );
   gpc1_1 gpc3212 (
      {stage0_20[457]},
      {stage1_20[239]}
   );
   gpc1_1 gpc3213 (
      {stage0_20[458]},
      {stage1_20[240]}
   );
   gpc1_1 gpc3214 (
      {stage0_20[459]},
      {stage1_20[241]}
   );
   gpc1_1 gpc3215 (
      {stage0_20[460]},
      {stage1_20[242]}
   );
   gpc1_1 gpc3216 (
      {stage0_20[461]},
      {stage1_20[243]}
   );
   gpc1_1 gpc3217 (
      {stage0_20[462]},
      {stage1_20[244]}
   );
   gpc1_1 gpc3218 (
      {stage0_20[463]},
      {stage1_20[245]}
   );
   gpc1_1 gpc3219 (
      {stage0_20[464]},
      {stage1_20[246]}
   );
   gpc1_1 gpc3220 (
      {stage0_20[465]},
      {stage1_20[247]}
   );
   gpc1_1 gpc3221 (
      {stage0_20[466]},
      {stage1_20[248]}
   );
   gpc1_1 gpc3222 (
      {stage0_20[467]},
      {stage1_20[249]}
   );
   gpc1_1 gpc3223 (
      {stage0_20[468]},
      {stage1_20[250]}
   );
   gpc1_1 gpc3224 (
      {stage0_20[469]},
      {stage1_20[251]}
   );
   gpc1_1 gpc3225 (
      {stage0_20[470]},
      {stage1_20[252]}
   );
   gpc1_1 gpc3226 (
      {stage0_20[471]},
      {stage1_20[253]}
   );
   gpc1_1 gpc3227 (
      {stage0_20[472]},
      {stage1_20[254]}
   );
   gpc1_1 gpc3228 (
      {stage0_20[473]},
      {stage1_20[255]}
   );
   gpc1_1 gpc3229 (
      {stage0_20[474]},
      {stage1_20[256]}
   );
   gpc1_1 gpc3230 (
      {stage0_20[475]},
      {stage1_20[257]}
   );
   gpc1_1 gpc3231 (
      {stage0_20[476]},
      {stage1_20[258]}
   );
   gpc1_1 gpc3232 (
      {stage0_20[477]},
      {stage1_20[259]}
   );
   gpc1_1 gpc3233 (
      {stage0_20[478]},
      {stage1_20[260]}
   );
   gpc1_1 gpc3234 (
      {stage0_20[479]},
      {stage1_20[261]}
   );
   gpc1_1 gpc3235 (
      {stage0_20[480]},
      {stage1_20[262]}
   );
   gpc1_1 gpc3236 (
      {stage0_20[481]},
      {stage1_20[263]}
   );
   gpc1_1 gpc3237 (
      {stage0_20[482]},
      {stage1_20[264]}
   );
   gpc1_1 gpc3238 (
      {stage0_20[483]},
      {stage1_20[265]}
   );
   gpc1_1 gpc3239 (
      {stage0_20[484]},
      {stage1_20[266]}
   );
   gpc1_1 gpc3240 (
      {stage0_20[485]},
      {stage1_20[267]}
   );
   gpc1_1 gpc3241 (
      {stage0_21[468]},
      {stage1_21[172]}
   );
   gpc1_1 gpc3242 (
      {stage0_21[469]},
      {stage1_21[173]}
   );
   gpc1_1 gpc3243 (
      {stage0_21[470]},
      {stage1_21[174]}
   );
   gpc1_1 gpc3244 (
      {stage0_21[471]},
      {stage1_21[175]}
   );
   gpc1_1 gpc3245 (
      {stage0_21[472]},
      {stage1_21[176]}
   );
   gpc1_1 gpc3246 (
      {stage0_21[473]},
      {stage1_21[177]}
   );
   gpc1_1 gpc3247 (
      {stage0_21[474]},
      {stage1_21[178]}
   );
   gpc1_1 gpc3248 (
      {stage0_21[475]},
      {stage1_21[179]}
   );
   gpc1_1 gpc3249 (
      {stage0_21[476]},
      {stage1_21[180]}
   );
   gpc1_1 gpc3250 (
      {stage0_21[477]},
      {stage1_21[181]}
   );
   gpc1_1 gpc3251 (
      {stage0_21[478]},
      {stage1_21[182]}
   );
   gpc1_1 gpc3252 (
      {stage0_21[479]},
      {stage1_21[183]}
   );
   gpc1_1 gpc3253 (
      {stage0_21[480]},
      {stage1_21[184]}
   );
   gpc1_1 gpc3254 (
      {stage0_21[481]},
      {stage1_21[185]}
   );
   gpc1_1 gpc3255 (
      {stage0_21[482]},
      {stage1_21[186]}
   );
   gpc1_1 gpc3256 (
      {stage0_21[483]},
      {stage1_21[187]}
   );
   gpc1_1 gpc3257 (
      {stage0_21[484]},
      {stage1_21[188]}
   );
   gpc1_1 gpc3258 (
      {stage0_21[485]},
      {stage1_21[189]}
   );
   gpc1_1 gpc3259 (
      {stage0_22[472]},
      {stage1_22[157]}
   );
   gpc1_1 gpc3260 (
      {stage0_22[473]},
      {stage1_22[158]}
   );
   gpc1_1 gpc3261 (
      {stage0_22[474]},
      {stage1_22[159]}
   );
   gpc1_1 gpc3262 (
      {stage0_22[475]},
      {stage1_22[160]}
   );
   gpc1_1 gpc3263 (
      {stage0_22[476]},
      {stage1_22[161]}
   );
   gpc1_1 gpc3264 (
      {stage0_22[477]},
      {stage1_22[162]}
   );
   gpc1_1 gpc3265 (
      {stage0_22[478]},
      {stage1_22[163]}
   );
   gpc1_1 gpc3266 (
      {stage0_22[479]},
      {stage1_22[164]}
   );
   gpc1_1 gpc3267 (
      {stage0_22[480]},
      {stage1_22[165]}
   );
   gpc1_1 gpc3268 (
      {stage0_22[481]},
      {stage1_22[166]}
   );
   gpc1_1 gpc3269 (
      {stage0_22[482]},
      {stage1_22[167]}
   );
   gpc1_1 gpc3270 (
      {stage0_22[483]},
      {stage1_22[168]}
   );
   gpc1_1 gpc3271 (
      {stage0_22[484]},
      {stage1_22[169]}
   );
   gpc1_1 gpc3272 (
      {stage0_22[485]},
      {stage1_22[170]}
   );
   gpc1_1 gpc3273 (
      {stage0_23[396]},
      {stage1_23[197]}
   );
   gpc1_1 gpc3274 (
      {stage0_23[397]},
      {stage1_23[198]}
   );
   gpc1_1 gpc3275 (
      {stage0_23[398]},
      {stage1_23[199]}
   );
   gpc1_1 gpc3276 (
      {stage0_23[399]},
      {stage1_23[200]}
   );
   gpc1_1 gpc3277 (
      {stage0_23[400]},
      {stage1_23[201]}
   );
   gpc1_1 gpc3278 (
      {stage0_23[401]},
      {stage1_23[202]}
   );
   gpc1_1 gpc3279 (
      {stage0_23[402]},
      {stage1_23[203]}
   );
   gpc1_1 gpc3280 (
      {stage0_23[403]},
      {stage1_23[204]}
   );
   gpc1_1 gpc3281 (
      {stage0_23[404]},
      {stage1_23[205]}
   );
   gpc1_1 gpc3282 (
      {stage0_23[405]},
      {stage1_23[206]}
   );
   gpc1_1 gpc3283 (
      {stage0_23[406]},
      {stage1_23[207]}
   );
   gpc1_1 gpc3284 (
      {stage0_23[407]},
      {stage1_23[208]}
   );
   gpc1_1 gpc3285 (
      {stage0_23[408]},
      {stage1_23[209]}
   );
   gpc1_1 gpc3286 (
      {stage0_23[409]},
      {stage1_23[210]}
   );
   gpc1_1 gpc3287 (
      {stage0_23[410]},
      {stage1_23[211]}
   );
   gpc1_1 gpc3288 (
      {stage0_23[411]},
      {stage1_23[212]}
   );
   gpc1_1 gpc3289 (
      {stage0_23[412]},
      {stage1_23[213]}
   );
   gpc1_1 gpc3290 (
      {stage0_23[413]},
      {stage1_23[214]}
   );
   gpc1_1 gpc3291 (
      {stage0_23[414]},
      {stage1_23[215]}
   );
   gpc1_1 gpc3292 (
      {stage0_23[415]},
      {stage1_23[216]}
   );
   gpc1_1 gpc3293 (
      {stage0_23[416]},
      {stage1_23[217]}
   );
   gpc1_1 gpc3294 (
      {stage0_23[417]},
      {stage1_23[218]}
   );
   gpc1_1 gpc3295 (
      {stage0_23[418]},
      {stage1_23[219]}
   );
   gpc1_1 gpc3296 (
      {stage0_23[419]},
      {stage1_23[220]}
   );
   gpc1_1 gpc3297 (
      {stage0_23[420]},
      {stage1_23[221]}
   );
   gpc1_1 gpc3298 (
      {stage0_23[421]},
      {stage1_23[222]}
   );
   gpc1_1 gpc3299 (
      {stage0_23[422]},
      {stage1_23[223]}
   );
   gpc1_1 gpc3300 (
      {stage0_23[423]},
      {stage1_23[224]}
   );
   gpc1_1 gpc3301 (
      {stage0_23[424]},
      {stage1_23[225]}
   );
   gpc1_1 gpc3302 (
      {stage0_23[425]},
      {stage1_23[226]}
   );
   gpc1_1 gpc3303 (
      {stage0_23[426]},
      {stage1_23[227]}
   );
   gpc1_1 gpc3304 (
      {stage0_23[427]},
      {stage1_23[228]}
   );
   gpc1_1 gpc3305 (
      {stage0_23[428]},
      {stage1_23[229]}
   );
   gpc1_1 gpc3306 (
      {stage0_23[429]},
      {stage1_23[230]}
   );
   gpc1_1 gpc3307 (
      {stage0_23[430]},
      {stage1_23[231]}
   );
   gpc1_1 gpc3308 (
      {stage0_23[431]},
      {stage1_23[232]}
   );
   gpc1_1 gpc3309 (
      {stage0_23[432]},
      {stage1_23[233]}
   );
   gpc1_1 gpc3310 (
      {stage0_23[433]},
      {stage1_23[234]}
   );
   gpc1_1 gpc3311 (
      {stage0_23[434]},
      {stage1_23[235]}
   );
   gpc1_1 gpc3312 (
      {stage0_23[435]},
      {stage1_23[236]}
   );
   gpc1_1 gpc3313 (
      {stage0_23[436]},
      {stage1_23[237]}
   );
   gpc1_1 gpc3314 (
      {stage0_23[437]},
      {stage1_23[238]}
   );
   gpc1_1 gpc3315 (
      {stage0_23[438]},
      {stage1_23[239]}
   );
   gpc1_1 gpc3316 (
      {stage0_23[439]},
      {stage1_23[240]}
   );
   gpc1_1 gpc3317 (
      {stage0_23[440]},
      {stage1_23[241]}
   );
   gpc1_1 gpc3318 (
      {stage0_23[441]},
      {stage1_23[242]}
   );
   gpc1_1 gpc3319 (
      {stage0_23[442]},
      {stage1_23[243]}
   );
   gpc1_1 gpc3320 (
      {stage0_23[443]},
      {stage1_23[244]}
   );
   gpc1_1 gpc3321 (
      {stage0_23[444]},
      {stage1_23[245]}
   );
   gpc1_1 gpc3322 (
      {stage0_23[445]},
      {stage1_23[246]}
   );
   gpc1_1 gpc3323 (
      {stage0_23[446]},
      {stage1_23[247]}
   );
   gpc1_1 gpc3324 (
      {stage0_23[447]},
      {stage1_23[248]}
   );
   gpc1_1 gpc3325 (
      {stage0_23[448]},
      {stage1_23[249]}
   );
   gpc1_1 gpc3326 (
      {stage0_23[449]},
      {stage1_23[250]}
   );
   gpc1_1 gpc3327 (
      {stage0_23[450]},
      {stage1_23[251]}
   );
   gpc1_1 gpc3328 (
      {stage0_23[451]},
      {stage1_23[252]}
   );
   gpc1_1 gpc3329 (
      {stage0_23[452]},
      {stage1_23[253]}
   );
   gpc1_1 gpc3330 (
      {stage0_23[453]},
      {stage1_23[254]}
   );
   gpc1_1 gpc3331 (
      {stage0_23[454]},
      {stage1_23[255]}
   );
   gpc1_1 gpc3332 (
      {stage0_23[455]},
      {stage1_23[256]}
   );
   gpc1_1 gpc3333 (
      {stage0_23[456]},
      {stage1_23[257]}
   );
   gpc1_1 gpc3334 (
      {stage0_23[457]},
      {stage1_23[258]}
   );
   gpc1_1 gpc3335 (
      {stage0_23[458]},
      {stage1_23[259]}
   );
   gpc1_1 gpc3336 (
      {stage0_23[459]},
      {stage1_23[260]}
   );
   gpc1_1 gpc3337 (
      {stage0_23[460]},
      {stage1_23[261]}
   );
   gpc1_1 gpc3338 (
      {stage0_23[461]},
      {stage1_23[262]}
   );
   gpc1_1 gpc3339 (
      {stage0_23[462]},
      {stage1_23[263]}
   );
   gpc1_1 gpc3340 (
      {stage0_23[463]},
      {stage1_23[264]}
   );
   gpc1_1 gpc3341 (
      {stage0_23[464]},
      {stage1_23[265]}
   );
   gpc1_1 gpc3342 (
      {stage0_23[465]},
      {stage1_23[266]}
   );
   gpc1_1 gpc3343 (
      {stage0_23[466]},
      {stage1_23[267]}
   );
   gpc1_1 gpc3344 (
      {stage0_23[467]},
      {stage1_23[268]}
   );
   gpc1_1 gpc3345 (
      {stage0_23[468]},
      {stage1_23[269]}
   );
   gpc1_1 gpc3346 (
      {stage0_23[469]},
      {stage1_23[270]}
   );
   gpc1_1 gpc3347 (
      {stage0_23[470]},
      {stage1_23[271]}
   );
   gpc1_1 gpc3348 (
      {stage0_23[471]},
      {stage1_23[272]}
   );
   gpc1_1 gpc3349 (
      {stage0_23[472]},
      {stage1_23[273]}
   );
   gpc1_1 gpc3350 (
      {stage0_23[473]},
      {stage1_23[274]}
   );
   gpc1_1 gpc3351 (
      {stage0_23[474]},
      {stage1_23[275]}
   );
   gpc1_1 gpc3352 (
      {stage0_23[475]},
      {stage1_23[276]}
   );
   gpc1_1 gpc3353 (
      {stage0_23[476]},
      {stage1_23[277]}
   );
   gpc1_1 gpc3354 (
      {stage0_23[477]},
      {stage1_23[278]}
   );
   gpc1_1 gpc3355 (
      {stage0_23[478]},
      {stage1_23[279]}
   );
   gpc1_1 gpc3356 (
      {stage0_23[479]},
      {stage1_23[280]}
   );
   gpc1_1 gpc3357 (
      {stage0_23[480]},
      {stage1_23[281]}
   );
   gpc1_1 gpc3358 (
      {stage0_23[481]},
      {stage1_23[282]}
   );
   gpc1_1 gpc3359 (
      {stage0_23[482]},
      {stage1_23[283]}
   );
   gpc1_1 gpc3360 (
      {stage0_23[483]},
      {stage1_23[284]}
   );
   gpc1_1 gpc3361 (
      {stage0_23[484]},
      {stage1_23[285]}
   );
   gpc1_1 gpc3362 (
      {stage0_23[485]},
      {stage1_23[286]}
   );
   gpc1_1 gpc3363 (
      {stage0_24[485]},
      {stage1_24[213]}
   );
   gpc1_1 gpc3364 (
      {stage0_26[402]},
      {stage1_26[167]}
   );
   gpc1_1 gpc3365 (
      {stage0_26[403]},
      {stage1_26[168]}
   );
   gpc1_1 gpc3366 (
      {stage0_26[404]},
      {stage1_26[169]}
   );
   gpc1_1 gpc3367 (
      {stage0_26[405]},
      {stage1_26[170]}
   );
   gpc1_1 gpc3368 (
      {stage0_26[406]},
      {stage1_26[171]}
   );
   gpc1_1 gpc3369 (
      {stage0_26[407]},
      {stage1_26[172]}
   );
   gpc1_1 gpc3370 (
      {stage0_26[408]},
      {stage1_26[173]}
   );
   gpc1_1 gpc3371 (
      {stage0_26[409]},
      {stage1_26[174]}
   );
   gpc1_1 gpc3372 (
      {stage0_26[410]},
      {stage1_26[175]}
   );
   gpc1_1 gpc3373 (
      {stage0_26[411]},
      {stage1_26[176]}
   );
   gpc1_1 gpc3374 (
      {stage0_26[412]},
      {stage1_26[177]}
   );
   gpc1_1 gpc3375 (
      {stage0_26[413]},
      {stage1_26[178]}
   );
   gpc1_1 gpc3376 (
      {stage0_26[414]},
      {stage1_26[179]}
   );
   gpc1_1 gpc3377 (
      {stage0_26[415]},
      {stage1_26[180]}
   );
   gpc1_1 gpc3378 (
      {stage0_26[416]},
      {stage1_26[181]}
   );
   gpc1_1 gpc3379 (
      {stage0_26[417]},
      {stage1_26[182]}
   );
   gpc1_1 gpc3380 (
      {stage0_26[418]},
      {stage1_26[183]}
   );
   gpc1_1 gpc3381 (
      {stage0_26[419]},
      {stage1_26[184]}
   );
   gpc1_1 gpc3382 (
      {stage0_26[420]},
      {stage1_26[185]}
   );
   gpc1_1 gpc3383 (
      {stage0_26[421]},
      {stage1_26[186]}
   );
   gpc1_1 gpc3384 (
      {stage0_26[422]},
      {stage1_26[187]}
   );
   gpc1_1 gpc3385 (
      {stage0_26[423]},
      {stage1_26[188]}
   );
   gpc1_1 gpc3386 (
      {stage0_26[424]},
      {stage1_26[189]}
   );
   gpc1_1 gpc3387 (
      {stage0_26[425]},
      {stage1_26[190]}
   );
   gpc1_1 gpc3388 (
      {stage0_26[426]},
      {stage1_26[191]}
   );
   gpc1_1 gpc3389 (
      {stage0_26[427]},
      {stage1_26[192]}
   );
   gpc1_1 gpc3390 (
      {stage0_26[428]},
      {stage1_26[193]}
   );
   gpc1_1 gpc3391 (
      {stage0_26[429]},
      {stage1_26[194]}
   );
   gpc1_1 gpc3392 (
      {stage0_26[430]},
      {stage1_26[195]}
   );
   gpc1_1 gpc3393 (
      {stage0_26[431]},
      {stage1_26[196]}
   );
   gpc1_1 gpc3394 (
      {stage0_26[432]},
      {stage1_26[197]}
   );
   gpc1_1 gpc3395 (
      {stage0_26[433]},
      {stage1_26[198]}
   );
   gpc1_1 gpc3396 (
      {stage0_26[434]},
      {stage1_26[199]}
   );
   gpc1_1 gpc3397 (
      {stage0_26[435]},
      {stage1_26[200]}
   );
   gpc1_1 gpc3398 (
      {stage0_26[436]},
      {stage1_26[201]}
   );
   gpc1_1 gpc3399 (
      {stage0_26[437]},
      {stage1_26[202]}
   );
   gpc1_1 gpc3400 (
      {stage0_26[438]},
      {stage1_26[203]}
   );
   gpc1_1 gpc3401 (
      {stage0_26[439]},
      {stage1_26[204]}
   );
   gpc1_1 gpc3402 (
      {stage0_26[440]},
      {stage1_26[205]}
   );
   gpc1_1 gpc3403 (
      {stage0_26[441]},
      {stage1_26[206]}
   );
   gpc1_1 gpc3404 (
      {stage0_26[442]},
      {stage1_26[207]}
   );
   gpc1_1 gpc3405 (
      {stage0_26[443]},
      {stage1_26[208]}
   );
   gpc1_1 gpc3406 (
      {stage0_26[444]},
      {stage1_26[209]}
   );
   gpc1_1 gpc3407 (
      {stage0_26[445]},
      {stage1_26[210]}
   );
   gpc1_1 gpc3408 (
      {stage0_26[446]},
      {stage1_26[211]}
   );
   gpc1_1 gpc3409 (
      {stage0_26[447]},
      {stage1_26[212]}
   );
   gpc1_1 gpc3410 (
      {stage0_26[448]},
      {stage1_26[213]}
   );
   gpc1_1 gpc3411 (
      {stage0_26[449]},
      {stage1_26[214]}
   );
   gpc1_1 gpc3412 (
      {stage0_26[450]},
      {stage1_26[215]}
   );
   gpc1_1 gpc3413 (
      {stage0_26[451]},
      {stage1_26[216]}
   );
   gpc1_1 gpc3414 (
      {stage0_26[452]},
      {stage1_26[217]}
   );
   gpc1_1 gpc3415 (
      {stage0_26[453]},
      {stage1_26[218]}
   );
   gpc1_1 gpc3416 (
      {stage0_26[454]},
      {stage1_26[219]}
   );
   gpc1_1 gpc3417 (
      {stage0_26[455]},
      {stage1_26[220]}
   );
   gpc1_1 gpc3418 (
      {stage0_26[456]},
      {stage1_26[221]}
   );
   gpc1_1 gpc3419 (
      {stage0_26[457]},
      {stage1_26[222]}
   );
   gpc1_1 gpc3420 (
      {stage0_26[458]},
      {stage1_26[223]}
   );
   gpc1_1 gpc3421 (
      {stage0_26[459]},
      {stage1_26[224]}
   );
   gpc1_1 gpc3422 (
      {stage0_26[460]},
      {stage1_26[225]}
   );
   gpc1_1 gpc3423 (
      {stage0_26[461]},
      {stage1_26[226]}
   );
   gpc1_1 gpc3424 (
      {stage0_26[462]},
      {stage1_26[227]}
   );
   gpc1_1 gpc3425 (
      {stage0_26[463]},
      {stage1_26[228]}
   );
   gpc1_1 gpc3426 (
      {stage0_26[464]},
      {stage1_26[229]}
   );
   gpc1_1 gpc3427 (
      {stage0_26[465]},
      {stage1_26[230]}
   );
   gpc1_1 gpc3428 (
      {stage0_26[466]},
      {stage1_26[231]}
   );
   gpc1_1 gpc3429 (
      {stage0_26[467]},
      {stage1_26[232]}
   );
   gpc1_1 gpc3430 (
      {stage0_26[468]},
      {stage1_26[233]}
   );
   gpc1_1 gpc3431 (
      {stage0_26[469]},
      {stage1_26[234]}
   );
   gpc1_1 gpc3432 (
      {stage0_26[470]},
      {stage1_26[235]}
   );
   gpc1_1 gpc3433 (
      {stage0_26[471]},
      {stage1_26[236]}
   );
   gpc1_1 gpc3434 (
      {stage0_26[472]},
      {stage1_26[237]}
   );
   gpc1_1 gpc3435 (
      {stage0_26[473]},
      {stage1_26[238]}
   );
   gpc1_1 gpc3436 (
      {stage0_26[474]},
      {stage1_26[239]}
   );
   gpc1_1 gpc3437 (
      {stage0_26[475]},
      {stage1_26[240]}
   );
   gpc1_1 gpc3438 (
      {stage0_26[476]},
      {stage1_26[241]}
   );
   gpc1_1 gpc3439 (
      {stage0_26[477]},
      {stage1_26[242]}
   );
   gpc1_1 gpc3440 (
      {stage0_26[478]},
      {stage1_26[243]}
   );
   gpc1_1 gpc3441 (
      {stage0_26[479]},
      {stage1_26[244]}
   );
   gpc1_1 gpc3442 (
      {stage0_26[480]},
      {stage1_26[245]}
   );
   gpc1_1 gpc3443 (
      {stage0_26[481]},
      {stage1_26[246]}
   );
   gpc1_1 gpc3444 (
      {stage0_26[482]},
      {stage1_26[247]}
   );
   gpc1_1 gpc3445 (
      {stage0_26[483]},
      {stage1_26[248]}
   );
   gpc1_1 gpc3446 (
      {stage0_26[484]},
      {stage1_26[249]}
   );
   gpc1_1 gpc3447 (
      {stage0_26[485]},
      {stage1_26[250]}
   );
   gpc1_1 gpc3448 (
      {stage0_27[473]},
      {stage1_27[193]}
   );
   gpc1_1 gpc3449 (
      {stage0_27[474]},
      {stage1_27[194]}
   );
   gpc1_1 gpc3450 (
      {stage0_27[475]},
      {stage1_27[195]}
   );
   gpc1_1 gpc3451 (
      {stage0_27[476]},
      {stage1_27[196]}
   );
   gpc1_1 gpc3452 (
      {stage0_27[477]},
      {stage1_27[197]}
   );
   gpc1_1 gpc3453 (
      {stage0_27[478]},
      {stage1_27[198]}
   );
   gpc1_1 gpc3454 (
      {stage0_27[479]},
      {stage1_27[199]}
   );
   gpc1_1 gpc3455 (
      {stage0_27[480]},
      {stage1_27[200]}
   );
   gpc1_1 gpc3456 (
      {stage0_27[481]},
      {stage1_27[201]}
   );
   gpc1_1 gpc3457 (
      {stage0_27[482]},
      {stage1_27[202]}
   );
   gpc1_1 gpc3458 (
      {stage0_27[483]},
      {stage1_27[203]}
   );
   gpc1_1 gpc3459 (
      {stage0_27[484]},
      {stage1_27[204]}
   );
   gpc1_1 gpc3460 (
      {stage0_27[485]},
      {stage1_27[205]}
   );
   gpc1_1 gpc3461 (
      {stage0_28[475]},
      {stage1_28[213]}
   );
   gpc1_1 gpc3462 (
      {stage0_28[476]},
      {stage1_28[214]}
   );
   gpc1_1 gpc3463 (
      {stage0_28[477]},
      {stage1_28[215]}
   );
   gpc1_1 gpc3464 (
      {stage0_28[478]},
      {stage1_28[216]}
   );
   gpc1_1 gpc3465 (
      {stage0_28[479]},
      {stage1_28[217]}
   );
   gpc1_1 gpc3466 (
      {stage0_28[480]},
      {stage1_28[218]}
   );
   gpc1_1 gpc3467 (
      {stage0_28[481]},
      {stage1_28[219]}
   );
   gpc1_1 gpc3468 (
      {stage0_28[482]},
      {stage1_28[220]}
   );
   gpc1_1 gpc3469 (
      {stage0_28[483]},
      {stage1_28[221]}
   );
   gpc1_1 gpc3470 (
      {stage0_28[484]},
      {stage1_28[222]}
   );
   gpc1_1 gpc3471 (
      {stage0_28[485]},
      {stage1_28[223]}
   );
   gpc1_1 gpc3472 (
      {stage0_29[444]},
      {stage1_29[187]}
   );
   gpc1_1 gpc3473 (
      {stage0_29[445]},
      {stage1_29[188]}
   );
   gpc1_1 gpc3474 (
      {stage0_29[446]},
      {stage1_29[189]}
   );
   gpc1_1 gpc3475 (
      {stage0_29[447]},
      {stage1_29[190]}
   );
   gpc1_1 gpc3476 (
      {stage0_29[448]},
      {stage1_29[191]}
   );
   gpc1_1 gpc3477 (
      {stage0_29[449]},
      {stage1_29[192]}
   );
   gpc1_1 gpc3478 (
      {stage0_29[450]},
      {stage1_29[193]}
   );
   gpc1_1 gpc3479 (
      {stage0_29[451]},
      {stage1_29[194]}
   );
   gpc1_1 gpc3480 (
      {stage0_29[452]},
      {stage1_29[195]}
   );
   gpc1_1 gpc3481 (
      {stage0_29[453]},
      {stage1_29[196]}
   );
   gpc1_1 gpc3482 (
      {stage0_29[454]},
      {stage1_29[197]}
   );
   gpc1_1 gpc3483 (
      {stage0_29[455]},
      {stage1_29[198]}
   );
   gpc1_1 gpc3484 (
      {stage0_29[456]},
      {stage1_29[199]}
   );
   gpc1_1 gpc3485 (
      {stage0_29[457]},
      {stage1_29[200]}
   );
   gpc1_1 gpc3486 (
      {stage0_29[458]},
      {stage1_29[201]}
   );
   gpc1_1 gpc3487 (
      {stage0_29[459]},
      {stage1_29[202]}
   );
   gpc1_1 gpc3488 (
      {stage0_29[460]},
      {stage1_29[203]}
   );
   gpc1_1 gpc3489 (
      {stage0_29[461]},
      {stage1_29[204]}
   );
   gpc1_1 gpc3490 (
      {stage0_29[462]},
      {stage1_29[205]}
   );
   gpc1_1 gpc3491 (
      {stage0_29[463]},
      {stage1_29[206]}
   );
   gpc1_1 gpc3492 (
      {stage0_29[464]},
      {stage1_29[207]}
   );
   gpc1_1 gpc3493 (
      {stage0_29[465]},
      {stage1_29[208]}
   );
   gpc1_1 gpc3494 (
      {stage0_29[466]},
      {stage1_29[209]}
   );
   gpc1_1 gpc3495 (
      {stage0_29[467]},
      {stage1_29[210]}
   );
   gpc1_1 gpc3496 (
      {stage0_29[468]},
      {stage1_29[211]}
   );
   gpc1_1 gpc3497 (
      {stage0_29[469]},
      {stage1_29[212]}
   );
   gpc1_1 gpc3498 (
      {stage0_29[470]},
      {stage1_29[213]}
   );
   gpc1_1 gpc3499 (
      {stage0_29[471]},
      {stage1_29[214]}
   );
   gpc1_1 gpc3500 (
      {stage0_29[472]},
      {stage1_29[215]}
   );
   gpc1_1 gpc3501 (
      {stage0_29[473]},
      {stage1_29[216]}
   );
   gpc1_1 gpc3502 (
      {stage0_29[474]},
      {stage1_29[217]}
   );
   gpc1_1 gpc3503 (
      {stage0_29[475]},
      {stage1_29[218]}
   );
   gpc1_1 gpc3504 (
      {stage0_29[476]},
      {stage1_29[219]}
   );
   gpc1_1 gpc3505 (
      {stage0_29[477]},
      {stage1_29[220]}
   );
   gpc1_1 gpc3506 (
      {stage0_29[478]},
      {stage1_29[221]}
   );
   gpc1_1 gpc3507 (
      {stage0_29[479]},
      {stage1_29[222]}
   );
   gpc1_1 gpc3508 (
      {stage0_29[480]},
      {stage1_29[223]}
   );
   gpc1_1 gpc3509 (
      {stage0_29[481]},
      {stage1_29[224]}
   );
   gpc1_1 gpc3510 (
      {stage0_29[482]},
      {stage1_29[225]}
   );
   gpc1_1 gpc3511 (
      {stage0_29[483]},
      {stage1_29[226]}
   );
   gpc1_1 gpc3512 (
      {stage0_29[484]},
      {stage1_29[227]}
   );
   gpc1_1 gpc3513 (
      {stage0_29[485]},
      {stage1_29[228]}
   );
   gpc1_1 gpc3514 (
      {stage0_30[460]},
      {stage1_30[166]}
   );
   gpc1_1 gpc3515 (
      {stage0_30[461]},
      {stage1_30[167]}
   );
   gpc1_1 gpc3516 (
      {stage0_30[462]},
      {stage1_30[168]}
   );
   gpc1_1 gpc3517 (
      {stage0_30[463]},
      {stage1_30[169]}
   );
   gpc1_1 gpc3518 (
      {stage0_30[464]},
      {stage1_30[170]}
   );
   gpc1_1 gpc3519 (
      {stage0_30[465]},
      {stage1_30[171]}
   );
   gpc1_1 gpc3520 (
      {stage0_30[466]},
      {stage1_30[172]}
   );
   gpc1_1 gpc3521 (
      {stage0_30[467]},
      {stage1_30[173]}
   );
   gpc1_1 gpc3522 (
      {stage0_30[468]},
      {stage1_30[174]}
   );
   gpc1_1 gpc3523 (
      {stage0_30[469]},
      {stage1_30[175]}
   );
   gpc1_1 gpc3524 (
      {stage0_30[470]},
      {stage1_30[176]}
   );
   gpc1_1 gpc3525 (
      {stage0_30[471]},
      {stage1_30[177]}
   );
   gpc1_1 gpc3526 (
      {stage0_30[472]},
      {stage1_30[178]}
   );
   gpc1_1 gpc3527 (
      {stage0_30[473]},
      {stage1_30[179]}
   );
   gpc1_1 gpc3528 (
      {stage0_30[474]},
      {stage1_30[180]}
   );
   gpc1_1 gpc3529 (
      {stage0_30[475]},
      {stage1_30[181]}
   );
   gpc1_1 gpc3530 (
      {stage0_30[476]},
      {stage1_30[182]}
   );
   gpc1_1 gpc3531 (
      {stage0_30[477]},
      {stage1_30[183]}
   );
   gpc1_1 gpc3532 (
      {stage0_30[478]},
      {stage1_30[184]}
   );
   gpc1_1 gpc3533 (
      {stage0_30[479]},
      {stage1_30[185]}
   );
   gpc1_1 gpc3534 (
      {stage0_30[480]},
      {stage1_30[186]}
   );
   gpc1_1 gpc3535 (
      {stage0_30[481]},
      {stage1_30[187]}
   );
   gpc1_1 gpc3536 (
      {stage0_30[482]},
      {stage1_30[188]}
   );
   gpc1_1 gpc3537 (
      {stage0_30[483]},
      {stage1_30[189]}
   );
   gpc1_1 gpc3538 (
      {stage0_30[484]},
      {stage1_30[190]}
   );
   gpc1_1 gpc3539 (
      {stage0_30[485]},
      {stage1_30[191]}
   );
   gpc1_1 gpc3540 (
      {stage0_31[476]},
      {stage1_31[208]}
   );
   gpc1_1 gpc3541 (
      {stage0_31[477]},
      {stage1_31[209]}
   );
   gpc1_1 gpc3542 (
      {stage0_31[478]},
      {stage1_31[210]}
   );
   gpc1_1 gpc3543 (
      {stage0_31[479]},
      {stage1_31[211]}
   );
   gpc1_1 gpc3544 (
      {stage0_31[480]},
      {stage1_31[212]}
   );
   gpc1_1 gpc3545 (
      {stage0_31[481]},
      {stage1_31[213]}
   );
   gpc1_1 gpc3546 (
      {stage0_31[482]},
      {stage1_31[214]}
   );
   gpc1_1 gpc3547 (
      {stage0_31[483]},
      {stage1_31[215]}
   );
   gpc1_1 gpc3548 (
      {stage0_31[484]},
      {stage1_31[216]}
   );
   gpc1_1 gpc3549 (
      {stage0_31[485]},
      {stage1_31[217]}
   );
   gpc1_1 gpc3550 (
      {stage0_33[396]},
      {stage1_33[169]}
   );
   gpc1_1 gpc3551 (
      {stage0_33[397]},
      {stage1_33[170]}
   );
   gpc1_1 gpc3552 (
      {stage0_33[398]},
      {stage1_33[171]}
   );
   gpc1_1 gpc3553 (
      {stage0_33[399]},
      {stage1_33[172]}
   );
   gpc1_1 gpc3554 (
      {stage0_33[400]},
      {stage1_33[173]}
   );
   gpc1_1 gpc3555 (
      {stage0_33[401]},
      {stage1_33[174]}
   );
   gpc1_1 gpc3556 (
      {stage0_33[402]},
      {stage1_33[175]}
   );
   gpc1_1 gpc3557 (
      {stage0_33[403]},
      {stage1_33[176]}
   );
   gpc1_1 gpc3558 (
      {stage0_33[404]},
      {stage1_33[177]}
   );
   gpc1_1 gpc3559 (
      {stage0_33[405]},
      {stage1_33[178]}
   );
   gpc1_1 gpc3560 (
      {stage0_33[406]},
      {stage1_33[179]}
   );
   gpc1_1 gpc3561 (
      {stage0_33[407]},
      {stage1_33[180]}
   );
   gpc1_1 gpc3562 (
      {stage0_33[408]},
      {stage1_33[181]}
   );
   gpc1_1 gpc3563 (
      {stage0_33[409]},
      {stage1_33[182]}
   );
   gpc1_1 gpc3564 (
      {stage0_33[410]},
      {stage1_33[183]}
   );
   gpc1_1 gpc3565 (
      {stage0_33[411]},
      {stage1_33[184]}
   );
   gpc1_1 gpc3566 (
      {stage0_33[412]},
      {stage1_33[185]}
   );
   gpc1_1 gpc3567 (
      {stage0_33[413]},
      {stage1_33[186]}
   );
   gpc1_1 gpc3568 (
      {stage0_33[414]},
      {stage1_33[187]}
   );
   gpc1_1 gpc3569 (
      {stage0_33[415]},
      {stage1_33[188]}
   );
   gpc1_1 gpc3570 (
      {stage0_33[416]},
      {stage1_33[189]}
   );
   gpc1_1 gpc3571 (
      {stage0_33[417]},
      {stage1_33[190]}
   );
   gpc1_1 gpc3572 (
      {stage0_33[418]},
      {stage1_33[191]}
   );
   gpc1_1 gpc3573 (
      {stage0_33[419]},
      {stage1_33[192]}
   );
   gpc1_1 gpc3574 (
      {stage0_33[420]},
      {stage1_33[193]}
   );
   gpc1_1 gpc3575 (
      {stage0_33[421]},
      {stage1_33[194]}
   );
   gpc1_1 gpc3576 (
      {stage0_33[422]},
      {stage1_33[195]}
   );
   gpc1_1 gpc3577 (
      {stage0_33[423]},
      {stage1_33[196]}
   );
   gpc1_1 gpc3578 (
      {stage0_33[424]},
      {stage1_33[197]}
   );
   gpc1_1 gpc3579 (
      {stage0_33[425]},
      {stage1_33[198]}
   );
   gpc1_1 gpc3580 (
      {stage0_33[426]},
      {stage1_33[199]}
   );
   gpc1_1 gpc3581 (
      {stage0_33[427]},
      {stage1_33[200]}
   );
   gpc1_1 gpc3582 (
      {stage0_33[428]},
      {stage1_33[201]}
   );
   gpc1_1 gpc3583 (
      {stage0_33[429]},
      {stage1_33[202]}
   );
   gpc1_1 gpc3584 (
      {stage0_33[430]},
      {stage1_33[203]}
   );
   gpc1_1 gpc3585 (
      {stage0_33[431]},
      {stage1_33[204]}
   );
   gpc1_1 gpc3586 (
      {stage0_33[432]},
      {stage1_33[205]}
   );
   gpc1_1 gpc3587 (
      {stage0_33[433]},
      {stage1_33[206]}
   );
   gpc1_1 gpc3588 (
      {stage0_33[434]},
      {stage1_33[207]}
   );
   gpc1_1 gpc3589 (
      {stage0_33[435]},
      {stage1_33[208]}
   );
   gpc1_1 gpc3590 (
      {stage0_33[436]},
      {stage1_33[209]}
   );
   gpc1_1 gpc3591 (
      {stage0_33[437]},
      {stage1_33[210]}
   );
   gpc1_1 gpc3592 (
      {stage0_33[438]},
      {stage1_33[211]}
   );
   gpc1_1 gpc3593 (
      {stage0_33[439]},
      {stage1_33[212]}
   );
   gpc1_1 gpc3594 (
      {stage0_33[440]},
      {stage1_33[213]}
   );
   gpc1_1 gpc3595 (
      {stage0_33[441]},
      {stage1_33[214]}
   );
   gpc1_1 gpc3596 (
      {stage0_33[442]},
      {stage1_33[215]}
   );
   gpc1_1 gpc3597 (
      {stage0_33[443]},
      {stage1_33[216]}
   );
   gpc1_1 gpc3598 (
      {stage0_33[444]},
      {stage1_33[217]}
   );
   gpc1_1 gpc3599 (
      {stage0_33[445]},
      {stage1_33[218]}
   );
   gpc1_1 gpc3600 (
      {stage0_33[446]},
      {stage1_33[219]}
   );
   gpc1_1 gpc3601 (
      {stage0_33[447]},
      {stage1_33[220]}
   );
   gpc1_1 gpc3602 (
      {stage0_33[448]},
      {stage1_33[221]}
   );
   gpc1_1 gpc3603 (
      {stage0_33[449]},
      {stage1_33[222]}
   );
   gpc1_1 gpc3604 (
      {stage0_33[450]},
      {stage1_33[223]}
   );
   gpc1_1 gpc3605 (
      {stage0_33[451]},
      {stage1_33[224]}
   );
   gpc1_1 gpc3606 (
      {stage0_33[452]},
      {stage1_33[225]}
   );
   gpc1_1 gpc3607 (
      {stage0_33[453]},
      {stage1_33[226]}
   );
   gpc1_1 gpc3608 (
      {stage0_33[454]},
      {stage1_33[227]}
   );
   gpc1_1 gpc3609 (
      {stage0_33[455]},
      {stage1_33[228]}
   );
   gpc1_1 gpc3610 (
      {stage0_33[456]},
      {stage1_33[229]}
   );
   gpc1_1 gpc3611 (
      {stage0_33[457]},
      {stage1_33[230]}
   );
   gpc1_1 gpc3612 (
      {stage0_33[458]},
      {stage1_33[231]}
   );
   gpc1_1 gpc3613 (
      {stage0_33[459]},
      {stage1_33[232]}
   );
   gpc1_1 gpc3614 (
      {stage0_33[460]},
      {stage1_33[233]}
   );
   gpc1_1 gpc3615 (
      {stage0_33[461]},
      {stage1_33[234]}
   );
   gpc1_1 gpc3616 (
      {stage0_33[462]},
      {stage1_33[235]}
   );
   gpc1_1 gpc3617 (
      {stage0_33[463]},
      {stage1_33[236]}
   );
   gpc1_1 gpc3618 (
      {stage0_33[464]},
      {stage1_33[237]}
   );
   gpc1_1 gpc3619 (
      {stage0_33[465]},
      {stage1_33[238]}
   );
   gpc1_1 gpc3620 (
      {stage0_33[466]},
      {stage1_33[239]}
   );
   gpc1_1 gpc3621 (
      {stage0_33[467]},
      {stage1_33[240]}
   );
   gpc1_1 gpc3622 (
      {stage0_33[468]},
      {stage1_33[241]}
   );
   gpc1_1 gpc3623 (
      {stage0_33[469]},
      {stage1_33[242]}
   );
   gpc1_1 gpc3624 (
      {stage0_33[470]},
      {stage1_33[243]}
   );
   gpc1_1 gpc3625 (
      {stage0_33[471]},
      {stage1_33[244]}
   );
   gpc1_1 gpc3626 (
      {stage0_33[472]},
      {stage1_33[245]}
   );
   gpc1_1 gpc3627 (
      {stage0_33[473]},
      {stage1_33[246]}
   );
   gpc1_1 gpc3628 (
      {stage0_33[474]},
      {stage1_33[247]}
   );
   gpc1_1 gpc3629 (
      {stage0_33[475]},
      {stage1_33[248]}
   );
   gpc1_1 gpc3630 (
      {stage0_33[476]},
      {stage1_33[249]}
   );
   gpc1_1 gpc3631 (
      {stage0_33[477]},
      {stage1_33[250]}
   );
   gpc1_1 gpc3632 (
      {stage0_33[478]},
      {stage1_33[251]}
   );
   gpc1_1 gpc3633 (
      {stage0_33[479]},
      {stage1_33[252]}
   );
   gpc1_1 gpc3634 (
      {stage0_33[480]},
      {stage1_33[253]}
   );
   gpc1_1 gpc3635 (
      {stage0_33[481]},
      {stage1_33[254]}
   );
   gpc1_1 gpc3636 (
      {stage0_33[482]},
      {stage1_33[255]}
   );
   gpc1_1 gpc3637 (
      {stage0_33[483]},
      {stage1_33[256]}
   );
   gpc1_1 gpc3638 (
      {stage0_33[484]},
      {stage1_33[257]}
   );
   gpc1_1 gpc3639 (
      {stage0_33[485]},
      {stage1_33[258]}
   );
   gpc1_1 gpc3640 (
      {stage0_35[464]},
      {stage1_35[195]}
   );
   gpc1_1 gpc3641 (
      {stage0_35[465]},
      {stage1_35[196]}
   );
   gpc1_1 gpc3642 (
      {stage0_35[466]},
      {stage1_35[197]}
   );
   gpc1_1 gpc3643 (
      {stage0_35[467]},
      {stage1_35[198]}
   );
   gpc1_1 gpc3644 (
      {stage0_35[468]},
      {stage1_35[199]}
   );
   gpc1_1 gpc3645 (
      {stage0_35[469]},
      {stage1_35[200]}
   );
   gpc1_1 gpc3646 (
      {stage0_35[470]},
      {stage1_35[201]}
   );
   gpc1_1 gpc3647 (
      {stage0_35[471]},
      {stage1_35[202]}
   );
   gpc1_1 gpc3648 (
      {stage0_35[472]},
      {stage1_35[203]}
   );
   gpc1_1 gpc3649 (
      {stage0_35[473]},
      {stage1_35[204]}
   );
   gpc1_1 gpc3650 (
      {stage0_35[474]},
      {stage1_35[205]}
   );
   gpc1_1 gpc3651 (
      {stage0_35[475]},
      {stage1_35[206]}
   );
   gpc1_1 gpc3652 (
      {stage0_35[476]},
      {stage1_35[207]}
   );
   gpc1_1 gpc3653 (
      {stage0_35[477]},
      {stage1_35[208]}
   );
   gpc1_1 gpc3654 (
      {stage0_35[478]},
      {stage1_35[209]}
   );
   gpc1_1 gpc3655 (
      {stage0_35[479]},
      {stage1_35[210]}
   );
   gpc1_1 gpc3656 (
      {stage0_35[480]},
      {stage1_35[211]}
   );
   gpc1_1 gpc3657 (
      {stage0_35[481]},
      {stage1_35[212]}
   );
   gpc1_1 gpc3658 (
      {stage0_35[482]},
      {stage1_35[213]}
   );
   gpc1_1 gpc3659 (
      {stage0_35[483]},
      {stage1_35[214]}
   );
   gpc1_1 gpc3660 (
      {stage0_35[484]},
      {stage1_35[215]}
   );
   gpc1_1 gpc3661 (
      {stage0_35[485]},
      {stage1_35[216]}
   );
   gpc1_1 gpc3662 (
      {stage0_37[355]},
      {stage1_37[177]}
   );
   gpc1_1 gpc3663 (
      {stage0_37[356]},
      {stage1_37[178]}
   );
   gpc1_1 gpc3664 (
      {stage0_37[357]},
      {stage1_37[179]}
   );
   gpc1_1 gpc3665 (
      {stage0_37[358]},
      {stage1_37[180]}
   );
   gpc1_1 gpc3666 (
      {stage0_37[359]},
      {stage1_37[181]}
   );
   gpc1_1 gpc3667 (
      {stage0_37[360]},
      {stage1_37[182]}
   );
   gpc1_1 gpc3668 (
      {stage0_37[361]},
      {stage1_37[183]}
   );
   gpc1_1 gpc3669 (
      {stage0_37[362]},
      {stage1_37[184]}
   );
   gpc1_1 gpc3670 (
      {stage0_37[363]},
      {stage1_37[185]}
   );
   gpc1_1 gpc3671 (
      {stage0_37[364]},
      {stage1_37[186]}
   );
   gpc1_1 gpc3672 (
      {stage0_37[365]},
      {stage1_37[187]}
   );
   gpc1_1 gpc3673 (
      {stage0_37[366]},
      {stage1_37[188]}
   );
   gpc1_1 gpc3674 (
      {stage0_37[367]},
      {stage1_37[189]}
   );
   gpc1_1 gpc3675 (
      {stage0_37[368]},
      {stage1_37[190]}
   );
   gpc1_1 gpc3676 (
      {stage0_37[369]},
      {stage1_37[191]}
   );
   gpc1_1 gpc3677 (
      {stage0_37[370]},
      {stage1_37[192]}
   );
   gpc1_1 gpc3678 (
      {stage0_37[371]},
      {stage1_37[193]}
   );
   gpc1_1 gpc3679 (
      {stage0_37[372]},
      {stage1_37[194]}
   );
   gpc1_1 gpc3680 (
      {stage0_37[373]},
      {stage1_37[195]}
   );
   gpc1_1 gpc3681 (
      {stage0_37[374]},
      {stage1_37[196]}
   );
   gpc1_1 gpc3682 (
      {stage0_37[375]},
      {stage1_37[197]}
   );
   gpc1_1 gpc3683 (
      {stage0_37[376]},
      {stage1_37[198]}
   );
   gpc1_1 gpc3684 (
      {stage0_37[377]},
      {stage1_37[199]}
   );
   gpc1_1 gpc3685 (
      {stage0_37[378]},
      {stage1_37[200]}
   );
   gpc1_1 gpc3686 (
      {stage0_37[379]},
      {stage1_37[201]}
   );
   gpc1_1 gpc3687 (
      {stage0_37[380]},
      {stage1_37[202]}
   );
   gpc1_1 gpc3688 (
      {stage0_37[381]},
      {stage1_37[203]}
   );
   gpc1_1 gpc3689 (
      {stage0_37[382]},
      {stage1_37[204]}
   );
   gpc1_1 gpc3690 (
      {stage0_37[383]},
      {stage1_37[205]}
   );
   gpc1_1 gpc3691 (
      {stage0_37[384]},
      {stage1_37[206]}
   );
   gpc1_1 gpc3692 (
      {stage0_37[385]},
      {stage1_37[207]}
   );
   gpc1_1 gpc3693 (
      {stage0_37[386]},
      {stage1_37[208]}
   );
   gpc1_1 gpc3694 (
      {stage0_37[387]},
      {stage1_37[209]}
   );
   gpc1_1 gpc3695 (
      {stage0_37[388]},
      {stage1_37[210]}
   );
   gpc1_1 gpc3696 (
      {stage0_37[389]},
      {stage1_37[211]}
   );
   gpc1_1 gpc3697 (
      {stage0_37[390]},
      {stage1_37[212]}
   );
   gpc1_1 gpc3698 (
      {stage0_37[391]},
      {stage1_37[213]}
   );
   gpc1_1 gpc3699 (
      {stage0_37[392]},
      {stage1_37[214]}
   );
   gpc1_1 gpc3700 (
      {stage0_37[393]},
      {stage1_37[215]}
   );
   gpc1_1 gpc3701 (
      {stage0_37[394]},
      {stage1_37[216]}
   );
   gpc1_1 gpc3702 (
      {stage0_37[395]},
      {stage1_37[217]}
   );
   gpc1_1 gpc3703 (
      {stage0_37[396]},
      {stage1_37[218]}
   );
   gpc1_1 gpc3704 (
      {stage0_37[397]},
      {stage1_37[219]}
   );
   gpc1_1 gpc3705 (
      {stage0_37[398]},
      {stage1_37[220]}
   );
   gpc1_1 gpc3706 (
      {stage0_37[399]},
      {stage1_37[221]}
   );
   gpc1_1 gpc3707 (
      {stage0_37[400]},
      {stage1_37[222]}
   );
   gpc1_1 gpc3708 (
      {stage0_37[401]},
      {stage1_37[223]}
   );
   gpc1_1 gpc3709 (
      {stage0_37[402]},
      {stage1_37[224]}
   );
   gpc1_1 gpc3710 (
      {stage0_37[403]},
      {stage1_37[225]}
   );
   gpc1_1 gpc3711 (
      {stage0_37[404]},
      {stage1_37[226]}
   );
   gpc1_1 gpc3712 (
      {stage0_37[405]},
      {stage1_37[227]}
   );
   gpc1_1 gpc3713 (
      {stage0_37[406]},
      {stage1_37[228]}
   );
   gpc1_1 gpc3714 (
      {stage0_37[407]},
      {stage1_37[229]}
   );
   gpc1_1 gpc3715 (
      {stage0_37[408]},
      {stage1_37[230]}
   );
   gpc1_1 gpc3716 (
      {stage0_37[409]},
      {stage1_37[231]}
   );
   gpc1_1 gpc3717 (
      {stage0_37[410]},
      {stage1_37[232]}
   );
   gpc1_1 gpc3718 (
      {stage0_37[411]},
      {stage1_37[233]}
   );
   gpc1_1 gpc3719 (
      {stage0_37[412]},
      {stage1_37[234]}
   );
   gpc1_1 gpc3720 (
      {stage0_37[413]},
      {stage1_37[235]}
   );
   gpc1_1 gpc3721 (
      {stage0_37[414]},
      {stage1_37[236]}
   );
   gpc1_1 gpc3722 (
      {stage0_37[415]},
      {stage1_37[237]}
   );
   gpc1_1 gpc3723 (
      {stage0_37[416]},
      {stage1_37[238]}
   );
   gpc1_1 gpc3724 (
      {stage0_37[417]},
      {stage1_37[239]}
   );
   gpc1_1 gpc3725 (
      {stage0_37[418]},
      {stage1_37[240]}
   );
   gpc1_1 gpc3726 (
      {stage0_37[419]},
      {stage1_37[241]}
   );
   gpc1_1 gpc3727 (
      {stage0_37[420]},
      {stage1_37[242]}
   );
   gpc1_1 gpc3728 (
      {stage0_37[421]},
      {stage1_37[243]}
   );
   gpc1_1 gpc3729 (
      {stage0_37[422]},
      {stage1_37[244]}
   );
   gpc1_1 gpc3730 (
      {stage0_37[423]},
      {stage1_37[245]}
   );
   gpc1_1 gpc3731 (
      {stage0_37[424]},
      {stage1_37[246]}
   );
   gpc1_1 gpc3732 (
      {stage0_37[425]},
      {stage1_37[247]}
   );
   gpc1_1 gpc3733 (
      {stage0_37[426]},
      {stage1_37[248]}
   );
   gpc1_1 gpc3734 (
      {stage0_37[427]},
      {stage1_37[249]}
   );
   gpc1_1 gpc3735 (
      {stage0_37[428]},
      {stage1_37[250]}
   );
   gpc1_1 gpc3736 (
      {stage0_37[429]},
      {stage1_37[251]}
   );
   gpc1_1 gpc3737 (
      {stage0_37[430]},
      {stage1_37[252]}
   );
   gpc1_1 gpc3738 (
      {stage0_37[431]},
      {stage1_37[253]}
   );
   gpc1_1 gpc3739 (
      {stage0_37[432]},
      {stage1_37[254]}
   );
   gpc1_1 gpc3740 (
      {stage0_37[433]},
      {stage1_37[255]}
   );
   gpc1_1 gpc3741 (
      {stage0_37[434]},
      {stage1_37[256]}
   );
   gpc1_1 gpc3742 (
      {stage0_37[435]},
      {stage1_37[257]}
   );
   gpc1_1 gpc3743 (
      {stage0_37[436]},
      {stage1_37[258]}
   );
   gpc1_1 gpc3744 (
      {stage0_37[437]},
      {stage1_37[259]}
   );
   gpc1_1 gpc3745 (
      {stage0_37[438]},
      {stage1_37[260]}
   );
   gpc1_1 gpc3746 (
      {stage0_37[439]},
      {stage1_37[261]}
   );
   gpc1_1 gpc3747 (
      {stage0_37[440]},
      {stage1_37[262]}
   );
   gpc1_1 gpc3748 (
      {stage0_37[441]},
      {stage1_37[263]}
   );
   gpc1_1 gpc3749 (
      {stage0_37[442]},
      {stage1_37[264]}
   );
   gpc1_1 gpc3750 (
      {stage0_37[443]},
      {stage1_37[265]}
   );
   gpc1_1 gpc3751 (
      {stage0_37[444]},
      {stage1_37[266]}
   );
   gpc1_1 gpc3752 (
      {stage0_37[445]},
      {stage1_37[267]}
   );
   gpc1_1 gpc3753 (
      {stage0_37[446]},
      {stage1_37[268]}
   );
   gpc1_1 gpc3754 (
      {stage0_37[447]},
      {stage1_37[269]}
   );
   gpc1_1 gpc3755 (
      {stage0_37[448]},
      {stage1_37[270]}
   );
   gpc1_1 gpc3756 (
      {stage0_37[449]},
      {stage1_37[271]}
   );
   gpc1_1 gpc3757 (
      {stage0_37[450]},
      {stage1_37[272]}
   );
   gpc1_1 gpc3758 (
      {stage0_37[451]},
      {stage1_37[273]}
   );
   gpc1_1 gpc3759 (
      {stage0_37[452]},
      {stage1_37[274]}
   );
   gpc1_1 gpc3760 (
      {stage0_37[453]},
      {stage1_37[275]}
   );
   gpc1_1 gpc3761 (
      {stage0_37[454]},
      {stage1_37[276]}
   );
   gpc1_1 gpc3762 (
      {stage0_37[455]},
      {stage1_37[277]}
   );
   gpc1_1 gpc3763 (
      {stage0_37[456]},
      {stage1_37[278]}
   );
   gpc1_1 gpc3764 (
      {stage0_37[457]},
      {stage1_37[279]}
   );
   gpc1_1 gpc3765 (
      {stage0_37[458]},
      {stage1_37[280]}
   );
   gpc1_1 gpc3766 (
      {stage0_37[459]},
      {stage1_37[281]}
   );
   gpc1_1 gpc3767 (
      {stage0_37[460]},
      {stage1_37[282]}
   );
   gpc1_1 gpc3768 (
      {stage0_37[461]},
      {stage1_37[283]}
   );
   gpc1_1 gpc3769 (
      {stage0_37[462]},
      {stage1_37[284]}
   );
   gpc1_1 gpc3770 (
      {stage0_37[463]},
      {stage1_37[285]}
   );
   gpc1_1 gpc3771 (
      {stage0_37[464]},
      {stage1_37[286]}
   );
   gpc1_1 gpc3772 (
      {stage0_37[465]},
      {stage1_37[287]}
   );
   gpc1_1 gpc3773 (
      {stage0_37[466]},
      {stage1_37[288]}
   );
   gpc1_1 gpc3774 (
      {stage0_37[467]},
      {stage1_37[289]}
   );
   gpc1_1 gpc3775 (
      {stage0_37[468]},
      {stage1_37[290]}
   );
   gpc1_1 gpc3776 (
      {stage0_37[469]},
      {stage1_37[291]}
   );
   gpc1_1 gpc3777 (
      {stage0_37[470]},
      {stage1_37[292]}
   );
   gpc1_1 gpc3778 (
      {stage0_37[471]},
      {stage1_37[293]}
   );
   gpc1_1 gpc3779 (
      {stage0_37[472]},
      {stage1_37[294]}
   );
   gpc1_1 gpc3780 (
      {stage0_37[473]},
      {stage1_37[295]}
   );
   gpc1_1 gpc3781 (
      {stage0_37[474]},
      {stage1_37[296]}
   );
   gpc1_1 gpc3782 (
      {stage0_37[475]},
      {stage1_37[297]}
   );
   gpc1_1 gpc3783 (
      {stage0_37[476]},
      {stage1_37[298]}
   );
   gpc1_1 gpc3784 (
      {stage0_37[477]},
      {stage1_37[299]}
   );
   gpc1_1 gpc3785 (
      {stage0_37[478]},
      {stage1_37[300]}
   );
   gpc1_1 gpc3786 (
      {stage0_37[479]},
      {stage1_37[301]}
   );
   gpc1_1 gpc3787 (
      {stage0_37[480]},
      {stage1_37[302]}
   );
   gpc1_1 gpc3788 (
      {stage0_37[481]},
      {stage1_37[303]}
   );
   gpc1_1 gpc3789 (
      {stage0_37[482]},
      {stage1_37[304]}
   );
   gpc1_1 gpc3790 (
      {stage0_37[483]},
      {stage1_37[305]}
   );
   gpc1_1 gpc3791 (
      {stage0_37[484]},
      {stage1_37[306]}
   );
   gpc1_1 gpc3792 (
      {stage0_37[485]},
      {stage1_37[307]}
   );
   gpc1_1 gpc3793 (
      {stage0_38[391]},
      {stage1_38[170]}
   );
   gpc1_1 gpc3794 (
      {stage0_38[392]},
      {stage1_38[171]}
   );
   gpc1_1 gpc3795 (
      {stage0_38[393]},
      {stage1_38[172]}
   );
   gpc1_1 gpc3796 (
      {stage0_38[394]},
      {stage1_38[173]}
   );
   gpc1_1 gpc3797 (
      {stage0_38[395]},
      {stage1_38[174]}
   );
   gpc1_1 gpc3798 (
      {stage0_38[396]},
      {stage1_38[175]}
   );
   gpc1_1 gpc3799 (
      {stage0_38[397]},
      {stage1_38[176]}
   );
   gpc1_1 gpc3800 (
      {stage0_38[398]},
      {stage1_38[177]}
   );
   gpc1_1 gpc3801 (
      {stage0_38[399]},
      {stage1_38[178]}
   );
   gpc1_1 gpc3802 (
      {stage0_38[400]},
      {stage1_38[179]}
   );
   gpc1_1 gpc3803 (
      {stage0_38[401]},
      {stage1_38[180]}
   );
   gpc1_1 gpc3804 (
      {stage0_38[402]},
      {stage1_38[181]}
   );
   gpc1_1 gpc3805 (
      {stage0_38[403]},
      {stage1_38[182]}
   );
   gpc1_1 gpc3806 (
      {stage0_38[404]},
      {stage1_38[183]}
   );
   gpc1_1 gpc3807 (
      {stage0_38[405]},
      {stage1_38[184]}
   );
   gpc1_1 gpc3808 (
      {stage0_38[406]},
      {stage1_38[185]}
   );
   gpc1_1 gpc3809 (
      {stage0_38[407]},
      {stage1_38[186]}
   );
   gpc1_1 gpc3810 (
      {stage0_38[408]},
      {stage1_38[187]}
   );
   gpc1_1 gpc3811 (
      {stage0_38[409]},
      {stage1_38[188]}
   );
   gpc1_1 gpc3812 (
      {stage0_38[410]},
      {stage1_38[189]}
   );
   gpc1_1 gpc3813 (
      {stage0_38[411]},
      {stage1_38[190]}
   );
   gpc1_1 gpc3814 (
      {stage0_38[412]},
      {stage1_38[191]}
   );
   gpc1_1 gpc3815 (
      {stage0_38[413]},
      {stage1_38[192]}
   );
   gpc1_1 gpc3816 (
      {stage0_38[414]},
      {stage1_38[193]}
   );
   gpc1_1 gpc3817 (
      {stage0_38[415]},
      {stage1_38[194]}
   );
   gpc1_1 gpc3818 (
      {stage0_38[416]},
      {stage1_38[195]}
   );
   gpc1_1 gpc3819 (
      {stage0_38[417]},
      {stage1_38[196]}
   );
   gpc1_1 gpc3820 (
      {stage0_38[418]},
      {stage1_38[197]}
   );
   gpc1_1 gpc3821 (
      {stage0_38[419]},
      {stage1_38[198]}
   );
   gpc1_1 gpc3822 (
      {stage0_38[420]},
      {stage1_38[199]}
   );
   gpc1_1 gpc3823 (
      {stage0_38[421]},
      {stage1_38[200]}
   );
   gpc1_1 gpc3824 (
      {stage0_38[422]},
      {stage1_38[201]}
   );
   gpc1_1 gpc3825 (
      {stage0_38[423]},
      {stage1_38[202]}
   );
   gpc1_1 gpc3826 (
      {stage0_38[424]},
      {stage1_38[203]}
   );
   gpc1_1 gpc3827 (
      {stage0_38[425]},
      {stage1_38[204]}
   );
   gpc1_1 gpc3828 (
      {stage0_38[426]},
      {stage1_38[205]}
   );
   gpc1_1 gpc3829 (
      {stage0_38[427]},
      {stage1_38[206]}
   );
   gpc1_1 gpc3830 (
      {stage0_38[428]},
      {stage1_38[207]}
   );
   gpc1_1 gpc3831 (
      {stage0_38[429]},
      {stage1_38[208]}
   );
   gpc1_1 gpc3832 (
      {stage0_38[430]},
      {stage1_38[209]}
   );
   gpc1_1 gpc3833 (
      {stage0_38[431]},
      {stage1_38[210]}
   );
   gpc1_1 gpc3834 (
      {stage0_38[432]},
      {stage1_38[211]}
   );
   gpc1_1 gpc3835 (
      {stage0_38[433]},
      {stage1_38[212]}
   );
   gpc1_1 gpc3836 (
      {stage0_38[434]},
      {stage1_38[213]}
   );
   gpc1_1 gpc3837 (
      {stage0_38[435]},
      {stage1_38[214]}
   );
   gpc1_1 gpc3838 (
      {stage0_38[436]},
      {stage1_38[215]}
   );
   gpc1_1 gpc3839 (
      {stage0_38[437]},
      {stage1_38[216]}
   );
   gpc1_1 gpc3840 (
      {stage0_38[438]},
      {stage1_38[217]}
   );
   gpc1_1 gpc3841 (
      {stage0_38[439]},
      {stage1_38[218]}
   );
   gpc1_1 gpc3842 (
      {stage0_38[440]},
      {stage1_38[219]}
   );
   gpc1_1 gpc3843 (
      {stage0_38[441]},
      {stage1_38[220]}
   );
   gpc1_1 gpc3844 (
      {stage0_38[442]},
      {stage1_38[221]}
   );
   gpc1_1 gpc3845 (
      {stage0_38[443]},
      {stage1_38[222]}
   );
   gpc1_1 gpc3846 (
      {stage0_38[444]},
      {stage1_38[223]}
   );
   gpc1_1 gpc3847 (
      {stage0_38[445]},
      {stage1_38[224]}
   );
   gpc1_1 gpc3848 (
      {stage0_38[446]},
      {stage1_38[225]}
   );
   gpc1_1 gpc3849 (
      {stage0_38[447]},
      {stage1_38[226]}
   );
   gpc1_1 gpc3850 (
      {stage0_38[448]},
      {stage1_38[227]}
   );
   gpc1_1 gpc3851 (
      {stage0_38[449]},
      {stage1_38[228]}
   );
   gpc1_1 gpc3852 (
      {stage0_38[450]},
      {stage1_38[229]}
   );
   gpc1_1 gpc3853 (
      {stage0_38[451]},
      {stage1_38[230]}
   );
   gpc1_1 gpc3854 (
      {stage0_38[452]},
      {stage1_38[231]}
   );
   gpc1_1 gpc3855 (
      {stage0_38[453]},
      {stage1_38[232]}
   );
   gpc1_1 gpc3856 (
      {stage0_38[454]},
      {stage1_38[233]}
   );
   gpc1_1 gpc3857 (
      {stage0_38[455]},
      {stage1_38[234]}
   );
   gpc1_1 gpc3858 (
      {stage0_38[456]},
      {stage1_38[235]}
   );
   gpc1_1 gpc3859 (
      {stage0_38[457]},
      {stage1_38[236]}
   );
   gpc1_1 gpc3860 (
      {stage0_38[458]},
      {stage1_38[237]}
   );
   gpc1_1 gpc3861 (
      {stage0_38[459]},
      {stage1_38[238]}
   );
   gpc1_1 gpc3862 (
      {stage0_38[460]},
      {stage1_38[239]}
   );
   gpc1_1 gpc3863 (
      {stage0_38[461]},
      {stage1_38[240]}
   );
   gpc1_1 gpc3864 (
      {stage0_38[462]},
      {stage1_38[241]}
   );
   gpc1_1 gpc3865 (
      {stage0_38[463]},
      {stage1_38[242]}
   );
   gpc1_1 gpc3866 (
      {stage0_38[464]},
      {stage1_38[243]}
   );
   gpc1_1 gpc3867 (
      {stage0_38[465]},
      {stage1_38[244]}
   );
   gpc1_1 gpc3868 (
      {stage0_38[466]},
      {stage1_38[245]}
   );
   gpc1_1 gpc3869 (
      {stage0_38[467]},
      {stage1_38[246]}
   );
   gpc1_1 gpc3870 (
      {stage0_38[468]},
      {stage1_38[247]}
   );
   gpc1_1 gpc3871 (
      {stage0_38[469]},
      {stage1_38[248]}
   );
   gpc1_1 gpc3872 (
      {stage0_38[470]},
      {stage1_38[249]}
   );
   gpc1_1 gpc3873 (
      {stage0_38[471]},
      {stage1_38[250]}
   );
   gpc1_1 gpc3874 (
      {stage0_38[472]},
      {stage1_38[251]}
   );
   gpc1_1 gpc3875 (
      {stage0_38[473]},
      {stage1_38[252]}
   );
   gpc1_1 gpc3876 (
      {stage0_38[474]},
      {stage1_38[253]}
   );
   gpc1_1 gpc3877 (
      {stage0_38[475]},
      {stage1_38[254]}
   );
   gpc1_1 gpc3878 (
      {stage0_38[476]},
      {stage1_38[255]}
   );
   gpc1_1 gpc3879 (
      {stage0_38[477]},
      {stage1_38[256]}
   );
   gpc1_1 gpc3880 (
      {stage0_38[478]},
      {stage1_38[257]}
   );
   gpc1_1 gpc3881 (
      {stage0_38[479]},
      {stage1_38[258]}
   );
   gpc1_1 gpc3882 (
      {stage0_38[480]},
      {stage1_38[259]}
   );
   gpc1_1 gpc3883 (
      {stage0_38[481]},
      {stage1_38[260]}
   );
   gpc1_1 gpc3884 (
      {stage0_38[482]},
      {stage1_38[261]}
   );
   gpc1_1 gpc3885 (
      {stage0_38[483]},
      {stage1_38[262]}
   );
   gpc1_1 gpc3886 (
      {stage0_38[484]},
      {stage1_38[263]}
   );
   gpc1_1 gpc3887 (
      {stage0_38[485]},
      {stage1_38[264]}
   );
   gpc1_1 gpc3888 (
      {stage0_39[447]},
      {stage1_39[174]}
   );
   gpc1_1 gpc3889 (
      {stage0_39[448]},
      {stage1_39[175]}
   );
   gpc1_1 gpc3890 (
      {stage0_39[449]},
      {stage1_39[176]}
   );
   gpc1_1 gpc3891 (
      {stage0_39[450]},
      {stage1_39[177]}
   );
   gpc1_1 gpc3892 (
      {stage0_39[451]},
      {stage1_39[178]}
   );
   gpc1_1 gpc3893 (
      {stage0_39[452]},
      {stage1_39[179]}
   );
   gpc1_1 gpc3894 (
      {stage0_39[453]},
      {stage1_39[180]}
   );
   gpc1_1 gpc3895 (
      {stage0_39[454]},
      {stage1_39[181]}
   );
   gpc1_1 gpc3896 (
      {stage0_39[455]},
      {stage1_39[182]}
   );
   gpc1_1 gpc3897 (
      {stage0_39[456]},
      {stage1_39[183]}
   );
   gpc1_1 gpc3898 (
      {stage0_39[457]},
      {stage1_39[184]}
   );
   gpc1_1 gpc3899 (
      {stage0_39[458]},
      {stage1_39[185]}
   );
   gpc1_1 gpc3900 (
      {stage0_39[459]},
      {stage1_39[186]}
   );
   gpc1_1 gpc3901 (
      {stage0_39[460]},
      {stage1_39[187]}
   );
   gpc1_1 gpc3902 (
      {stage0_39[461]},
      {stage1_39[188]}
   );
   gpc1_1 gpc3903 (
      {stage0_39[462]},
      {stage1_39[189]}
   );
   gpc1_1 gpc3904 (
      {stage0_39[463]},
      {stage1_39[190]}
   );
   gpc1_1 gpc3905 (
      {stage0_39[464]},
      {stage1_39[191]}
   );
   gpc1_1 gpc3906 (
      {stage0_39[465]},
      {stage1_39[192]}
   );
   gpc1_1 gpc3907 (
      {stage0_39[466]},
      {stage1_39[193]}
   );
   gpc1_1 gpc3908 (
      {stage0_39[467]},
      {stage1_39[194]}
   );
   gpc1_1 gpc3909 (
      {stage0_39[468]},
      {stage1_39[195]}
   );
   gpc1_1 gpc3910 (
      {stage0_39[469]},
      {stage1_39[196]}
   );
   gpc1_1 gpc3911 (
      {stage0_39[470]},
      {stage1_39[197]}
   );
   gpc1_1 gpc3912 (
      {stage0_39[471]},
      {stage1_39[198]}
   );
   gpc1_1 gpc3913 (
      {stage0_39[472]},
      {stage1_39[199]}
   );
   gpc1_1 gpc3914 (
      {stage0_39[473]},
      {stage1_39[200]}
   );
   gpc1_1 gpc3915 (
      {stage0_39[474]},
      {stage1_39[201]}
   );
   gpc1_1 gpc3916 (
      {stage0_39[475]},
      {stage1_39[202]}
   );
   gpc1_1 gpc3917 (
      {stage0_39[476]},
      {stage1_39[203]}
   );
   gpc1_1 gpc3918 (
      {stage0_39[477]},
      {stage1_39[204]}
   );
   gpc1_1 gpc3919 (
      {stage0_39[478]},
      {stage1_39[205]}
   );
   gpc1_1 gpc3920 (
      {stage0_39[479]},
      {stage1_39[206]}
   );
   gpc1_1 gpc3921 (
      {stage0_39[480]},
      {stage1_39[207]}
   );
   gpc1_1 gpc3922 (
      {stage0_39[481]},
      {stage1_39[208]}
   );
   gpc1_1 gpc3923 (
      {stage0_39[482]},
      {stage1_39[209]}
   );
   gpc1_1 gpc3924 (
      {stage0_39[483]},
      {stage1_39[210]}
   );
   gpc1_1 gpc3925 (
      {stage0_39[484]},
      {stage1_39[211]}
   );
   gpc1_1 gpc3926 (
      {stage0_39[485]},
      {stage1_39[212]}
   );
   gpc1_1 gpc3927 (
      {stage0_40[380]},
      {stage1_40[198]}
   );
   gpc1_1 gpc3928 (
      {stage0_40[381]},
      {stage1_40[199]}
   );
   gpc1_1 gpc3929 (
      {stage0_40[382]},
      {stage1_40[200]}
   );
   gpc1_1 gpc3930 (
      {stage0_40[383]},
      {stage1_40[201]}
   );
   gpc1_1 gpc3931 (
      {stage0_40[384]},
      {stage1_40[202]}
   );
   gpc1_1 gpc3932 (
      {stage0_40[385]},
      {stage1_40[203]}
   );
   gpc1_1 gpc3933 (
      {stage0_40[386]},
      {stage1_40[204]}
   );
   gpc1_1 gpc3934 (
      {stage0_40[387]},
      {stage1_40[205]}
   );
   gpc1_1 gpc3935 (
      {stage0_40[388]},
      {stage1_40[206]}
   );
   gpc1_1 gpc3936 (
      {stage0_40[389]},
      {stage1_40[207]}
   );
   gpc1_1 gpc3937 (
      {stage0_40[390]},
      {stage1_40[208]}
   );
   gpc1_1 gpc3938 (
      {stage0_40[391]},
      {stage1_40[209]}
   );
   gpc1_1 gpc3939 (
      {stage0_40[392]},
      {stage1_40[210]}
   );
   gpc1_1 gpc3940 (
      {stage0_40[393]},
      {stage1_40[211]}
   );
   gpc1_1 gpc3941 (
      {stage0_40[394]},
      {stage1_40[212]}
   );
   gpc1_1 gpc3942 (
      {stage0_40[395]},
      {stage1_40[213]}
   );
   gpc1_1 gpc3943 (
      {stage0_40[396]},
      {stage1_40[214]}
   );
   gpc1_1 gpc3944 (
      {stage0_40[397]},
      {stage1_40[215]}
   );
   gpc1_1 gpc3945 (
      {stage0_40[398]},
      {stage1_40[216]}
   );
   gpc1_1 gpc3946 (
      {stage0_40[399]},
      {stage1_40[217]}
   );
   gpc1_1 gpc3947 (
      {stage0_40[400]},
      {stage1_40[218]}
   );
   gpc1_1 gpc3948 (
      {stage0_40[401]},
      {stage1_40[219]}
   );
   gpc1_1 gpc3949 (
      {stage0_40[402]},
      {stage1_40[220]}
   );
   gpc1_1 gpc3950 (
      {stage0_40[403]},
      {stage1_40[221]}
   );
   gpc1_1 gpc3951 (
      {stage0_40[404]},
      {stage1_40[222]}
   );
   gpc1_1 gpc3952 (
      {stage0_40[405]},
      {stage1_40[223]}
   );
   gpc1_1 gpc3953 (
      {stage0_40[406]},
      {stage1_40[224]}
   );
   gpc1_1 gpc3954 (
      {stage0_40[407]},
      {stage1_40[225]}
   );
   gpc1_1 gpc3955 (
      {stage0_40[408]},
      {stage1_40[226]}
   );
   gpc1_1 gpc3956 (
      {stage0_40[409]},
      {stage1_40[227]}
   );
   gpc1_1 gpc3957 (
      {stage0_40[410]},
      {stage1_40[228]}
   );
   gpc1_1 gpc3958 (
      {stage0_40[411]},
      {stage1_40[229]}
   );
   gpc1_1 gpc3959 (
      {stage0_40[412]},
      {stage1_40[230]}
   );
   gpc1_1 gpc3960 (
      {stage0_40[413]},
      {stage1_40[231]}
   );
   gpc1_1 gpc3961 (
      {stage0_40[414]},
      {stage1_40[232]}
   );
   gpc1_1 gpc3962 (
      {stage0_40[415]},
      {stage1_40[233]}
   );
   gpc1_1 gpc3963 (
      {stage0_40[416]},
      {stage1_40[234]}
   );
   gpc1_1 gpc3964 (
      {stage0_40[417]},
      {stage1_40[235]}
   );
   gpc1_1 gpc3965 (
      {stage0_40[418]},
      {stage1_40[236]}
   );
   gpc1_1 gpc3966 (
      {stage0_40[419]},
      {stage1_40[237]}
   );
   gpc1_1 gpc3967 (
      {stage0_40[420]},
      {stage1_40[238]}
   );
   gpc1_1 gpc3968 (
      {stage0_40[421]},
      {stage1_40[239]}
   );
   gpc1_1 gpc3969 (
      {stage0_40[422]},
      {stage1_40[240]}
   );
   gpc1_1 gpc3970 (
      {stage0_40[423]},
      {stage1_40[241]}
   );
   gpc1_1 gpc3971 (
      {stage0_40[424]},
      {stage1_40[242]}
   );
   gpc1_1 gpc3972 (
      {stage0_40[425]},
      {stage1_40[243]}
   );
   gpc1_1 gpc3973 (
      {stage0_40[426]},
      {stage1_40[244]}
   );
   gpc1_1 gpc3974 (
      {stage0_40[427]},
      {stage1_40[245]}
   );
   gpc1_1 gpc3975 (
      {stage0_40[428]},
      {stage1_40[246]}
   );
   gpc1_1 gpc3976 (
      {stage0_40[429]},
      {stage1_40[247]}
   );
   gpc1_1 gpc3977 (
      {stage0_40[430]},
      {stage1_40[248]}
   );
   gpc1_1 gpc3978 (
      {stage0_40[431]},
      {stage1_40[249]}
   );
   gpc1_1 gpc3979 (
      {stage0_40[432]},
      {stage1_40[250]}
   );
   gpc1_1 gpc3980 (
      {stage0_40[433]},
      {stage1_40[251]}
   );
   gpc1_1 gpc3981 (
      {stage0_40[434]},
      {stage1_40[252]}
   );
   gpc1_1 gpc3982 (
      {stage0_40[435]},
      {stage1_40[253]}
   );
   gpc1_1 gpc3983 (
      {stage0_40[436]},
      {stage1_40[254]}
   );
   gpc1_1 gpc3984 (
      {stage0_40[437]},
      {stage1_40[255]}
   );
   gpc1_1 gpc3985 (
      {stage0_40[438]},
      {stage1_40[256]}
   );
   gpc1_1 gpc3986 (
      {stage0_40[439]},
      {stage1_40[257]}
   );
   gpc1_1 gpc3987 (
      {stage0_40[440]},
      {stage1_40[258]}
   );
   gpc1_1 gpc3988 (
      {stage0_40[441]},
      {stage1_40[259]}
   );
   gpc1_1 gpc3989 (
      {stage0_40[442]},
      {stage1_40[260]}
   );
   gpc1_1 gpc3990 (
      {stage0_40[443]},
      {stage1_40[261]}
   );
   gpc1_1 gpc3991 (
      {stage0_40[444]},
      {stage1_40[262]}
   );
   gpc1_1 gpc3992 (
      {stage0_40[445]},
      {stage1_40[263]}
   );
   gpc1_1 gpc3993 (
      {stage0_40[446]},
      {stage1_40[264]}
   );
   gpc1_1 gpc3994 (
      {stage0_40[447]},
      {stage1_40[265]}
   );
   gpc1_1 gpc3995 (
      {stage0_40[448]},
      {stage1_40[266]}
   );
   gpc1_1 gpc3996 (
      {stage0_40[449]},
      {stage1_40[267]}
   );
   gpc1_1 gpc3997 (
      {stage0_40[450]},
      {stage1_40[268]}
   );
   gpc1_1 gpc3998 (
      {stage0_40[451]},
      {stage1_40[269]}
   );
   gpc1_1 gpc3999 (
      {stage0_40[452]},
      {stage1_40[270]}
   );
   gpc1_1 gpc4000 (
      {stage0_40[453]},
      {stage1_40[271]}
   );
   gpc1_1 gpc4001 (
      {stage0_40[454]},
      {stage1_40[272]}
   );
   gpc1_1 gpc4002 (
      {stage0_40[455]},
      {stage1_40[273]}
   );
   gpc1_1 gpc4003 (
      {stage0_40[456]},
      {stage1_40[274]}
   );
   gpc1_1 gpc4004 (
      {stage0_40[457]},
      {stage1_40[275]}
   );
   gpc1_1 gpc4005 (
      {stage0_40[458]},
      {stage1_40[276]}
   );
   gpc1_1 gpc4006 (
      {stage0_40[459]},
      {stage1_40[277]}
   );
   gpc1_1 gpc4007 (
      {stage0_40[460]},
      {stage1_40[278]}
   );
   gpc1_1 gpc4008 (
      {stage0_40[461]},
      {stage1_40[279]}
   );
   gpc1_1 gpc4009 (
      {stage0_40[462]},
      {stage1_40[280]}
   );
   gpc1_1 gpc4010 (
      {stage0_40[463]},
      {stage1_40[281]}
   );
   gpc1_1 gpc4011 (
      {stage0_40[464]},
      {stage1_40[282]}
   );
   gpc1_1 gpc4012 (
      {stage0_40[465]},
      {stage1_40[283]}
   );
   gpc1_1 gpc4013 (
      {stage0_40[466]},
      {stage1_40[284]}
   );
   gpc1_1 gpc4014 (
      {stage0_40[467]},
      {stage1_40[285]}
   );
   gpc1_1 gpc4015 (
      {stage0_40[468]},
      {stage1_40[286]}
   );
   gpc1_1 gpc4016 (
      {stage0_40[469]},
      {stage1_40[287]}
   );
   gpc1_1 gpc4017 (
      {stage0_40[470]},
      {stage1_40[288]}
   );
   gpc1_1 gpc4018 (
      {stage0_40[471]},
      {stage1_40[289]}
   );
   gpc1_1 gpc4019 (
      {stage0_40[472]},
      {stage1_40[290]}
   );
   gpc1_1 gpc4020 (
      {stage0_40[473]},
      {stage1_40[291]}
   );
   gpc1_1 gpc4021 (
      {stage0_40[474]},
      {stage1_40[292]}
   );
   gpc1_1 gpc4022 (
      {stage0_40[475]},
      {stage1_40[293]}
   );
   gpc1_1 gpc4023 (
      {stage0_40[476]},
      {stage1_40[294]}
   );
   gpc1_1 gpc4024 (
      {stage0_40[477]},
      {stage1_40[295]}
   );
   gpc1_1 gpc4025 (
      {stage0_40[478]},
      {stage1_40[296]}
   );
   gpc1_1 gpc4026 (
      {stage0_40[479]},
      {stage1_40[297]}
   );
   gpc1_1 gpc4027 (
      {stage0_40[480]},
      {stage1_40[298]}
   );
   gpc1_1 gpc4028 (
      {stage0_40[481]},
      {stage1_40[299]}
   );
   gpc1_1 gpc4029 (
      {stage0_40[482]},
      {stage1_40[300]}
   );
   gpc1_1 gpc4030 (
      {stage0_40[483]},
      {stage1_40[301]}
   );
   gpc1_1 gpc4031 (
      {stage0_40[484]},
      {stage1_40[302]}
   );
   gpc1_1 gpc4032 (
      {stage0_40[485]},
      {stage1_40[303]}
   );
   gpc1_1 gpc4033 (
      {stage0_41[477]},
      {stage1_41[162]}
   );
   gpc1_1 gpc4034 (
      {stage0_41[478]},
      {stage1_41[163]}
   );
   gpc1_1 gpc4035 (
      {stage0_41[479]},
      {stage1_41[164]}
   );
   gpc1_1 gpc4036 (
      {stage0_41[480]},
      {stage1_41[165]}
   );
   gpc1_1 gpc4037 (
      {stage0_41[481]},
      {stage1_41[166]}
   );
   gpc1_1 gpc4038 (
      {stage0_41[482]},
      {stage1_41[167]}
   );
   gpc1_1 gpc4039 (
      {stage0_41[483]},
      {stage1_41[168]}
   );
   gpc1_1 gpc4040 (
      {stage0_41[484]},
      {stage1_41[169]}
   );
   gpc1_1 gpc4041 (
      {stage0_41[485]},
      {stage1_41[170]}
   );
   gpc1_1 gpc4042 (
      {stage0_42[483]},
      {stage1_42[171]}
   );
   gpc1_1 gpc4043 (
      {stage0_42[484]},
      {stage1_42[172]}
   );
   gpc1_1 gpc4044 (
      {stage0_42[485]},
      {stage1_42[173]}
   );
   gpc1_1 gpc4045 (
      {stage0_43[451]},
      {stage1_43[219]}
   );
   gpc1_1 gpc4046 (
      {stage0_43[452]},
      {stage1_43[220]}
   );
   gpc1_1 gpc4047 (
      {stage0_43[453]},
      {stage1_43[221]}
   );
   gpc1_1 gpc4048 (
      {stage0_43[454]},
      {stage1_43[222]}
   );
   gpc1_1 gpc4049 (
      {stage0_43[455]},
      {stage1_43[223]}
   );
   gpc1_1 gpc4050 (
      {stage0_43[456]},
      {stage1_43[224]}
   );
   gpc1_1 gpc4051 (
      {stage0_43[457]},
      {stage1_43[225]}
   );
   gpc1_1 gpc4052 (
      {stage0_43[458]},
      {stage1_43[226]}
   );
   gpc1_1 gpc4053 (
      {stage0_43[459]},
      {stage1_43[227]}
   );
   gpc1_1 gpc4054 (
      {stage0_43[460]},
      {stage1_43[228]}
   );
   gpc1_1 gpc4055 (
      {stage0_43[461]},
      {stage1_43[229]}
   );
   gpc1_1 gpc4056 (
      {stage0_43[462]},
      {stage1_43[230]}
   );
   gpc1_1 gpc4057 (
      {stage0_43[463]},
      {stage1_43[231]}
   );
   gpc1_1 gpc4058 (
      {stage0_43[464]},
      {stage1_43[232]}
   );
   gpc1_1 gpc4059 (
      {stage0_43[465]},
      {stage1_43[233]}
   );
   gpc1_1 gpc4060 (
      {stage0_43[466]},
      {stage1_43[234]}
   );
   gpc1_1 gpc4061 (
      {stage0_43[467]},
      {stage1_43[235]}
   );
   gpc1_1 gpc4062 (
      {stage0_43[468]},
      {stage1_43[236]}
   );
   gpc1_1 gpc4063 (
      {stage0_43[469]},
      {stage1_43[237]}
   );
   gpc1_1 gpc4064 (
      {stage0_43[470]},
      {stage1_43[238]}
   );
   gpc1_1 gpc4065 (
      {stage0_43[471]},
      {stage1_43[239]}
   );
   gpc1_1 gpc4066 (
      {stage0_43[472]},
      {stage1_43[240]}
   );
   gpc1_1 gpc4067 (
      {stage0_43[473]},
      {stage1_43[241]}
   );
   gpc1_1 gpc4068 (
      {stage0_43[474]},
      {stage1_43[242]}
   );
   gpc1_1 gpc4069 (
      {stage0_43[475]},
      {stage1_43[243]}
   );
   gpc1_1 gpc4070 (
      {stage0_43[476]},
      {stage1_43[244]}
   );
   gpc1_1 gpc4071 (
      {stage0_43[477]},
      {stage1_43[245]}
   );
   gpc1_1 gpc4072 (
      {stage0_43[478]},
      {stage1_43[246]}
   );
   gpc1_1 gpc4073 (
      {stage0_43[479]},
      {stage1_43[247]}
   );
   gpc1_1 gpc4074 (
      {stage0_43[480]},
      {stage1_43[248]}
   );
   gpc1_1 gpc4075 (
      {stage0_43[481]},
      {stage1_43[249]}
   );
   gpc1_1 gpc4076 (
      {stage0_43[482]},
      {stage1_43[250]}
   );
   gpc1_1 gpc4077 (
      {stage0_43[483]},
      {stage1_43[251]}
   );
   gpc1_1 gpc4078 (
      {stage0_43[484]},
      {stage1_43[252]}
   );
   gpc1_1 gpc4079 (
      {stage0_43[485]},
      {stage1_43[253]}
   );
   gpc1_1 gpc4080 (
      {stage0_44[424]},
      {stage1_44[194]}
   );
   gpc1_1 gpc4081 (
      {stage0_44[425]},
      {stage1_44[195]}
   );
   gpc1_1 gpc4082 (
      {stage0_44[426]},
      {stage1_44[196]}
   );
   gpc1_1 gpc4083 (
      {stage0_44[427]},
      {stage1_44[197]}
   );
   gpc1_1 gpc4084 (
      {stage0_44[428]},
      {stage1_44[198]}
   );
   gpc1_1 gpc4085 (
      {stage0_44[429]},
      {stage1_44[199]}
   );
   gpc1_1 gpc4086 (
      {stage0_44[430]},
      {stage1_44[200]}
   );
   gpc1_1 gpc4087 (
      {stage0_44[431]},
      {stage1_44[201]}
   );
   gpc1_1 gpc4088 (
      {stage0_44[432]},
      {stage1_44[202]}
   );
   gpc1_1 gpc4089 (
      {stage0_44[433]},
      {stage1_44[203]}
   );
   gpc1_1 gpc4090 (
      {stage0_44[434]},
      {stage1_44[204]}
   );
   gpc1_1 gpc4091 (
      {stage0_44[435]},
      {stage1_44[205]}
   );
   gpc1_1 gpc4092 (
      {stage0_44[436]},
      {stage1_44[206]}
   );
   gpc1_1 gpc4093 (
      {stage0_44[437]},
      {stage1_44[207]}
   );
   gpc1_1 gpc4094 (
      {stage0_44[438]},
      {stage1_44[208]}
   );
   gpc1_1 gpc4095 (
      {stage0_44[439]},
      {stage1_44[209]}
   );
   gpc1_1 gpc4096 (
      {stage0_44[440]},
      {stage1_44[210]}
   );
   gpc1_1 gpc4097 (
      {stage0_44[441]},
      {stage1_44[211]}
   );
   gpc1_1 gpc4098 (
      {stage0_44[442]},
      {stage1_44[212]}
   );
   gpc1_1 gpc4099 (
      {stage0_44[443]},
      {stage1_44[213]}
   );
   gpc1_1 gpc4100 (
      {stage0_44[444]},
      {stage1_44[214]}
   );
   gpc1_1 gpc4101 (
      {stage0_44[445]},
      {stage1_44[215]}
   );
   gpc1_1 gpc4102 (
      {stage0_44[446]},
      {stage1_44[216]}
   );
   gpc1_1 gpc4103 (
      {stage0_44[447]},
      {stage1_44[217]}
   );
   gpc1_1 gpc4104 (
      {stage0_44[448]},
      {stage1_44[218]}
   );
   gpc1_1 gpc4105 (
      {stage0_44[449]},
      {stage1_44[219]}
   );
   gpc1_1 gpc4106 (
      {stage0_44[450]},
      {stage1_44[220]}
   );
   gpc1_1 gpc4107 (
      {stage0_44[451]},
      {stage1_44[221]}
   );
   gpc1_1 gpc4108 (
      {stage0_44[452]},
      {stage1_44[222]}
   );
   gpc1_1 gpc4109 (
      {stage0_44[453]},
      {stage1_44[223]}
   );
   gpc1_1 gpc4110 (
      {stage0_44[454]},
      {stage1_44[224]}
   );
   gpc1_1 gpc4111 (
      {stage0_44[455]},
      {stage1_44[225]}
   );
   gpc1_1 gpc4112 (
      {stage0_44[456]},
      {stage1_44[226]}
   );
   gpc1_1 gpc4113 (
      {stage0_44[457]},
      {stage1_44[227]}
   );
   gpc1_1 gpc4114 (
      {stage0_44[458]},
      {stage1_44[228]}
   );
   gpc1_1 gpc4115 (
      {stage0_44[459]},
      {stage1_44[229]}
   );
   gpc1_1 gpc4116 (
      {stage0_44[460]},
      {stage1_44[230]}
   );
   gpc1_1 gpc4117 (
      {stage0_44[461]},
      {stage1_44[231]}
   );
   gpc1_1 gpc4118 (
      {stage0_44[462]},
      {stage1_44[232]}
   );
   gpc1_1 gpc4119 (
      {stage0_44[463]},
      {stage1_44[233]}
   );
   gpc1_1 gpc4120 (
      {stage0_44[464]},
      {stage1_44[234]}
   );
   gpc1_1 gpc4121 (
      {stage0_44[465]},
      {stage1_44[235]}
   );
   gpc1_1 gpc4122 (
      {stage0_44[466]},
      {stage1_44[236]}
   );
   gpc1_1 gpc4123 (
      {stage0_44[467]},
      {stage1_44[237]}
   );
   gpc1_1 gpc4124 (
      {stage0_44[468]},
      {stage1_44[238]}
   );
   gpc1_1 gpc4125 (
      {stage0_44[469]},
      {stage1_44[239]}
   );
   gpc1_1 gpc4126 (
      {stage0_44[470]},
      {stage1_44[240]}
   );
   gpc1_1 gpc4127 (
      {stage0_44[471]},
      {stage1_44[241]}
   );
   gpc1_1 gpc4128 (
      {stage0_44[472]},
      {stage1_44[242]}
   );
   gpc1_1 gpc4129 (
      {stage0_44[473]},
      {stage1_44[243]}
   );
   gpc1_1 gpc4130 (
      {stage0_44[474]},
      {stage1_44[244]}
   );
   gpc1_1 gpc4131 (
      {stage0_44[475]},
      {stage1_44[245]}
   );
   gpc1_1 gpc4132 (
      {stage0_44[476]},
      {stage1_44[246]}
   );
   gpc1_1 gpc4133 (
      {stage0_44[477]},
      {stage1_44[247]}
   );
   gpc1_1 gpc4134 (
      {stage0_44[478]},
      {stage1_44[248]}
   );
   gpc1_1 gpc4135 (
      {stage0_44[479]},
      {stage1_44[249]}
   );
   gpc1_1 gpc4136 (
      {stage0_44[480]},
      {stage1_44[250]}
   );
   gpc1_1 gpc4137 (
      {stage0_44[481]},
      {stage1_44[251]}
   );
   gpc1_1 gpc4138 (
      {stage0_44[482]},
      {stage1_44[252]}
   );
   gpc1_1 gpc4139 (
      {stage0_44[483]},
      {stage1_44[253]}
   );
   gpc1_1 gpc4140 (
      {stage0_44[484]},
      {stage1_44[254]}
   );
   gpc1_1 gpc4141 (
      {stage0_44[485]},
      {stage1_44[255]}
   );
   gpc1_1 gpc4142 (
      {stage0_45[433]},
      {stage1_45[159]}
   );
   gpc1_1 gpc4143 (
      {stage0_45[434]},
      {stage1_45[160]}
   );
   gpc1_1 gpc4144 (
      {stage0_45[435]},
      {stage1_45[161]}
   );
   gpc1_1 gpc4145 (
      {stage0_45[436]},
      {stage1_45[162]}
   );
   gpc1_1 gpc4146 (
      {stage0_45[437]},
      {stage1_45[163]}
   );
   gpc1_1 gpc4147 (
      {stage0_45[438]},
      {stage1_45[164]}
   );
   gpc1_1 gpc4148 (
      {stage0_45[439]},
      {stage1_45[165]}
   );
   gpc1_1 gpc4149 (
      {stage0_45[440]},
      {stage1_45[166]}
   );
   gpc1_1 gpc4150 (
      {stage0_45[441]},
      {stage1_45[167]}
   );
   gpc1_1 gpc4151 (
      {stage0_45[442]},
      {stage1_45[168]}
   );
   gpc1_1 gpc4152 (
      {stage0_45[443]},
      {stage1_45[169]}
   );
   gpc1_1 gpc4153 (
      {stage0_45[444]},
      {stage1_45[170]}
   );
   gpc1_1 gpc4154 (
      {stage0_45[445]},
      {stage1_45[171]}
   );
   gpc1_1 gpc4155 (
      {stage0_45[446]},
      {stage1_45[172]}
   );
   gpc1_1 gpc4156 (
      {stage0_45[447]},
      {stage1_45[173]}
   );
   gpc1_1 gpc4157 (
      {stage0_45[448]},
      {stage1_45[174]}
   );
   gpc1_1 gpc4158 (
      {stage0_45[449]},
      {stage1_45[175]}
   );
   gpc1_1 gpc4159 (
      {stage0_45[450]},
      {stage1_45[176]}
   );
   gpc1_1 gpc4160 (
      {stage0_45[451]},
      {stage1_45[177]}
   );
   gpc1_1 gpc4161 (
      {stage0_45[452]},
      {stage1_45[178]}
   );
   gpc1_1 gpc4162 (
      {stage0_45[453]},
      {stage1_45[179]}
   );
   gpc1_1 gpc4163 (
      {stage0_45[454]},
      {stage1_45[180]}
   );
   gpc1_1 gpc4164 (
      {stage0_45[455]},
      {stage1_45[181]}
   );
   gpc1_1 gpc4165 (
      {stage0_45[456]},
      {stage1_45[182]}
   );
   gpc1_1 gpc4166 (
      {stage0_45[457]},
      {stage1_45[183]}
   );
   gpc1_1 gpc4167 (
      {stage0_45[458]},
      {stage1_45[184]}
   );
   gpc1_1 gpc4168 (
      {stage0_45[459]},
      {stage1_45[185]}
   );
   gpc1_1 gpc4169 (
      {stage0_45[460]},
      {stage1_45[186]}
   );
   gpc1_1 gpc4170 (
      {stage0_45[461]},
      {stage1_45[187]}
   );
   gpc1_1 gpc4171 (
      {stage0_45[462]},
      {stage1_45[188]}
   );
   gpc1_1 gpc4172 (
      {stage0_45[463]},
      {stage1_45[189]}
   );
   gpc1_1 gpc4173 (
      {stage0_45[464]},
      {stage1_45[190]}
   );
   gpc1_1 gpc4174 (
      {stage0_45[465]},
      {stage1_45[191]}
   );
   gpc1_1 gpc4175 (
      {stage0_45[466]},
      {stage1_45[192]}
   );
   gpc1_1 gpc4176 (
      {stage0_45[467]},
      {stage1_45[193]}
   );
   gpc1_1 gpc4177 (
      {stage0_45[468]},
      {stage1_45[194]}
   );
   gpc1_1 gpc4178 (
      {stage0_45[469]},
      {stage1_45[195]}
   );
   gpc1_1 gpc4179 (
      {stage0_45[470]},
      {stage1_45[196]}
   );
   gpc1_1 gpc4180 (
      {stage0_45[471]},
      {stage1_45[197]}
   );
   gpc1_1 gpc4181 (
      {stage0_45[472]},
      {stage1_45[198]}
   );
   gpc1_1 gpc4182 (
      {stage0_45[473]},
      {stage1_45[199]}
   );
   gpc1_1 gpc4183 (
      {stage0_45[474]},
      {stage1_45[200]}
   );
   gpc1_1 gpc4184 (
      {stage0_45[475]},
      {stage1_45[201]}
   );
   gpc1_1 gpc4185 (
      {stage0_45[476]},
      {stage1_45[202]}
   );
   gpc1_1 gpc4186 (
      {stage0_45[477]},
      {stage1_45[203]}
   );
   gpc1_1 gpc4187 (
      {stage0_45[478]},
      {stage1_45[204]}
   );
   gpc1_1 gpc4188 (
      {stage0_45[479]},
      {stage1_45[205]}
   );
   gpc1_1 gpc4189 (
      {stage0_45[480]},
      {stage1_45[206]}
   );
   gpc1_1 gpc4190 (
      {stage0_45[481]},
      {stage1_45[207]}
   );
   gpc1_1 gpc4191 (
      {stage0_45[482]},
      {stage1_45[208]}
   );
   gpc1_1 gpc4192 (
      {stage0_45[483]},
      {stage1_45[209]}
   );
   gpc1_1 gpc4193 (
      {stage0_45[484]},
      {stage1_45[210]}
   );
   gpc1_1 gpc4194 (
      {stage0_45[485]},
      {stage1_45[211]}
   );
   gpc1_1 gpc4195 (
      {stage0_46[356]},
      {stage1_46[168]}
   );
   gpc1_1 gpc4196 (
      {stage0_46[357]},
      {stage1_46[169]}
   );
   gpc1_1 gpc4197 (
      {stage0_46[358]},
      {stage1_46[170]}
   );
   gpc1_1 gpc4198 (
      {stage0_46[359]},
      {stage1_46[171]}
   );
   gpc1_1 gpc4199 (
      {stage0_46[360]},
      {stage1_46[172]}
   );
   gpc1_1 gpc4200 (
      {stage0_46[361]},
      {stage1_46[173]}
   );
   gpc1_1 gpc4201 (
      {stage0_46[362]},
      {stage1_46[174]}
   );
   gpc1_1 gpc4202 (
      {stage0_46[363]},
      {stage1_46[175]}
   );
   gpc1_1 gpc4203 (
      {stage0_46[364]},
      {stage1_46[176]}
   );
   gpc1_1 gpc4204 (
      {stage0_46[365]},
      {stage1_46[177]}
   );
   gpc1_1 gpc4205 (
      {stage0_46[366]},
      {stage1_46[178]}
   );
   gpc1_1 gpc4206 (
      {stage0_46[367]},
      {stage1_46[179]}
   );
   gpc1_1 gpc4207 (
      {stage0_46[368]},
      {stage1_46[180]}
   );
   gpc1_1 gpc4208 (
      {stage0_46[369]},
      {stage1_46[181]}
   );
   gpc1_1 gpc4209 (
      {stage0_46[370]},
      {stage1_46[182]}
   );
   gpc1_1 gpc4210 (
      {stage0_46[371]},
      {stage1_46[183]}
   );
   gpc1_1 gpc4211 (
      {stage0_46[372]},
      {stage1_46[184]}
   );
   gpc1_1 gpc4212 (
      {stage0_46[373]},
      {stage1_46[185]}
   );
   gpc1_1 gpc4213 (
      {stage0_46[374]},
      {stage1_46[186]}
   );
   gpc1_1 gpc4214 (
      {stage0_46[375]},
      {stage1_46[187]}
   );
   gpc1_1 gpc4215 (
      {stage0_46[376]},
      {stage1_46[188]}
   );
   gpc1_1 gpc4216 (
      {stage0_46[377]},
      {stage1_46[189]}
   );
   gpc1_1 gpc4217 (
      {stage0_46[378]},
      {stage1_46[190]}
   );
   gpc1_1 gpc4218 (
      {stage0_46[379]},
      {stage1_46[191]}
   );
   gpc1_1 gpc4219 (
      {stage0_46[380]},
      {stage1_46[192]}
   );
   gpc1_1 gpc4220 (
      {stage0_46[381]},
      {stage1_46[193]}
   );
   gpc1_1 gpc4221 (
      {stage0_46[382]},
      {stage1_46[194]}
   );
   gpc1_1 gpc4222 (
      {stage0_46[383]},
      {stage1_46[195]}
   );
   gpc1_1 gpc4223 (
      {stage0_46[384]},
      {stage1_46[196]}
   );
   gpc1_1 gpc4224 (
      {stage0_46[385]},
      {stage1_46[197]}
   );
   gpc1_1 gpc4225 (
      {stage0_46[386]},
      {stage1_46[198]}
   );
   gpc1_1 gpc4226 (
      {stage0_46[387]},
      {stage1_46[199]}
   );
   gpc1_1 gpc4227 (
      {stage0_46[388]},
      {stage1_46[200]}
   );
   gpc1_1 gpc4228 (
      {stage0_46[389]},
      {stage1_46[201]}
   );
   gpc1_1 gpc4229 (
      {stage0_46[390]},
      {stage1_46[202]}
   );
   gpc1_1 gpc4230 (
      {stage0_46[391]},
      {stage1_46[203]}
   );
   gpc1_1 gpc4231 (
      {stage0_46[392]},
      {stage1_46[204]}
   );
   gpc1_1 gpc4232 (
      {stage0_46[393]},
      {stage1_46[205]}
   );
   gpc1_1 gpc4233 (
      {stage0_46[394]},
      {stage1_46[206]}
   );
   gpc1_1 gpc4234 (
      {stage0_46[395]},
      {stage1_46[207]}
   );
   gpc1_1 gpc4235 (
      {stage0_46[396]},
      {stage1_46[208]}
   );
   gpc1_1 gpc4236 (
      {stage0_46[397]},
      {stage1_46[209]}
   );
   gpc1_1 gpc4237 (
      {stage0_46[398]},
      {stage1_46[210]}
   );
   gpc1_1 gpc4238 (
      {stage0_46[399]},
      {stage1_46[211]}
   );
   gpc1_1 gpc4239 (
      {stage0_46[400]},
      {stage1_46[212]}
   );
   gpc1_1 gpc4240 (
      {stage0_46[401]},
      {stage1_46[213]}
   );
   gpc1_1 gpc4241 (
      {stage0_46[402]},
      {stage1_46[214]}
   );
   gpc1_1 gpc4242 (
      {stage0_46[403]},
      {stage1_46[215]}
   );
   gpc1_1 gpc4243 (
      {stage0_46[404]},
      {stage1_46[216]}
   );
   gpc1_1 gpc4244 (
      {stage0_46[405]},
      {stage1_46[217]}
   );
   gpc1_1 gpc4245 (
      {stage0_46[406]},
      {stage1_46[218]}
   );
   gpc1_1 gpc4246 (
      {stage0_46[407]},
      {stage1_46[219]}
   );
   gpc1_1 gpc4247 (
      {stage0_46[408]},
      {stage1_46[220]}
   );
   gpc1_1 gpc4248 (
      {stage0_46[409]},
      {stage1_46[221]}
   );
   gpc1_1 gpc4249 (
      {stage0_46[410]},
      {stage1_46[222]}
   );
   gpc1_1 gpc4250 (
      {stage0_46[411]},
      {stage1_46[223]}
   );
   gpc1_1 gpc4251 (
      {stage0_46[412]},
      {stage1_46[224]}
   );
   gpc1_1 gpc4252 (
      {stage0_46[413]},
      {stage1_46[225]}
   );
   gpc1_1 gpc4253 (
      {stage0_46[414]},
      {stage1_46[226]}
   );
   gpc1_1 gpc4254 (
      {stage0_46[415]},
      {stage1_46[227]}
   );
   gpc1_1 gpc4255 (
      {stage0_46[416]},
      {stage1_46[228]}
   );
   gpc1_1 gpc4256 (
      {stage0_46[417]},
      {stage1_46[229]}
   );
   gpc1_1 gpc4257 (
      {stage0_46[418]},
      {stage1_46[230]}
   );
   gpc1_1 gpc4258 (
      {stage0_46[419]},
      {stage1_46[231]}
   );
   gpc1_1 gpc4259 (
      {stage0_46[420]},
      {stage1_46[232]}
   );
   gpc1_1 gpc4260 (
      {stage0_46[421]},
      {stage1_46[233]}
   );
   gpc1_1 gpc4261 (
      {stage0_46[422]},
      {stage1_46[234]}
   );
   gpc1_1 gpc4262 (
      {stage0_46[423]},
      {stage1_46[235]}
   );
   gpc1_1 gpc4263 (
      {stage0_46[424]},
      {stage1_46[236]}
   );
   gpc1_1 gpc4264 (
      {stage0_46[425]},
      {stage1_46[237]}
   );
   gpc1_1 gpc4265 (
      {stage0_46[426]},
      {stage1_46[238]}
   );
   gpc1_1 gpc4266 (
      {stage0_46[427]},
      {stage1_46[239]}
   );
   gpc1_1 gpc4267 (
      {stage0_46[428]},
      {stage1_46[240]}
   );
   gpc1_1 gpc4268 (
      {stage0_46[429]},
      {stage1_46[241]}
   );
   gpc1_1 gpc4269 (
      {stage0_46[430]},
      {stage1_46[242]}
   );
   gpc1_1 gpc4270 (
      {stage0_46[431]},
      {stage1_46[243]}
   );
   gpc1_1 gpc4271 (
      {stage0_46[432]},
      {stage1_46[244]}
   );
   gpc1_1 gpc4272 (
      {stage0_46[433]},
      {stage1_46[245]}
   );
   gpc1_1 gpc4273 (
      {stage0_46[434]},
      {stage1_46[246]}
   );
   gpc1_1 gpc4274 (
      {stage0_46[435]},
      {stage1_46[247]}
   );
   gpc1_1 gpc4275 (
      {stage0_46[436]},
      {stage1_46[248]}
   );
   gpc1_1 gpc4276 (
      {stage0_46[437]},
      {stage1_46[249]}
   );
   gpc1_1 gpc4277 (
      {stage0_46[438]},
      {stage1_46[250]}
   );
   gpc1_1 gpc4278 (
      {stage0_46[439]},
      {stage1_46[251]}
   );
   gpc1_1 gpc4279 (
      {stage0_46[440]},
      {stage1_46[252]}
   );
   gpc1_1 gpc4280 (
      {stage0_46[441]},
      {stage1_46[253]}
   );
   gpc1_1 gpc4281 (
      {stage0_46[442]},
      {stage1_46[254]}
   );
   gpc1_1 gpc4282 (
      {stage0_46[443]},
      {stage1_46[255]}
   );
   gpc1_1 gpc4283 (
      {stage0_46[444]},
      {stage1_46[256]}
   );
   gpc1_1 gpc4284 (
      {stage0_46[445]},
      {stage1_46[257]}
   );
   gpc1_1 gpc4285 (
      {stage0_46[446]},
      {stage1_46[258]}
   );
   gpc1_1 gpc4286 (
      {stage0_46[447]},
      {stage1_46[259]}
   );
   gpc1_1 gpc4287 (
      {stage0_46[448]},
      {stage1_46[260]}
   );
   gpc1_1 gpc4288 (
      {stage0_46[449]},
      {stage1_46[261]}
   );
   gpc1_1 gpc4289 (
      {stage0_46[450]},
      {stage1_46[262]}
   );
   gpc1_1 gpc4290 (
      {stage0_46[451]},
      {stage1_46[263]}
   );
   gpc1_1 gpc4291 (
      {stage0_46[452]},
      {stage1_46[264]}
   );
   gpc1_1 gpc4292 (
      {stage0_46[453]},
      {stage1_46[265]}
   );
   gpc1_1 gpc4293 (
      {stage0_46[454]},
      {stage1_46[266]}
   );
   gpc1_1 gpc4294 (
      {stage0_46[455]},
      {stage1_46[267]}
   );
   gpc1_1 gpc4295 (
      {stage0_46[456]},
      {stage1_46[268]}
   );
   gpc1_1 gpc4296 (
      {stage0_46[457]},
      {stage1_46[269]}
   );
   gpc1_1 gpc4297 (
      {stage0_46[458]},
      {stage1_46[270]}
   );
   gpc1_1 gpc4298 (
      {stage0_46[459]},
      {stage1_46[271]}
   );
   gpc1_1 gpc4299 (
      {stage0_46[460]},
      {stage1_46[272]}
   );
   gpc1_1 gpc4300 (
      {stage0_46[461]},
      {stage1_46[273]}
   );
   gpc1_1 gpc4301 (
      {stage0_46[462]},
      {stage1_46[274]}
   );
   gpc1_1 gpc4302 (
      {stage0_46[463]},
      {stage1_46[275]}
   );
   gpc1_1 gpc4303 (
      {stage0_46[464]},
      {stage1_46[276]}
   );
   gpc1_1 gpc4304 (
      {stage0_46[465]},
      {stage1_46[277]}
   );
   gpc1_1 gpc4305 (
      {stage0_46[466]},
      {stage1_46[278]}
   );
   gpc1_1 gpc4306 (
      {stage0_46[467]},
      {stage1_46[279]}
   );
   gpc1_1 gpc4307 (
      {stage0_46[468]},
      {stage1_46[280]}
   );
   gpc1_1 gpc4308 (
      {stage0_46[469]},
      {stage1_46[281]}
   );
   gpc1_1 gpc4309 (
      {stage0_46[470]},
      {stage1_46[282]}
   );
   gpc1_1 gpc4310 (
      {stage0_46[471]},
      {stage1_46[283]}
   );
   gpc1_1 gpc4311 (
      {stage0_46[472]},
      {stage1_46[284]}
   );
   gpc1_1 gpc4312 (
      {stage0_46[473]},
      {stage1_46[285]}
   );
   gpc1_1 gpc4313 (
      {stage0_46[474]},
      {stage1_46[286]}
   );
   gpc1_1 gpc4314 (
      {stage0_46[475]},
      {stage1_46[287]}
   );
   gpc1_1 gpc4315 (
      {stage0_46[476]},
      {stage1_46[288]}
   );
   gpc1_1 gpc4316 (
      {stage0_46[477]},
      {stage1_46[289]}
   );
   gpc1_1 gpc4317 (
      {stage0_46[478]},
      {stage1_46[290]}
   );
   gpc1_1 gpc4318 (
      {stage0_46[479]},
      {stage1_46[291]}
   );
   gpc1_1 gpc4319 (
      {stage0_46[480]},
      {stage1_46[292]}
   );
   gpc1_1 gpc4320 (
      {stage0_46[481]},
      {stage1_46[293]}
   );
   gpc1_1 gpc4321 (
      {stage0_46[482]},
      {stage1_46[294]}
   );
   gpc1_1 gpc4322 (
      {stage0_46[483]},
      {stage1_46[295]}
   );
   gpc1_1 gpc4323 (
      {stage0_46[484]},
      {stage1_46[296]}
   );
   gpc1_1 gpc4324 (
      {stage0_46[485]},
      {stage1_46[297]}
   );
   gpc1_1 gpc4325 (
      {stage0_47[443]},
      {stage1_47[193]}
   );
   gpc1_1 gpc4326 (
      {stage0_47[444]},
      {stage1_47[194]}
   );
   gpc1_1 gpc4327 (
      {stage0_47[445]},
      {stage1_47[195]}
   );
   gpc1_1 gpc4328 (
      {stage0_47[446]},
      {stage1_47[196]}
   );
   gpc1_1 gpc4329 (
      {stage0_47[447]},
      {stage1_47[197]}
   );
   gpc1_1 gpc4330 (
      {stage0_47[448]},
      {stage1_47[198]}
   );
   gpc1_1 gpc4331 (
      {stage0_47[449]},
      {stage1_47[199]}
   );
   gpc1_1 gpc4332 (
      {stage0_47[450]},
      {stage1_47[200]}
   );
   gpc1_1 gpc4333 (
      {stage0_47[451]},
      {stage1_47[201]}
   );
   gpc1_1 gpc4334 (
      {stage0_47[452]},
      {stage1_47[202]}
   );
   gpc1_1 gpc4335 (
      {stage0_47[453]},
      {stage1_47[203]}
   );
   gpc1_1 gpc4336 (
      {stage0_47[454]},
      {stage1_47[204]}
   );
   gpc1_1 gpc4337 (
      {stage0_47[455]},
      {stage1_47[205]}
   );
   gpc1_1 gpc4338 (
      {stage0_47[456]},
      {stage1_47[206]}
   );
   gpc1_1 gpc4339 (
      {stage0_47[457]},
      {stage1_47[207]}
   );
   gpc1_1 gpc4340 (
      {stage0_47[458]},
      {stage1_47[208]}
   );
   gpc1_1 gpc4341 (
      {stage0_47[459]},
      {stage1_47[209]}
   );
   gpc1_1 gpc4342 (
      {stage0_47[460]},
      {stage1_47[210]}
   );
   gpc1_1 gpc4343 (
      {stage0_47[461]},
      {stage1_47[211]}
   );
   gpc1_1 gpc4344 (
      {stage0_47[462]},
      {stage1_47[212]}
   );
   gpc1_1 gpc4345 (
      {stage0_47[463]},
      {stage1_47[213]}
   );
   gpc1_1 gpc4346 (
      {stage0_47[464]},
      {stage1_47[214]}
   );
   gpc1_1 gpc4347 (
      {stage0_47[465]},
      {stage1_47[215]}
   );
   gpc1_1 gpc4348 (
      {stage0_47[466]},
      {stage1_47[216]}
   );
   gpc1_1 gpc4349 (
      {stage0_47[467]},
      {stage1_47[217]}
   );
   gpc1_1 gpc4350 (
      {stage0_47[468]},
      {stage1_47[218]}
   );
   gpc1_1 gpc4351 (
      {stage0_47[469]},
      {stage1_47[219]}
   );
   gpc1_1 gpc4352 (
      {stage0_47[470]},
      {stage1_47[220]}
   );
   gpc1_1 gpc4353 (
      {stage0_47[471]},
      {stage1_47[221]}
   );
   gpc1_1 gpc4354 (
      {stage0_47[472]},
      {stage1_47[222]}
   );
   gpc1_1 gpc4355 (
      {stage0_47[473]},
      {stage1_47[223]}
   );
   gpc1_1 gpc4356 (
      {stage0_47[474]},
      {stage1_47[224]}
   );
   gpc1_1 gpc4357 (
      {stage0_47[475]},
      {stage1_47[225]}
   );
   gpc1_1 gpc4358 (
      {stage0_47[476]},
      {stage1_47[226]}
   );
   gpc1_1 gpc4359 (
      {stage0_47[477]},
      {stage1_47[227]}
   );
   gpc1_1 gpc4360 (
      {stage0_47[478]},
      {stage1_47[228]}
   );
   gpc1_1 gpc4361 (
      {stage0_47[479]},
      {stage1_47[229]}
   );
   gpc1_1 gpc4362 (
      {stage0_47[480]},
      {stage1_47[230]}
   );
   gpc1_1 gpc4363 (
      {stage0_47[481]},
      {stage1_47[231]}
   );
   gpc1_1 gpc4364 (
      {stage0_47[482]},
      {stage1_47[232]}
   );
   gpc1_1 gpc4365 (
      {stage0_47[483]},
      {stage1_47[233]}
   );
   gpc1_1 gpc4366 (
      {stage0_47[484]},
      {stage1_47[234]}
   );
   gpc1_1 gpc4367 (
      {stage0_47[485]},
      {stage1_47[235]}
   );
   gpc1_1 gpc4368 (
      {stage0_48[478]},
      {stage1_48[190]}
   );
   gpc1_1 gpc4369 (
      {stage0_48[479]},
      {stage1_48[191]}
   );
   gpc1_1 gpc4370 (
      {stage0_48[480]},
      {stage1_48[192]}
   );
   gpc1_1 gpc4371 (
      {stage0_48[481]},
      {stage1_48[193]}
   );
   gpc1_1 gpc4372 (
      {stage0_48[482]},
      {stage1_48[194]}
   );
   gpc1_1 gpc4373 (
      {stage0_48[483]},
      {stage1_48[195]}
   );
   gpc1_1 gpc4374 (
      {stage0_48[484]},
      {stage1_48[196]}
   );
   gpc1_1 gpc4375 (
      {stage0_48[485]},
      {stage1_48[197]}
   );
   gpc1_1 gpc4376 (
      {stage0_50[481]},
      {stage1_50[185]}
   );
   gpc1_1 gpc4377 (
      {stage0_50[482]},
      {stage1_50[186]}
   );
   gpc1_1 gpc4378 (
      {stage0_50[483]},
      {stage1_50[187]}
   );
   gpc1_1 gpc4379 (
      {stage0_50[484]},
      {stage1_50[188]}
   );
   gpc1_1 gpc4380 (
      {stage0_50[485]},
      {stage1_50[189]}
   );
   gpc1_1 gpc4381 (
      {stage0_51[435]},
      {stage1_51[224]}
   );
   gpc1_1 gpc4382 (
      {stage0_51[436]},
      {stage1_51[225]}
   );
   gpc1_1 gpc4383 (
      {stage0_51[437]},
      {stage1_51[226]}
   );
   gpc1_1 gpc4384 (
      {stage0_51[438]},
      {stage1_51[227]}
   );
   gpc1_1 gpc4385 (
      {stage0_51[439]},
      {stage1_51[228]}
   );
   gpc1_1 gpc4386 (
      {stage0_51[440]},
      {stage1_51[229]}
   );
   gpc1_1 gpc4387 (
      {stage0_51[441]},
      {stage1_51[230]}
   );
   gpc1_1 gpc4388 (
      {stage0_51[442]},
      {stage1_51[231]}
   );
   gpc1_1 gpc4389 (
      {stage0_51[443]},
      {stage1_51[232]}
   );
   gpc1_1 gpc4390 (
      {stage0_51[444]},
      {stage1_51[233]}
   );
   gpc1_1 gpc4391 (
      {stage0_51[445]},
      {stage1_51[234]}
   );
   gpc1_1 gpc4392 (
      {stage0_51[446]},
      {stage1_51[235]}
   );
   gpc1_1 gpc4393 (
      {stage0_51[447]},
      {stage1_51[236]}
   );
   gpc1_1 gpc4394 (
      {stage0_51[448]},
      {stage1_51[237]}
   );
   gpc1_1 gpc4395 (
      {stage0_51[449]},
      {stage1_51[238]}
   );
   gpc1_1 gpc4396 (
      {stage0_51[450]},
      {stage1_51[239]}
   );
   gpc1_1 gpc4397 (
      {stage0_51[451]},
      {stage1_51[240]}
   );
   gpc1_1 gpc4398 (
      {stage0_51[452]},
      {stage1_51[241]}
   );
   gpc1_1 gpc4399 (
      {stage0_51[453]},
      {stage1_51[242]}
   );
   gpc1_1 gpc4400 (
      {stage0_51[454]},
      {stage1_51[243]}
   );
   gpc1_1 gpc4401 (
      {stage0_51[455]},
      {stage1_51[244]}
   );
   gpc1_1 gpc4402 (
      {stage0_51[456]},
      {stage1_51[245]}
   );
   gpc1_1 gpc4403 (
      {stage0_51[457]},
      {stage1_51[246]}
   );
   gpc1_1 gpc4404 (
      {stage0_51[458]},
      {stage1_51[247]}
   );
   gpc1_1 gpc4405 (
      {stage0_51[459]},
      {stage1_51[248]}
   );
   gpc1_1 gpc4406 (
      {stage0_51[460]},
      {stage1_51[249]}
   );
   gpc1_1 gpc4407 (
      {stage0_51[461]},
      {stage1_51[250]}
   );
   gpc1_1 gpc4408 (
      {stage0_51[462]},
      {stage1_51[251]}
   );
   gpc1_1 gpc4409 (
      {stage0_51[463]},
      {stage1_51[252]}
   );
   gpc1_1 gpc4410 (
      {stage0_51[464]},
      {stage1_51[253]}
   );
   gpc1_1 gpc4411 (
      {stage0_51[465]},
      {stage1_51[254]}
   );
   gpc1_1 gpc4412 (
      {stage0_51[466]},
      {stage1_51[255]}
   );
   gpc1_1 gpc4413 (
      {stage0_51[467]},
      {stage1_51[256]}
   );
   gpc1_1 gpc4414 (
      {stage0_51[468]},
      {stage1_51[257]}
   );
   gpc1_1 gpc4415 (
      {stage0_51[469]},
      {stage1_51[258]}
   );
   gpc1_1 gpc4416 (
      {stage0_51[470]},
      {stage1_51[259]}
   );
   gpc1_1 gpc4417 (
      {stage0_51[471]},
      {stage1_51[260]}
   );
   gpc1_1 gpc4418 (
      {stage0_51[472]},
      {stage1_51[261]}
   );
   gpc1_1 gpc4419 (
      {stage0_51[473]},
      {stage1_51[262]}
   );
   gpc1_1 gpc4420 (
      {stage0_51[474]},
      {stage1_51[263]}
   );
   gpc1_1 gpc4421 (
      {stage0_51[475]},
      {stage1_51[264]}
   );
   gpc1_1 gpc4422 (
      {stage0_51[476]},
      {stage1_51[265]}
   );
   gpc1_1 gpc4423 (
      {stage0_51[477]},
      {stage1_51[266]}
   );
   gpc1_1 gpc4424 (
      {stage0_51[478]},
      {stage1_51[267]}
   );
   gpc1_1 gpc4425 (
      {stage0_51[479]},
      {stage1_51[268]}
   );
   gpc1_1 gpc4426 (
      {stage0_51[480]},
      {stage1_51[269]}
   );
   gpc1_1 gpc4427 (
      {stage0_51[481]},
      {stage1_51[270]}
   );
   gpc1_1 gpc4428 (
      {stage0_51[482]},
      {stage1_51[271]}
   );
   gpc1_1 gpc4429 (
      {stage0_51[483]},
      {stage1_51[272]}
   );
   gpc1_1 gpc4430 (
      {stage0_51[484]},
      {stage1_51[273]}
   );
   gpc1_1 gpc4431 (
      {stage0_51[485]},
      {stage1_51[274]}
   );
   gpc1_1 gpc4432 (
      {stage0_54[453]},
      {stage1_54[198]}
   );
   gpc1_1 gpc4433 (
      {stage0_54[454]},
      {stage1_54[199]}
   );
   gpc1_1 gpc4434 (
      {stage0_54[455]},
      {stage1_54[200]}
   );
   gpc1_1 gpc4435 (
      {stage0_54[456]},
      {stage1_54[201]}
   );
   gpc1_1 gpc4436 (
      {stage0_54[457]},
      {stage1_54[202]}
   );
   gpc1_1 gpc4437 (
      {stage0_54[458]},
      {stage1_54[203]}
   );
   gpc1_1 gpc4438 (
      {stage0_54[459]},
      {stage1_54[204]}
   );
   gpc1_1 gpc4439 (
      {stage0_54[460]},
      {stage1_54[205]}
   );
   gpc1_1 gpc4440 (
      {stage0_54[461]},
      {stage1_54[206]}
   );
   gpc1_1 gpc4441 (
      {stage0_54[462]},
      {stage1_54[207]}
   );
   gpc1_1 gpc4442 (
      {stage0_54[463]},
      {stage1_54[208]}
   );
   gpc1_1 gpc4443 (
      {stage0_54[464]},
      {stage1_54[209]}
   );
   gpc1_1 gpc4444 (
      {stage0_54[465]},
      {stage1_54[210]}
   );
   gpc1_1 gpc4445 (
      {stage0_54[466]},
      {stage1_54[211]}
   );
   gpc1_1 gpc4446 (
      {stage0_54[467]},
      {stage1_54[212]}
   );
   gpc1_1 gpc4447 (
      {stage0_54[468]},
      {stage1_54[213]}
   );
   gpc1_1 gpc4448 (
      {stage0_54[469]},
      {stage1_54[214]}
   );
   gpc1_1 gpc4449 (
      {stage0_54[470]},
      {stage1_54[215]}
   );
   gpc1_1 gpc4450 (
      {stage0_54[471]},
      {stage1_54[216]}
   );
   gpc1_1 gpc4451 (
      {stage0_54[472]},
      {stage1_54[217]}
   );
   gpc1_1 gpc4452 (
      {stage0_54[473]},
      {stage1_54[218]}
   );
   gpc1_1 gpc4453 (
      {stage0_54[474]},
      {stage1_54[219]}
   );
   gpc1_1 gpc4454 (
      {stage0_54[475]},
      {stage1_54[220]}
   );
   gpc1_1 gpc4455 (
      {stage0_54[476]},
      {stage1_54[221]}
   );
   gpc1_1 gpc4456 (
      {stage0_54[477]},
      {stage1_54[222]}
   );
   gpc1_1 gpc4457 (
      {stage0_54[478]},
      {stage1_54[223]}
   );
   gpc1_1 gpc4458 (
      {stage0_54[479]},
      {stage1_54[224]}
   );
   gpc1_1 gpc4459 (
      {stage0_54[480]},
      {stage1_54[225]}
   );
   gpc1_1 gpc4460 (
      {stage0_54[481]},
      {stage1_54[226]}
   );
   gpc1_1 gpc4461 (
      {stage0_54[482]},
      {stage1_54[227]}
   );
   gpc1_1 gpc4462 (
      {stage0_54[483]},
      {stage1_54[228]}
   );
   gpc1_1 gpc4463 (
      {stage0_54[484]},
      {stage1_54[229]}
   );
   gpc1_1 gpc4464 (
      {stage0_54[485]},
      {stage1_54[230]}
   );
   gpc1_1 gpc4465 (
      {stage0_55[425]},
      {stage1_55[206]}
   );
   gpc1_1 gpc4466 (
      {stage0_55[426]},
      {stage1_55[207]}
   );
   gpc1_1 gpc4467 (
      {stage0_55[427]},
      {stage1_55[208]}
   );
   gpc1_1 gpc4468 (
      {stage0_55[428]},
      {stage1_55[209]}
   );
   gpc1_1 gpc4469 (
      {stage0_55[429]},
      {stage1_55[210]}
   );
   gpc1_1 gpc4470 (
      {stage0_55[430]},
      {stage1_55[211]}
   );
   gpc1_1 gpc4471 (
      {stage0_55[431]},
      {stage1_55[212]}
   );
   gpc1_1 gpc4472 (
      {stage0_55[432]},
      {stage1_55[213]}
   );
   gpc1_1 gpc4473 (
      {stage0_55[433]},
      {stage1_55[214]}
   );
   gpc1_1 gpc4474 (
      {stage0_55[434]},
      {stage1_55[215]}
   );
   gpc1_1 gpc4475 (
      {stage0_55[435]},
      {stage1_55[216]}
   );
   gpc1_1 gpc4476 (
      {stage0_55[436]},
      {stage1_55[217]}
   );
   gpc1_1 gpc4477 (
      {stage0_55[437]},
      {stage1_55[218]}
   );
   gpc1_1 gpc4478 (
      {stage0_55[438]},
      {stage1_55[219]}
   );
   gpc1_1 gpc4479 (
      {stage0_55[439]},
      {stage1_55[220]}
   );
   gpc1_1 gpc4480 (
      {stage0_55[440]},
      {stage1_55[221]}
   );
   gpc1_1 gpc4481 (
      {stage0_55[441]},
      {stage1_55[222]}
   );
   gpc1_1 gpc4482 (
      {stage0_55[442]},
      {stage1_55[223]}
   );
   gpc1_1 gpc4483 (
      {stage0_55[443]},
      {stage1_55[224]}
   );
   gpc1_1 gpc4484 (
      {stage0_55[444]},
      {stage1_55[225]}
   );
   gpc1_1 gpc4485 (
      {stage0_55[445]},
      {stage1_55[226]}
   );
   gpc1_1 gpc4486 (
      {stage0_55[446]},
      {stage1_55[227]}
   );
   gpc1_1 gpc4487 (
      {stage0_55[447]},
      {stage1_55[228]}
   );
   gpc1_1 gpc4488 (
      {stage0_55[448]},
      {stage1_55[229]}
   );
   gpc1_1 gpc4489 (
      {stage0_55[449]},
      {stage1_55[230]}
   );
   gpc1_1 gpc4490 (
      {stage0_55[450]},
      {stage1_55[231]}
   );
   gpc1_1 gpc4491 (
      {stage0_55[451]},
      {stage1_55[232]}
   );
   gpc1_1 gpc4492 (
      {stage0_55[452]},
      {stage1_55[233]}
   );
   gpc1_1 gpc4493 (
      {stage0_55[453]},
      {stage1_55[234]}
   );
   gpc1_1 gpc4494 (
      {stage0_55[454]},
      {stage1_55[235]}
   );
   gpc1_1 gpc4495 (
      {stage0_55[455]},
      {stage1_55[236]}
   );
   gpc1_1 gpc4496 (
      {stage0_55[456]},
      {stage1_55[237]}
   );
   gpc1_1 gpc4497 (
      {stage0_55[457]},
      {stage1_55[238]}
   );
   gpc1_1 gpc4498 (
      {stage0_55[458]},
      {stage1_55[239]}
   );
   gpc1_1 gpc4499 (
      {stage0_55[459]},
      {stage1_55[240]}
   );
   gpc1_1 gpc4500 (
      {stage0_55[460]},
      {stage1_55[241]}
   );
   gpc1_1 gpc4501 (
      {stage0_55[461]},
      {stage1_55[242]}
   );
   gpc1_1 gpc4502 (
      {stage0_55[462]},
      {stage1_55[243]}
   );
   gpc1_1 gpc4503 (
      {stage0_55[463]},
      {stage1_55[244]}
   );
   gpc1_1 gpc4504 (
      {stage0_55[464]},
      {stage1_55[245]}
   );
   gpc1_1 gpc4505 (
      {stage0_55[465]},
      {stage1_55[246]}
   );
   gpc1_1 gpc4506 (
      {stage0_55[466]},
      {stage1_55[247]}
   );
   gpc1_1 gpc4507 (
      {stage0_55[467]},
      {stage1_55[248]}
   );
   gpc1_1 gpc4508 (
      {stage0_55[468]},
      {stage1_55[249]}
   );
   gpc1_1 gpc4509 (
      {stage0_55[469]},
      {stage1_55[250]}
   );
   gpc1_1 gpc4510 (
      {stage0_55[470]},
      {stage1_55[251]}
   );
   gpc1_1 gpc4511 (
      {stage0_55[471]},
      {stage1_55[252]}
   );
   gpc1_1 gpc4512 (
      {stage0_55[472]},
      {stage1_55[253]}
   );
   gpc1_1 gpc4513 (
      {stage0_55[473]},
      {stage1_55[254]}
   );
   gpc1_1 gpc4514 (
      {stage0_55[474]},
      {stage1_55[255]}
   );
   gpc1_1 gpc4515 (
      {stage0_55[475]},
      {stage1_55[256]}
   );
   gpc1_1 gpc4516 (
      {stage0_55[476]},
      {stage1_55[257]}
   );
   gpc1_1 gpc4517 (
      {stage0_55[477]},
      {stage1_55[258]}
   );
   gpc1_1 gpc4518 (
      {stage0_55[478]},
      {stage1_55[259]}
   );
   gpc1_1 gpc4519 (
      {stage0_55[479]},
      {stage1_55[260]}
   );
   gpc1_1 gpc4520 (
      {stage0_55[480]},
      {stage1_55[261]}
   );
   gpc1_1 gpc4521 (
      {stage0_55[481]},
      {stage1_55[262]}
   );
   gpc1_1 gpc4522 (
      {stage0_55[482]},
      {stage1_55[263]}
   );
   gpc1_1 gpc4523 (
      {stage0_55[483]},
      {stage1_55[264]}
   );
   gpc1_1 gpc4524 (
      {stage0_55[484]},
      {stage1_55[265]}
   );
   gpc1_1 gpc4525 (
      {stage0_55[485]},
      {stage1_55[266]}
   );
   gpc1_1 gpc4526 (
      {stage0_58[460]},
      {stage1_58[194]}
   );
   gpc1_1 gpc4527 (
      {stage0_58[461]},
      {stage1_58[195]}
   );
   gpc1_1 gpc4528 (
      {stage0_58[462]},
      {stage1_58[196]}
   );
   gpc1_1 gpc4529 (
      {stage0_58[463]},
      {stage1_58[197]}
   );
   gpc1_1 gpc4530 (
      {stage0_58[464]},
      {stage1_58[198]}
   );
   gpc1_1 gpc4531 (
      {stage0_58[465]},
      {stage1_58[199]}
   );
   gpc1_1 gpc4532 (
      {stage0_58[466]},
      {stage1_58[200]}
   );
   gpc1_1 gpc4533 (
      {stage0_58[467]},
      {stage1_58[201]}
   );
   gpc1_1 gpc4534 (
      {stage0_58[468]},
      {stage1_58[202]}
   );
   gpc1_1 gpc4535 (
      {stage0_58[469]},
      {stage1_58[203]}
   );
   gpc1_1 gpc4536 (
      {stage0_58[470]},
      {stage1_58[204]}
   );
   gpc1_1 gpc4537 (
      {stage0_58[471]},
      {stage1_58[205]}
   );
   gpc1_1 gpc4538 (
      {stage0_58[472]},
      {stage1_58[206]}
   );
   gpc1_1 gpc4539 (
      {stage0_58[473]},
      {stage1_58[207]}
   );
   gpc1_1 gpc4540 (
      {stage0_58[474]},
      {stage1_58[208]}
   );
   gpc1_1 gpc4541 (
      {stage0_58[475]},
      {stage1_58[209]}
   );
   gpc1_1 gpc4542 (
      {stage0_58[476]},
      {stage1_58[210]}
   );
   gpc1_1 gpc4543 (
      {stage0_58[477]},
      {stage1_58[211]}
   );
   gpc1_1 gpc4544 (
      {stage0_58[478]},
      {stage1_58[212]}
   );
   gpc1_1 gpc4545 (
      {stage0_58[479]},
      {stage1_58[213]}
   );
   gpc1_1 gpc4546 (
      {stage0_58[480]},
      {stage1_58[214]}
   );
   gpc1_1 gpc4547 (
      {stage0_58[481]},
      {stage1_58[215]}
   );
   gpc1_1 gpc4548 (
      {stage0_58[482]},
      {stage1_58[216]}
   );
   gpc1_1 gpc4549 (
      {stage0_58[483]},
      {stage1_58[217]}
   );
   gpc1_1 gpc4550 (
      {stage0_58[484]},
      {stage1_58[218]}
   );
   gpc1_1 gpc4551 (
      {stage0_58[485]},
      {stage1_58[219]}
   );
   gpc1_1 gpc4552 (
      {stage0_59[469]},
      {stage1_59[189]}
   );
   gpc1_1 gpc4553 (
      {stage0_59[470]},
      {stage1_59[190]}
   );
   gpc1_1 gpc4554 (
      {stage0_59[471]},
      {stage1_59[191]}
   );
   gpc1_1 gpc4555 (
      {stage0_59[472]},
      {stage1_59[192]}
   );
   gpc1_1 gpc4556 (
      {stage0_59[473]},
      {stage1_59[193]}
   );
   gpc1_1 gpc4557 (
      {stage0_59[474]},
      {stage1_59[194]}
   );
   gpc1_1 gpc4558 (
      {stage0_59[475]},
      {stage1_59[195]}
   );
   gpc1_1 gpc4559 (
      {stage0_59[476]},
      {stage1_59[196]}
   );
   gpc1_1 gpc4560 (
      {stage0_59[477]},
      {stage1_59[197]}
   );
   gpc1_1 gpc4561 (
      {stage0_59[478]},
      {stage1_59[198]}
   );
   gpc1_1 gpc4562 (
      {stage0_59[479]},
      {stage1_59[199]}
   );
   gpc1_1 gpc4563 (
      {stage0_59[480]},
      {stage1_59[200]}
   );
   gpc1_1 gpc4564 (
      {stage0_59[481]},
      {stage1_59[201]}
   );
   gpc1_1 gpc4565 (
      {stage0_59[482]},
      {stage1_59[202]}
   );
   gpc1_1 gpc4566 (
      {stage0_59[483]},
      {stage1_59[203]}
   );
   gpc1_1 gpc4567 (
      {stage0_59[484]},
      {stage1_59[204]}
   );
   gpc1_1 gpc4568 (
      {stage0_59[485]},
      {stage1_59[205]}
   );
   gpc1_1 gpc4569 (
      {stage0_62[474]},
      {stage1_62[181]}
   );
   gpc1_1 gpc4570 (
      {stage0_62[475]},
      {stage1_62[182]}
   );
   gpc1_1 gpc4571 (
      {stage0_62[476]},
      {stage1_62[183]}
   );
   gpc1_1 gpc4572 (
      {stage0_62[477]},
      {stage1_62[184]}
   );
   gpc1_1 gpc4573 (
      {stage0_62[478]},
      {stage1_62[185]}
   );
   gpc1_1 gpc4574 (
      {stage0_62[479]},
      {stage1_62[186]}
   );
   gpc1_1 gpc4575 (
      {stage0_62[480]},
      {stage1_62[187]}
   );
   gpc1_1 gpc4576 (
      {stage0_62[481]},
      {stage1_62[188]}
   );
   gpc1_1 gpc4577 (
      {stage0_62[482]},
      {stage1_62[189]}
   );
   gpc1_1 gpc4578 (
      {stage0_62[483]},
      {stage1_62[190]}
   );
   gpc1_1 gpc4579 (
      {stage0_62[484]},
      {stage1_62[191]}
   );
   gpc1_1 gpc4580 (
      {stage0_62[485]},
      {stage1_62[192]}
   );
   gpc1_1 gpc4581 (
      {stage0_63[324]},
      {stage1_63[146]}
   );
   gpc1_1 gpc4582 (
      {stage0_63[325]},
      {stage1_63[147]}
   );
   gpc1_1 gpc4583 (
      {stage0_63[326]},
      {stage1_63[148]}
   );
   gpc1_1 gpc4584 (
      {stage0_63[327]},
      {stage1_63[149]}
   );
   gpc1_1 gpc4585 (
      {stage0_63[328]},
      {stage1_63[150]}
   );
   gpc1_1 gpc4586 (
      {stage0_63[329]},
      {stage1_63[151]}
   );
   gpc1_1 gpc4587 (
      {stage0_63[330]},
      {stage1_63[152]}
   );
   gpc1_1 gpc4588 (
      {stage0_63[331]},
      {stage1_63[153]}
   );
   gpc1_1 gpc4589 (
      {stage0_63[332]},
      {stage1_63[154]}
   );
   gpc1_1 gpc4590 (
      {stage0_63[333]},
      {stage1_63[155]}
   );
   gpc1_1 gpc4591 (
      {stage0_63[334]},
      {stage1_63[156]}
   );
   gpc1_1 gpc4592 (
      {stage0_63[335]},
      {stage1_63[157]}
   );
   gpc1_1 gpc4593 (
      {stage0_63[336]},
      {stage1_63[158]}
   );
   gpc1_1 gpc4594 (
      {stage0_63[337]},
      {stage1_63[159]}
   );
   gpc1_1 gpc4595 (
      {stage0_63[338]},
      {stage1_63[160]}
   );
   gpc1_1 gpc4596 (
      {stage0_63[339]},
      {stage1_63[161]}
   );
   gpc1_1 gpc4597 (
      {stage0_63[340]},
      {stage1_63[162]}
   );
   gpc1_1 gpc4598 (
      {stage0_63[341]},
      {stage1_63[163]}
   );
   gpc1_1 gpc4599 (
      {stage0_63[342]},
      {stage1_63[164]}
   );
   gpc1_1 gpc4600 (
      {stage0_63[343]},
      {stage1_63[165]}
   );
   gpc1_1 gpc4601 (
      {stage0_63[344]},
      {stage1_63[166]}
   );
   gpc1_1 gpc4602 (
      {stage0_63[345]},
      {stage1_63[167]}
   );
   gpc1_1 gpc4603 (
      {stage0_63[346]},
      {stage1_63[168]}
   );
   gpc1_1 gpc4604 (
      {stage0_63[347]},
      {stage1_63[169]}
   );
   gpc1_1 gpc4605 (
      {stage0_63[348]},
      {stage1_63[170]}
   );
   gpc1_1 gpc4606 (
      {stage0_63[349]},
      {stage1_63[171]}
   );
   gpc1_1 gpc4607 (
      {stage0_63[350]},
      {stage1_63[172]}
   );
   gpc1_1 gpc4608 (
      {stage0_63[351]},
      {stage1_63[173]}
   );
   gpc1_1 gpc4609 (
      {stage0_63[352]},
      {stage1_63[174]}
   );
   gpc1_1 gpc4610 (
      {stage0_63[353]},
      {stage1_63[175]}
   );
   gpc1_1 gpc4611 (
      {stage0_63[354]},
      {stage1_63[176]}
   );
   gpc1_1 gpc4612 (
      {stage0_63[355]},
      {stage1_63[177]}
   );
   gpc1_1 gpc4613 (
      {stage0_63[356]},
      {stage1_63[178]}
   );
   gpc1_1 gpc4614 (
      {stage0_63[357]},
      {stage1_63[179]}
   );
   gpc1_1 gpc4615 (
      {stage0_63[358]},
      {stage1_63[180]}
   );
   gpc1_1 gpc4616 (
      {stage0_63[359]},
      {stage1_63[181]}
   );
   gpc1_1 gpc4617 (
      {stage0_63[360]},
      {stage1_63[182]}
   );
   gpc1_1 gpc4618 (
      {stage0_63[361]},
      {stage1_63[183]}
   );
   gpc1_1 gpc4619 (
      {stage0_63[362]},
      {stage1_63[184]}
   );
   gpc1_1 gpc4620 (
      {stage0_63[363]},
      {stage1_63[185]}
   );
   gpc1_1 gpc4621 (
      {stage0_63[364]},
      {stage1_63[186]}
   );
   gpc1_1 gpc4622 (
      {stage0_63[365]},
      {stage1_63[187]}
   );
   gpc1_1 gpc4623 (
      {stage0_63[366]},
      {stage1_63[188]}
   );
   gpc1_1 gpc4624 (
      {stage0_63[367]},
      {stage1_63[189]}
   );
   gpc1_1 gpc4625 (
      {stage0_63[368]},
      {stage1_63[190]}
   );
   gpc1_1 gpc4626 (
      {stage0_63[369]},
      {stage1_63[191]}
   );
   gpc1_1 gpc4627 (
      {stage0_63[370]},
      {stage1_63[192]}
   );
   gpc1_1 gpc4628 (
      {stage0_63[371]},
      {stage1_63[193]}
   );
   gpc1_1 gpc4629 (
      {stage0_63[372]},
      {stage1_63[194]}
   );
   gpc1_1 gpc4630 (
      {stage0_63[373]},
      {stage1_63[195]}
   );
   gpc1_1 gpc4631 (
      {stage0_63[374]},
      {stage1_63[196]}
   );
   gpc1_1 gpc4632 (
      {stage0_63[375]},
      {stage1_63[197]}
   );
   gpc1_1 gpc4633 (
      {stage0_63[376]},
      {stage1_63[198]}
   );
   gpc1_1 gpc4634 (
      {stage0_63[377]},
      {stage1_63[199]}
   );
   gpc1_1 gpc4635 (
      {stage0_63[378]},
      {stage1_63[200]}
   );
   gpc1_1 gpc4636 (
      {stage0_63[379]},
      {stage1_63[201]}
   );
   gpc1_1 gpc4637 (
      {stage0_63[380]},
      {stage1_63[202]}
   );
   gpc1_1 gpc4638 (
      {stage0_63[381]},
      {stage1_63[203]}
   );
   gpc1_1 gpc4639 (
      {stage0_63[382]},
      {stage1_63[204]}
   );
   gpc1_1 gpc4640 (
      {stage0_63[383]},
      {stage1_63[205]}
   );
   gpc1_1 gpc4641 (
      {stage0_63[384]},
      {stage1_63[206]}
   );
   gpc1_1 gpc4642 (
      {stage0_63[385]},
      {stage1_63[207]}
   );
   gpc1_1 gpc4643 (
      {stage0_63[386]},
      {stage1_63[208]}
   );
   gpc1_1 gpc4644 (
      {stage0_63[387]},
      {stage1_63[209]}
   );
   gpc1_1 gpc4645 (
      {stage0_63[388]},
      {stage1_63[210]}
   );
   gpc1_1 gpc4646 (
      {stage0_63[389]},
      {stage1_63[211]}
   );
   gpc1_1 gpc4647 (
      {stage0_63[390]},
      {stage1_63[212]}
   );
   gpc1_1 gpc4648 (
      {stage0_63[391]},
      {stage1_63[213]}
   );
   gpc1_1 gpc4649 (
      {stage0_63[392]},
      {stage1_63[214]}
   );
   gpc1_1 gpc4650 (
      {stage0_63[393]},
      {stage1_63[215]}
   );
   gpc1_1 gpc4651 (
      {stage0_63[394]},
      {stage1_63[216]}
   );
   gpc1_1 gpc4652 (
      {stage0_63[395]},
      {stage1_63[217]}
   );
   gpc1_1 gpc4653 (
      {stage0_63[396]},
      {stage1_63[218]}
   );
   gpc1_1 gpc4654 (
      {stage0_63[397]},
      {stage1_63[219]}
   );
   gpc1_1 gpc4655 (
      {stage0_63[398]},
      {stage1_63[220]}
   );
   gpc1_1 gpc4656 (
      {stage0_63[399]},
      {stage1_63[221]}
   );
   gpc1_1 gpc4657 (
      {stage0_63[400]},
      {stage1_63[222]}
   );
   gpc1_1 gpc4658 (
      {stage0_63[401]},
      {stage1_63[223]}
   );
   gpc1_1 gpc4659 (
      {stage0_63[402]},
      {stage1_63[224]}
   );
   gpc1_1 gpc4660 (
      {stage0_63[403]},
      {stage1_63[225]}
   );
   gpc1_1 gpc4661 (
      {stage0_63[404]},
      {stage1_63[226]}
   );
   gpc1_1 gpc4662 (
      {stage0_63[405]},
      {stage1_63[227]}
   );
   gpc1_1 gpc4663 (
      {stage0_63[406]},
      {stage1_63[228]}
   );
   gpc1_1 gpc4664 (
      {stage0_63[407]},
      {stage1_63[229]}
   );
   gpc1_1 gpc4665 (
      {stage0_63[408]},
      {stage1_63[230]}
   );
   gpc1_1 gpc4666 (
      {stage0_63[409]},
      {stage1_63[231]}
   );
   gpc1_1 gpc4667 (
      {stage0_63[410]},
      {stage1_63[232]}
   );
   gpc1_1 gpc4668 (
      {stage0_63[411]},
      {stage1_63[233]}
   );
   gpc1_1 gpc4669 (
      {stage0_63[412]},
      {stage1_63[234]}
   );
   gpc1_1 gpc4670 (
      {stage0_63[413]},
      {stage1_63[235]}
   );
   gpc1_1 gpc4671 (
      {stage0_63[414]},
      {stage1_63[236]}
   );
   gpc1_1 gpc4672 (
      {stage0_63[415]},
      {stage1_63[237]}
   );
   gpc1_1 gpc4673 (
      {stage0_63[416]},
      {stage1_63[238]}
   );
   gpc1_1 gpc4674 (
      {stage0_63[417]},
      {stage1_63[239]}
   );
   gpc1_1 gpc4675 (
      {stage0_63[418]},
      {stage1_63[240]}
   );
   gpc1_1 gpc4676 (
      {stage0_63[419]},
      {stage1_63[241]}
   );
   gpc1_1 gpc4677 (
      {stage0_63[420]},
      {stage1_63[242]}
   );
   gpc1_1 gpc4678 (
      {stage0_63[421]},
      {stage1_63[243]}
   );
   gpc1_1 gpc4679 (
      {stage0_63[422]},
      {stage1_63[244]}
   );
   gpc1_1 gpc4680 (
      {stage0_63[423]},
      {stage1_63[245]}
   );
   gpc1_1 gpc4681 (
      {stage0_63[424]},
      {stage1_63[246]}
   );
   gpc1_1 gpc4682 (
      {stage0_63[425]},
      {stage1_63[247]}
   );
   gpc1_1 gpc4683 (
      {stage0_63[426]},
      {stage1_63[248]}
   );
   gpc1_1 gpc4684 (
      {stage0_63[427]},
      {stage1_63[249]}
   );
   gpc1_1 gpc4685 (
      {stage0_63[428]},
      {stage1_63[250]}
   );
   gpc1_1 gpc4686 (
      {stage0_63[429]},
      {stage1_63[251]}
   );
   gpc1_1 gpc4687 (
      {stage0_63[430]},
      {stage1_63[252]}
   );
   gpc1_1 gpc4688 (
      {stage0_63[431]},
      {stage1_63[253]}
   );
   gpc1_1 gpc4689 (
      {stage0_63[432]},
      {stage1_63[254]}
   );
   gpc1_1 gpc4690 (
      {stage0_63[433]},
      {stage1_63[255]}
   );
   gpc1_1 gpc4691 (
      {stage0_63[434]},
      {stage1_63[256]}
   );
   gpc1_1 gpc4692 (
      {stage0_63[435]},
      {stage1_63[257]}
   );
   gpc1_1 gpc4693 (
      {stage0_63[436]},
      {stage1_63[258]}
   );
   gpc1_1 gpc4694 (
      {stage0_63[437]},
      {stage1_63[259]}
   );
   gpc1_1 gpc4695 (
      {stage0_63[438]},
      {stage1_63[260]}
   );
   gpc1_1 gpc4696 (
      {stage0_63[439]},
      {stage1_63[261]}
   );
   gpc1_1 gpc4697 (
      {stage0_63[440]},
      {stage1_63[262]}
   );
   gpc1_1 gpc4698 (
      {stage0_63[441]},
      {stage1_63[263]}
   );
   gpc1_1 gpc4699 (
      {stage0_63[442]},
      {stage1_63[264]}
   );
   gpc1_1 gpc4700 (
      {stage0_63[443]},
      {stage1_63[265]}
   );
   gpc1_1 gpc4701 (
      {stage0_63[444]},
      {stage1_63[266]}
   );
   gpc1_1 gpc4702 (
      {stage0_63[445]},
      {stage1_63[267]}
   );
   gpc1_1 gpc4703 (
      {stage0_63[446]},
      {stage1_63[268]}
   );
   gpc1_1 gpc4704 (
      {stage0_63[447]},
      {stage1_63[269]}
   );
   gpc1_1 gpc4705 (
      {stage0_63[448]},
      {stage1_63[270]}
   );
   gpc1_1 gpc4706 (
      {stage0_63[449]},
      {stage1_63[271]}
   );
   gpc1_1 gpc4707 (
      {stage0_63[450]},
      {stage1_63[272]}
   );
   gpc1_1 gpc4708 (
      {stage0_63[451]},
      {stage1_63[273]}
   );
   gpc1_1 gpc4709 (
      {stage0_63[452]},
      {stage1_63[274]}
   );
   gpc1_1 gpc4710 (
      {stage0_63[453]},
      {stage1_63[275]}
   );
   gpc1_1 gpc4711 (
      {stage0_63[454]},
      {stage1_63[276]}
   );
   gpc1_1 gpc4712 (
      {stage0_63[455]},
      {stage1_63[277]}
   );
   gpc1_1 gpc4713 (
      {stage0_63[456]},
      {stage1_63[278]}
   );
   gpc1_1 gpc4714 (
      {stage0_63[457]},
      {stage1_63[279]}
   );
   gpc1_1 gpc4715 (
      {stage0_63[458]},
      {stage1_63[280]}
   );
   gpc1_1 gpc4716 (
      {stage0_63[459]},
      {stage1_63[281]}
   );
   gpc1_1 gpc4717 (
      {stage0_63[460]},
      {stage1_63[282]}
   );
   gpc1_1 gpc4718 (
      {stage0_63[461]},
      {stage1_63[283]}
   );
   gpc1_1 gpc4719 (
      {stage0_63[462]},
      {stage1_63[284]}
   );
   gpc1_1 gpc4720 (
      {stage0_63[463]},
      {stage1_63[285]}
   );
   gpc1_1 gpc4721 (
      {stage0_63[464]},
      {stage1_63[286]}
   );
   gpc1_1 gpc4722 (
      {stage0_63[465]},
      {stage1_63[287]}
   );
   gpc1_1 gpc4723 (
      {stage0_63[466]},
      {stage1_63[288]}
   );
   gpc1_1 gpc4724 (
      {stage0_63[467]},
      {stage1_63[289]}
   );
   gpc1_1 gpc4725 (
      {stage0_63[468]},
      {stage1_63[290]}
   );
   gpc1_1 gpc4726 (
      {stage0_63[469]},
      {stage1_63[291]}
   );
   gpc1_1 gpc4727 (
      {stage0_63[470]},
      {stage1_63[292]}
   );
   gpc1_1 gpc4728 (
      {stage0_63[471]},
      {stage1_63[293]}
   );
   gpc1_1 gpc4729 (
      {stage0_63[472]},
      {stage1_63[294]}
   );
   gpc1_1 gpc4730 (
      {stage0_63[473]},
      {stage1_63[295]}
   );
   gpc1_1 gpc4731 (
      {stage0_63[474]},
      {stage1_63[296]}
   );
   gpc1_1 gpc4732 (
      {stage0_63[475]},
      {stage1_63[297]}
   );
   gpc1_1 gpc4733 (
      {stage0_63[476]},
      {stage1_63[298]}
   );
   gpc1_1 gpc4734 (
      {stage0_63[477]},
      {stage1_63[299]}
   );
   gpc1_1 gpc4735 (
      {stage0_63[478]},
      {stage1_63[300]}
   );
   gpc1_1 gpc4736 (
      {stage0_63[479]},
      {stage1_63[301]}
   );
   gpc1_1 gpc4737 (
      {stage0_63[480]},
      {stage1_63[302]}
   );
   gpc1_1 gpc4738 (
      {stage0_63[481]},
      {stage1_63[303]}
   );
   gpc1_1 gpc4739 (
      {stage0_63[482]},
      {stage1_63[304]}
   );
   gpc1_1 gpc4740 (
      {stage0_63[483]},
      {stage1_63[305]}
   );
   gpc1_1 gpc4741 (
      {stage0_63[484]},
      {stage1_63[306]}
   );
   gpc1_1 gpc4742 (
      {stage0_63[485]},
      {stage1_63[307]}
   );
   gpc606_5 gpc4743 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc4744 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc4745 (
      {stage1_0[12], stage1_0[13], stage1_0[14], stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc4746 (
      {stage1_0[18], stage1_0[19], stage1_0[20], stage1_0[21], stage1_0[22]},
      {stage1_1[0]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc4747 (
      {stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27]},
      {stage1_1[1]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc4748 (
      {stage1_0[28], stage1_0[29], stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[2]},
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc4749 (
      {stage1_0[33], stage1_0[34], stage1_0[35], stage1_0[36], stage1_0[37]},
      {stage1_1[3]},
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc615_5 gpc4750 (
      {stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41], stage1_0[42]},
      {stage1_1[4]},
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc615_5 gpc4751 (
      {stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_1[5]},
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc615_5 gpc4752 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52]},
      {stage1_1[6]},
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc615_5 gpc4753 (
      {stage1_0[53], stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57]},
      {stage1_1[7]},
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc615_5 gpc4754 (
      {stage1_0[58], stage1_0[59], stage1_0[60], stage1_0[61], stage1_0[62]},
      {stage1_1[8]},
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc615_5 gpc4755 (
      {stage1_0[63], stage1_0[64], stage1_0[65], stage1_0[66], stage1_0[67]},
      {stage1_1[9]},
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc615_5 gpc4756 (
      {stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71], stage1_0[72]},
      {stage1_1[10]},
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc615_5 gpc4757 (
      {stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_1[11]},
      {stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87], stage1_2[88], stage1_2[89]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc615_5 gpc4758 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82]},
      {stage1_1[12]},
      {stage1_2[90], stage1_2[91], stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc615_5 gpc4759 (
      {stage1_0[83], stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87]},
      {stage1_1[13]},
      {stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc615_5 gpc4760 (
      {stage1_0[88], stage1_0[89], stage1_0[90], stage1_0[91], stage1_0[92]},
      {stage1_1[14]},
      {stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc615_5 gpc4761 (
      {stage1_0[93], stage1_0[94], stage1_0[95], stage1_0[96], stage1_0[97]},
      {stage1_1[15]},
      {stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112], stage1_2[113]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc615_5 gpc4762 (
      {stage1_0[98], stage1_0[99], stage1_0[100], stage1_0[101], stage1_0[102]},
      {stage1_1[16]},
      {stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117], stage1_2[118], stage1_2[119]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc615_5 gpc4763 (
      {stage1_0[103], stage1_0[104], stage1_0[105], stage1_0[106], stage1_0[107]},
      {stage1_1[17]},
      {stage1_2[120], stage1_2[121], stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc4764 (
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc606_5 gpc4765 (
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc4766 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc4767 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc4768 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29]},
      {stage2_5[4],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc4769 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage2_5[5],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc4770 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage2_5[6],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc4771 (
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage2_5[7],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc4772 (
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage2_5[8],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc4773 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59]},
      {stage2_5[9],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc4774 (
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage2_5[10],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc4775 (
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage2_5[11],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc4776 (
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77]},
      {stage2_5[12],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc4777 (
      {stage1_1[96], stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101]},
      {stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage2_5[13],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc4778 (
      {stage1_1[102], stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107]},
      {stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89]},
      {stage2_5[14],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc4779 (
      {stage1_1[108], stage1_1[109], stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113]},
      {stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage2_5[15],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc4780 (
      {stage1_1[114], stage1_1[115], stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119]},
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101]},
      {stage2_5[16],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc4781 (
      {stage1_1[120], stage1_1[121], stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125]},
      {stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage2_5[17],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc606_5 gpc4782 (
      {stage1_1[126], stage1_1[127], stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131]},
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113]},
      {stage2_5[18],stage2_4[39],stage2_3[39],stage2_2[39],stage2_1[39]}
   );
   gpc606_5 gpc4783 (
      {stage1_1[132], stage1_1[133], stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137]},
      {stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119]},
      {stage2_5[19],stage2_4[40],stage2_3[40],stage2_2[40],stage2_1[40]}
   );
   gpc606_5 gpc4784 (
      {stage1_1[138], stage1_1[139], stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143]},
      {stage1_3[120], stage1_3[121], stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125]},
      {stage2_5[20],stage2_4[41],stage2_3[41],stage2_2[41],stage2_1[41]}
   );
   gpc606_5 gpc4785 (
      {stage1_1[144], stage1_1[145], stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149]},
      {stage1_3[126], stage1_3[127], stage1_3[128], stage1_3[129], stage1_3[130], stage1_3[131]},
      {stage2_5[21],stage2_4[42],stage2_3[42],stage2_2[42],stage2_1[42]}
   );
   gpc606_5 gpc4786 (
      {stage1_1[150], stage1_1[151], stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155]},
      {stage1_3[132], stage1_3[133], stage1_3[134], stage1_3[135], stage1_3[136], stage1_3[137]},
      {stage2_5[22],stage2_4[43],stage2_3[43],stage2_2[43],stage2_1[43]}
   );
   gpc606_5 gpc4787 (
      {stage1_1[156], stage1_1[157], stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161]},
      {stage1_3[138], stage1_3[139], stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143]},
      {stage2_5[23],stage2_4[44],stage2_3[44],stage2_2[44],stage2_1[44]}
   );
   gpc606_5 gpc4788 (
      {stage1_1[162], stage1_1[163], stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167]},
      {stage1_3[144], stage1_3[145], stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149]},
      {stage2_5[24],stage2_4[45],stage2_3[45],stage2_2[45],stage2_1[45]}
   );
   gpc606_5 gpc4789 (
      {stage1_2[126], stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[25],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc606_5 gpc4790 (
      {stage1_2[132], stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[26],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc606_5 gpc4791 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142], stage1_2[143]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[27],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc1343_5 gpc4792 (
      {stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3]},
      {stage1_6[0], stage1_6[1], stage1_6[2]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[0],stage2_6[3],stage2_5[28],stage2_4[49]}
   );
   gpc1406_5 gpc4793 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage1_7[1]},
      {stage2_8[1],stage2_7[1],stage2_6[4],stage2_5[29],stage2_4[50]}
   );
   gpc606_5 gpc4794 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[2],stage2_6[5],stage2_5[30],stage2_4[51]}
   );
   gpc606_5 gpc4795 (
      {stage1_4[33], stage1_4[34], stage1_4[35], stage1_4[36], stage1_4[37], stage1_4[38]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[3],stage2_7[3],stage2_6[6],stage2_5[31],stage2_4[52]}
   );
   gpc606_5 gpc4796 (
      {stage1_4[39], stage1_4[40], stage1_4[41], stage1_4[42], stage1_4[43], stage1_4[44]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[4],stage2_7[4],stage2_6[7],stage2_5[32],stage2_4[53]}
   );
   gpc606_5 gpc4797 (
      {stage1_4[45], stage1_4[46], stage1_4[47], stage1_4[48], stage1_4[49], stage1_4[50]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[5],stage2_7[5],stage2_6[8],stage2_5[33],stage2_4[54]}
   );
   gpc606_5 gpc4798 (
      {stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[6],stage2_7[6],stage2_6[9],stage2_5[34],stage2_4[55]}
   );
   gpc606_5 gpc4799 (
      {stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[7],stage2_7[7],stage2_6[10],stage2_5[35],stage2_4[56]}
   );
   gpc606_5 gpc4800 (
      {stage1_4[63], stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67], stage1_4[68]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[8],stage2_7[8],stage2_6[11],stage2_5[36],stage2_4[57]}
   );
   gpc606_5 gpc4801 (
      {stage1_4[69], stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73], stage1_4[74]},
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage2_8[9],stage2_7[9],stage2_6[12],stage2_5[37],stage2_4[58]}
   );
   gpc606_5 gpc4802 (
      {stage1_4[75], stage1_4[76], stage1_4[77], stage1_4[78], stage1_4[79], stage1_4[80]},
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage2_8[10],stage2_7[10],stage2_6[13],stage2_5[38],stage2_4[59]}
   );
   gpc606_5 gpc4803 (
      {stage1_4[81], stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86]},
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage2_8[11],stage2_7[11],stage2_6[14],stage2_5[39],stage2_4[60]}
   );
   gpc606_5 gpc4804 (
      {stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91], stage1_4[92]},
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72]},
      {stage2_8[12],stage2_7[12],stage2_6[15],stage2_5[40],stage2_4[61]}
   );
   gpc606_5 gpc4805 (
      {stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96], stage1_4[97], stage1_4[98]},
      {stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78]},
      {stage2_8[13],stage2_7[13],stage2_6[16],stage2_5[41],stage2_4[62]}
   );
   gpc606_5 gpc4806 (
      {stage1_4[99], stage1_4[100], stage1_4[101], stage1_4[102], stage1_4[103], stage1_4[104]},
      {stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage2_8[14],stage2_7[14],stage2_6[17],stage2_5[42],stage2_4[63]}
   );
   gpc606_5 gpc4807 (
      {stage1_4[105], stage1_4[106], stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110]},
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage2_8[15],stage2_7[15],stage2_6[18],stage2_5[43],stage2_4[64]}
   );
   gpc606_5 gpc4808 (
      {stage1_4[111], stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116]},
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage2_8[16],stage2_7[16],stage2_6[19],stage2_5[44],stage2_4[65]}
   );
   gpc606_5 gpc4809 (
      {stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121], stage1_4[122]},
      {stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102]},
      {stage2_8[17],stage2_7[17],stage2_6[20],stage2_5[45],stage2_4[66]}
   );
   gpc606_5 gpc4810 (
      {stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126], stage1_4[127], stage1_4[128]},
      {stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108]},
      {stage2_8[18],stage2_7[18],stage2_6[21],stage2_5[46],stage2_4[67]}
   );
   gpc606_5 gpc4811 (
      {stage1_4[129], stage1_4[130], stage1_4[131], stage1_4[132], stage1_4[133], stage1_4[134]},
      {stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage2_8[19],stage2_7[19],stage2_6[22],stage2_5[47],stage2_4[68]}
   );
   gpc606_5 gpc4812 (
      {stage1_4[135], stage1_4[136], stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140]},
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119], stage1_6[120]},
      {stage2_8[20],stage2_7[20],stage2_6[23],stage2_5[48],stage2_4[69]}
   );
   gpc606_5 gpc4813 (
      {stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146]},
      {stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125], stage1_6[126]},
      {stage2_8[21],stage2_7[21],stage2_6[24],stage2_5[49],stage2_4[70]}
   );
   gpc606_5 gpc4814 (
      {stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151], stage1_4[152]},
      {stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131], stage1_6[132]},
      {stage2_8[22],stage2_7[22],stage2_6[25],stage2_5[50],stage2_4[71]}
   );
   gpc606_5 gpc4815 (
      {stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156], stage1_4[157], stage1_4[158]},
      {stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137], stage1_6[138]},
      {stage2_8[23],stage2_7[23],stage2_6[26],stage2_5[51],stage2_4[72]}
   );
   gpc606_5 gpc4816 (
      {stage1_4[159], stage1_4[160], stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164]},
      {stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143], stage1_6[144]},
      {stage2_8[24],stage2_7[24],stage2_6[27],stage2_5[52],stage2_4[73]}
   );
   gpc606_5 gpc4817 (
      {stage1_4[165], stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170]},
      {stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149], stage1_6[150]},
      {stage2_8[25],stage2_7[25],stage2_6[28],stage2_5[53],stage2_4[74]}
   );
   gpc606_5 gpc4818 (
      {stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176]},
      {stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155], stage1_6[156]},
      {stage2_8[26],stage2_7[26],stage2_6[29],stage2_5[54],stage2_4[75]}
   );
   gpc606_5 gpc4819 (
      {stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181], stage1_4[182]},
      {stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161], stage1_6[162]},
      {stage2_8[27],stage2_7[27],stage2_6[30],stage2_5[55],stage2_4[76]}
   );
   gpc606_5 gpc4820 (
      {stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186], stage1_4[187], stage1_4[188]},
      {stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167], stage1_6[168]},
      {stage2_8[28],stage2_7[28],stage2_6[31],stage2_5[56],stage2_4[77]}
   );
   gpc606_5 gpc4821 (
      {stage1_4[189], stage1_4[190], stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194]},
      {stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173], stage1_6[174]},
      {stage2_8[29],stage2_7[29],stage2_6[32],stage2_5[57],stage2_4[78]}
   );
   gpc606_5 gpc4822 (
      {stage1_5[4], stage1_5[5], stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9]},
      {stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage2_9[0],stage2_8[30],stage2_7[30],stage2_6[33],stage2_5[58]}
   );
   gpc606_5 gpc4823 (
      {stage1_5[10], stage1_5[11], stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15]},
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[31],stage2_7[31],stage2_6[34],stage2_5[59]}
   );
   gpc606_5 gpc4824 (
      {stage1_5[16], stage1_5[17], stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21]},
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19]},
      {stage2_9[2],stage2_8[32],stage2_7[32],stage2_6[35],stage2_5[60]}
   );
   gpc606_5 gpc4825 (
      {stage1_5[22], stage1_5[23], stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27]},
      {stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24], stage1_7[25]},
      {stage2_9[3],stage2_8[33],stage2_7[33],stage2_6[36],stage2_5[61]}
   );
   gpc606_5 gpc4826 (
      {stage1_5[28], stage1_5[29], stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33]},
      {stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31]},
      {stage2_9[4],stage2_8[34],stage2_7[34],stage2_6[37],stage2_5[62]}
   );
   gpc606_5 gpc4827 (
      {stage1_5[34], stage1_5[35], stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39]},
      {stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37]},
      {stage2_9[5],stage2_8[35],stage2_7[35],stage2_6[38],stage2_5[63]}
   );
   gpc606_5 gpc4828 (
      {stage1_5[40], stage1_5[41], stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45]},
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage2_9[6],stage2_8[36],stage2_7[36],stage2_6[39],stage2_5[64]}
   );
   gpc606_5 gpc4829 (
      {stage1_5[46], stage1_5[47], stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51]},
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48], stage1_7[49]},
      {stage2_9[7],stage2_8[37],stage2_7[37],stage2_6[40],stage2_5[65]}
   );
   gpc606_5 gpc4830 (
      {stage1_5[52], stage1_5[53], stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57]},
      {stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54], stage1_7[55]},
      {stage2_9[8],stage2_8[38],stage2_7[38],stage2_6[41],stage2_5[66]}
   );
   gpc606_5 gpc4831 (
      {stage1_5[58], stage1_5[59], stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63]},
      {stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61]},
      {stage2_9[9],stage2_8[39],stage2_7[39],stage2_6[42],stage2_5[67]}
   );
   gpc606_5 gpc4832 (
      {stage1_5[64], stage1_5[65], stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69]},
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66], stage1_7[67]},
      {stage2_9[10],stage2_8[40],stage2_7[40],stage2_6[43],stage2_5[68]}
   );
   gpc606_5 gpc4833 (
      {stage1_5[70], stage1_5[71], stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75]},
      {stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71], stage1_7[72], stage1_7[73]},
      {stage2_9[11],stage2_8[41],stage2_7[41],stage2_6[44],stage2_5[69]}
   );
   gpc606_5 gpc4834 (
      {stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81]},
      {stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77], stage1_7[78], stage1_7[79]},
      {stage2_9[12],stage2_8[42],stage2_7[42],stage2_6[45],stage2_5[70]}
   );
   gpc606_5 gpc4835 (
      {stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87]},
      {stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85]},
      {stage2_9[13],stage2_8[43],stage2_7[43],stage2_6[46],stage2_5[71]}
   );
   gpc606_5 gpc4836 (
      {stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93]},
      {stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage2_9[14],stage2_8[44],stage2_7[44],stage2_6[47],stage2_5[72]}
   );
   gpc606_5 gpc4837 (
      {stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99]},
      {stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95], stage1_7[96], stage1_7[97]},
      {stage2_9[15],stage2_8[45],stage2_7[45],stage2_6[48],stage2_5[73]}
   );
   gpc606_5 gpc4838 (
      {stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105]},
      {stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101], stage1_7[102], stage1_7[103]},
      {stage2_9[16],stage2_8[46],stage2_7[46],stage2_6[49],stage2_5[74]}
   );
   gpc606_5 gpc4839 (
      {stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111]},
      {stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107], stage1_7[108], stage1_7[109]},
      {stage2_9[17],stage2_8[47],stage2_7[47],stage2_6[50],stage2_5[75]}
   );
   gpc606_5 gpc4840 (
      {stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117]},
      {stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114], stage1_7[115]},
      {stage2_9[18],stage2_8[48],stage2_7[48],stage2_6[51],stage2_5[76]}
   );
   gpc606_5 gpc4841 (
      {stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123]},
      {stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120], stage1_7[121]},
      {stage2_9[19],stage2_8[49],stage2_7[49],stage2_6[52],stage2_5[77]}
   );
   gpc615_5 gpc4842 (
      {stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[20],stage2_8[50],stage2_7[50]}
   );
   gpc615_5 gpc4843 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[21],stage2_8[51],stage2_7[51]}
   );
   gpc615_5 gpc4844 (
      {stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136]},
      {stage1_8[2]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[2],stage2_9[22],stage2_8[52],stage2_7[52]}
   );
   gpc615_5 gpc4845 (
      {stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140], stage1_7[141]},
      {stage1_8[3]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[3],stage2_9[23],stage2_8[53],stage2_7[53]}
   );
   gpc615_5 gpc4846 (
      {stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145], stage1_7[146]},
      {stage1_8[4]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[4],stage2_9[24],stage2_8[54],stage2_7[54]}
   );
   gpc615_5 gpc4847 (
      {stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150], stage1_7[151]},
      {stage1_8[5]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[5],stage2_9[25],stage2_8[55],stage2_7[55]}
   );
   gpc615_5 gpc4848 (
      {stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_8[6]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[6],stage2_9[26],stage2_8[56],stage2_7[56]}
   );
   gpc615_5 gpc4849 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161]},
      {stage1_8[7]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[7],stage2_9[27],stage2_8[57],stage2_7[57]}
   );
   gpc615_5 gpc4850 (
      {stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165], stage1_7[166]},
      {stage1_8[8]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[8],stage2_9[28],stage2_8[58],stage2_7[58]}
   );
   gpc615_5 gpc4851 (
      {stage1_7[167], stage1_7[168], stage1_7[169], stage1_7[170], stage1_7[171]},
      {stage1_8[9]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[9],stage2_9[29],stage2_8[59],stage2_7[59]}
   );
   gpc615_5 gpc4852 (
      {stage1_7[172], stage1_7[173], stage1_7[174], stage1_7[175], stage1_7[176]},
      {stage1_8[10]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[10],stage2_9[30],stage2_8[60],stage2_7[60]}
   );
   gpc615_5 gpc4853 (
      {stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180], stage1_7[181]},
      {stage1_8[11]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[11],stage2_9[31],stage2_8[61],stage2_7[61]}
   );
   gpc615_5 gpc4854 (
      {stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185], stage1_7[186]},
      {stage1_8[12]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[12],stage2_9[32],stage2_8[62],stage2_7[62]}
   );
   gpc615_5 gpc4855 (
      {stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190], stage1_7[191]},
      {stage1_8[13]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[13],stage2_9[33],stage2_8[63],stage2_7[63]}
   );
   gpc615_5 gpc4856 (
      {stage1_7[192], stage1_7[193], stage1_7[194], stage1_7[195], stage1_7[196]},
      {stage1_8[14]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[14],stage2_9[34],stage2_8[64],stage2_7[64]}
   );
   gpc615_5 gpc4857 (
      {stage1_7[197], stage1_7[198], stage1_7[199], stage1_7[200], stage1_7[201]},
      {stage1_8[15]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[15],stage2_9[35],stage2_8[65],stage2_7[65]}
   );
   gpc615_5 gpc4858 (
      {stage1_7[202], stage1_7[203], stage1_7[204], stage1_7[205], stage1_7[206]},
      {stage1_8[16]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[16],stage2_9[36],stage2_8[66],stage2_7[66]}
   );
   gpc615_5 gpc4859 (
      {stage1_7[207], stage1_7[208], stage1_7[209], stage1_7[210], stage1_7[211]},
      {stage1_8[17]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[17],stage2_9[37],stage2_8[67],stage2_7[67]}
   );
   gpc615_5 gpc4860 (
      {stage1_7[212], stage1_7[213], stage1_7[214], stage1_7[215], stage1_7[216]},
      {stage1_8[18]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[18],stage2_9[38],stage2_8[68],stage2_7[68]}
   );
   gpc207_4 gpc4861 (
      {stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25]},
      {stage1_10[0], stage1_10[1]},
      {stage2_11[19],stage2_10[19],stage2_9[39],stage2_8[69]}
   );
   gpc606_5 gpc4862 (
      {stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31]},
      {stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6], stage1_10[7]},
      {stage2_12[0],stage2_11[20],stage2_10[20],stage2_9[40],stage2_8[70]}
   );
   gpc606_5 gpc4863 (
      {stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37]},
      {stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12], stage1_10[13]},
      {stage2_12[1],stage2_11[21],stage2_10[21],stage2_9[41],stage2_8[71]}
   );
   gpc606_5 gpc4864 (
      {stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43]},
      {stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19]},
      {stage2_12[2],stage2_11[22],stage2_10[22],stage2_9[42],stage2_8[72]}
   );
   gpc606_5 gpc4865 (
      {stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49]},
      {stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25]},
      {stage2_12[3],stage2_11[23],stage2_10[23],stage2_9[43],stage2_8[73]}
   );
   gpc606_5 gpc4866 (
      {stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54], stage1_8[55]},
      {stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30], stage1_10[31]},
      {stage2_12[4],stage2_11[24],stage2_10[24],stage2_9[44],stage2_8[74]}
   );
   gpc606_5 gpc4867 (
      {stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59], stage1_8[60], stage1_8[61]},
      {stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36], stage1_10[37]},
      {stage2_12[5],stage2_11[25],stage2_10[25],stage2_9[45],stage2_8[75]}
   );
   gpc606_5 gpc4868 (
      {stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66], stage1_8[67]},
      {stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42], stage1_10[43]},
      {stage2_12[6],stage2_11[26],stage2_10[26],stage2_9[46],stage2_8[76]}
   );
   gpc606_5 gpc4869 (
      {stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71], stage1_8[72], stage1_8[73]},
      {stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49]},
      {stage2_12[7],stage2_11[27],stage2_10[27],stage2_9[47],stage2_8[77]}
   );
   gpc606_5 gpc4870 (
      {stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77], stage1_8[78], stage1_8[79]},
      {stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55]},
      {stage2_12[8],stage2_11[28],stage2_10[28],stage2_9[48],stage2_8[78]}
   );
   gpc606_5 gpc4871 (
      {stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83], stage1_8[84], stage1_8[85]},
      {stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61]},
      {stage2_12[9],stage2_11[29],stage2_10[29],stage2_9[49],stage2_8[79]}
   );
   gpc606_5 gpc4872 (
      {stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89], stage1_8[90], stage1_8[91]},
      {stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67]},
      {stage2_12[10],stage2_11[30],stage2_10[30],stage2_9[50],stage2_8[80]}
   );
   gpc606_5 gpc4873 (
      {stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95], stage1_8[96], stage1_8[97]},
      {stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72], stage1_10[73]},
      {stage2_12[11],stage2_11[31],stage2_10[31],stage2_9[51],stage2_8[81]}
   );
   gpc606_5 gpc4874 (
      {stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101], stage1_8[102], stage1_8[103]},
      {stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78], stage1_10[79]},
      {stage2_12[12],stage2_11[32],stage2_10[32],stage2_9[52],stage2_8[82]}
   );
   gpc606_5 gpc4875 (
      {stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107], stage1_8[108], stage1_8[109]},
      {stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83], stage1_10[84], stage1_10[85]},
      {stage2_12[13],stage2_11[33],stage2_10[33],stage2_9[53],stage2_8[83]}
   );
   gpc606_5 gpc4876 (
      {stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113], stage1_8[114], stage1_8[115]},
      {stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90], stage1_10[91]},
      {stage2_12[14],stage2_11[34],stage2_10[34],stage2_9[54],stage2_8[84]}
   );
   gpc606_5 gpc4877 (
      {stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119], stage1_8[120], stage1_8[121]},
      {stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96], stage1_10[97]},
      {stage2_12[15],stage2_11[35],stage2_10[35],stage2_9[55],stage2_8[85]}
   );
   gpc606_5 gpc4878 (
      {stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125], stage1_8[126], stage1_8[127]},
      {stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101], stage1_10[102], stage1_10[103]},
      {stage2_12[16],stage2_11[36],stage2_10[36],stage2_9[56],stage2_8[86]}
   );
   gpc606_5 gpc4879 (
      {stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131], stage1_8[132], stage1_8[133]},
      {stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107], stage1_10[108], stage1_10[109]},
      {stage2_12[17],stage2_11[37],stage2_10[37],stage2_9[57],stage2_8[87]}
   );
   gpc606_5 gpc4880 (
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[18],stage2_11[38],stage2_10[38],stage2_9[58]}
   );
   gpc606_5 gpc4881 (
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[19],stage2_11[39],stage2_10[39],stage2_9[59]}
   );
   gpc606_5 gpc4882 (
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[20],stage2_11[40],stage2_10[40],stage2_9[60]}
   );
   gpc615_5 gpc4883 (
      {stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113], stage1_10[114]},
      {stage1_11[18]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[3],stage2_12[21],stage2_11[41],stage2_10[41]}
   );
   gpc615_5 gpc4884 (
      {stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage1_11[19]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[4],stage2_12[22],stage2_11[42],stage2_10[42]}
   );
   gpc615_5 gpc4885 (
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124]},
      {stage1_11[20]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[5],stage2_12[23],stage2_11[43],stage2_10[43]}
   );
   gpc615_5 gpc4886 (
      {stage1_10[125], stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129]},
      {stage1_11[21]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[6],stage2_12[24],stage2_11[44],stage2_10[44]}
   );
   gpc615_5 gpc4887 (
      {stage1_10[130], stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134]},
      {stage1_11[22]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[7],stage2_12[25],stage2_11[45],stage2_10[45]}
   );
   gpc615_5 gpc4888 (
      {stage1_10[135], stage1_10[136], stage1_10[137], stage1_10[138], stage1_10[139]},
      {stage1_11[23]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[8],stage2_12[26],stage2_11[46],stage2_10[46]}
   );
   gpc615_5 gpc4889 (
      {stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143], stage1_10[144]},
      {stage1_11[24]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[9],stage2_12[27],stage2_11[47],stage2_10[47]}
   );
   gpc615_5 gpc4890 (
      {stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage1_11[25]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[10],stage2_12[28],stage2_11[48],stage2_10[48]}
   );
   gpc615_5 gpc4891 (
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154]},
      {stage1_11[26]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[11],stage2_12[29],stage2_11[49],stage2_10[49]}
   );
   gpc615_5 gpc4892 (
      {stage1_10[155], stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159]},
      {stage1_11[27]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[12],stage2_12[30],stage2_11[50],stage2_10[50]}
   );
   gpc615_5 gpc4893 (
      {stage1_10[160], stage1_10[161], stage1_10[162], stage1_10[163], stage1_10[164]},
      {stage1_11[28]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[13],stage2_12[31],stage2_11[51],stage2_10[51]}
   );
   gpc615_5 gpc4894 (
      {stage1_10[165], stage1_10[166], stage1_10[167], stage1_10[168], stage1_10[169]},
      {stage1_11[29]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[14],stage2_12[32],stage2_11[52],stage2_10[52]}
   );
   gpc615_5 gpc4895 (
      {stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173], stage1_10[174]},
      {stage1_11[30]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[15],stage2_12[33],stage2_11[53],stage2_10[53]}
   );
   gpc606_5 gpc4896 (
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[13],stage2_13[16],stage2_12[34],stage2_11[54]}
   );
   gpc606_5 gpc4897 (
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[14],stage2_13[17],stage2_12[35],stage2_11[55]}
   );
   gpc606_5 gpc4898 (
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[15],stage2_13[18],stage2_12[36],stage2_11[56]}
   );
   gpc606_5 gpc4899 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[16],stage2_13[19],stage2_12[37],stage2_11[57]}
   );
   gpc606_5 gpc4900 (
      {stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59], stage1_11[60]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[17],stage2_13[20],stage2_12[38],stage2_11[58]}
   );
   gpc606_5 gpc4901 (
      {stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65], stage1_11[66]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[18],stage2_13[21],stage2_12[39],stage2_11[59]}
   );
   gpc606_5 gpc4902 (
      {stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[19],stage2_13[22],stage2_12[40],stage2_11[60]}
   );
   gpc606_5 gpc4903 (
      {stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77], stage1_11[78]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[20],stage2_13[23],stage2_12[41],stage2_11[61]}
   );
   gpc606_5 gpc4904 (
      {stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83], stage1_11[84]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[21],stage2_13[24],stage2_12[42],stage2_11[62]}
   );
   gpc606_5 gpc4905 (
      {stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89], stage1_11[90]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[22],stage2_13[25],stage2_12[43],stage2_11[63]}
   );
   gpc606_5 gpc4906 (
      {stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95], stage1_11[96]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[23],stage2_13[26],stage2_12[44],stage2_11[64]}
   );
   gpc606_5 gpc4907 (
      {stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101], stage1_11[102]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[24],stage2_13[27],stage2_12[45],stage2_11[65]}
   );
   gpc606_5 gpc4908 (
      {stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108]},
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage2_15[12],stage2_14[25],stage2_13[28],stage2_12[46],stage2_11[66]}
   );
   gpc606_5 gpc4909 (
      {stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage2_15[13],stage2_14[26],stage2_13[29],stage2_12[47],stage2_11[67]}
   );
   gpc606_5 gpc4910 (
      {stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119], stage1_11[120]},
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage2_15[14],stage2_14[27],stage2_13[30],stage2_12[48],stage2_11[68]}
   );
   gpc606_5 gpc4911 (
      {stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125], stage1_11[126]},
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage2_15[15],stage2_14[28],stage2_13[31],stage2_12[49],stage2_11[69]}
   );
   gpc606_5 gpc4912 (
      {stage1_11[127], stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131], stage1_11[132]},
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage2_15[16],stage2_14[29],stage2_13[32],stage2_12[50],stage2_11[70]}
   );
   gpc615_5 gpc4913 (
      {stage1_11[133], stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137]},
      {stage1_12[78]},
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage2_15[17],stage2_14[30],stage2_13[33],stage2_12[51],stage2_11[71]}
   );
   gpc615_5 gpc4914 (
      {stage1_11[138], stage1_11[139], stage1_11[140], stage1_11[141], stage1_11[142]},
      {stage1_12[79]},
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage2_15[18],stage2_14[31],stage2_13[34],stage2_12[52],stage2_11[72]}
   );
   gpc615_5 gpc4915 (
      {stage1_11[143], stage1_11[144], stage1_11[145], stage1_11[146], stage1_11[147]},
      {stage1_12[80]},
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage2_15[19],stage2_14[32],stage2_13[35],stage2_12[53],stage2_11[73]}
   );
   gpc615_5 gpc4916 (
      {stage1_11[148], stage1_11[149], stage1_11[150], stage1_11[151], stage1_11[152]},
      {stage1_12[81]},
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage2_15[20],stage2_14[33],stage2_13[36],stage2_12[54],stage2_11[74]}
   );
   gpc615_5 gpc4917 (
      {stage1_11[153], stage1_11[154], stage1_11[155], stage1_11[156], stage1_11[157]},
      {stage1_12[82]},
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage2_15[21],stage2_14[34],stage2_13[37],stage2_12[55],stage2_11[75]}
   );
   gpc615_5 gpc4918 (
      {stage1_11[158], stage1_11[159], stage1_11[160], stage1_11[161], stage1_11[162]},
      {stage1_12[83]},
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage2_15[22],stage2_14[35],stage2_13[38],stage2_12[56],stage2_11[76]}
   );
   gpc615_5 gpc4919 (
      {stage1_11[163], stage1_11[164], stage1_11[165], stage1_11[166], stage1_11[167]},
      {stage1_12[84]},
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage2_15[23],stage2_14[36],stage2_13[39],stage2_12[57],stage2_11[77]}
   );
   gpc615_5 gpc4920 (
      {stage1_11[168], stage1_11[169], stage1_11[170], stage1_11[171], stage1_11[172]},
      {stage1_12[85]},
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage2_15[24],stage2_14[37],stage2_13[40],stage2_12[58],stage2_11[78]}
   );
   gpc615_5 gpc4921 (
      {stage1_11[173], stage1_11[174], stage1_11[175], stage1_11[176], stage1_11[177]},
      {stage1_12[86]},
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155]},
      {stage2_15[25],stage2_14[38],stage2_13[41],stage2_12[59],stage2_11[79]}
   );
   gpc615_5 gpc4922 (
      {stage1_11[178], stage1_11[179], stage1_11[180], stage1_11[181], stage1_11[182]},
      {stage1_12[87]},
      {stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage2_15[26],stage2_14[39],stage2_13[42],stage2_12[60],stage2_11[80]}
   );
   gpc615_5 gpc4923 (
      {stage1_11[183], stage1_11[184], stage1_11[185], stage1_11[186], stage1_11[187]},
      {stage1_12[88]},
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166], stage1_13[167]},
      {stage2_15[27],stage2_14[40],stage2_13[43],stage2_12[61],stage2_11[81]}
   );
   gpc615_5 gpc4924 (
      {stage1_11[188], stage1_11[189], stage1_11[190], stage1_11[191], stage1_11[192]},
      {stage1_12[89]},
      {stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173]},
      {stage2_15[28],stage2_14[41],stage2_13[44],stage2_12[62],stage2_11[82]}
   );
   gpc615_5 gpc4925 (
      {stage1_11[193], stage1_11[194], stage1_11[195], stage1_11[196], stage1_11[197]},
      {stage1_12[90]},
      {stage1_13[174], stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage2_15[29],stage2_14[42],stage2_13[45],stage2_12[63],stage2_11[83]}
   );
   gpc615_5 gpc4926 (
      {stage1_11[198], stage1_11[199], stage1_11[200], stage1_11[201], stage1_11[202]},
      {stage1_12[91]},
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184], stage1_13[185]},
      {stage2_15[30],stage2_14[43],stage2_13[46],stage2_12[64],stage2_11[84]}
   );
   gpc615_5 gpc4927 (
      {stage1_11[203], stage1_11[204], stage1_11[205], stage1_11[206], stage1_11[207]},
      {stage1_12[92]},
      {stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189], stage1_13[190], stage1_13[191]},
      {stage2_15[31],stage2_14[44],stage2_13[47],stage2_12[65],stage2_11[85]}
   );
   gpc615_5 gpc4928 (
      {stage1_11[208], stage1_11[209], stage1_11[210], stage1_11[211], stage1_11[212]},
      {stage1_12[93]},
      {stage1_13[192], stage1_13[193], stage1_13[194], stage1_13[195], stage1_13[196], stage1_13[197]},
      {stage2_15[32],stage2_14[45],stage2_13[48],stage2_12[66],stage2_11[86]}
   );
   gpc615_5 gpc4929 (
      {stage1_11[213], stage1_11[214], stage1_11[215], stage1_11[216], stage1_11[217]},
      {stage1_12[94]},
      {stage1_13[198], stage1_13[199], stage1_13[200], stage1_13[201], stage1_13[202], stage1_13[203]},
      {stage2_15[33],stage2_14[46],stage2_13[49],stage2_12[67],stage2_11[87]}
   );
   gpc615_5 gpc4930 (
      {stage1_11[218], stage1_11[219], stage1_11[220], stage1_11[221], stage1_11[222]},
      {stage1_12[95]},
      {stage1_13[204], stage1_13[205], stage1_13[206], stage1_13[207], stage1_13[208], stage1_13[209]},
      {stage2_15[34],stage2_14[47],stage2_13[50],stage2_12[68],stage2_11[88]}
   );
   gpc1325_5 gpc4931 (
      {stage1_11[223], stage1_11[224], stage1_11[225], stage1_11[226], stage1_11[227]},
      {stage1_12[96], stage1_12[97]},
      {stage1_13[210], stage1_13[211], stage1_13[212]},
      {stage1_14[0]},
      {stage2_15[35],stage2_14[48],stage2_13[51],stage2_12[69],stage2_11[89]}
   );
   gpc2135_5 gpc4932 (
      {stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101], stage1_12[102]},
      {stage1_13[213], stage1_13[214], stage1_13[215]},
      {stage1_14[1]},
      {stage1_15[0], stage1_15[1]},
      {stage2_16[0],stage2_15[36],stage2_14[49],stage2_13[52],stage2_12[70]}
   );
   gpc606_5 gpc4933 (
      {stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107], stage1_12[108]},
      {stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage2_16[1],stage2_15[37],stage2_14[50],stage2_13[53],stage2_12[71]}
   );
   gpc606_5 gpc4934 (
      {stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113], stage1_12[114]},
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage2_16[2],stage2_15[38],stage2_14[51],stage2_13[54],stage2_12[72]}
   );
   gpc606_5 gpc4935 (
      {stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119], stage1_12[120]},
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18], stage1_14[19]},
      {stage2_16[3],stage2_15[39],stage2_14[52],stage2_13[55],stage2_12[73]}
   );
   gpc606_5 gpc4936 (
      {stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125], stage1_12[126]},
      {stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage2_16[4],stage2_15[40],stage2_14[53],stage2_13[56],stage2_12[74]}
   );
   gpc606_5 gpc4937 (
      {stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131], stage1_12[132]},
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31]},
      {stage2_16[5],stage2_15[41],stage2_14[54],stage2_13[57],stage2_12[75]}
   );
   gpc606_5 gpc4938 (
      {stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137], stage1_12[138]},
      {stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37]},
      {stage2_16[6],stage2_15[42],stage2_14[55],stage2_13[58],stage2_12[76]}
   );
   gpc606_5 gpc4939 (
      {stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143], stage1_12[144]},
      {stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42], stage1_14[43]},
      {stage2_16[7],stage2_15[43],stage2_14[56],stage2_13[59],stage2_12[77]}
   );
   gpc606_5 gpc4940 (
      {stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149], stage1_12[150]},
      {stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48], stage1_14[49]},
      {stage2_16[8],stage2_15[44],stage2_14[57],stage2_13[60],stage2_12[78]}
   );
   gpc606_5 gpc4941 (
      {stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154], stage1_12[155], stage1_12[156]},
      {stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54], stage1_14[55]},
      {stage2_16[9],stage2_15[45],stage2_14[58],stage2_13[61],stage2_12[79]}
   );
   gpc606_5 gpc4942 (
      {stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162]},
      {stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59], stage1_14[60], stage1_14[61]},
      {stage2_16[10],stage2_15[46],stage2_14[59],stage2_13[62],stage2_12[80]}
   );
   gpc606_5 gpc4943 (
      {stage1_13[216], stage1_13[217], stage1_13[218], stage1_13[219], stage1_13[220], stage1_13[221]},
      {stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7]},
      {stage2_17[0],stage2_16[11],stage2_15[47],stage2_14[60],stage2_13[63]}
   );
   gpc606_5 gpc4944 (
      {stage1_13[222], stage1_13[223], stage1_13[224], stage1_13[225], stage1_13[226], stage1_13[227]},
      {stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11], stage1_15[12], stage1_15[13]},
      {stage2_17[1],stage2_16[12],stage2_15[48],stage2_14[61],stage2_13[64]}
   );
   gpc606_5 gpc4945 (
      {stage1_13[228], stage1_13[229], stage1_13[230], stage1_13[231], stage1_13[232], stage1_13[233]},
      {stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19]},
      {stage2_17[2],stage2_16[13],stage2_15[49],stage2_14[62],stage2_13[65]}
   );
   gpc606_5 gpc4946 (
      {stage1_13[234], stage1_13[235], stage1_13[236], stage1_13[237], stage1_13[238], stage1_13[239]},
      {stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25]},
      {stage2_17[3],stage2_16[14],stage2_15[50],stage2_14[63],stage2_13[66]}
   );
   gpc606_5 gpc4947 (
      {stage1_13[240], stage1_13[241], stage1_13[242], stage1_13[243], stage1_13[244], stage1_13[245]},
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31]},
      {stage2_17[4],stage2_16[15],stage2_15[51],stage2_14[64],stage2_13[67]}
   );
   gpc606_5 gpc4948 (
      {stage1_13[246], stage1_13[247], stage1_13[248], stage1_13[249], stage1_13[250], stage1_13[251]},
      {stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage2_17[5],stage2_16[16],stage2_15[52],stage2_14[65],stage2_13[68]}
   );
   gpc606_5 gpc4949 (
      {stage1_13[252], stage1_13[253], stage1_13[254], stage1_13[255], stage1_13[256], stage1_13[257]},
      {stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage2_17[6],stage2_16[17],stage2_15[53],stage2_14[66],stage2_13[69]}
   );
   gpc606_5 gpc4950 (
      {stage1_13[258], stage1_13[259], stage1_13[260], stage1_13[261], stage1_13[262], stage1_13[263]},
      {stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48], stage1_15[49]},
      {stage2_17[7],stage2_16[18],stage2_15[54],stage2_14[67],stage2_13[70]}
   );
   gpc606_5 gpc4951 (
      {stage1_13[264], stage1_13[265], stage1_13[266], stage1_13[267], stage1_13[268], stage1_13[269]},
      {stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55]},
      {stage2_17[8],stage2_16[19],stage2_15[55],stage2_14[68],stage2_13[71]}
   );
   gpc606_5 gpc4952 (
      {stage1_13[270], stage1_13[271], stage1_13[272], stage1_13[273], stage1_13[274], stage1_13[275]},
      {stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61]},
      {stage2_17[9],stage2_16[20],stage2_15[56],stage2_14[69],stage2_13[72]}
   );
   gpc606_5 gpc4953 (
      {stage1_13[276], stage1_13[277], stage1_13[278], stage1_13[279], stage1_13[280], stage1_13[281]},
      {stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67]},
      {stage2_17[10],stage2_16[21],stage2_15[57],stage2_14[70],stage2_13[73]}
   );
   gpc606_5 gpc4954 (
      {stage1_13[282], stage1_13[283], stage1_13[284], stage1_13[285], stage1_13[286], stage1_13[287]},
      {stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72], stage1_15[73]},
      {stage2_17[11],stage2_16[22],stage2_15[58],stage2_14[71],stage2_13[74]}
   );
   gpc606_5 gpc4955 (
      {stage1_13[288], stage1_13[289], stage1_13[290], stage1_13[291], stage1_13[292], stage1_13[293]},
      {stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77], stage1_15[78], stage1_15[79]},
      {stage2_17[12],stage2_16[23],stage2_15[59],stage2_14[72],stage2_13[75]}
   );
   gpc606_5 gpc4956 (
      {stage1_13[294], stage1_13[295], stage1_13[296], stage1_13[297], stage1_13[298], stage1_13[299]},
      {stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83], stage1_15[84], stage1_15[85]},
      {stage2_17[13],stage2_16[24],stage2_15[60],stage2_14[73],stage2_13[76]}
   );
   gpc606_5 gpc4957 (
      {stage1_13[300], stage1_13[301], stage1_13[302], stage1_13[303], stage1_13[304], 1'b0},
      {stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89], stage1_15[90], stage1_15[91]},
      {stage2_17[14],stage2_16[25],stage2_15[61],stage2_14[74],stage2_13[77]}
   );
   gpc615_5 gpc4958 (
      {stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65], stage1_14[66]},
      {stage1_15[92]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[15],stage2_16[26],stage2_15[62],stage2_14[75]}
   );
   gpc615_5 gpc4959 (
      {stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage1_15[93]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[16],stage2_16[27],stage2_15[63],stage2_14[76]}
   );
   gpc615_5 gpc4960 (
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76]},
      {stage1_15[94]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[17],stage2_16[28],stage2_15[64],stage2_14[77]}
   );
   gpc615_5 gpc4961 (
      {stage1_14[77], stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81]},
      {stage1_15[95]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[18],stage2_16[29],stage2_15[65],stage2_14[78]}
   );
   gpc615_5 gpc4962 (
      {stage1_14[82], stage1_14[83], stage1_14[84], stage1_14[85], stage1_14[86]},
      {stage1_15[96]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[19],stage2_16[30],stage2_15[66],stage2_14[79]}
   );
   gpc615_5 gpc4963 (
      {stage1_14[87], stage1_14[88], stage1_14[89], stage1_14[90], stage1_14[91]},
      {stage1_15[97]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[20],stage2_16[31],stage2_15[67],stage2_14[80]}
   );
   gpc615_5 gpc4964 (
      {stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95], stage1_14[96]},
      {stage1_15[98]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[21],stage2_16[32],stage2_15[68],stage2_14[81]}
   );
   gpc615_5 gpc4965 (
      {stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage1_15[99]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[22],stage2_16[33],stage2_15[69],stage2_14[82]}
   );
   gpc615_5 gpc4966 (
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106]},
      {stage1_15[100]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[23],stage2_16[34],stage2_15[70],stage2_14[83]}
   );
   gpc615_5 gpc4967 (
      {stage1_14[107], stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111]},
      {stage1_15[101]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[24],stage2_16[35],stage2_15[71],stage2_14[84]}
   );
   gpc615_5 gpc4968 (
      {stage1_14[112], stage1_14[113], stage1_14[114], stage1_14[115], stage1_14[116]},
      {stage1_15[102]},
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage2_18[10],stage2_17[25],stage2_16[36],stage2_15[72],stage2_14[85]}
   );
   gpc615_5 gpc4969 (
      {stage1_14[117], stage1_14[118], stage1_14[119], stage1_14[120], stage1_14[121]},
      {stage1_15[103]},
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage2_18[11],stage2_17[26],stage2_16[37],stage2_15[73],stage2_14[86]}
   );
   gpc615_5 gpc4970 (
      {stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125], stage1_14[126]},
      {stage1_15[104]},
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage2_18[12],stage2_17[27],stage2_16[38],stage2_15[74],stage2_14[87]}
   );
   gpc615_5 gpc4971 (
      {stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage1_15[105]},
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage2_18[13],stage2_17[28],stage2_16[39],stage2_15[75],stage2_14[88]}
   );
   gpc615_5 gpc4972 (
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136]},
      {stage1_15[106]},
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage2_18[14],stage2_17[29],stage2_16[40],stage2_15[76],stage2_14[89]}
   );
   gpc615_5 gpc4973 (
      {stage1_14[137], stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141]},
      {stage1_15[107]},
      {stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95]},
      {stage2_18[15],stage2_17[30],stage2_16[41],stage2_15[77],stage2_14[90]}
   );
   gpc615_5 gpc4974 (
      {stage1_14[142], stage1_14[143], stage1_14[144], stage1_14[145], stage1_14[146]},
      {stage1_15[108]},
      {stage1_16[96], stage1_16[97], stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101]},
      {stage2_18[16],stage2_17[31],stage2_16[42],stage2_15[78],stage2_14[91]}
   );
   gpc615_5 gpc4975 (
      {stage1_14[147], stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151]},
      {stage1_15[109]},
      {stage1_16[102], stage1_16[103], stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107]},
      {stage2_18[17],stage2_17[32],stage2_16[43],stage2_15[79],stage2_14[92]}
   );
   gpc615_5 gpc4976 (
      {stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155], stage1_14[156]},
      {stage1_15[110]},
      {stage1_16[108], stage1_16[109], stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113]},
      {stage2_18[18],stage2_17[33],stage2_16[44],stage2_15[80],stage2_14[93]}
   );
   gpc615_5 gpc4977 (
      {stage1_14[157], stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161]},
      {stage1_15[111]},
      {stage1_16[114], stage1_16[115], stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119]},
      {stage2_18[19],stage2_17[34],stage2_16[45],stage2_15[81],stage2_14[94]}
   );
   gpc615_5 gpc4978 (
      {stage1_14[162], stage1_14[163], stage1_14[164], stage1_14[165], stage1_14[166]},
      {stage1_15[112]},
      {stage1_16[120], stage1_16[121], stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125]},
      {stage2_18[20],stage2_17[35],stage2_16[46],stage2_15[82],stage2_14[95]}
   );
   gpc615_5 gpc4979 (
      {stage1_14[167], stage1_14[168], stage1_14[169], stage1_14[170], stage1_14[171]},
      {stage1_15[113]},
      {stage1_16[126], stage1_16[127], stage1_16[128], stage1_16[129], stage1_16[130], stage1_16[131]},
      {stage2_18[21],stage2_17[36],stage2_16[47],stage2_15[83],stage2_14[96]}
   );
   gpc615_5 gpc4980 (
      {stage1_14[172], stage1_14[173], stage1_14[174], stage1_14[175], stage1_14[176]},
      {stage1_15[114]},
      {stage1_16[132], stage1_16[133], stage1_16[134], stage1_16[135], stage1_16[136], stage1_16[137]},
      {stage2_18[22],stage2_17[37],stage2_16[48],stage2_15[84],stage2_14[97]}
   );
   gpc615_5 gpc4981 (
      {stage1_14[177], stage1_14[178], stage1_14[179], stage1_14[180], stage1_14[181]},
      {stage1_15[115]},
      {stage1_16[138], stage1_16[139], stage1_16[140], stage1_16[141], stage1_16[142], stage1_16[143]},
      {stage2_18[23],stage2_17[38],stage2_16[49],stage2_15[85],stage2_14[98]}
   );
   gpc615_5 gpc4982 (
      {stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185], stage1_14[186]},
      {stage1_15[116]},
      {stage1_16[144], stage1_16[145], stage1_16[146], stage1_16[147], stage1_16[148], stage1_16[149]},
      {stage2_18[24],stage2_17[39],stage2_16[50],stage2_15[86],stage2_14[99]}
   );
   gpc615_5 gpc4983 (
      {stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191]},
      {stage1_15[117]},
      {stage1_16[150], stage1_16[151], stage1_16[152], stage1_16[153], stage1_16[154], stage1_16[155]},
      {stage2_18[25],stage2_17[40],stage2_16[51],stage2_15[87],stage2_14[100]}
   );
   gpc615_5 gpc4984 (
      {stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195], stage1_14[196]},
      {stage1_15[118]},
      {stage1_16[156], stage1_16[157], stage1_16[158], stage1_16[159], stage1_16[160], stage1_16[161]},
      {stage2_18[26],stage2_17[41],stage2_16[52],stage2_15[88],stage2_14[101]}
   );
   gpc615_5 gpc4985 (
      {stage1_14[197], stage1_14[198], stage1_14[199], stage1_14[200], stage1_14[201]},
      {stage1_15[119]},
      {stage1_16[162], stage1_16[163], stage1_16[164], stage1_16[165], stage1_16[166], stage1_16[167]},
      {stage2_18[27],stage2_17[42],stage2_16[53],stage2_15[89],stage2_14[102]}
   );
   gpc615_5 gpc4986 (
      {stage1_14[202], stage1_14[203], stage1_14[204], stage1_14[205], stage1_14[206]},
      {stage1_15[120]},
      {stage1_16[168], stage1_16[169], stage1_16[170], stage1_16[171], stage1_16[172], stage1_16[173]},
      {stage2_18[28],stage2_17[43],stage2_16[54],stage2_15[90],stage2_14[103]}
   );
   gpc615_5 gpc4987 (
      {stage1_14[207], stage1_14[208], stage1_14[209], stage1_14[210], stage1_14[211]},
      {stage1_15[121]},
      {stage1_16[174], stage1_16[175], stage1_16[176], stage1_16[177], stage1_16[178], stage1_16[179]},
      {stage2_18[29],stage2_17[44],stage2_16[55],stage2_15[91],stage2_14[104]}
   );
   gpc615_5 gpc4988 (
      {stage1_14[212], stage1_14[213], stage1_14[214], stage1_14[215], stage1_14[216]},
      {stage1_15[122]},
      {stage1_16[180], stage1_16[181], stage1_16[182], stage1_16[183], stage1_16[184], stage1_16[185]},
      {stage2_18[30],stage2_17[45],stage2_16[56],stage2_15[92],stage2_14[105]}
   );
   gpc606_5 gpc4989 (
      {stage1_16[186], stage1_16[187], stage1_16[188], stage1_16[189], stage1_16[190], stage1_16[191]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[31],stage2_17[46],stage2_16[57]}
   );
   gpc606_5 gpc4990 (
      {stage1_16[192], stage1_16[193], stage1_16[194], stage1_16[195], stage1_16[196], stage1_16[197]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[1],stage2_18[32],stage2_17[47],stage2_16[58]}
   );
   gpc606_5 gpc4991 (
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[33],stage2_17[48]}
   );
   gpc606_5 gpc4992 (
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[34],stage2_17[49]}
   );
   gpc606_5 gpc4993 (
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[35],stage2_17[50]}
   );
   gpc606_5 gpc4994 (
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[5],stage2_19[5],stage2_18[36],stage2_17[51]}
   );
   gpc606_5 gpc4995 (
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[6],stage2_19[6],stage2_18[37],stage2_17[52]}
   );
   gpc606_5 gpc4996 (
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[7],stage2_19[7],stage2_18[38],stage2_17[53]}
   );
   gpc606_5 gpc4997 (
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[8],stage2_19[8],stage2_18[39],stage2_17[54]}
   );
   gpc606_5 gpc4998 (
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[9],stage2_19[9],stage2_18[40],stage2_17[55]}
   );
   gpc606_5 gpc4999 (
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[10],stage2_19[10],stage2_18[41],stage2_17[56]}
   );
   gpc606_5 gpc5000 (
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[11],stage2_19[11],stage2_18[42],stage2_17[57]}
   );
   gpc606_5 gpc5001 (
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[12],stage2_19[12],stage2_18[43],stage2_17[58]}
   );
   gpc606_5 gpc5002 (
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[13],stage2_19[13],stage2_18[44],stage2_17[59]}
   );
   gpc606_5 gpc5003 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[14],stage2_19[14],stage2_18[45],stage2_17[60]}
   );
   gpc606_5 gpc5004 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[15],stage2_19[15],stage2_18[46],stage2_17[61]}
   );
   gpc606_5 gpc5005 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[16],stage2_19[16],stage2_18[47],stage2_17[62]}
   );
   gpc606_5 gpc5006 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[17],stage2_19[17],stage2_18[48],stage2_17[63]}
   );
   gpc606_5 gpc5007 (
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99], stage1_19[100], stage1_19[101]},
      {stage2_21[16],stage2_20[18],stage2_19[18],stage2_18[49],stage2_17[64]}
   );
   gpc606_5 gpc5008 (
      {stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105], stage1_17[106], stage1_17[107]},
      {stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107]},
      {stage2_21[17],stage2_20[19],stage2_19[19],stage2_18[50],stage2_17[65]}
   );
   gpc606_5 gpc5009 (
      {stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111], stage1_17[112], stage1_17[113]},
      {stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage2_21[18],stage2_20[20],stage2_19[20],stage2_18[51],stage2_17[66]}
   );
   gpc606_5 gpc5010 (
      {stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117], stage1_17[118], stage1_17[119]},
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118], stage1_19[119]},
      {stage2_21[19],stage2_20[21],stage2_19[21],stage2_18[52],stage2_17[67]}
   );
   gpc606_5 gpc5011 (
      {stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123], stage1_17[124], stage1_17[125]},
      {stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123], stage1_19[124], stage1_19[125]},
      {stage2_21[20],stage2_20[22],stage2_19[22],stage2_18[53],stage2_17[68]}
   );
   gpc606_5 gpc5012 (
      {stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129], stage1_17[130], stage1_17[131]},
      {stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129], stage1_19[130], stage1_19[131]},
      {stage2_21[21],stage2_20[23],stage2_19[23],stage2_18[54],stage2_17[69]}
   );
   gpc606_5 gpc5013 (
      {stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135], stage1_17[136], stage1_17[137]},
      {stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135], stage1_19[136], stage1_19[137]},
      {stage2_21[22],stage2_20[24],stage2_19[24],stage2_18[55],stage2_17[70]}
   );
   gpc606_5 gpc5014 (
      {stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141], stage1_17[142], stage1_17[143]},
      {stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141], stage1_19[142], stage1_19[143]},
      {stage2_21[23],stage2_20[25],stage2_19[25],stage2_18[56],stage2_17[71]}
   );
   gpc606_5 gpc5015 (
      {stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147], stage1_17[148], stage1_17[149]},
      {stage1_19[144], stage1_19[145], stage1_19[146], stage1_19[147], stage1_19[148], stage1_19[149]},
      {stage2_21[24],stage2_20[26],stage2_19[26],stage2_18[57],stage2_17[72]}
   );
   gpc606_5 gpc5016 (
      {stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153], stage1_17[154], stage1_17[155]},
      {stage1_19[150], stage1_19[151], stage1_19[152], stage1_19[153], stage1_19[154], stage1_19[155]},
      {stage2_21[25],stage2_20[27],stage2_19[27],stage2_18[58],stage2_17[73]}
   );
   gpc606_5 gpc5017 (
      {stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159], stage1_17[160], stage1_17[161]},
      {stage1_19[156], stage1_19[157], stage1_19[158], stage1_19[159], stage1_19[160], stage1_19[161]},
      {stage2_21[26],stage2_20[28],stage2_19[28],stage2_18[59],stage2_17[74]}
   );
   gpc606_5 gpc5018 (
      {stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165], stage1_17[166], stage1_17[167]},
      {stage1_19[162], stage1_19[163], stage1_19[164], stage1_19[165], stage1_19[166], stage1_19[167]},
      {stage2_21[27],stage2_20[29],stage2_19[29],stage2_18[60],stage2_17[75]}
   );
   gpc606_5 gpc5019 (
      {stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171], stage1_17[172], stage1_17[173]},
      {stage1_19[168], stage1_19[169], stage1_19[170], stage1_19[171], stage1_19[172], stage1_19[173]},
      {stage2_21[28],stage2_20[30],stage2_19[30],stage2_18[61],stage2_17[76]}
   );
   gpc606_5 gpc5020 (
      {stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177], stage1_17[178], stage1_17[179]},
      {stage1_19[174], stage1_19[175], stage1_19[176], stage1_19[177], stage1_19[178], stage1_19[179]},
      {stage2_21[29],stage2_20[31],stage2_19[31],stage2_18[62],stage2_17[77]}
   );
   gpc606_5 gpc5021 (
      {stage1_17[180], stage1_17[181], stage1_17[182], stage1_17[183], stage1_17[184], stage1_17[185]},
      {stage1_19[180], stage1_19[181], stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185]},
      {stage2_21[30],stage2_20[32],stage2_19[32],stage2_18[63],stage2_17[78]}
   );
   gpc606_5 gpc5022 (
      {stage1_17[186], stage1_17[187], stage1_17[188], stage1_17[189], stage1_17[190], stage1_17[191]},
      {stage1_19[186], stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190], stage1_19[191]},
      {stage2_21[31],stage2_20[33],stage2_19[33],stage2_18[64],stage2_17[79]}
   );
   gpc606_5 gpc5023 (
      {stage1_17[192], stage1_17[193], stage1_17[194], stage1_17[195], stage1_17[196], stage1_17[197]},
      {stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195], stage1_19[196], stage1_19[197]},
      {stage2_21[32],stage2_20[34],stage2_19[34],stage2_18[65],stage2_17[80]}
   );
   gpc606_5 gpc5024 (
      {stage1_17[198], stage1_17[199], stage1_17[200], stage1_17[201], stage1_17[202], stage1_17[203]},
      {stage1_19[198], stage1_19[199], stage1_19[200], stage1_19[201], stage1_19[202], stage1_19[203]},
      {stage2_21[33],stage2_20[35],stage2_19[35],stage2_18[66],stage2_17[81]}
   );
   gpc606_5 gpc5025 (
      {stage1_17[204], stage1_17[205], stage1_17[206], stage1_17[207], stage1_17[208], stage1_17[209]},
      {stage1_19[204], stage1_19[205], stage1_19[206], stage1_19[207], stage1_19[208], stage1_19[209]},
      {stage2_21[34],stage2_20[36],stage2_19[36],stage2_18[67],stage2_17[82]}
   );
   gpc606_5 gpc5026 (
      {stage1_17[210], stage1_17[211], stage1_17[212], stage1_17[213], stage1_17[214], stage1_17[215]},
      {stage1_19[210], stage1_19[211], stage1_19[212], stage1_19[213], stage1_19[214], stage1_19[215]},
      {stage2_21[35],stage2_20[37],stage2_19[37],stage2_18[68],stage2_17[83]}
   );
   gpc606_5 gpc5027 (
      {stage1_17[216], stage1_17[217], stage1_17[218], stage1_17[219], stage1_17[220], stage1_17[221]},
      {stage1_19[216], stage1_19[217], stage1_19[218], stage1_19[219], stage1_19[220], stage1_19[221]},
      {stage2_21[36],stage2_20[38],stage2_19[38],stage2_18[69],stage2_17[84]}
   );
   gpc606_5 gpc5028 (
      {stage1_17[222], stage1_17[223], stage1_17[224], stage1_17[225], stage1_17[226], stage1_17[227]},
      {stage1_19[222], stage1_19[223], stage1_19[224], stage1_19[225], stage1_19[226], stage1_19[227]},
      {stage2_21[37],stage2_20[39],stage2_19[39],stage2_18[70],stage2_17[85]}
   );
   gpc606_5 gpc5029 (
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[38],stage2_20[40],stage2_19[40],stage2_18[71]}
   );
   gpc606_5 gpc5030 (
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[39],stage2_20[41],stage2_19[41],stage2_18[72]}
   );
   gpc606_5 gpc5031 (
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[40],stage2_20[42],stage2_19[42],stage2_18[73]}
   );
   gpc606_5 gpc5032 (
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[41],stage2_20[43],stage2_19[43],stage2_18[74]}
   );
   gpc606_5 gpc5033 (
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage2_22[4],stage2_21[42],stage2_20[44],stage2_19[44],stage2_18[75]}
   );
   gpc606_5 gpc5034 (
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34], stage1_20[35]},
      {stage2_22[5],stage2_21[43],stage2_20[45],stage2_19[45],stage2_18[76]}
   );
   gpc606_5 gpc5035 (
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40], stage1_20[41]},
      {stage2_22[6],stage2_21[44],stage2_20[46],stage2_19[46],stage2_18[77]}
   );
   gpc606_5 gpc5036 (
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46], stage1_20[47]},
      {stage2_22[7],stage2_21[45],stage2_20[47],stage2_19[47],stage2_18[78]}
   );
   gpc606_5 gpc5037 (
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52], stage1_20[53]},
      {stage2_22[8],stage2_21[46],stage2_20[48],stage2_19[48],stage2_18[79]}
   );
   gpc606_5 gpc5038 (
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58], stage1_20[59]},
      {stage2_22[9],stage2_21[47],stage2_20[49],stage2_19[49],stage2_18[80]}
   );
   gpc606_5 gpc5039 (
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64], stage1_20[65]},
      {stage2_22[10],stage2_21[48],stage2_20[50],stage2_19[50],stage2_18[81]}
   );
   gpc606_5 gpc5040 (
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70], stage1_20[71]},
      {stage2_22[11],stage2_21[49],stage2_20[51],stage2_19[51],stage2_18[82]}
   );
   gpc606_5 gpc5041 (
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88], stage1_18[89]},
      {stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76], stage1_20[77]},
      {stage2_22[12],stage2_21[50],stage2_20[52],stage2_19[52],stage2_18[83]}
   );
   gpc606_5 gpc5042 (
      {stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93], stage1_18[94], stage1_18[95]},
      {stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82], stage1_20[83]},
      {stage2_22[13],stage2_21[51],stage2_20[53],stage2_19[53],stage2_18[84]}
   );
   gpc606_5 gpc5043 (
      {stage1_18[96], stage1_18[97], stage1_18[98], stage1_18[99], stage1_18[100], stage1_18[101]},
      {stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88], stage1_20[89]},
      {stage2_22[14],stage2_21[52],stage2_20[54],stage2_19[54],stage2_18[85]}
   );
   gpc606_5 gpc5044 (
      {stage1_18[102], stage1_18[103], stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107]},
      {stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94], stage1_20[95]},
      {stage2_22[15],stage2_21[53],stage2_20[55],stage2_19[55],stage2_18[86]}
   );
   gpc606_5 gpc5045 (
      {stage1_18[108], stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage1_20[96], stage1_20[97], stage1_20[98], stage1_20[99], stage1_20[100], stage1_20[101]},
      {stage2_22[16],stage2_21[54],stage2_20[56],stage2_19[56],stage2_18[87]}
   );
   gpc606_5 gpc5046 (
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118], stage1_18[119]},
      {stage1_20[102], stage1_20[103], stage1_20[104], stage1_20[105], stage1_20[106], stage1_20[107]},
      {stage2_22[17],stage2_21[55],stage2_20[57],stage2_19[57],stage2_18[88]}
   );
   gpc606_5 gpc5047 (
      {stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123], stage1_18[124], stage1_18[125]},
      {stage1_20[108], stage1_20[109], stage1_20[110], stage1_20[111], stage1_20[112], stage1_20[113]},
      {stage2_22[18],stage2_21[56],stage2_20[58],stage2_19[58],stage2_18[89]}
   );
   gpc606_5 gpc5048 (
      {stage1_18[126], stage1_18[127], stage1_18[128], stage1_18[129], stage1_18[130], stage1_18[131]},
      {stage1_20[114], stage1_20[115], stage1_20[116], stage1_20[117], stage1_20[118], stage1_20[119]},
      {stage2_22[19],stage2_21[57],stage2_20[59],stage2_19[59],stage2_18[90]}
   );
   gpc606_5 gpc5049 (
      {stage1_18[132], stage1_18[133], stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137]},
      {stage1_20[120], stage1_20[121], stage1_20[122], stage1_20[123], stage1_20[124], stage1_20[125]},
      {stage2_22[20],stage2_21[58],stage2_20[60],stage2_19[60],stage2_18[91]}
   );
   gpc606_5 gpc5050 (
      {stage1_18[138], stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage1_20[126], stage1_20[127], stage1_20[128], stage1_20[129], stage1_20[130], stage1_20[131]},
      {stage2_22[21],stage2_21[59],stage2_20[61],stage2_19[61],stage2_18[92]}
   );
   gpc606_5 gpc5051 (
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148], stage1_18[149]},
      {stage1_20[132], stage1_20[133], stage1_20[134], stage1_20[135], stage1_20[136], stage1_20[137]},
      {stage2_22[22],stage2_21[60],stage2_20[62],stage2_19[62],stage2_18[93]}
   );
   gpc606_5 gpc5052 (
      {stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153], stage1_18[154], stage1_18[155]},
      {stage1_20[138], stage1_20[139], stage1_20[140], stage1_20[141], stage1_20[142], stage1_20[143]},
      {stage2_22[23],stage2_21[61],stage2_20[63],stage2_19[63],stage2_18[94]}
   );
   gpc606_5 gpc5053 (
      {stage1_18[156], stage1_18[157], stage1_18[158], stage1_18[159], stage1_18[160], stage1_18[161]},
      {stage1_20[144], stage1_20[145], stage1_20[146], stage1_20[147], stage1_20[148], stage1_20[149]},
      {stage2_22[24],stage2_21[62],stage2_20[64],stage2_19[64],stage2_18[95]}
   );
   gpc606_5 gpc5054 (
      {stage1_18[162], stage1_18[163], stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167]},
      {stage1_20[150], stage1_20[151], stage1_20[152], stage1_20[153], stage1_20[154], stage1_20[155]},
      {stage2_22[25],stage2_21[63],stage2_20[65],stage2_19[65],stage2_18[96]}
   );
   gpc606_5 gpc5055 (
      {stage1_18[168], stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage1_20[156], stage1_20[157], stage1_20[158], stage1_20[159], stage1_20[160], stage1_20[161]},
      {stage2_22[26],stage2_21[64],stage2_20[66],stage2_19[66],stage2_18[97]}
   );
   gpc606_5 gpc5056 (
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178], stage1_18[179]},
      {stage1_20[162], stage1_20[163], stage1_20[164], stage1_20[165], stage1_20[166], stage1_20[167]},
      {stage2_22[27],stage2_21[65],stage2_20[67],stage2_19[67],stage2_18[98]}
   );
   gpc606_5 gpc5057 (
      {stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183], stage1_18[184], stage1_18[185]},
      {stage1_20[168], stage1_20[169], stage1_20[170], stage1_20[171], stage1_20[172], stage1_20[173]},
      {stage2_22[28],stage2_21[66],stage2_20[68],stage2_19[68],stage2_18[99]}
   );
   gpc615_5 gpc5058 (
      {stage1_18[186], stage1_18[187], stage1_18[188], stage1_18[189], stage1_18[190]},
      {stage1_19[228]},
      {stage1_20[174], stage1_20[175], stage1_20[176], stage1_20[177], stage1_20[178], stage1_20[179]},
      {stage2_22[29],stage2_21[67],stage2_20[69],stage2_19[69],stage2_18[100]}
   );
   gpc615_5 gpc5059 (
      {stage1_19[229], stage1_19[230], stage1_19[231], stage1_19[232], stage1_19[233]},
      {stage1_20[180]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[30],stage2_21[68],stage2_20[70],stage2_19[70]}
   );
   gpc606_5 gpc5060 (
      {stage1_20[181], stage1_20[182], stage1_20[183], stage1_20[184], stage1_20[185], stage1_20[186]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[1],stage2_22[31],stage2_21[69],stage2_20[71]}
   );
   gpc615_5 gpc5061 (
      {stage1_20[187], stage1_20[188], stage1_20[189], stage1_20[190], stage1_20[191]},
      {stage1_21[6]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[2],stage2_22[32],stage2_21[70],stage2_20[72]}
   );
   gpc615_5 gpc5062 (
      {stage1_20[192], stage1_20[193], stage1_20[194], stage1_20[195], stage1_20[196]},
      {stage1_21[7]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[3],stage2_22[33],stage2_21[71],stage2_20[73]}
   );
   gpc615_5 gpc5063 (
      {stage1_20[197], stage1_20[198], stage1_20[199], stage1_20[200], stage1_20[201]},
      {stage1_21[8]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[4],stage2_22[34],stage2_21[72],stage2_20[74]}
   );
   gpc615_5 gpc5064 (
      {stage1_20[202], stage1_20[203], stage1_20[204], stage1_20[205], stage1_20[206]},
      {stage1_21[9]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[5],stage2_22[35],stage2_21[73],stage2_20[75]}
   );
   gpc615_5 gpc5065 (
      {stage1_20[207], stage1_20[208], stage1_20[209], stage1_20[210], stage1_20[211]},
      {stage1_21[10]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[6],stage2_22[36],stage2_21[74],stage2_20[76]}
   );
   gpc615_5 gpc5066 (
      {stage1_20[212], stage1_20[213], stage1_20[214], stage1_20[215], stage1_20[216]},
      {stage1_21[11]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[7],stage2_22[37],stage2_21[75],stage2_20[77]}
   );
   gpc615_5 gpc5067 (
      {stage1_20[217], stage1_20[218], stage1_20[219], stage1_20[220], stage1_20[221]},
      {stage1_21[12]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[8],stage2_22[38],stage2_21[76],stage2_20[78]}
   );
   gpc615_5 gpc5068 (
      {stage1_20[222], stage1_20[223], stage1_20[224], stage1_20[225], stage1_20[226]},
      {stage1_21[13]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[9],stage2_22[39],stage2_21[77],stage2_20[79]}
   );
   gpc615_5 gpc5069 (
      {stage1_20[227], stage1_20[228], stage1_20[229], stage1_20[230], stage1_20[231]},
      {stage1_21[14]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[10],stage2_22[40],stage2_21[78],stage2_20[80]}
   );
   gpc615_5 gpc5070 (
      {stage1_20[232], stage1_20[233], stage1_20[234], stage1_20[235], stage1_20[236]},
      {stage1_21[15]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[11],stage2_22[41],stage2_21[79],stage2_20[81]}
   );
   gpc615_5 gpc5071 (
      {stage1_20[237], stage1_20[238], stage1_20[239], stage1_20[240], stage1_20[241]},
      {stage1_21[16]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[12],stage2_22[42],stage2_21[80],stage2_20[82]}
   );
   gpc615_5 gpc5072 (
      {stage1_20[242], stage1_20[243], stage1_20[244], stage1_20[245], stage1_20[246]},
      {stage1_21[17]},
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage2_24[12],stage2_23[13],stage2_22[43],stage2_21[81],stage2_20[83]}
   );
   gpc615_5 gpc5073 (
      {stage1_20[247], stage1_20[248], stage1_20[249], stage1_20[250], stage1_20[251]},
      {stage1_21[18]},
      {stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage2_24[13],stage2_23[14],stage2_22[44],stage2_21[82],stage2_20[84]}
   );
   gpc615_5 gpc5074 (
      {stage1_20[252], stage1_20[253], stage1_20[254], stage1_20[255], stage1_20[256]},
      {stage1_21[19]},
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88], stage1_22[89]},
      {stage2_24[14],stage2_23[15],stage2_22[45],stage2_21[83],stage2_20[85]}
   );
   gpc615_5 gpc5075 (
      {stage1_20[257], stage1_20[258], stage1_20[259], stage1_20[260], stage1_20[261]},
      {stage1_21[20]},
      {stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93], stage1_22[94], stage1_22[95]},
      {stage2_24[15],stage2_23[16],stage2_22[46],stage2_21[84],stage2_20[86]}
   );
   gpc606_5 gpc5076 (
      {stage1_21[21], stage1_21[22], stage1_21[23], stage1_21[24], stage1_21[25], stage1_21[26]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[16],stage2_23[17],stage2_22[47],stage2_21[85]}
   );
   gpc606_5 gpc5077 (
      {stage1_21[27], stage1_21[28], stage1_21[29], stage1_21[30], stage1_21[31], stage1_21[32]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[17],stage2_23[18],stage2_22[48],stage2_21[86]}
   );
   gpc606_5 gpc5078 (
      {stage1_21[33], stage1_21[34], stage1_21[35], stage1_21[36], stage1_21[37], stage1_21[38]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[18],stage2_23[19],stage2_22[49],stage2_21[87]}
   );
   gpc606_5 gpc5079 (
      {stage1_21[39], stage1_21[40], stage1_21[41], stage1_21[42], stage1_21[43], stage1_21[44]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[19],stage2_23[20],stage2_22[50],stage2_21[88]}
   );
   gpc606_5 gpc5080 (
      {stage1_21[45], stage1_21[46], stage1_21[47], stage1_21[48], stage1_21[49], stage1_21[50]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[20],stage2_23[21],stage2_22[51],stage2_21[89]}
   );
   gpc606_5 gpc5081 (
      {stage1_21[51], stage1_21[52], stage1_21[53], stage1_21[54], stage1_21[55], stage1_21[56]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[21],stage2_23[22],stage2_22[52],stage2_21[90]}
   );
   gpc606_5 gpc5082 (
      {stage1_21[57], stage1_21[58], stage1_21[59], stage1_21[60], stage1_21[61], stage1_21[62]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[22],stage2_23[23],stage2_22[53],stage2_21[91]}
   );
   gpc606_5 gpc5083 (
      {stage1_21[63], stage1_21[64], stage1_21[65], stage1_21[66], stage1_21[67], stage1_21[68]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[23],stage2_23[24],stage2_22[54],stage2_21[92]}
   );
   gpc606_5 gpc5084 (
      {stage1_21[69], stage1_21[70], stage1_21[71], stage1_21[72], stage1_21[73], stage1_21[74]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage2_25[8],stage2_24[24],stage2_23[25],stage2_22[55],stage2_21[93]}
   );
   gpc606_5 gpc5085 (
      {stage1_21[75], stage1_21[76], stage1_21[77], stage1_21[78], stage1_21[79], stage1_21[80]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage2_25[9],stage2_24[25],stage2_23[26],stage2_22[56],stage2_21[94]}
   );
   gpc606_5 gpc5086 (
      {stage1_21[81], stage1_21[82], stage1_21[83], stage1_21[84], stage1_21[85], stage1_21[86]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage2_25[10],stage2_24[26],stage2_23[27],stage2_22[57],stage2_21[95]}
   );
   gpc606_5 gpc5087 (
      {stage1_21[87], stage1_21[88], stage1_21[89], stage1_21[90], stage1_21[91], stage1_21[92]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage2_25[11],stage2_24[27],stage2_23[28],stage2_22[58],stage2_21[96]}
   );
   gpc606_5 gpc5088 (
      {stage1_21[93], stage1_21[94], stage1_21[95], stage1_21[96], stage1_21[97], stage1_21[98]},
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage2_25[12],stage2_24[28],stage2_23[29],stage2_22[59],stage2_21[97]}
   );
   gpc606_5 gpc5089 (
      {stage1_21[99], stage1_21[100], stage1_21[101], stage1_21[102], stage1_21[103], stage1_21[104]},
      {stage1_23[78], stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82], stage1_23[83]},
      {stage2_25[13],stage2_24[29],stage2_23[30],stage2_22[60],stage2_21[98]}
   );
   gpc606_5 gpc5090 (
      {stage1_21[105], stage1_21[106], stage1_21[107], stage1_21[108], stage1_21[109], stage1_21[110]},
      {stage1_23[84], stage1_23[85], stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89]},
      {stage2_25[14],stage2_24[30],stage2_23[31],stage2_22[61],stage2_21[99]}
   );
   gpc606_5 gpc5091 (
      {stage1_21[111], stage1_21[112], stage1_21[113], stage1_21[114], stage1_21[115], stage1_21[116]},
      {stage1_23[90], stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95]},
      {stage2_25[15],stage2_24[31],stage2_23[32],stage2_22[62],stage2_21[100]}
   );
   gpc606_5 gpc5092 (
      {stage1_21[117], stage1_21[118], stage1_21[119], stage1_21[120], stage1_21[121], stage1_21[122]},
      {stage1_23[96], stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101]},
      {stage2_25[16],stage2_24[32],stage2_23[33],stage2_22[63],stage2_21[101]}
   );
   gpc606_5 gpc5093 (
      {stage1_21[123], stage1_21[124], stage1_21[125], stage1_21[126], stage1_21[127], stage1_21[128]},
      {stage1_23[102], stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107]},
      {stage2_25[17],stage2_24[33],stage2_23[34],stage2_22[64],stage2_21[102]}
   );
   gpc615_5 gpc5094 (
      {stage1_21[129], stage1_21[130], stage1_21[131], stage1_21[132], stage1_21[133]},
      {stage1_22[96]},
      {stage1_23[108], stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112], stage1_23[113]},
      {stage2_25[18],stage2_24[34],stage2_23[35],stage2_22[65],stage2_21[103]}
   );
   gpc615_5 gpc5095 (
      {stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137], stage1_21[138]},
      {stage1_22[97]},
      {stage1_23[114], stage1_23[115], stage1_23[116], stage1_23[117], stage1_23[118], stage1_23[119]},
      {stage2_25[19],stage2_24[35],stage2_23[36],stage2_22[66],stage2_21[104]}
   );
   gpc615_5 gpc5096 (
      {stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage1_22[98]},
      {stage1_23[120], stage1_23[121], stage1_23[122], stage1_23[123], stage1_23[124], stage1_23[125]},
      {stage2_25[20],stage2_24[36],stage2_23[37],stage2_22[67],stage2_21[105]}
   );
   gpc615_5 gpc5097 (
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148]},
      {stage1_22[99]},
      {stage1_23[126], stage1_23[127], stage1_23[128], stage1_23[129], stage1_23[130], stage1_23[131]},
      {stage2_25[21],stage2_24[37],stage2_23[38],stage2_22[68],stage2_21[106]}
   );
   gpc615_5 gpc5098 (
      {stage1_21[149], stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153]},
      {stage1_22[100]},
      {stage1_23[132], stage1_23[133], stage1_23[134], stage1_23[135], stage1_23[136], stage1_23[137]},
      {stage2_25[22],stage2_24[38],stage2_23[39],stage2_22[69],stage2_21[107]}
   );
   gpc615_5 gpc5099 (
      {stage1_21[154], stage1_21[155], stage1_21[156], stage1_21[157], stage1_21[158]},
      {stage1_22[101]},
      {stage1_23[138], stage1_23[139], stage1_23[140], stage1_23[141], stage1_23[142], stage1_23[143]},
      {stage2_25[23],stage2_24[39],stage2_23[40],stage2_22[70],stage2_21[108]}
   );
   gpc615_5 gpc5100 (
      {stage1_21[159], stage1_21[160], stage1_21[161], stage1_21[162], stage1_21[163]},
      {stage1_22[102]},
      {stage1_23[144], stage1_23[145], stage1_23[146], stage1_23[147], stage1_23[148], stage1_23[149]},
      {stage2_25[24],stage2_24[40],stage2_23[41],stage2_22[71],stage2_21[109]}
   );
   gpc615_5 gpc5101 (
      {stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167], stage1_21[168]},
      {stage1_22[103]},
      {stage1_23[150], stage1_23[151], stage1_23[152], stage1_23[153], stage1_23[154], stage1_23[155]},
      {stage2_25[25],stage2_24[41],stage2_23[42],stage2_22[72],stage2_21[110]}
   );
   gpc615_5 gpc5102 (
      {stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage1_22[104]},
      {stage1_23[156], stage1_23[157], stage1_23[158], stage1_23[159], stage1_23[160], stage1_23[161]},
      {stage2_25[26],stage2_24[42],stage2_23[43],stage2_22[73],stage2_21[111]}
   );
   gpc615_5 gpc5103 (
      {stage1_22[105], stage1_22[106], stage1_22[107], stage1_22[108], stage1_22[109]},
      {stage1_23[162]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[27],stage2_24[43],stage2_23[44],stage2_22[74]}
   );
   gpc615_5 gpc5104 (
      {stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113], stage1_22[114]},
      {stage1_23[163]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[28],stage2_24[44],stage2_23[45],stage2_22[75]}
   );
   gpc615_5 gpc5105 (
      {stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118], stage1_22[119]},
      {stage1_23[164]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[29],stage2_24[45],stage2_23[46],stage2_22[76]}
   );
   gpc615_5 gpc5106 (
      {stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123], stage1_22[124]},
      {stage1_23[165]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[30],stage2_24[46],stage2_23[47],stage2_22[77]}
   );
   gpc615_5 gpc5107 (
      {stage1_22[125], stage1_22[126], stage1_22[127], stage1_22[128], stage1_22[129]},
      {stage1_23[166]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[31],stage2_24[47],stage2_23[48],stage2_22[78]}
   );
   gpc615_5 gpc5108 (
      {stage1_22[130], stage1_22[131], stage1_22[132], stage1_22[133], stage1_22[134]},
      {stage1_23[167]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[32],stage2_24[48],stage2_23[49],stage2_22[79]}
   );
   gpc615_5 gpc5109 (
      {stage1_22[135], stage1_22[136], stage1_22[137], stage1_22[138], stage1_22[139]},
      {stage1_23[168]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[33],stage2_24[49],stage2_23[50],stage2_22[80]}
   );
   gpc615_5 gpc5110 (
      {stage1_22[140], stage1_22[141], stage1_22[142], stage1_22[143], stage1_22[144]},
      {stage1_23[169]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[34],stage2_24[50],stage2_23[51],stage2_22[81]}
   );
   gpc615_5 gpc5111 (
      {stage1_23[170], stage1_23[171], stage1_23[172], stage1_23[173], stage1_23[174]},
      {stage1_24[48]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[8],stage2_25[35],stage2_24[51],stage2_23[52]}
   );
   gpc615_5 gpc5112 (
      {stage1_23[175], stage1_23[176], stage1_23[177], stage1_23[178], stage1_23[179]},
      {stage1_24[49]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[9],stage2_25[36],stage2_24[52],stage2_23[53]}
   );
   gpc615_5 gpc5113 (
      {stage1_23[180], stage1_23[181], stage1_23[182], stage1_23[183], stage1_23[184]},
      {stage1_24[50]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[10],stage2_25[37],stage2_24[53],stage2_23[54]}
   );
   gpc615_5 gpc5114 (
      {stage1_23[185], stage1_23[186], stage1_23[187], stage1_23[188], stage1_23[189]},
      {stage1_24[51]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[11],stage2_25[38],stage2_24[54],stage2_23[55]}
   );
   gpc615_5 gpc5115 (
      {stage1_23[190], stage1_23[191], stage1_23[192], stage1_23[193], stage1_23[194]},
      {stage1_24[52]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[12],stage2_25[39],stage2_24[55],stage2_23[56]}
   );
   gpc615_5 gpc5116 (
      {stage1_23[195], stage1_23[196], stage1_23[197], stage1_23[198], stage1_23[199]},
      {stage1_24[53]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[13],stage2_25[40],stage2_24[56],stage2_23[57]}
   );
   gpc615_5 gpc5117 (
      {stage1_23[200], stage1_23[201], stage1_23[202], stage1_23[203], stage1_23[204]},
      {stage1_24[54]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[14],stage2_25[41],stage2_24[57],stage2_23[58]}
   );
   gpc615_5 gpc5118 (
      {stage1_23[205], stage1_23[206], stage1_23[207], stage1_23[208], stage1_23[209]},
      {stage1_24[55]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[15],stage2_25[42],stage2_24[58],stage2_23[59]}
   );
   gpc615_5 gpc5119 (
      {stage1_23[210], stage1_23[211], stage1_23[212], stage1_23[213], stage1_23[214]},
      {stage1_24[56]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[16],stage2_25[43],stage2_24[59],stage2_23[60]}
   );
   gpc615_5 gpc5120 (
      {stage1_23[215], stage1_23[216], stage1_23[217], stage1_23[218], stage1_23[219]},
      {stage1_24[57]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[17],stage2_25[44],stage2_24[60],stage2_23[61]}
   );
   gpc615_5 gpc5121 (
      {stage1_23[220], stage1_23[221], stage1_23[222], stage1_23[223], stage1_23[224]},
      {stage1_24[58]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[18],stage2_25[45],stage2_24[61],stage2_23[62]}
   );
   gpc615_5 gpc5122 (
      {stage1_23[225], stage1_23[226], stage1_23[227], stage1_23[228], stage1_23[229]},
      {stage1_24[59]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[19],stage2_25[46],stage2_24[62],stage2_23[63]}
   );
   gpc615_5 gpc5123 (
      {stage1_23[230], stage1_23[231], stage1_23[232], stage1_23[233], stage1_23[234]},
      {stage1_24[60]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[20],stage2_25[47],stage2_24[63],stage2_23[64]}
   );
   gpc615_5 gpc5124 (
      {stage1_23[235], stage1_23[236], stage1_23[237], stage1_23[238], stage1_23[239]},
      {stage1_24[61]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[21],stage2_25[48],stage2_24[64],stage2_23[65]}
   );
   gpc615_5 gpc5125 (
      {stage1_23[240], stage1_23[241], stage1_23[242], stage1_23[243], stage1_23[244]},
      {stage1_24[62]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[22],stage2_25[49],stage2_24[65],stage2_23[66]}
   );
   gpc615_5 gpc5126 (
      {stage1_23[245], stage1_23[246], stage1_23[247], stage1_23[248], stage1_23[249]},
      {stage1_24[63]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[23],stage2_25[50],stage2_24[66],stage2_23[67]}
   );
   gpc615_5 gpc5127 (
      {stage1_23[250], stage1_23[251], stage1_23[252], stage1_23[253], stage1_23[254]},
      {stage1_24[64]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[24],stage2_25[51],stage2_24[67],stage2_23[68]}
   );
   gpc615_5 gpc5128 (
      {stage1_23[255], stage1_23[256], stage1_23[257], stage1_23[258], stage1_23[259]},
      {stage1_24[65]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[25],stage2_25[52],stage2_24[68],stage2_23[69]}
   );
   gpc615_5 gpc5129 (
      {stage1_23[260], stage1_23[261], stage1_23[262], stage1_23[263], stage1_23[264]},
      {stage1_24[66]},
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage2_27[18],stage2_26[26],stage2_25[53],stage2_24[69],stage2_23[70]}
   );
   gpc615_5 gpc5130 (
      {stage1_23[265], stage1_23[266], stage1_23[267], stage1_23[268], stage1_23[269]},
      {stage1_24[67]},
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage2_27[19],stage2_26[27],stage2_25[54],stage2_24[70],stage2_23[71]}
   );
   gpc615_5 gpc5131 (
      {stage1_23[270], stage1_23[271], stage1_23[272], stage1_23[273], stage1_23[274]},
      {stage1_24[68]},
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage2_27[20],stage2_26[28],stage2_25[55],stage2_24[71],stage2_23[72]}
   );
   gpc615_5 gpc5132 (
      {stage1_23[275], stage1_23[276], stage1_23[277], stage1_23[278], stage1_23[279]},
      {stage1_24[69]},
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage2_27[21],stage2_26[29],stage2_25[56],stage2_24[72],stage2_23[73]}
   );
   gpc615_5 gpc5133 (
      {stage1_23[280], stage1_23[281], stage1_23[282], stage1_23[283], stage1_23[284]},
      {stage1_24[70]},
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage2_27[22],stage2_26[30],stage2_25[57],stage2_24[73],stage2_23[74]}
   );
   gpc615_5 gpc5134 (
      {stage1_23[285], stage1_23[286], 1'b0, 1'b0, 1'b0},
      {stage1_24[71]},
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage2_27[23],stage2_26[31],stage2_25[58],stage2_24[74],stage2_23[75]}
   );
   gpc606_5 gpc5135 (
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[24],stage2_26[32],stage2_25[59],stage2_24[75]}
   );
   gpc606_5 gpc5136 (
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[25],stage2_26[33],stage2_25[60],stage2_24[76]}
   );
   gpc606_5 gpc5137 (
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[26],stage2_26[34],stage2_25[61],stage2_24[77]}
   );
   gpc606_5 gpc5138 (
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[27],stage2_26[35],stage2_25[62],stage2_24[78]}
   );
   gpc606_5 gpc5139 (
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[28],stage2_26[36],stage2_25[63],stage2_24[79]}
   );
   gpc606_5 gpc5140 (
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[29],stage2_26[37],stage2_25[64],stage2_24[80]}
   );
   gpc606_5 gpc5141 (
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[30],stage2_26[38],stage2_25[65],stage2_24[81]}
   );
   gpc606_5 gpc5142 (
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[31],stage2_26[39],stage2_25[66],stage2_24[82]}
   );
   gpc606_5 gpc5143 (
      {stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[32],stage2_26[40],stage2_25[67],stage2_24[83]}
   );
   gpc606_5 gpc5144 (
      {stage1_24[126], stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131]},
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage2_28[9],stage2_27[33],stage2_26[41],stage2_25[68],stage2_24[84]}
   );
   gpc606_5 gpc5145 (
      {stage1_24[132], stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137]},
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage2_28[10],stage2_27[34],stage2_26[42],stage2_25[69],stage2_24[85]}
   );
   gpc606_5 gpc5146 (
      {stage1_24[138], stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143]},
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70], stage1_26[71]},
      {stage2_28[11],stage2_27[35],stage2_26[43],stage2_25[70],stage2_24[86]}
   );
   gpc606_5 gpc5147 (
      {stage1_24[144], stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148], stage1_24[149]},
      {stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77]},
      {stage2_28[12],stage2_27[36],stage2_26[44],stage2_25[71],stage2_24[87]}
   );
   gpc606_5 gpc5148 (
      {stage1_24[150], stage1_24[151], stage1_24[152], stage1_24[153], stage1_24[154], stage1_24[155]},
      {stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83]},
      {stage2_28[13],stage2_27[37],stage2_26[45],stage2_25[72],stage2_24[88]}
   );
   gpc606_5 gpc5149 (
      {stage1_24[156], stage1_24[157], stage1_24[158], stage1_24[159], stage1_24[160], stage1_24[161]},
      {stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage2_28[14],stage2_27[38],stage2_26[46],stage2_25[73],stage2_24[89]}
   );
   gpc606_5 gpc5150 (
      {stage1_24[162], stage1_24[163], stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167]},
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage2_28[15],stage2_27[39],stage2_26[47],stage2_25[74],stage2_24[90]}
   );
   gpc606_5 gpc5151 (
      {stage1_24[168], stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100], stage1_26[101]},
      {stage2_28[16],stage2_27[40],stage2_26[48],stage2_25[75],stage2_24[91]}
   );
   gpc606_5 gpc5152 (
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178], stage1_24[179]},
      {stage1_26[102], stage1_26[103], stage1_26[104], stage1_26[105], stage1_26[106], stage1_26[107]},
      {stage2_28[17],stage2_27[41],stage2_26[49],stage2_25[76],stage2_24[92]}
   );
   gpc606_5 gpc5153 (
      {stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183], stage1_24[184], stage1_24[185]},
      {stage1_26[108], stage1_26[109], stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113]},
      {stage2_28[18],stage2_27[42],stage2_26[50],stage2_25[77],stage2_24[93]}
   );
   gpc606_5 gpc5154 (
      {stage1_24[186], stage1_24[187], stage1_24[188], stage1_24[189], stage1_24[190], stage1_24[191]},
      {stage1_26[114], stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119]},
      {stage2_28[19],stage2_27[43],stage2_26[51],stage2_25[78],stage2_24[94]}
   );
   gpc606_5 gpc5155 (
      {stage1_24[192], stage1_24[193], stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197]},
      {stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage2_28[20],stage2_27[44],stage2_26[52],stage2_25[79],stage2_24[95]}
   );
   gpc606_5 gpc5156 (
      {stage1_24[198], stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203]},
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130], stage1_26[131]},
      {stage2_28[21],stage2_27[45],stage2_26[53],stage2_25[80],stage2_24[96]}
   );
   gpc606_5 gpc5157 (
      {stage1_24[204], stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208], stage1_24[209]},
      {stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135], stage1_26[136], stage1_26[137]},
      {stage2_28[22],stage2_27[46],stage2_26[54],stage2_25[81],stage2_24[97]}
   );
   gpc207_4 gpc5158 (
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149], stage1_25[150]},
      {stage1_27[0], stage1_27[1]},
      {stage2_28[23],stage2_27[47],stage2_26[55],stage2_25[82]}
   );
   gpc606_5 gpc5159 (
      {stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155], stage1_25[156]},
      {stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5], stage1_27[6], stage1_27[7]},
      {stage2_29[0],stage2_28[24],stage2_27[48],stage2_26[56],stage2_25[83]}
   );
   gpc606_5 gpc5160 (
      {stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161], stage1_25[162]},
      {stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13]},
      {stage2_29[1],stage2_28[25],stage2_27[49],stage2_26[57],stage2_25[84]}
   );
   gpc606_5 gpc5161 (
      {stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167], stage1_25[168]},
      {stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19]},
      {stage2_29[2],stage2_28[26],stage2_27[50],stage2_26[58],stage2_25[85]}
   );
   gpc606_5 gpc5162 (
      {stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173], stage1_25[174]},
      {stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23], stage1_27[24], stage1_27[25]},
      {stage2_29[3],stage2_28[27],stage2_27[51],stage2_26[59],stage2_25[86]}
   );
   gpc615_5 gpc5163 (
      {stage1_26[138], stage1_26[139], stage1_26[140], stage1_26[141], stage1_26[142]},
      {stage1_27[26]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[4],stage2_28[28],stage2_27[52],stage2_26[60]}
   );
   gpc615_5 gpc5164 (
      {stage1_26[143], stage1_26[144], stage1_26[145], stage1_26[146], stage1_26[147]},
      {stage1_27[27]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[5],stage2_28[29],stage2_27[53],stage2_26[61]}
   );
   gpc615_5 gpc5165 (
      {stage1_26[148], stage1_26[149], stage1_26[150], stage1_26[151], stage1_26[152]},
      {stage1_27[28]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[6],stage2_28[30],stage2_27[54],stage2_26[62]}
   );
   gpc615_5 gpc5166 (
      {stage1_26[153], stage1_26[154], stage1_26[155], stage1_26[156], stage1_26[157]},
      {stage1_27[29]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[7],stage2_28[31],stage2_27[55],stage2_26[63]}
   );
   gpc615_5 gpc5167 (
      {stage1_26[158], stage1_26[159], stage1_26[160], stage1_26[161], stage1_26[162]},
      {stage1_27[30]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[8],stage2_28[32],stage2_27[56],stage2_26[64]}
   );
   gpc615_5 gpc5168 (
      {stage1_26[163], stage1_26[164], stage1_26[165], stage1_26[166], stage1_26[167]},
      {stage1_27[31]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[9],stage2_28[33],stage2_27[57],stage2_26[65]}
   );
   gpc615_5 gpc5169 (
      {stage1_26[168], stage1_26[169], stage1_26[170], stage1_26[171], stage1_26[172]},
      {stage1_27[32]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[10],stage2_28[34],stage2_27[58],stage2_26[66]}
   );
   gpc615_5 gpc5170 (
      {stage1_26[173], stage1_26[174], stage1_26[175], stage1_26[176], stage1_26[177]},
      {stage1_27[33]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[11],stage2_28[35],stage2_27[59],stage2_26[67]}
   );
   gpc615_5 gpc5171 (
      {stage1_26[178], stage1_26[179], stage1_26[180], stage1_26[181], stage1_26[182]},
      {stage1_27[34]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[12],stage2_28[36],stage2_27[60],stage2_26[68]}
   );
   gpc615_5 gpc5172 (
      {stage1_26[183], stage1_26[184], stage1_26[185], stage1_26[186], stage1_26[187]},
      {stage1_27[35]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[13],stage2_28[37],stage2_27[61],stage2_26[69]}
   );
   gpc615_5 gpc5173 (
      {stage1_26[188], stage1_26[189], stage1_26[190], stage1_26[191], stage1_26[192]},
      {stage1_27[36]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[14],stage2_28[38],stage2_27[62],stage2_26[70]}
   );
   gpc615_5 gpc5174 (
      {stage1_26[193], stage1_26[194], stage1_26[195], stage1_26[196], stage1_26[197]},
      {stage1_27[37]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[15],stage2_28[39],stage2_27[63],stage2_26[71]}
   );
   gpc615_5 gpc5175 (
      {stage1_26[198], stage1_26[199], stage1_26[200], stage1_26[201], stage1_26[202]},
      {stage1_27[38]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[16],stage2_28[40],stage2_27[64],stage2_26[72]}
   );
   gpc615_5 gpc5176 (
      {stage1_26[203], stage1_26[204], stage1_26[205], stage1_26[206], stage1_26[207]},
      {stage1_27[39]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[17],stage2_28[41],stage2_27[65],stage2_26[73]}
   );
   gpc615_5 gpc5177 (
      {stage1_26[208], stage1_26[209], stage1_26[210], stage1_26[211], stage1_26[212]},
      {stage1_27[40]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[18],stage2_28[42],stage2_27[66],stage2_26[74]}
   );
   gpc615_5 gpc5178 (
      {stage1_26[213], stage1_26[214], stage1_26[215], stage1_26[216], stage1_26[217]},
      {stage1_27[41]},
      {stage1_28[90], stage1_28[91], stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95]},
      {stage2_30[15],stage2_29[19],stage2_28[43],stage2_27[67],stage2_26[75]}
   );
   gpc615_5 gpc5179 (
      {stage1_26[218], stage1_26[219], stage1_26[220], stage1_26[221], stage1_26[222]},
      {stage1_27[42]},
      {stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101]},
      {stage2_30[16],stage2_29[20],stage2_28[44],stage2_27[68],stage2_26[76]}
   );
   gpc615_5 gpc5180 (
      {stage1_26[223], stage1_26[224], stage1_26[225], stage1_26[226], stage1_26[227]},
      {stage1_27[43]},
      {stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106], stage1_28[107]},
      {stage2_30[17],stage2_29[21],stage2_28[45],stage2_27[69],stage2_26[77]}
   );
   gpc615_5 gpc5181 (
      {stage1_26[228], stage1_26[229], stage1_26[230], stage1_26[231], stage1_26[232]},
      {stage1_27[44]},
      {stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112], stage1_28[113]},
      {stage2_30[18],stage2_29[22],stage2_28[46],stage2_27[70],stage2_26[78]}
   );
   gpc615_5 gpc5182 (
      {stage1_26[233], stage1_26[234], stage1_26[235], stage1_26[236], stage1_26[237]},
      {stage1_27[45]},
      {stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118], stage1_28[119]},
      {stage2_30[19],stage2_29[23],stage2_28[47],stage2_27[71],stage2_26[79]}
   );
   gpc615_5 gpc5183 (
      {stage1_26[238], stage1_26[239], stage1_26[240], stage1_26[241], stage1_26[242]},
      {stage1_27[46]},
      {stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124], stage1_28[125]},
      {stage2_30[20],stage2_29[24],stage2_28[48],stage2_27[72],stage2_26[80]}
   );
   gpc615_5 gpc5184 (
      {stage1_26[243], stage1_26[244], stage1_26[245], stage1_26[246], stage1_26[247]},
      {stage1_27[47]},
      {stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130], stage1_28[131]},
      {stage2_30[21],stage2_29[25],stage2_28[49],stage2_27[73],stage2_26[81]}
   );
   gpc615_5 gpc5185 (
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_28[132]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[22],stage2_29[26],stage2_28[50],stage2_27[74]}
   );
   gpc615_5 gpc5186 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[133]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[23],stage2_29[27],stage2_28[51],stage2_27[75]}
   );
   gpc615_5 gpc5187 (
      {stage1_27[58], stage1_27[59], stage1_27[60], stage1_27[61], stage1_27[62]},
      {stage1_28[134]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[24],stage2_29[28],stage2_28[52],stage2_27[76]}
   );
   gpc615_5 gpc5188 (
      {stage1_27[63], stage1_27[64], stage1_27[65], stage1_27[66], stage1_27[67]},
      {stage1_28[135]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[25],stage2_29[29],stage2_28[53],stage2_27[77]}
   );
   gpc615_5 gpc5189 (
      {stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71], stage1_27[72]},
      {stage1_28[136]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[26],stage2_29[30],stage2_28[54],stage2_27[78]}
   );
   gpc615_5 gpc5190 (
      {stage1_27[73], stage1_27[74], stage1_27[75], stage1_27[76], stage1_27[77]},
      {stage1_28[137]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[27],stage2_29[31],stage2_28[55],stage2_27[79]}
   );
   gpc615_5 gpc5191 (
      {stage1_27[78], stage1_27[79], stage1_27[80], stage1_27[81], stage1_27[82]},
      {stage1_28[138]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[28],stage2_29[32],stage2_28[56],stage2_27[80]}
   );
   gpc615_5 gpc5192 (
      {stage1_27[83], stage1_27[84], stage1_27[85], stage1_27[86], stage1_27[87]},
      {stage1_28[139]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[29],stage2_29[33],stage2_28[57],stage2_27[81]}
   );
   gpc615_5 gpc5193 (
      {stage1_27[88], stage1_27[89], stage1_27[90], stage1_27[91], stage1_27[92]},
      {stage1_28[140]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[30],stage2_29[34],stage2_28[58],stage2_27[82]}
   );
   gpc615_5 gpc5194 (
      {stage1_27[93], stage1_27[94], stage1_27[95], stage1_27[96], stage1_27[97]},
      {stage1_28[141]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[31],stage2_29[35],stage2_28[59],stage2_27[83]}
   );
   gpc615_5 gpc5195 (
      {stage1_27[98], stage1_27[99], stage1_27[100], stage1_27[101], stage1_27[102]},
      {stage1_28[142]},
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage2_31[10],stage2_30[32],stage2_29[36],stage2_28[60],stage2_27[84]}
   );
   gpc615_5 gpc5196 (
      {stage1_27[103], stage1_27[104], stage1_27[105], stage1_27[106], stage1_27[107]},
      {stage1_28[143]},
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage2_31[11],stage2_30[33],stage2_29[37],stage2_28[61],stage2_27[85]}
   );
   gpc615_5 gpc5197 (
      {stage1_27[108], stage1_27[109], stage1_27[110], stage1_27[111], stage1_27[112]},
      {stage1_28[144]},
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage2_31[12],stage2_30[34],stage2_29[38],stage2_28[62],stage2_27[86]}
   );
   gpc615_5 gpc5198 (
      {stage1_27[113], stage1_27[114], stage1_27[115], stage1_27[116], stage1_27[117]},
      {stage1_28[145]},
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage2_31[13],stage2_30[35],stage2_29[39],stage2_28[63],stage2_27[87]}
   );
   gpc615_5 gpc5199 (
      {stage1_27[118], stage1_27[119], stage1_27[120], stage1_27[121], stage1_27[122]},
      {stage1_28[146]},
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage2_31[14],stage2_30[36],stage2_29[40],stage2_28[64],stage2_27[88]}
   );
   gpc615_5 gpc5200 (
      {stage1_27[123], stage1_27[124], stage1_27[125], stage1_27[126], stage1_27[127]},
      {stage1_28[147]},
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage2_31[15],stage2_30[37],stage2_29[41],stage2_28[65],stage2_27[89]}
   );
   gpc615_5 gpc5201 (
      {stage1_27[128], stage1_27[129], stage1_27[130], stage1_27[131], stage1_27[132]},
      {stage1_28[148]},
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage2_31[16],stage2_30[38],stage2_29[42],stage2_28[66],stage2_27[90]}
   );
   gpc615_5 gpc5202 (
      {stage1_27[133], stage1_27[134], stage1_27[135], stage1_27[136], stage1_27[137]},
      {stage1_28[149]},
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage2_31[17],stage2_30[39],stage2_29[43],stage2_28[67],stage2_27[91]}
   );
   gpc615_5 gpc5203 (
      {stage1_27[138], stage1_27[139], stage1_27[140], stage1_27[141], stage1_27[142]},
      {stage1_28[150]},
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage2_31[18],stage2_30[40],stage2_29[44],stage2_28[68],stage2_27[92]}
   );
   gpc615_5 gpc5204 (
      {stage1_27[143], stage1_27[144], stage1_27[145], stage1_27[146], stage1_27[147]},
      {stage1_28[151]},
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage2_31[19],stage2_30[41],stage2_29[45],stage2_28[69],stage2_27[93]}
   );
   gpc615_5 gpc5205 (
      {stage1_27[148], stage1_27[149], stage1_27[150], stage1_27[151], stage1_27[152]},
      {stage1_28[152]},
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage2_31[20],stage2_30[42],stage2_29[46],stage2_28[70],stage2_27[94]}
   );
   gpc615_5 gpc5206 (
      {stage1_27[153], stage1_27[154], stage1_27[155], stage1_27[156], stage1_27[157]},
      {stage1_28[153]},
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage2_31[21],stage2_30[43],stage2_29[47],stage2_28[71],stage2_27[95]}
   );
   gpc615_5 gpc5207 (
      {stage1_27[158], stage1_27[159], stage1_27[160], stage1_27[161], stage1_27[162]},
      {stage1_28[154]},
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage2_31[22],stage2_30[44],stage2_29[48],stage2_28[72],stage2_27[96]}
   );
   gpc615_5 gpc5208 (
      {stage1_27[163], stage1_27[164], stage1_27[165], stage1_27[166], stage1_27[167]},
      {stage1_28[155]},
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage2_31[23],stage2_30[45],stage2_29[49],stage2_28[73],stage2_27[97]}
   );
   gpc615_5 gpc5209 (
      {stage1_27[168], stage1_27[169], stage1_27[170], stage1_27[171], stage1_27[172]},
      {stage1_28[156]},
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage2_31[24],stage2_30[46],stage2_29[50],stage2_28[74],stage2_27[98]}
   );
   gpc615_5 gpc5210 (
      {stage1_27[173], stage1_27[174], stage1_27[175], stage1_27[176], stage1_27[177]},
      {stage1_28[157]},
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage2_31[25],stage2_30[47],stage2_29[51],stage2_28[75],stage2_27[99]}
   );
   gpc615_5 gpc5211 (
      {stage1_27[178], stage1_27[179], stage1_27[180], stage1_27[181], stage1_27[182]},
      {stage1_28[158]},
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage2_31[26],stage2_30[48],stage2_29[52],stage2_28[76],stage2_27[100]}
   );
   gpc615_5 gpc5212 (
      {stage1_27[183], stage1_27[184], stage1_27[185], stage1_27[186], stage1_27[187]},
      {stage1_28[159]},
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage2_31[27],stage2_30[49],stage2_29[53],stage2_28[77],stage2_27[101]}
   );
   gpc615_5 gpc5213 (
      {stage1_27[188], stage1_27[189], stage1_27[190], stage1_27[191], stage1_27[192]},
      {stage1_28[160]},
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage2_31[28],stage2_30[50],stage2_29[54],stage2_28[78],stage2_27[102]}
   );
   gpc615_5 gpc5214 (
      {stage1_27[193], stage1_27[194], stage1_27[195], stage1_27[196], stage1_27[197]},
      {stage1_28[161]},
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage2_31[29],stage2_30[51],stage2_29[55],stage2_28[79],stage2_27[103]}
   );
   gpc615_5 gpc5215 (
      {stage1_27[198], stage1_27[199], stage1_27[200], stage1_27[201], stage1_27[202]},
      {stage1_28[162]},
      {stage1_29[180], stage1_29[181], stage1_29[182], stage1_29[183], stage1_29[184], stage1_29[185]},
      {stage2_31[30],stage2_30[52],stage2_29[56],stage2_28[80],stage2_27[104]}
   );
   gpc615_5 gpc5216 (
      {stage1_27[203], stage1_27[204], stage1_27[205], 1'b0, 1'b0},
      {stage1_28[163]},
      {stage1_29[186], stage1_29[187], stage1_29[188], stage1_29[189], stage1_29[190], stage1_29[191]},
      {stage2_31[31],stage2_30[53],stage2_29[57],stage2_28[81],stage2_27[105]}
   );
   gpc606_5 gpc5217 (
      {stage1_28[164], stage1_28[165], stage1_28[166], stage1_28[167], stage1_28[168], stage1_28[169]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[32],stage2_30[54],stage2_29[58],stage2_28[82]}
   );
   gpc606_5 gpc5218 (
      {stage1_28[170], stage1_28[171], stage1_28[172], stage1_28[173], stage1_28[174], stage1_28[175]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[33],stage2_30[55],stage2_29[59],stage2_28[83]}
   );
   gpc606_5 gpc5219 (
      {stage1_28[176], stage1_28[177], stage1_28[178], stage1_28[179], stage1_28[180], stage1_28[181]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[34],stage2_30[56],stage2_29[60],stage2_28[84]}
   );
   gpc606_5 gpc5220 (
      {stage1_28[182], stage1_28[183], stage1_28[184], stage1_28[185], stage1_28[186], stage1_28[187]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[35],stage2_30[57],stage2_29[61],stage2_28[85]}
   );
   gpc606_5 gpc5221 (
      {stage1_28[188], stage1_28[189], stage1_28[190], stage1_28[191], stage1_28[192], stage1_28[193]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[36],stage2_30[58],stage2_29[62],stage2_28[86]}
   );
   gpc606_5 gpc5222 (
      {stage1_28[194], stage1_28[195], stage1_28[196], stage1_28[197], stage1_28[198], stage1_28[199]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[37],stage2_30[59],stage2_29[63],stage2_28[87]}
   );
   gpc606_5 gpc5223 (
      {stage1_28[200], stage1_28[201], stage1_28[202], stage1_28[203], stage1_28[204], stage1_28[205]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[38],stage2_30[60],stage2_29[64],stage2_28[88]}
   );
   gpc606_5 gpc5224 (
      {stage1_28[206], stage1_28[207], stage1_28[208], stage1_28[209], stage1_28[210], stage1_28[211]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[39],stage2_30[61],stage2_29[65],stage2_28[89]}
   );
   gpc606_5 gpc5225 (
      {stage1_28[212], stage1_28[213], stage1_28[214], stage1_28[215], stage1_28[216], stage1_28[217]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[40],stage2_30[62],stage2_29[66],stage2_28[90]}
   );
   gpc606_5 gpc5226 (
      {stage1_28[218], stage1_28[219], stage1_28[220], stage1_28[221], stage1_28[222], stage1_28[223]},
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage2_32[9],stage2_31[41],stage2_30[63],stage2_29[67],stage2_28[91]}
   );
   gpc1163_5 gpc5227 (
      {stage1_29[192], stage1_29[193], stage1_29[194]},
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_31[0]},
      {stage1_32[0]},
      {stage2_33[0],stage2_32[10],stage2_31[42],stage2_30[64],stage2_29[68]}
   );
   gpc1163_5 gpc5228 (
      {stage1_29[195], stage1_29[196], stage1_29[197]},
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_31[1]},
      {stage1_32[1]},
      {stage2_33[1],stage2_32[11],stage2_31[43],stage2_30[65],stage2_29[69]}
   );
   gpc1163_5 gpc5229 (
      {stage1_29[198], stage1_29[199], stage1_29[200]},
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_31[2]},
      {stage1_32[2]},
      {stage2_33[2],stage2_32[12],stage2_31[44],stage2_30[66],stage2_29[70]}
   );
   gpc1163_5 gpc5230 (
      {stage1_29[201], stage1_29[202], stage1_29[203]},
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_31[3]},
      {stage1_32[3]},
      {stage2_33[3],stage2_32[13],stage2_31[45],stage2_30[67],stage2_29[71]}
   );
   gpc606_5 gpc5231 (
      {stage1_29[204], stage1_29[205], stage1_29[206], stage1_29[207], stage1_29[208], stage1_29[209]},
      {stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9]},
      {stage2_33[4],stage2_32[14],stage2_31[46],stage2_30[68],stage2_29[72]}
   );
   gpc606_5 gpc5232 (
      {stage1_29[210], stage1_29[211], stage1_29[212], stage1_29[213], stage1_29[214], stage1_29[215]},
      {stage1_31[10], stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage2_33[5],stage2_32[15],stage2_31[47],stage2_30[69],stage2_29[73]}
   );
   gpc606_5 gpc5233 (
      {stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87], stage1_30[88], stage1_30[89]},
      {stage1_32[4], stage1_32[5], stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9]},
      {stage2_34[0],stage2_33[6],stage2_32[16],stage2_31[48],stage2_30[70]}
   );
   gpc615_5 gpc5234 (
      {stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93], stage1_30[94]},
      {stage1_31[16]},
      {stage1_32[10], stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15]},
      {stage2_34[1],stage2_33[7],stage2_32[17],stage2_31[49],stage2_30[71]}
   );
   gpc615_5 gpc5235 (
      {stage1_30[95], stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99]},
      {stage1_31[17]},
      {stage1_32[16], stage1_32[17], stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21]},
      {stage2_34[2],stage2_33[8],stage2_32[18],stage2_31[50],stage2_30[72]}
   );
   gpc615_5 gpc5236 (
      {stage1_30[100], stage1_30[101], stage1_30[102], stage1_30[103], stage1_30[104]},
      {stage1_31[18]},
      {stage1_32[22], stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27]},
      {stage2_34[3],stage2_33[9],stage2_32[19],stage2_31[51],stage2_30[73]}
   );
   gpc615_5 gpc5237 (
      {stage1_30[105], stage1_30[106], stage1_30[107], stage1_30[108], stage1_30[109]},
      {stage1_31[19]},
      {stage1_32[28], stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33]},
      {stage2_34[4],stage2_33[10],stage2_32[20],stage2_31[52],stage2_30[74]}
   );
   gpc615_5 gpc5238 (
      {stage1_30[110], stage1_30[111], stage1_30[112], stage1_30[113], stage1_30[114]},
      {stage1_31[20]},
      {stage1_32[34], stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39]},
      {stage2_34[5],stage2_33[11],stage2_32[21],stage2_31[53],stage2_30[75]}
   );
   gpc615_5 gpc5239 (
      {stage1_30[115], stage1_30[116], stage1_30[117], stage1_30[118], stage1_30[119]},
      {stage1_31[21]},
      {stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45]},
      {stage2_34[6],stage2_33[12],stage2_32[22],stage2_31[54],stage2_30[76]}
   );
   gpc615_5 gpc5240 (
      {stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123], stage1_30[124]},
      {stage1_31[22]},
      {stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51]},
      {stage2_34[7],stage2_33[13],stage2_32[23],stage2_31[55],stage2_30[77]}
   );
   gpc615_5 gpc5241 (
      {stage1_30[125], stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129]},
      {stage1_31[23]},
      {stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57]},
      {stage2_34[8],stage2_33[14],stage2_32[24],stage2_31[56],stage2_30[78]}
   );
   gpc615_5 gpc5242 (
      {stage1_30[130], stage1_30[131], stage1_30[132], stage1_30[133], stage1_30[134]},
      {stage1_31[24]},
      {stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63]},
      {stage2_34[9],stage2_33[15],stage2_32[25],stage2_31[57],stage2_30[79]}
   );
   gpc615_5 gpc5243 (
      {stage1_30[135], stage1_30[136], stage1_30[137], stage1_30[138], stage1_30[139]},
      {stage1_31[25]},
      {stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69]},
      {stage2_34[10],stage2_33[16],stage2_32[26],stage2_31[58],stage2_30[80]}
   );
   gpc615_5 gpc5244 (
      {stage1_30[140], stage1_30[141], stage1_30[142], stage1_30[143], stage1_30[144]},
      {stage1_31[26]},
      {stage1_32[70], stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75]},
      {stage2_34[11],stage2_33[17],stage2_32[27],stage2_31[59],stage2_30[81]}
   );
   gpc615_5 gpc5245 (
      {stage1_30[145], stage1_30[146], stage1_30[147], stage1_30[148], stage1_30[149]},
      {stage1_31[27]},
      {stage1_32[76], stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81]},
      {stage2_34[12],stage2_33[18],stage2_32[28],stage2_31[60],stage2_30[82]}
   );
   gpc615_5 gpc5246 (
      {stage1_30[150], stage1_30[151], stage1_30[152], stage1_30[153], stage1_30[154]},
      {stage1_31[28]},
      {stage1_32[82], stage1_32[83], stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87]},
      {stage2_34[13],stage2_33[19],stage2_32[29],stage2_31[61],stage2_30[83]}
   );
   gpc615_5 gpc5247 (
      {stage1_30[155], stage1_30[156], stage1_30[157], stage1_30[158], stage1_30[159]},
      {stage1_31[29]},
      {stage1_32[88], stage1_32[89], stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93]},
      {stage2_34[14],stage2_33[20],stage2_32[30],stage2_31[62],stage2_30[84]}
   );
   gpc1163_5 gpc5248 (
      {stage1_31[30], stage1_31[31], stage1_31[32]},
      {stage1_32[94], stage1_32[95], stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99]},
      {stage1_33[0]},
      {stage1_34[0]},
      {stage2_35[0],stage2_34[15],stage2_33[21],stage2_32[31],stage2_31[63]}
   );
   gpc606_5 gpc5249 (
      {stage1_31[33], stage1_31[34], stage1_31[35], stage1_31[36], stage1_31[37], stage1_31[38]},
      {stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6]},
      {stage2_35[1],stage2_34[16],stage2_33[22],stage2_32[32],stage2_31[64]}
   );
   gpc606_5 gpc5250 (
      {stage1_31[39], stage1_31[40], stage1_31[41], stage1_31[42], stage1_31[43], stage1_31[44]},
      {stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12]},
      {stage2_35[2],stage2_34[17],stage2_33[23],stage2_32[33],stage2_31[65]}
   );
   gpc606_5 gpc5251 (
      {stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49], stage1_31[50]},
      {stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17], stage1_33[18]},
      {stage2_35[3],stage2_34[18],stage2_33[24],stage2_32[34],stage2_31[66]}
   );
   gpc606_5 gpc5252 (
      {stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54], stage1_31[55], stage1_31[56]},
      {stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23], stage1_33[24]},
      {stage2_35[4],stage2_34[19],stage2_33[25],stage2_32[35],stage2_31[67]}
   );
   gpc606_5 gpc5253 (
      {stage1_31[57], stage1_31[58], stage1_31[59], stage1_31[60], stage1_31[61], stage1_31[62]},
      {stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29], stage1_33[30]},
      {stage2_35[5],stage2_34[20],stage2_33[26],stage2_32[36],stage2_31[68]}
   );
   gpc606_5 gpc5254 (
      {stage1_31[63], stage1_31[64], stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68]},
      {stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35], stage1_33[36]},
      {stage2_35[6],stage2_34[21],stage2_33[27],stage2_32[37],stage2_31[69]}
   );
   gpc606_5 gpc5255 (
      {stage1_31[69], stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73], stage1_31[74]},
      {stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41], stage1_33[42]},
      {stage2_35[7],stage2_34[22],stage2_33[28],stage2_32[38],stage2_31[70]}
   );
   gpc606_5 gpc5256 (
      {stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78], stage1_31[79], stage1_31[80]},
      {stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47], stage1_33[48]},
      {stage2_35[8],stage2_34[23],stage2_33[29],stage2_32[39],stage2_31[71]}
   );
   gpc606_5 gpc5257 (
      {stage1_31[81], stage1_31[82], stage1_31[83], stage1_31[84], stage1_31[85], stage1_31[86]},
      {stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53], stage1_33[54]},
      {stage2_35[9],stage2_34[24],stage2_33[30],stage2_32[40],stage2_31[72]}
   );
   gpc606_5 gpc5258 (
      {stage1_31[87], stage1_31[88], stage1_31[89], stage1_31[90], stage1_31[91], stage1_31[92]},
      {stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59], stage1_33[60]},
      {stage2_35[10],stage2_34[25],stage2_33[31],stage2_32[41],stage2_31[73]}
   );
   gpc606_5 gpc5259 (
      {stage1_31[93], stage1_31[94], stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98]},
      {stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65], stage1_33[66]},
      {stage2_35[11],stage2_34[26],stage2_33[32],stage2_32[42],stage2_31[74]}
   );
   gpc606_5 gpc5260 (
      {stage1_31[99], stage1_31[100], stage1_31[101], stage1_31[102], stage1_31[103], stage1_31[104]},
      {stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71], stage1_33[72]},
      {stage2_35[12],stage2_34[27],stage2_33[33],stage2_32[43],stage2_31[75]}
   );
   gpc615_5 gpc5261 (
      {stage1_31[105], stage1_31[106], stage1_31[107], stage1_31[108], stage1_31[109]},
      {stage1_32[100]},
      {stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77], stage1_33[78]},
      {stage2_35[13],stage2_34[28],stage2_33[34],stage2_32[44],stage2_31[76]}
   );
   gpc615_5 gpc5262 (
      {stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113], stage1_31[114]},
      {stage1_32[101]},
      {stage1_33[79], stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83], stage1_33[84]},
      {stage2_35[14],stage2_34[29],stage2_33[35],stage2_32[45],stage2_31[77]}
   );
   gpc615_5 gpc5263 (
      {stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage1_32[102]},
      {stage1_33[85], stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89], stage1_33[90]},
      {stage2_35[15],stage2_34[30],stage2_33[36],stage2_32[46],stage2_31[78]}
   );
   gpc615_5 gpc5264 (
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124]},
      {stage1_32[103]},
      {stage1_33[91], stage1_33[92], stage1_33[93], stage1_33[94], stage1_33[95], stage1_33[96]},
      {stage2_35[16],stage2_34[31],stage2_33[37],stage2_32[47],stage2_31[79]}
   );
   gpc615_5 gpc5265 (
      {stage1_31[125], stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129]},
      {stage1_32[104]},
      {stage1_33[97], stage1_33[98], stage1_33[99], stage1_33[100], stage1_33[101], stage1_33[102]},
      {stage2_35[17],stage2_34[32],stage2_33[38],stage2_32[48],stage2_31[80]}
   );
   gpc615_5 gpc5266 (
      {stage1_31[130], stage1_31[131], stage1_31[132], stage1_31[133], stage1_31[134]},
      {stage1_32[105]},
      {stage1_33[103], stage1_33[104], stage1_33[105], stage1_33[106], stage1_33[107], stage1_33[108]},
      {stage2_35[18],stage2_34[33],stage2_33[39],stage2_32[49],stage2_31[81]}
   );
   gpc615_5 gpc5267 (
      {stage1_31[135], stage1_31[136], stage1_31[137], stage1_31[138], stage1_31[139]},
      {stage1_32[106]},
      {stage1_33[109], stage1_33[110], stage1_33[111], stage1_33[112], stage1_33[113], stage1_33[114]},
      {stage2_35[19],stage2_34[34],stage2_33[40],stage2_32[50],stage2_31[82]}
   );
   gpc615_5 gpc5268 (
      {stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143], stage1_31[144]},
      {stage1_32[107]},
      {stage1_33[115], stage1_33[116], stage1_33[117], stage1_33[118], stage1_33[119], stage1_33[120]},
      {stage2_35[20],stage2_34[35],stage2_33[41],stage2_32[51],stage2_31[83]}
   );
   gpc615_5 gpc5269 (
      {stage1_31[145], stage1_31[146], stage1_31[147], stage1_31[148], stage1_31[149]},
      {stage1_32[108]},
      {stage1_33[121], stage1_33[122], stage1_33[123], stage1_33[124], stage1_33[125], stage1_33[126]},
      {stage2_35[21],stage2_34[36],stage2_33[42],stage2_32[52],stage2_31[84]}
   );
   gpc615_5 gpc5270 (
      {stage1_31[150], stage1_31[151], stage1_31[152], stage1_31[153], stage1_31[154]},
      {stage1_32[109]},
      {stage1_33[127], stage1_33[128], stage1_33[129], stage1_33[130], stage1_33[131], stage1_33[132]},
      {stage2_35[22],stage2_34[37],stage2_33[43],stage2_32[53],stage2_31[85]}
   );
   gpc615_5 gpc5271 (
      {stage1_31[155], stage1_31[156], stage1_31[157], stage1_31[158], stage1_31[159]},
      {stage1_32[110]},
      {stage1_33[133], stage1_33[134], stage1_33[135], stage1_33[136], stage1_33[137], stage1_33[138]},
      {stage2_35[23],stage2_34[38],stage2_33[44],stage2_32[54],stage2_31[86]}
   );
   gpc615_5 gpc5272 (
      {stage1_31[160], stage1_31[161], stage1_31[162], stage1_31[163], stage1_31[164]},
      {stage1_32[111]},
      {stage1_33[139], stage1_33[140], stage1_33[141], stage1_33[142], stage1_33[143], stage1_33[144]},
      {stage2_35[24],stage2_34[39],stage2_33[45],stage2_32[55],stage2_31[87]}
   );
   gpc615_5 gpc5273 (
      {stage1_31[165], stage1_31[166], stage1_31[167], stage1_31[168], stage1_31[169]},
      {stage1_32[112]},
      {stage1_33[145], stage1_33[146], stage1_33[147], stage1_33[148], stage1_33[149], stage1_33[150]},
      {stage2_35[25],stage2_34[40],stage2_33[46],stage2_32[56],stage2_31[88]}
   );
   gpc615_5 gpc5274 (
      {stage1_31[170], stage1_31[171], stage1_31[172], stage1_31[173], stage1_31[174]},
      {stage1_32[113]},
      {stage1_33[151], stage1_33[152], stage1_33[153], stage1_33[154], stage1_33[155], stage1_33[156]},
      {stage2_35[26],stage2_34[41],stage2_33[47],stage2_32[57],stage2_31[89]}
   );
   gpc615_5 gpc5275 (
      {stage1_31[175], stage1_31[176], stage1_31[177], stage1_31[178], stage1_31[179]},
      {stage1_32[114]},
      {stage1_33[157], stage1_33[158], stage1_33[159], stage1_33[160], stage1_33[161], stage1_33[162]},
      {stage2_35[27],stage2_34[42],stage2_33[48],stage2_32[58],stage2_31[90]}
   );
   gpc615_5 gpc5276 (
      {stage1_31[180], stage1_31[181], stage1_31[182], stage1_31[183], stage1_31[184]},
      {stage1_32[115]},
      {stage1_33[163], stage1_33[164], stage1_33[165], stage1_33[166], stage1_33[167], stage1_33[168]},
      {stage2_35[28],stage2_34[43],stage2_33[49],stage2_32[59],stage2_31[91]}
   );
   gpc615_5 gpc5277 (
      {stage1_31[185], stage1_31[186], stage1_31[187], stage1_31[188], stage1_31[189]},
      {stage1_32[116]},
      {stage1_33[169], stage1_33[170], stage1_33[171], stage1_33[172], stage1_33[173], stage1_33[174]},
      {stage2_35[29],stage2_34[44],stage2_33[50],stage2_32[60],stage2_31[92]}
   );
   gpc615_5 gpc5278 (
      {stage1_31[190], stage1_31[191], stage1_31[192], stage1_31[193], stage1_31[194]},
      {stage1_32[117]},
      {stage1_33[175], stage1_33[176], stage1_33[177], stage1_33[178], stage1_33[179], stage1_33[180]},
      {stage2_35[30],stage2_34[45],stage2_33[51],stage2_32[61],stage2_31[93]}
   );
   gpc615_5 gpc5279 (
      {stage1_31[195], stage1_31[196], stage1_31[197], stage1_31[198], stage1_31[199]},
      {stage1_32[118]},
      {stage1_33[181], stage1_33[182], stage1_33[183], stage1_33[184], stage1_33[185], stage1_33[186]},
      {stage2_35[31],stage2_34[46],stage2_33[52],stage2_32[62],stage2_31[94]}
   );
   gpc615_5 gpc5280 (
      {stage1_31[200], stage1_31[201], stage1_31[202], stage1_31[203], stage1_31[204]},
      {stage1_32[119]},
      {stage1_33[187], stage1_33[188], stage1_33[189], stage1_33[190], stage1_33[191], stage1_33[192]},
      {stage2_35[32],stage2_34[47],stage2_33[53],stage2_32[63],stage2_31[95]}
   );
   gpc615_5 gpc5281 (
      {stage1_31[205], stage1_31[206], stage1_31[207], stage1_31[208], stage1_31[209]},
      {stage1_32[120]},
      {stage1_33[193], stage1_33[194], stage1_33[195], stage1_33[196], stage1_33[197], stage1_33[198]},
      {stage2_35[33],stage2_34[48],stage2_33[54],stage2_32[64],stage2_31[96]}
   );
   gpc615_5 gpc5282 (
      {stage1_31[210], stage1_31[211], stage1_31[212], stage1_31[213], stage1_31[214]},
      {stage1_32[121]},
      {stage1_33[199], stage1_33[200], stage1_33[201], stage1_33[202], stage1_33[203], stage1_33[204]},
      {stage2_35[34],stage2_34[49],stage2_33[55],stage2_32[65],stage2_31[97]}
   );
   gpc615_5 gpc5283 (
      {stage1_31[215], stage1_31[216], stage1_31[217], 1'b0, 1'b0},
      {stage1_32[122]},
      {stage1_33[205], stage1_33[206], stage1_33[207], stage1_33[208], stage1_33[209], stage1_33[210]},
      {stage2_35[35],stage2_34[50],stage2_33[56],stage2_32[66],stage2_31[98]}
   );
   gpc606_5 gpc5284 (
      {stage1_32[123], stage1_32[124], stage1_32[125], stage1_32[126], stage1_32[127], stage1_32[128]},
      {stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5], stage1_34[6]},
      {stage2_36[0],stage2_35[36],stage2_34[51],stage2_33[57],stage2_32[67]}
   );
   gpc606_5 gpc5285 (
      {stage1_32[129], stage1_32[130], stage1_32[131], stage1_32[132], stage1_32[133], stage1_32[134]},
      {stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11], stage1_34[12]},
      {stage2_36[1],stage2_35[37],stage2_34[52],stage2_33[58],stage2_32[68]}
   );
   gpc606_5 gpc5286 (
      {stage1_32[135], stage1_32[136], stage1_32[137], stage1_32[138], stage1_32[139], stage1_32[140]},
      {stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17], stage1_34[18]},
      {stage2_36[2],stage2_35[38],stage2_34[53],stage2_33[59],stage2_32[69]}
   );
   gpc606_5 gpc5287 (
      {stage1_32[141], stage1_32[142], stage1_32[143], stage1_32[144], stage1_32[145], stage1_32[146]},
      {stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23], stage1_34[24]},
      {stage2_36[3],stage2_35[39],stage2_34[54],stage2_33[60],stage2_32[70]}
   );
   gpc606_5 gpc5288 (
      {stage1_32[147], stage1_32[148], stage1_32[149], stage1_32[150], stage1_32[151], stage1_32[152]},
      {stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29], stage1_34[30]},
      {stage2_36[4],stage2_35[40],stage2_34[55],stage2_33[61],stage2_32[71]}
   );
   gpc606_5 gpc5289 (
      {stage1_32[153], stage1_32[154], stage1_32[155], stage1_32[156], stage1_32[157], stage1_32[158]},
      {stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35], stage1_34[36]},
      {stage2_36[5],stage2_35[41],stage2_34[56],stage2_33[62],stage2_32[72]}
   );
   gpc606_5 gpc5290 (
      {stage1_32[159], stage1_32[160], stage1_32[161], stage1_32[162], stage1_32[163], stage1_32[164]},
      {stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41], stage1_34[42]},
      {stage2_36[6],stage2_35[42],stage2_34[57],stage2_33[63],stage2_32[73]}
   );
   gpc606_5 gpc5291 (
      {stage1_32[165], stage1_32[166], stage1_32[167], stage1_32[168], stage1_32[169], stage1_32[170]},
      {stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47], stage1_34[48]},
      {stage2_36[7],stage2_35[43],stage2_34[58],stage2_33[64],stage2_32[74]}
   );
   gpc606_5 gpc5292 (
      {stage1_32[171], stage1_32[172], stage1_32[173], stage1_32[174], stage1_32[175], stage1_32[176]},
      {stage1_34[49], stage1_34[50], stage1_34[51], stage1_34[52], stage1_34[53], stage1_34[54]},
      {stage2_36[8],stage2_35[44],stage2_34[59],stage2_33[65],stage2_32[75]}
   );
   gpc606_5 gpc5293 (
      {stage1_32[177], stage1_32[178], stage1_32[179], stage1_32[180], stage1_32[181], stage1_32[182]},
      {stage1_34[55], stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59], stage1_34[60]},
      {stage2_36[9],stage2_35[45],stage2_34[60],stage2_33[66],stage2_32[76]}
   );
   gpc606_5 gpc5294 (
      {stage1_32[183], stage1_32[184], stage1_32[185], stage1_32[186], stage1_32[187], stage1_32[188]},
      {stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65], stage1_34[66]},
      {stage2_36[10],stage2_35[46],stage2_34[61],stage2_33[67],stage2_32[77]}
   );
   gpc2116_5 gpc5295 (
      {stage1_33[211], stage1_33[212], stage1_33[213], stage1_33[214], stage1_33[215], stage1_33[216]},
      {stage1_34[67]},
      {stage1_35[0]},
      {stage1_36[0], stage1_36[1]},
      {stage2_37[0],stage2_36[11],stage2_35[47],stage2_34[62],stage2_33[68]}
   );
   gpc606_5 gpc5296 (
      {stage1_33[217], stage1_33[218], stage1_33[219], stage1_33[220], stage1_33[221], stage1_33[222]},
      {stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5], stage1_35[6]},
      {stage2_37[1],stage2_36[12],stage2_35[48],stage2_34[63],stage2_33[69]}
   );
   gpc606_5 gpc5297 (
      {stage1_33[223], stage1_33[224], stage1_33[225], stage1_33[226], stage1_33[227], stage1_33[228]},
      {stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11], stage1_35[12]},
      {stage2_37[2],stage2_36[13],stage2_35[49],stage2_34[64],stage2_33[70]}
   );
   gpc606_5 gpc5298 (
      {stage1_33[229], stage1_33[230], stage1_33[231], stage1_33[232], stage1_33[233], stage1_33[234]},
      {stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17], stage1_35[18]},
      {stage2_37[3],stage2_36[14],stage2_35[50],stage2_34[65],stage2_33[71]}
   );
   gpc606_5 gpc5299 (
      {stage1_33[235], stage1_33[236], stage1_33[237], stage1_33[238], stage1_33[239], stage1_33[240]},
      {stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23], stage1_35[24]},
      {stage2_37[4],stage2_36[15],stage2_35[51],stage2_34[66],stage2_33[72]}
   );
   gpc606_5 gpc5300 (
      {stage1_33[241], stage1_33[242], stage1_33[243], stage1_33[244], stage1_33[245], stage1_33[246]},
      {stage1_35[25], stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29], stage1_35[30]},
      {stage2_37[5],stage2_36[16],stage2_35[52],stage2_34[67],stage2_33[73]}
   );
   gpc606_5 gpc5301 (
      {stage1_33[247], stage1_33[248], stage1_33[249], stage1_33[250], stage1_33[251], stage1_33[252]},
      {stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35], stage1_35[36]},
      {stage2_37[6],stage2_36[17],stage2_35[53],stage2_34[68],stage2_33[74]}
   );
   gpc606_5 gpc5302 (
      {stage1_33[253], stage1_33[254], stage1_33[255], stage1_33[256], stage1_33[257], stage1_33[258]},
      {stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41], stage1_35[42]},
      {stage2_37[7],stage2_36[18],stage2_35[54],stage2_34[69],stage2_33[75]}
   );
   gpc606_5 gpc5303 (
      {stage1_34[68], stage1_34[69], stage1_34[70], stage1_34[71], stage1_34[72], stage1_34[73]},
      {stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5], stage1_36[6], stage1_36[7]},
      {stage2_38[0],stage2_37[8],stage2_36[19],stage2_35[55],stage2_34[70]}
   );
   gpc606_5 gpc5304 (
      {stage1_34[74], stage1_34[75], stage1_34[76], stage1_34[77], stage1_34[78], stage1_34[79]},
      {stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11], stage1_36[12], stage1_36[13]},
      {stage2_38[1],stage2_37[9],stage2_36[20],stage2_35[56],stage2_34[71]}
   );
   gpc606_5 gpc5305 (
      {stage1_34[80], stage1_34[81], stage1_34[82], stage1_34[83], stage1_34[84], stage1_34[85]},
      {stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17], stage1_36[18], stage1_36[19]},
      {stage2_38[2],stage2_37[10],stage2_36[21],stage2_35[57],stage2_34[72]}
   );
   gpc606_5 gpc5306 (
      {stage1_34[86], stage1_34[87], stage1_34[88], stage1_34[89], stage1_34[90], stage1_34[91]},
      {stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23], stage1_36[24], stage1_36[25]},
      {stage2_38[3],stage2_37[11],stage2_36[22],stage2_35[58],stage2_34[73]}
   );
   gpc606_5 gpc5307 (
      {stage1_34[92], stage1_34[93], stage1_34[94], stage1_34[95], stage1_34[96], stage1_34[97]},
      {stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29], stage1_36[30], stage1_36[31]},
      {stage2_38[4],stage2_37[12],stage2_36[23],stage2_35[59],stage2_34[74]}
   );
   gpc606_5 gpc5308 (
      {stage1_34[98], stage1_34[99], stage1_34[100], stage1_34[101], stage1_34[102], stage1_34[103]},
      {stage1_36[32], stage1_36[33], stage1_36[34], stage1_36[35], stage1_36[36], stage1_36[37]},
      {stage2_38[5],stage2_37[13],stage2_36[24],stage2_35[60],stage2_34[75]}
   );
   gpc606_5 gpc5309 (
      {stage1_34[104], stage1_34[105], stage1_34[106], stage1_34[107], stage1_34[108], stage1_34[109]},
      {stage1_36[38], stage1_36[39], stage1_36[40], stage1_36[41], stage1_36[42], stage1_36[43]},
      {stage2_38[6],stage2_37[14],stage2_36[25],stage2_35[61],stage2_34[76]}
   );
   gpc606_5 gpc5310 (
      {stage1_34[110], stage1_34[111], stage1_34[112], stage1_34[113], stage1_34[114], stage1_34[115]},
      {stage1_36[44], stage1_36[45], stage1_36[46], stage1_36[47], stage1_36[48], stage1_36[49]},
      {stage2_38[7],stage2_37[15],stage2_36[26],stage2_35[62],stage2_34[77]}
   );
   gpc606_5 gpc5311 (
      {stage1_34[116], stage1_34[117], stage1_34[118], stage1_34[119], stage1_34[120], stage1_34[121]},
      {stage1_36[50], stage1_36[51], stage1_36[52], stage1_36[53], stage1_36[54], stage1_36[55]},
      {stage2_38[8],stage2_37[16],stage2_36[27],stage2_35[63],stage2_34[78]}
   );
   gpc606_5 gpc5312 (
      {stage1_34[122], stage1_34[123], stage1_34[124], stage1_34[125], stage1_34[126], stage1_34[127]},
      {stage1_36[56], stage1_36[57], stage1_36[58], stage1_36[59], stage1_36[60], stage1_36[61]},
      {stage2_38[9],stage2_37[17],stage2_36[28],stage2_35[64],stage2_34[79]}
   );
   gpc606_5 gpc5313 (
      {stage1_34[128], stage1_34[129], stage1_34[130], stage1_34[131], stage1_34[132], stage1_34[133]},
      {stage1_36[62], stage1_36[63], stage1_36[64], stage1_36[65], stage1_36[66], stage1_36[67]},
      {stage2_38[10],stage2_37[18],stage2_36[29],stage2_35[65],stage2_34[80]}
   );
   gpc606_5 gpc5314 (
      {stage1_34[134], stage1_34[135], stage1_34[136], stage1_34[137], stage1_34[138], stage1_34[139]},
      {stage1_36[68], stage1_36[69], stage1_36[70], stage1_36[71], stage1_36[72], stage1_36[73]},
      {stage2_38[11],stage2_37[19],stage2_36[30],stage2_35[66],stage2_34[81]}
   );
   gpc615_5 gpc5315 (
      {stage1_35[43], stage1_35[44], stage1_35[45], stage1_35[46], stage1_35[47]},
      {stage1_36[74]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[12],stage2_37[20],stage2_36[31],stage2_35[67]}
   );
   gpc615_5 gpc5316 (
      {stage1_35[48], stage1_35[49], stage1_35[50], stage1_35[51], stage1_35[52]},
      {stage1_36[75]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[13],stage2_37[21],stage2_36[32],stage2_35[68]}
   );
   gpc615_5 gpc5317 (
      {stage1_35[53], stage1_35[54], stage1_35[55], stage1_35[56], stage1_35[57]},
      {stage1_36[76]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[14],stage2_37[22],stage2_36[33],stage2_35[69]}
   );
   gpc615_5 gpc5318 (
      {stage1_35[58], stage1_35[59], stage1_35[60], stage1_35[61], stage1_35[62]},
      {stage1_36[77]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[15],stage2_37[23],stage2_36[34],stage2_35[70]}
   );
   gpc615_5 gpc5319 (
      {stage1_35[63], stage1_35[64], stage1_35[65], stage1_35[66], stage1_35[67]},
      {stage1_36[78]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[16],stage2_37[24],stage2_36[35],stage2_35[71]}
   );
   gpc615_5 gpc5320 (
      {stage1_35[68], stage1_35[69], stage1_35[70], stage1_35[71], stage1_35[72]},
      {stage1_36[79]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[17],stage2_37[25],stage2_36[36],stage2_35[72]}
   );
   gpc615_5 gpc5321 (
      {stage1_35[73], stage1_35[74], stage1_35[75], stage1_35[76], stage1_35[77]},
      {stage1_36[80]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[18],stage2_37[26],stage2_36[37],stage2_35[73]}
   );
   gpc615_5 gpc5322 (
      {stage1_35[78], stage1_35[79], stage1_35[80], stage1_35[81], stage1_35[82]},
      {stage1_36[81]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[19],stage2_37[27],stage2_36[38],stage2_35[74]}
   );
   gpc615_5 gpc5323 (
      {stage1_35[83], stage1_35[84], stage1_35[85], stage1_35[86], stage1_35[87]},
      {stage1_36[82]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage2_39[8],stage2_38[20],stage2_37[28],stage2_36[39],stage2_35[75]}
   );
   gpc615_5 gpc5324 (
      {stage1_35[88], stage1_35[89], stage1_35[90], stage1_35[91], stage1_35[92]},
      {stage1_36[83]},
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58], stage1_37[59]},
      {stage2_39[9],stage2_38[21],stage2_37[29],stage2_36[40],stage2_35[76]}
   );
   gpc615_5 gpc5325 (
      {stage1_35[93], stage1_35[94], stage1_35[95], stage1_35[96], stage1_35[97]},
      {stage1_36[84]},
      {stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63], stage1_37[64], stage1_37[65]},
      {stage2_39[10],stage2_38[22],stage2_37[30],stage2_36[41],stage2_35[77]}
   );
   gpc615_5 gpc5326 (
      {stage1_35[98], stage1_35[99], stage1_35[100], stage1_35[101], stage1_35[102]},
      {stage1_36[85]},
      {stage1_37[66], stage1_37[67], stage1_37[68], stage1_37[69], stage1_37[70], stage1_37[71]},
      {stage2_39[11],stage2_38[23],stage2_37[31],stage2_36[42],stage2_35[78]}
   );
   gpc615_5 gpc5327 (
      {stage1_35[103], stage1_35[104], stage1_35[105], stage1_35[106], stage1_35[107]},
      {stage1_36[86]},
      {stage1_37[72], stage1_37[73], stage1_37[74], stage1_37[75], stage1_37[76], stage1_37[77]},
      {stage2_39[12],stage2_38[24],stage2_37[32],stage2_36[43],stage2_35[79]}
   );
   gpc615_5 gpc5328 (
      {stage1_35[108], stage1_35[109], stage1_35[110], stage1_35[111], stage1_35[112]},
      {stage1_36[87]},
      {stage1_37[78], stage1_37[79], stage1_37[80], stage1_37[81], stage1_37[82], stage1_37[83]},
      {stage2_39[13],stage2_38[25],stage2_37[33],stage2_36[44],stage2_35[80]}
   );
   gpc615_5 gpc5329 (
      {stage1_35[113], stage1_35[114], stage1_35[115], stage1_35[116], stage1_35[117]},
      {stage1_36[88]},
      {stage1_37[84], stage1_37[85], stage1_37[86], stage1_37[87], stage1_37[88], stage1_37[89]},
      {stage2_39[14],stage2_38[26],stage2_37[34],stage2_36[45],stage2_35[81]}
   );
   gpc615_5 gpc5330 (
      {stage1_35[118], stage1_35[119], stage1_35[120], stage1_35[121], stage1_35[122]},
      {stage1_36[89]},
      {stage1_37[90], stage1_37[91], stage1_37[92], stage1_37[93], stage1_37[94], stage1_37[95]},
      {stage2_39[15],stage2_38[27],stage2_37[35],stage2_36[46],stage2_35[82]}
   );
   gpc615_5 gpc5331 (
      {stage1_35[123], stage1_35[124], stage1_35[125], stage1_35[126], stage1_35[127]},
      {stage1_36[90]},
      {stage1_37[96], stage1_37[97], stage1_37[98], stage1_37[99], stage1_37[100], stage1_37[101]},
      {stage2_39[16],stage2_38[28],stage2_37[36],stage2_36[47],stage2_35[83]}
   );
   gpc615_5 gpc5332 (
      {stage1_35[128], stage1_35[129], stage1_35[130], stage1_35[131], stage1_35[132]},
      {stage1_36[91]},
      {stage1_37[102], stage1_37[103], stage1_37[104], stage1_37[105], stage1_37[106], stage1_37[107]},
      {stage2_39[17],stage2_38[29],stage2_37[37],stage2_36[48],stage2_35[84]}
   );
   gpc615_5 gpc5333 (
      {stage1_35[133], stage1_35[134], stage1_35[135], stage1_35[136], stage1_35[137]},
      {stage1_36[92]},
      {stage1_37[108], stage1_37[109], stage1_37[110], stage1_37[111], stage1_37[112], stage1_37[113]},
      {stage2_39[18],stage2_38[30],stage2_37[38],stage2_36[49],stage2_35[85]}
   );
   gpc615_5 gpc5334 (
      {stage1_35[138], stage1_35[139], stage1_35[140], stage1_35[141], stage1_35[142]},
      {stage1_36[93]},
      {stage1_37[114], stage1_37[115], stage1_37[116], stage1_37[117], stage1_37[118], stage1_37[119]},
      {stage2_39[19],stage2_38[31],stage2_37[39],stage2_36[50],stage2_35[86]}
   );
   gpc615_5 gpc5335 (
      {stage1_35[143], stage1_35[144], stage1_35[145], stage1_35[146], stage1_35[147]},
      {stage1_36[94]},
      {stage1_37[120], stage1_37[121], stage1_37[122], stage1_37[123], stage1_37[124], stage1_37[125]},
      {stage2_39[20],stage2_38[32],stage2_37[40],stage2_36[51],stage2_35[87]}
   );
   gpc615_5 gpc5336 (
      {stage1_35[148], stage1_35[149], stage1_35[150], stage1_35[151], stage1_35[152]},
      {stage1_36[95]},
      {stage1_37[126], stage1_37[127], stage1_37[128], stage1_37[129], stage1_37[130], stage1_37[131]},
      {stage2_39[21],stage2_38[33],stage2_37[41],stage2_36[52],stage2_35[88]}
   );
   gpc615_5 gpc5337 (
      {stage1_35[153], stage1_35[154], stage1_35[155], stage1_35[156], stage1_35[157]},
      {stage1_36[96]},
      {stage1_37[132], stage1_37[133], stage1_37[134], stage1_37[135], stage1_37[136], stage1_37[137]},
      {stage2_39[22],stage2_38[34],stage2_37[42],stage2_36[53],stage2_35[89]}
   );
   gpc615_5 gpc5338 (
      {stage1_35[158], stage1_35[159], stage1_35[160], stage1_35[161], stage1_35[162]},
      {stage1_36[97]},
      {stage1_37[138], stage1_37[139], stage1_37[140], stage1_37[141], stage1_37[142], stage1_37[143]},
      {stage2_39[23],stage2_38[35],stage2_37[43],stage2_36[54],stage2_35[90]}
   );
   gpc615_5 gpc5339 (
      {stage1_35[163], stage1_35[164], stage1_35[165], stage1_35[166], stage1_35[167]},
      {stage1_36[98]},
      {stage1_37[144], stage1_37[145], stage1_37[146], stage1_37[147], stage1_37[148], stage1_37[149]},
      {stage2_39[24],stage2_38[36],stage2_37[44],stage2_36[55],stage2_35[91]}
   );
   gpc615_5 gpc5340 (
      {stage1_35[168], stage1_35[169], stage1_35[170], stage1_35[171], stage1_35[172]},
      {stage1_36[99]},
      {stage1_37[150], stage1_37[151], stage1_37[152], stage1_37[153], stage1_37[154], stage1_37[155]},
      {stage2_39[25],stage2_38[37],stage2_37[45],stage2_36[56],stage2_35[92]}
   );
   gpc615_5 gpc5341 (
      {stage1_35[173], stage1_35[174], stage1_35[175], stage1_35[176], stage1_35[177]},
      {stage1_36[100]},
      {stage1_37[156], stage1_37[157], stage1_37[158], stage1_37[159], stage1_37[160], stage1_37[161]},
      {stage2_39[26],stage2_38[38],stage2_37[46],stage2_36[57],stage2_35[93]}
   );
   gpc1406_5 gpc5342 (
      {stage1_36[101], stage1_36[102], stage1_36[103], stage1_36[104], stage1_36[105], stage1_36[106]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[27],stage2_38[39],stage2_37[47],stage2_36[58]}
   );
   gpc606_5 gpc5343 (
      {stage1_36[107], stage1_36[108], stage1_36[109], stage1_36[110], stage1_36[111], stage1_36[112]},
      {stage1_38[4], stage1_38[5], stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9]},
      {stage2_40[1],stage2_39[28],stage2_38[40],stage2_37[48],stage2_36[59]}
   );
   gpc606_5 gpc5344 (
      {stage1_36[113], stage1_36[114], stage1_36[115], stage1_36[116], stage1_36[117], stage1_36[118]},
      {stage1_38[10], stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15]},
      {stage2_40[2],stage2_39[29],stage2_38[41],stage2_37[49],stage2_36[60]}
   );
   gpc606_5 gpc5345 (
      {stage1_36[119], stage1_36[120], stage1_36[121], stage1_36[122], stage1_36[123], stage1_36[124]},
      {stage1_38[16], stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20], stage1_38[21]},
      {stage2_40[3],stage2_39[30],stage2_38[42],stage2_37[50],stage2_36[61]}
   );
   gpc606_5 gpc5346 (
      {stage1_36[125], stage1_36[126], stage1_36[127], stage1_36[128], stage1_36[129], stage1_36[130]},
      {stage1_38[22], stage1_38[23], stage1_38[24], stage1_38[25], stage1_38[26], stage1_38[27]},
      {stage2_40[4],stage2_39[31],stage2_38[43],stage2_37[51],stage2_36[62]}
   );
   gpc606_5 gpc5347 (
      {stage1_36[131], stage1_36[132], stage1_36[133], stage1_36[134], stage1_36[135], stage1_36[136]},
      {stage1_38[28], stage1_38[29], stage1_38[30], stage1_38[31], stage1_38[32], stage1_38[33]},
      {stage2_40[5],stage2_39[32],stage2_38[44],stage2_37[52],stage2_36[63]}
   );
   gpc606_5 gpc5348 (
      {stage1_36[137], stage1_36[138], stage1_36[139], stage1_36[140], stage1_36[141], stage1_36[142]},
      {stage1_38[34], stage1_38[35], stage1_38[36], stage1_38[37], stage1_38[38], stage1_38[39]},
      {stage2_40[6],stage2_39[33],stage2_38[45],stage2_37[53],stage2_36[64]}
   );
   gpc606_5 gpc5349 (
      {stage1_36[143], stage1_36[144], stage1_36[145], stage1_36[146], stage1_36[147], stage1_36[148]},
      {stage1_38[40], stage1_38[41], stage1_38[42], stage1_38[43], stage1_38[44], stage1_38[45]},
      {stage2_40[7],stage2_39[34],stage2_38[46],stage2_37[54],stage2_36[65]}
   );
   gpc606_5 gpc5350 (
      {stage1_36[149], stage1_36[150], stage1_36[151], stage1_36[152], stage1_36[153], stage1_36[154]},
      {stage1_38[46], stage1_38[47], stage1_38[48], stage1_38[49], stage1_38[50], stage1_38[51]},
      {stage2_40[8],stage2_39[35],stage2_38[47],stage2_37[55],stage2_36[66]}
   );
   gpc606_5 gpc5351 (
      {stage1_36[155], stage1_36[156], stage1_36[157], stage1_36[158], stage1_36[159], stage1_36[160]},
      {stage1_38[52], stage1_38[53], stage1_38[54], stage1_38[55], stage1_38[56], stage1_38[57]},
      {stage2_40[9],stage2_39[36],stage2_38[48],stage2_37[56],stage2_36[67]}
   );
   gpc606_5 gpc5352 (
      {stage1_36[161], stage1_36[162], stage1_36[163], stage1_36[164], stage1_36[165], stage1_36[166]},
      {stage1_38[58], stage1_38[59], stage1_38[60], stage1_38[61], stage1_38[62], stage1_38[63]},
      {stage2_40[10],stage2_39[37],stage2_38[49],stage2_37[57],stage2_36[68]}
   );
   gpc606_5 gpc5353 (
      {stage1_36[167], stage1_36[168], stage1_36[169], stage1_36[170], stage1_36[171], stage1_36[172]},
      {stage1_38[64], stage1_38[65], stage1_38[66], stage1_38[67], stage1_38[68], stage1_38[69]},
      {stage2_40[11],stage2_39[38],stage2_38[50],stage2_37[58],stage2_36[69]}
   );
   gpc606_5 gpc5354 (
      {stage1_36[173], stage1_36[174], stage1_36[175], stage1_36[176], stage1_36[177], stage1_36[178]},
      {stage1_38[70], stage1_38[71], stage1_38[72], stage1_38[73], stage1_38[74], stage1_38[75]},
      {stage2_40[12],stage2_39[39],stage2_38[51],stage2_37[59],stage2_36[70]}
   );
   gpc606_5 gpc5355 (
      {stage1_36[179], stage1_36[180], stage1_36[181], stage1_36[182], stage1_36[183], stage1_36[184]},
      {stage1_38[76], stage1_38[77], stage1_38[78], stage1_38[79], stage1_38[80], stage1_38[81]},
      {stage2_40[13],stage2_39[40],stage2_38[52],stage2_37[60],stage2_36[71]}
   );
   gpc606_5 gpc5356 (
      {stage1_36[185], stage1_36[186], stage1_36[187], stage1_36[188], stage1_36[189], stage1_36[190]},
      {stage1_38[82], stage1_38[83], stage1_38[84], stage1_38[85], stage1_38[86], stage1_38[87]},
      {stage2_40[14],stage2_39[41],stage2_38[53],stage2_37[61],stage2_36[72]}
   );
   gpc606_5 gpc5357 (
      {stage1_36[191], stage1_36[192], stage1_36[193], stage1_36[194], stage1_36[195], stage1_36[196]},
      {stage1_38[88], stage1_38[89], stage1_38[90], stage1_38[91], stage1_38[92], stage1_38[93]},
      {stage2_40[15],stage2_39[42],stage2_38[54],stage2_37[62],stage2_36[73]}
   );
   gpc606_5 gpc5358 (
      {stage1_36[197], stage1_36[198], stage1_36[199], stage1_36[200], stage1_36[201], 1'b0},
      {stage1_38[94], stage1_38[95], stage1_38[96], stage1_38[97], stage1_38[98], stage1_38[99]},
      {stage2_40[16],stage2_39[43],stage2_38[55],stage2_37[63],stage2_36[74]}
   );
   gpc606_5 gpc5359 (
      {stage1_37[162], stage1_37[163], stage1_37[164], stage1_37[165], stage1_37[166], stage1_37[167]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[17],stage2_39[44],stage2_38[56],stage2_37[64]}
   );
   gpc606_5 gpc5360 (
      {stage1_37[168], stage1_37[169], stage1_37[170], stage1_37[171], stage1_37[172], stage1_37[173]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[18],stage2_39[45],stage2_38[57],stage2_37[65]}
   );
   gpc606_5 gpc5361 (
      {stage1_37[174], stage1_37[175], stage1_37[176], stage1_37[177], stage1_37[178], stage1_37[179]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[19],stage2_39[46],stage2_38[58],stage2_37[66]}
   );
   gpc606_5 gpc5362 (
      {stage1_37[180], stage1_37[181], stage1_37[182], stage1_37[183], stage1_37[184], stage1_37[185]},
      {stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24]},
      {stage2_41[3],stage2_40[20],stage2_39[47],stage2_38[59],stage2_37[67]}
   );
   gpc606_5 gpc5363 (
      {stage1_37[186], stage1_37[187], stage1_37[188], stage1_37[189], stage1_37[190], stage1_37[191]},
      {stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30]},
      {stage2_41[4],stage2_40[21],stage2_39[48],stage2_38[60],stage2_37[68]}
   );
   gpc606_5 gpc5364 (
      {stage1_37[192], stage1_37[193], stage1_37[194], stage1_37[195], stage1_37[196], stage1_37[197]},
      {stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36]},
      {stage2_41[5],stage2_40[22],stage2_39[49],stage2_38[61],stage2_37[69]}
   );
   gpc606_5 gpc5365 (
      {stage1_37[198], stage1_37[199], stage1_37[200], stage1_37[201], stage1_37[202], stage1_37[203]},
      {stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42]},
      {stage2_41[6],stage2_40[23],stage2_39[50],stage2_38[62],stage2_37[70]}
   );
   gpc606_5 gpc5366 (
      {stage1_37[204], stage1_37[205], stage1_37[206], stage1_37[207], stage1_37[208], stage1_37[209]},
      {stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48]},
      {stage2_41[7],stage2_40[24],stage2_39[51],stage2_38[63],stage2_37[71]}
   );
   gpc606_5 gpc5367 (
      {stage1_37[210], stage1_37[211], stage1_37[212], stage1_37[213], stage1_37[214], stage1_37[215]},
      {stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54]},
      {stage2_41[8],stage2_40[25],stage2_39[52],stage2_38[64],stage2_37[72]}
   );
   gpc606_5 gpc5368 (
      {stage1_37[216], stage1_37[217], stage1_37[218], stage1_37[219], stage1_37[220], stage1_37[221]},
      {stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60]},
      {stage2_41[9],stage2_40[26],stage2_39[53],stage2_38[65],stage2_37[73]}
   );
   gpc606_5 gpc5369 (
      {stage1_37[222], stage1_37[223], stage1_37[224], stage1_37[225], stage1_37[226], stage1_37[227]},
      {stage1_39[61], stage1_39[62], stage1_39[63], stage1_39[64], stage1_39[65], stage1_39[66]},
      {stage2_41[10],stage2_40[27],stage2_39[54],stage2_38[66],stage2_37[74]}
   );
   gpc606_5 gpc5370 (
      {stage1_37[228], stage1_37[229], stage1_37[230], stage1_37[231], stage1_37[232], stage1_37[233]},
      {stage1_39[67], stage1_39[68], stage1_39[69], stage1_39[70], stage1_39[71], stage1_39[72]},
      {stage2_41[11],stage2_40[28],stage2_39[55],stage2_38[67],stage2_37[75]}
   );
   gpc606_5 gpc5371 (
      {stage1_37[234], stage1_37[235], stage1_37[236], stage1_37[237], stage1_37[238], stage1_37[239]},
      {stage1_39[73], stage1_39[74], stage1_39[75], stage1_39[76], stage1_39[77], stage1_39[78]},
      {stage2_41[12],stage2_40[29],stage2_39[56],stage2_38[68],stage2_37[76]}
   );
   gpc606_5 gpc5372 (
      {stage1_37[240], stage1_37[241], stage1_37[242], stage1_37[243], stage1_37[244], stage1_37[245]},
      {stage1_39[79], stage1_39[80], stage1_39[81], stage1_39[82], stage1_39[83], stage1_39[84]},
      {stage2_41[13],stage2_40[30],stage2_39[57],stage2_38[69],stage2_37[77]}
   );
   gpc606_5 gpc5373 (
      {stage1_37[246], stage1_37[247], stage1_37[248], stage1_37[249], stage1_37[250], stage1_37[251]},
      {stage1_39[85], stage1_39[86], stage1_39[87], stage1_39[88], stage1_39[89], stage1_39[90]},
      {stage2_41[14],stage2_40[31],stage2_39[58],stage2_38[70],stage2_37[78]}
   );
   gpc606_5 gpc5374 (
      {stage1_37[252], stage1_37[253], stage1_37[254], stage1_37[255], stage1_37[256], stage1_37[257]},
      {stage1_39[91], stage1_39[92], stage1_39[93], stage1_39[94], stage1_39[95], stage1_39[96]},
      {stage2_41[15],stage2_40[32],stage2_39[59],stage2_38[71],stage2_37[79]}
   );
   gpc606_5 gpc5375 (
      {stage1_37[258], stage1_37[259], stage1_37[260], stage1_37[261], stage1_37[262], stage1_37[263]},
      {stage1_39[97], stage1_39[98], stage1_39[99], stage1_39[100], stage1_39[101], stage1_39[102]},
      {stage2_41[16],stage2_40[33],stage2_39[60],stage2_38[72],stage2_37[80]}
   );
   gpc606_5 gpc5376 (
      {stage1_37[264], stage1_37[265], stage1_37[266], stage1_37[267], stage1_37[268], stage1_37[269]},
      {stage1_39[103], stage1_39[104], stage1_39[105], stage1_39[106], stage1_39[107], stage1_39[108]},
      {stage2_41[17],stage2_40[34],stage2_39[61],stage2_38[73],stage2_37[81]}
   );
   gpc606_5 gpc5377 (
      {stage1_37[270], stage1_37[271], stage1_37[272], stage1_37[273], stage1_37[274], stage1_37[275]},
      {stage1_39[109], stage1_39[110], stage1_39[111], stage1_39[112], stage1_39[113], stage1_39[114]},
      {stage2_41[18],stage2_40[35],stage2_39[62],stage2_38[74],stage2_37[82]}
   );
   gpc606_5 gpc5378 (
      {stage1_37[276], stage1_37[277], stage1_37[278], stage1_37[279], stage1_37[280], stage1_37[281]},
      {stage1_39[115], stage1_39[116], stage1_39[117], stage1_39[118], stage1_39[119], stage1_39[120]},
      {stage2_41[19],stage2_40[36],stage2_39[63],stage2_38[75],stage2_37[83]}
   );
   gpc606_5 gpc5379 (
      {stage1_37[282], stage1_37[283], stage1_37[284], stage1_37[285], stage1_37[286], stage1_37[287]},
      {stage1_39[121], stage1_39[122], stage1_39[123], stage1_39[124], stage1_39[125], stage1_39[126]},
      {stage2_41[20],stage2_40[37],stage2_39[64],stage2_38[76],stage2_37[84]}
   );
   gpc606_5 gpc5380 (
      {stage1_37[288], stage1_37[289], stage1_37[290], stage1_37[291], stage1_37[292], stage1_37[293]},
      {stage1_39[127], stage1_39[128], stage1_39[129], stage1_39[130], stage1_39[131], stage1_39[132]},
      {stage2_41[21],stage2_40[38],stage2_39[65],stage2_38[77],stage2_37[85]}
   );
   gpc606_5 gpc5381 (
      {stage1_37[294], stage1_37[295], stage1_37[296], stage1_37[297], stage1_37[298], stage1_37[299]},
      {stage1_39[133], stage1_39[134], stage1_39[135], stage1_39[136], stage1_39[137], stage1_39[138]},
      {stage2_41[22],stage2_40[39],stage2_39[66],stage2_38[78],stage2_37[86]}
   );
   gpc606_5 gpc5382 (
      {stage1_37[300], stage1_37[301], stage1_37[302], stage1_37[303], stage1_37[304], stage1_37[305]},
      {stage1_39[139], stage1_39[140], stage1_39[141], stage1_39[142], stage1_39[143], stage1_39[144]},
      {stage2_41[23],stage2_40[40],stage2_39[67],stage2_38[79],stage2_37[87]}
   );
   gpc606_5 gpc5383 (
      {stage1_38[100], stage1_38[101], stage1_38[102], stage1_38[103], stage1_38[104], stage1_38[105]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[24],stage2_40[41],stage2_39[68],stage2_38[80]}
   );
   gpc615_5 gpc5384 (
      {stage1_38[106], stage1_38[107], stage1_38[108], stage1_38[109], stage1_38[110]},
      {stage1_39[145]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[25],stage2_40[42],stage2_39[69],stage2_38[81]}
   );
   gpc615_5 gpc5385 (
      {stage1_38[111], stage1_38[112], stage1_38[113], stage1_38[114], stage1_38[115]},
      {stage1_39[146]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[26],stage2_40[43],stage2_39[70],stage2_38[82]}
   );
   gpc615_5 gpc5386 (
      {stage1_38[116], stage1_38[117], stage1_38[118], stage1_38[119], stage1_38[120]},
      {stage1_39[147]},
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage2_42[3],stage2_41[27],stage2_40[44],stage2_39[71],stage2_38[83]}
   );
   gpc615_5 gpc5387 (
      {stage1_38[121], stage1_38[122], stage1_38[123], stage1_38[124], stage1_38[125]},
      {stage1_39[148]},
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage2_42[4],stage2_41[28],stage2_40[45],stage2_39[72],stage2_38[84]}
   );
   gpc615_5 gpc5388 (
      {stage1_38[126], stage1_38[127], stage1_38[128], stage1_38[129], stage1_38[130]},
      {stage1_39[149]},
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage2_42[5],stage2_41[29],stage2_40[46],stage2_39[73],stage2_38[85]}
   );
   gpc615_5 gpc5389 (
      {stage1_38[131], stage1_38[132], stage1_38[133], stage1_38[134], stage1_38[135]},
      {stage1_39[150]},
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage2_42[6],stage2_41[30],stage2_40[47],stage2_39[74],stage2_38[86]}
   );
   gpc615_5 gpc5390 (
      {stage1_38[136], stage1_38[137], stage1_38[138], stage1_38[139], stage1_38[140]},
      {stage1_39[151]},
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage2_42[7],stage2_41[31],stage2_40[48],stage2_39[75],stage2_38[87]}
   );
   gpc615_5 gpc5391 (
      {stage1_38[141], stage1_38[142], stage1_38[143], stage1_38[144], stage1_38[145]},
      {stage1_39[152]},
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage2_42[8],stage2_41[32],stage2_40[49],stage2_39[76],stage2_38[88]}
   );
   gpc615_5 gpc5392 (
      {stage1_38[146], stage1_38[147], stage1_38[148], stage1_38[149], stage1_38[150]},
      {stage1_39[153]},
      {stage1_40[54], stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58], stage1_40[59]},
      {stage2_42[9],stage2_41[33],stage2_40[50],stage2_39[77],stage2_38[89]}
   );
   gpc615_5 gpc5393 (
      {stage1_38[151], stage1_38[152], stage1_38[153], stage1_38[154], stage1_38[155]},
      {stage1_39[154]},
      {stage1_40[60], stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64], stage1_40[65]},
      {stage2_42[10],stage2_41[34],stage2_40[51],stage2_39[78],stage2_38[90]}
   );
   gpc615_5 gpc5394 (
      {stage1_38[156], stage1_38[157], stage1_38[158], stage1_38[159], stage1_38[160]},
      {stage1_39[155]},
      {stage1_40[66], stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70], stage1_40[71]},
      {stage2_42[11],stage2_41[35],stage2_40[52],stage2_39[79],stage2_38[91]}
   );
   gpc615_5 gpc5395 (
      {stage1_38[161], stage1_38[162], stage1_38[163], stage1_38[164], stage1_38[165]},
      {stage1_39[156]},
      {stage1_40[72], stage1_40[73], stage1_40[74], stage1_40[75], stage1_40[76], stage1_40[77]},
      {stage2_42[12],stage2_41[36],stage2_40[53],stage2_39[80],stage2_38[92]}
   );
   gpc615_5 gpc5396 (
      {stage1_38[166], stage1_38[167], stage1_38[168], stage1_38[169], stage1_38[170]},
      {stage1_39[157]},
      {stage1_40[78], stage1_40[79], stage1_40[80], stage1_40[81], stage1_40[82], stage1_40[83]},
      {stage2_42[13],stage2_41[37],stage2_40[54],stage2_39[81],stage2_38[93]}
   );
   gpc615_5 gpc5397 (
      {stage1_38[171], stage1_38[172], stage1_38[173], stage1_38[174], stage1_38[175]},
      {stage1_39[158]},
      {stage1_40[84], stage1_40[85], stage1_40[86], stage1_40[87], stage1_40[88], stage1_40[89]},
      {stage2_42[14],stage2_41[38],stage2_40[55],stage2_39[82],stage2_38[94]}
   );
   gpc615_5 gpc5398 (
      {stage1_38[176], stage1_38[177], stage1_38[178], stage1_38[179], stage1_38[180]},
      {stage1_39[159]},
      {stage1_40[90], stage1_40[91], stage1_40[92], stage1_40[93], stage1_40[94], stage1_40[95]},
      {stage2_42[15],stage2_41[39],stage2_40[56],stage2_39[83],stage2_38[95]}
   );
   gpc615_5 gpc5399 (
      {stage1_38[181], stage1_38[182], stage1_38[183], stage1_38[184], stage1_38[185]},
      {stage1_39[160]},
      {stage1_40[96], stage1_40[97], stage1_40[98], stage1_40[99], stage1_40[100], stage1_40[101]},
      {stage2_42[16],stage2_41[40],stage2_40[57],stage2_39[84],stage2_38[96]}
   );
   gpc615_5 gpc5400 (
      {stage1_38[186], stage1_38[187], stage1_38[188], stage1_38[189], stage1_38[190]},
      {stage1_39[161]},
      {stage1_40[102], stage1_40[103], stage1_40[104], stage1_40[105], stage1_40[106], stage1_40[107]},
      {stage2_42[17],stage2_41[41],stage2_40[58],stage2_39[85],stage2_38[97]}
   );
   gpc615_5 gpc5401 (
      {stage1_38[191], stage1_38[192], stage1_38[193], stage1_38[194], stage1_38[195]},
      {stage1_39[162]},
      {stage1_40[108], stage1_40[109], stage1_40[110], stage1_40[111], stage1_40[112], stage1_40[113]},
      {stage2_42[18],stage2_41[42],stage2_40[59],stage2_39[86],stage2_38[98]}
   );
   gpc615_5 gpc5402 (
      {stage1_38[196], stage1_38[197], stage1_38[198], stage1_38[199], stage1_38[200]},
      {stage1_39[163]},
      {stage1_40[114], stage1_40[115], stage1_40[116], stage1_40[117], stage1_40[118], stage1_40[119]},
      {stage2_42[19],stage2_41[43],stage2_40[60],stage2_39[87],stage2_38[99]}
   );
   gpc615_5 gpc5403 (
      {stage1_38[201], stage1_38[202], stage1_38[203], stage1_38[204], stage1_38[205]},
      {stage1_39[164]},
      {stage1_40[120], stage1_40[121], stage1_40[122], stage1_40[123], stage1_40[124], stage1_40[125]},
      {stage2_42[20],stage2_41[44],stage2_40[61],stage2_39[88],stage2_38[100]}
   );
   gpc615_5 gpc5404 (
      {stage1_38[206], stage1_38[207], stage1_38[208], stage1_38[209], stage1_38[210]},
      {stage1_39[165]},
      {stage1_40[126], stage1_40[127], stage1_40[128], stage1_40[129], stage1_40[130], stage1_40[131]},
      {stage2_42[21],stage2_41[45],stage2_40[62],stage2_39[89],stage2_38[101]}
   );
   gpc615_5 gpc5405 (
      {stage1_38[211], stage1_38[212], stage1_38[213], stage1_38[214], stage1_38[215]},
      {stage1_39[166]},
      {stage1_40[132], stage1_40[133], stage1_40[134], stage1_40[135], stage1_40[136], stage1_40[137]},
      {stage2_42[22],stage2_41[46],stage2_40[63],stage2_39[90],stage2_38[102]}
   );
   gpc615_5 gpc5406 (
      {stage1_38[216], stage1_38[217], stage1_38[218], stage1_38[219], stage1_38[220]},
      {stage1_39[167]},
      {stage1_40[138], stage1_40[139], stage1_40[140], stage1_40[141], stage1_40[142], stage1_40[143]},
      {stage2_42[23],stage2_41[47],stage2_40[64],stage2_39[91],stage2_38[103]}
   );
   gpc615_5 gpc5407 (
      {stage1_38[221], stage1_38[222], stage1_38[223], stage1_38[224], stage1_38[225]},
      {stage1_39[168]},
      {stage1_40[144], stage1_40[145], stage1_40[146], stage1_40[147], stage1_40[148], stage1_40[149]},
      {stage2_42[24],stage2_41[48],stage2_40[65],stage2_39[92],stage2_38[104]}
   );
   gpc615_5 gpc5408 (
      {stage1_38[226], stage1_38[227], stage1_38[228], stage1_38[229], stage1_38[230]},
      {stage1_39[169]},
      {stage1_40[150], stage1_40[151], stage1_40[152], stage1_40[153], stage1_40[154], stage1_40[155]},
      {stage2_42[25],stage2_41[49],stage2_40[66],stage2_39[93],stage2_38[105]}
   );
   gpc606_5 gpc5409 (
      {stage1_40[156], stage1_40[157], stage1_40[158], stage1_40[159], stage1_40[160], stage1_40[161]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[26],stage2_41[50],stage2_40[67]}
   );
   gpc606_5 gpc5410 (
      {stage1_40[162], stage1_40[163], stage1_40[164], stage1_40[165], stage1_40[166], stage1_40[167]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[1],stage2_42[27],stage2_41[51],stage2_40[68]}
   );
   gpc606_5 gpc5411 (
      {stage1_40[168], stage1_40[169], stage1_40[170], stage1_40[171], stage1_40[172], stage1_40[173]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[2],stage2_42[28],stage2_41[52],stage2_40[69]}
   );
   gpc606_5 gpc5412 (
      {stage1_40[174], stage1_40[175], stage1_40[176], stage1_40[177], stage1_40[178], stage1_40[179]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[3],stage2_42[29],stage2_41[53],stage2_40[70]}
   );
   gpc606_5 gpc5413 (
      {stage1_40[180], stage1_40[181], stage1_40[182], stage1_40[183], stage1_40[184], stage1_40[185]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[4],stage2_42[30],stage2_41[54],stage2_40[71]}
   );
   gpc606_5 gpc5414 (
      {stage1_40[186], stage1_40[187], stage1_40[188], stage1_40[189], stage1_40[190], stage1_40[191]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[5],stage2_42[31],stage2_41[55],stage2_40[72]}
   );
   gpc606_5 gpc5415 (
      {stage1_40[192], stage1_40[193], stage1_40[194], stage1_40[195], stage1_40[196], stage1_40[197]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[6],stage2_42[32],stage2_41[56],stage2_40[73]}
   );
   gpc606_5 gpc5416 (
      {stage1_40[198], stage1_40[199], stage1_40[200], stage1_40[201], stage1_40[202], stage1_40[203]},
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage2_44[7],stage2_43[7],stage2_42[33],stage2_41[57],stage2_40[74]}
   );
   gpc606_5 gpc5417 (
      {stage1_40[204], stage1_40[205], stage1_40[206], stage1_40[207], stage1_40[208], stage1_40[209]},
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage2_44[8],stage2_43[8],stage2_42[34],stage2_41[58],stage2_40[75]}
   );
   gpc606_5 gpc5418 (
      {stage1_40[210], stage1_40[211], stage1_40[212], stage1_40[213], stage1_40[214], stage1_40[215]},
      {stage1_42[54], stage1_42[55], stage1_42[56], stage1_42[57], stage1_42[58], stage1_42[59]},
      {stage2_44[9],stage2_43[9],stage2_42[35],stage2_41[59],stage2_40[76]}
   );
   gpc615_5 gpc5419 (
      {stage1_40[216], stage1_40[217], stage1_40[218], stage1_40[219], stage1_40[220]},
      {stage1_41[0]},
      {stage1_42[60], stage1_42[61], stage1_42[62], stage1_42[63], stage1_42[64], stage1_42[65]},
      {stage2_44[10],stage2_43[10],stage2_42[36],stage2_41[60],stage2_40[77]}
   );
   gpc615_5 gpc5420 (
      {stage1_40[221], stage1_40[222], stage1_40[223], stage1_40[224], stage1_40[225]},
      {stage1_41[1]},
      {stage1_42[66], stage1_42[67], stage1_42[68], stage1_42[69], stage1_42[70], stage1_42[71]},
      {stage2_44[11],stage2_43[11],stage2_42[37],stage2_41[61],stage2_40[78]}
   );
   gpc615_5 gpc5421 (
      {stage1_40[226], stage1_40[227], stage1_40[228], stage1_40[229], stage1_40[230]},
      {stage1_41[2]},
      {stage1_42[72], stage1_42[73], stage1_42[74], stage1_42[75], stage1_42[76], stage1_42[77]},
      {stage2_44[12],stage2_43[12],stage2_42[38],stage2_41[62],stage2_40[79]}
   );
   gpc615_5 gpc5422 (
      {stage1_40[231], stage1_40[232], stage1_40[233], stage1_40[234], stage1_40[235]},
      {stage1_41[3]},
      {stage1_42[78], stage1_42[79], stage1_42[80], stage1_42[81], stage1_42[82], stage1_42[83]},
      {stage2_44[13],stage2_43[13],stage2_42[39],stage2_41[63],stage2_40[80]}
   );
   gpc615_5 gpc5423 (
      {stage1_40[236], stage1_40[237], stage1_40[238], stage1_40[239], stage1_40[240]},
      {stage1_41[4]},
      {stage1_42[84], stage1_42[85], stage1_42[86], stage1_42[87], stage1_42[88], stage1_42[89]},
      {stage2_44[14],stage2_43[14],stage2_42[40],stage2_41[64],stage2_40[81]}
   );
   gpc615_5 gpc5424 (
      {stage1_40[241], stage1_40[242], stage1_40[243], stage1_40[244], stage1_40[245]},
      {stage1_41[5]},
      {stage1_42[90], stage1_42[91], stage1_42[92], stage1_42[93], stage1_42[94], stage1_42[95]},
      {stage2_44[15],stage2_43[15],stage2_42[41],stage2_41[65],stage2_40[82]}
   );
   gpc615_5 gpc5425 (
      {stage1_40[246], stage1_40[247], stage1_40[248], stage1_40[249], stage1_40[250]},
      {stage1_41[6]},
      {stage1_42[96], stage1_42[97], stage1_42[98], stage1_42[99], stage1_42[100], stage1_42[101]},
      {stage2_44[16],stage2_43[16],stage2_42[42],stage2_41[66],stage2_40[83]}
   );
   gpc615_5 gpc5426 (
      {stage1_40[251], stage1_40[252], stage1_40[253], stage1_40[254], stage1_40[255]},
      {stage1_41[7]},
      {stage1_42[102], stage1_42[103], stage1_42[104], stage1_42[105], stage1_42[106], stage1_42[107]},
      {stage2_44[17],stage2_43[17],stage2_42[43],stage2_41[67],stage2_40[84]}
   );
   gpc615_5 gpc5427 (
      {stage1_40[256], stage1_40[257], stage1_40[258], stage1_40[259], stage1_40[260]},
      {stage1_41[8]},
      {stage1_42[108], stage1_42[109], stage1_42[110], stage1_42[111], stage1_42[112], stage1_42[113]},
      {stage2_44[18],stage2_43[18],stage2_42[44],stage2_41[68],stage2_40[85]}
   );
   gpc615_5 gpc5428 (
      {stage1_40[261], stage1_40[262], stage1_40[263], stage1_40[264], stage1_40[265]},
      {stage1_41[9]},
      {stage1_42[114], stage1_42[115], stage1_42[116], stage1_42[117], stage1_42[118], stage1_42[119]},
      {stage2_44[19],stage2_43[19],stage2_42[45],stage2_41[69],stage2_40[86]}
   );
   gpc615_5 gpc5429 (
      {stage1_40[266], stage1_40[267], stage1_40[268], stage1_40[269], stage1_40[270]},
      {stage1_41[10]},
      {stage1_42[120], stage1_42[121], stage1_42[122], stage1_42[123], stage1_42[124], stage1_42[125]},
      {stage2_44[20],stage2_43[20],stage2_42[46],stage2_41[70],stage2_40[87]}
   );
   gpc615_5 gpc5430 (
      {stage1_40[271], stage1_40[272], stage1_40[273], stage1_40[274], stage1_40[275]},
      {stage1_41[11]},
      {stage1_42[126], stage1_42[127], stage1_42[128], stage1_42[129], stage1_42[130], stage1_42[131]},
      {stage2_44[21],stage2_43[21],stage2_42[47],stage2_41[71],stage2_40[88]}
   );
   gpc615_5 gpc5431 (
      {stage1_40[276], stage1_40[277], stage1_40[278], stage1_40[279], stage1_40[280]},
      {stage1_41[12]},
      {stage1_42[132], stage1_42[133], stage1_42[134], stage1_42[135], stage1_42[136], stage1_42[137]},
      {stage2_44[22],stage2_43[22],stage2_42[48],stage2_41[72],stage2_40[89]}
   );
   gpc606_5 gpc5432 (
      {stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[23],stage2_43[23],stage2_42[49],stage2_41[73]}
   );
   gpc606_5 gpc5433 (
      {stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23], stage1_41[24]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[24],stage2_43[24],stage2_42[50],stage2_41[74]}
   );
   gpc606_5 gpc5434 (
      {stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29], stage1_41[30]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[25],stage2_43[25],stage2_42[51],stage2_41[75]}
   );
   gpc606_5 gpc5435 (
      {stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35], stage1_41[36]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[26],stage2_43[26],stage2_42[52],stage2_41[76]}
   );
   gpc606_5 gpc5436 (
      {stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41], stage1_41[42]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[27],stage2_43[27],stage2_42[53],stage2_41[77]}
   );
   gpc615_5 gpc5437 (
      {stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage1_42[138]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[28],stage2_43[28],stage2_42[54],stage2_41[78]}
   );
   gpc615_5 gpc5438 (
      {stage1_41[48], stage1_41[49], stage1_41[50], stage1_41[51], stage1_41[52]},
      {stage1_42[139]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[29],stage2_43[29],stage2_42[55],stage2_41[79]}
   );
   gpc615_5 gpc5439 (
      {stage1_41[53], stage1_41[54], stage1_41[55], stage1_41[56], stage1_41[57]},
      {stage1_42[140]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[30],stage2_43[30],stage2_42[56],stage2_41[80]}
   );
   gpc615_5 gpc5440 (
      {stage1_41[58], stage1_41[59], stage1_41[60], stage1_41[61], stage1_41[62]},
      {stage1_42[141]},
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage2_45[8],stage2_44[31],stage2_43[31],stage2_42[57],stage2_41[81]}
   );
   gpc615_5 gpc5441 (
      {stage1_41[63], stage1_41[64], stage1_41[65], stage1_41[66], stage1_41[67]},
      {stage1_42[142]},
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage2_45[9],stage2_44[32],stage2_43[32],stage2_42[58],stage2_41[82]}
   );
   gpc615_5 gpc5442 (
      {stage1_41[68], stage1_41[69], stage1_41[70], stage1_41[71], stage1_41[72]},
      {stage1_42[143]},
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage2_45[10],stage2_44[33],stage2_43[33],stage2_42[59],stage2_41[83]}
   );
   gpc615_5 gpc5443 (
      {stage1_41[73], stage1_41[74], stage1_41[75], stage1_41[76], stage1_41[77]},
      {stage1_42[144]},
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage2_45[11],stage2_44[34],stage2_43[34],stage2_42[60],stage2_41[84]}
   );
   gpc615_5 gpc5444 (
      {stage1_41[78], stage1_41[79], stage1_41[80], stage1_41[81], stage1_41[82]},
      {stage1_42[145]},
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage2_45[12],stage2_44[35],stage2_43[35],stage2_42[61],stage2_41[85]}
   );
   gpc615_5 gpc5445 (
      {stage1_41[83], stage1_41[84], stage1_41[85], stage1_41[86], stage1_41[87]},
      {stage1_42[146]},
      {stage1_43[78], stage1_43[79], stage1_43[80], stage1_43[81], stage1_43[82], stage1_43[83]},
      {stage2_45[13],stage2_44[36],stage2_43[36],stage2_42[62],stage2_41[86]}
   );
   gpc615_5 gpc5446 (
      {stage1_41[88], stage1_41[89], stage1_41[90], stage1_41[91], stage1_41[92]},
      {stage1_42[147]},
      {stage1_43[84], stage1_43[85], stage1_43[86], stage1_43[87], stage1_43[88], stage1_43[89]},
      {stage2_45[14],stage2_44[37],stage2_43[37],stage2_42[63],stage2_41[87]}
   );
   gpc615_5 gpc5447 (
      {stage1_41[93], stage1_41[94], stage1_41[95], stage1_41[96], stage1_41[97]},
      {stage1_42[148]},
      {stage1_43[90], stage1_43[91], stage1_43[92], stage1_43[93], stage1_43[94], stage1_43[95]},
      {stage2_45[15],stage2_44[38],stage2_43[38],stage2_42[64],stage2_41[88]}
   );
   gpc615_5 gpc5448 (
      {stage1_41[98], stage1_41[99], stage1_41[100], stage1_41[101], stage1_41[102]},
      {stage1_42[149]},
      {stage1_43[96], stage1_43[97], stage1_43[98], stage1_43[99], stage1_43[100], stage1_43[101]},
      {stage2_45[16],stage2_44[39],stage2_43[39],stage2_42[65],stage2_41[89]}
   );
   gpc615_5 gpc5449 (
      {stage1_41[103], stage1_41[104], stage1_41[105], stage1_41[106], stage1_41[107]},
      {stage1_42[150]},
      {stage1_43[102], stage1_43[103], stage1_43[104], stage1_43[105], stage1_43[106], stage1_43[107]},
      {stage2_45[17],stage2_44[40],stage2_43[40],stage2_42[66],stage2_41[90]}
   );
   gpc615_5 gpc5450 (
      {stage1_41[108], stage1_41[109], stage1_41[110], stage1_41[111], stage1_41[112]},
      {stage1_42[151]},
      {stage1_43[108], stage1_43[109], stage1_43[110], stage1_43[111], stage1_43[112], stage1_43[113]},
      {stage2_45[18],stage2_44[41],stage2_43[41],stage2_42[67],stage2_41[91]}
   );
   gpc615_5 gpc5451 (
      {stage1_41[113], stage1_41[114], stage1_41[115], stage1_41[116], stage1_41[117]},
      {stage1_42[152]},
      {stage1_43[114], stage1_43[115], stage1_43[116], stage1_43[117], stage1_43[118], stage1_43[119]},
      {stage2_45[19],stage2_44[42],stage2_43[42],stage2_42[68],stage2_41[92]}
   );
   gpc615_5 gpc5452 (
      {stage1_41[118], stage1_41[119], stage1_41[120], stage1_41[121], stage1_41[122]},
      {stage1_42[153]},
      {stage1_43[120], stage1_43[121], stage1_43[122], stage1_43[123], stage1_43[124], stage1_43[125]},
      {stage2_45[20],stage2_44[43],stage2_43[43],stage2_42[69],stage2_41[93]}
   );
   gpc615_5 gpc5453 (
      {stage1_41[123], stage1_41[124], stage1_41[125], stage1_41[126], stage1_41[127]},
      {stage1_42[154]},
      {stage1_43[126], stage1_43[127], stage1_43[128], stage1_43[129], stage1_43[130], stage1_43[131]},
      {stage2_45[21],stage2_44[44],stage2_43[44],stage2_42[70],stage2_41[94]}
   );
   gpc615_5 gpc5454 (
      {stage1_41[128], stage1_41[129], stage1_41[130], stage1_41[131], stage1_41[132]},
      {stage1_42[155]},
      {stage1_43[132], stage1_43[133], stage1_43[134], stage1_43[135], stage1_43[136], stage1_43[137]},
      {stage2_45[22],stage2_44[45],stage2_43[45],stage2_42[71],stage2_41[95]}
   );
   gpc615_5 gpc5455 (
      {stage1_41[133], stage1_41[134], stage1_41[135], stage1_41[136], stage1_41[137]},
      {stage1_42[156]},
      {stage1_43[138], stage1_43[139], stage1_43[140], stage1_43[141], stage1_43[142], stage1_43[143]},
      {stage2_45[23],stage2_44[46],stage2_43[46],stage2_42[72],stage2_41[96]}
   );
   gpc615_5 gpc5456 (
      {stage1_41[138], stage1_41[139], stage1_41[140], stage1_41[141], stage1_41[142]},
      {stage1_42[157]},
      {stage1_43[144], stage1_43[145], stage1_43[146], stage1_43[147], stage1_43[148], stage1_43[149]},
      {stage2_45[24],stage2_44[47],stage2_43[47],stage2_42[73],stage2_41[97]}
   );
   gpc615_5 gpc5457 (
      {stage1_41[143], stage1_41[144], stage1_41[145], stage1_41[146], stage1_41[147]},
      {stage1_42[158]},
      {stage1_43[150], stage1_43[151], stage1_43[152], stage1_43[153], stage1_43[154], stage1_43[155]},
      {stage2_45[25],stage2_44[48],stage2_43[48],stage2_42[74],stage2_41[98]}
   );
   gpc615_5 gpc5458 (
      {stage1_41[148], stage1_41[149], stage1_41[150], stage1_41[151], stage1_41[152]},
      {stage1_42[159]},
      {stage1_43[156], stage1_43[157], stage1_43[158], stage1_43[159], stage1_43[160], stage1_43[161]},
      {stage2_45[26],stage2_44[49],stage2_43[49],stage2_42[75],stage2_41[99]}
   );
   gpc615_5 gpc5459 (
      {stage1_41[153], stage1_41[154], stage1_41[155], stage1_41[156], stage1_41[157]},
      {stage1_42[160]},
      {stage1_43[162], stage1_43[163], stage1_43[164], stage1_43[165], stage1_43[166], stage1_43[167]},
      {stage2_45[27],stage2_44[50],stage2_43[50],stage2_42[76],stage2_41[100]}
   );
   gpc615_5 gpc5460 (
      {stage1_41[158], stage1_41[159], stage1_41[160], stage1_41[161], stage1_41[162]},
      {stage1_42[161]},
      {stage1_43[168], stage1_43[169], stage1_43[170], stage1_43[171], stage1_43[172], stage1_43[173]},
      {stage2_45[28],stage2_44[51],stage2_43[51],stage2_42[77],stage2_41[101]}
   );
   gpc615_5 gpc5461 (
      {stage1_41[163], stage1_41[164], stage1_41[165], stage1_41[166], stage1_41[167]},
      {stage1_42[162]},
      {stage1_43[174], stage1_43[175], stage1_43[176], stage1_43[177], stage1_43[178], stage1_43[179]},
      {stage2_45[29],stage2_44[52],stage2_43[52],stage2_42[78],stage2_41[102]}
   );
   gpc615_5 gpc5462 (
      {stage1_42[163], stage1_42[164], stage1_42[165], stage1_42[166], stage1_42[167]},
      {stage1_43[180]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[30],stage2_44[53],stage2_43[53],stage2_42[79]}
   );
   gpc615_5 gpc5463 (
      {stage1_43[181], stage1_43[182], stage1_43[183], stage1_43[184], stage1_43[185]},
      {stage1_44[6]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[1],stage2_45[31],stage2_44[54],stage2_43[54]}
   );
   gpc615_5 gpc5464 (
      {stage1_43[186], stage1_43[187], stage1_43[188], stage1_43[189], stage1_43[190]},
      {stage1_44[7]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[2],stage2_45[32],stage2_44[55],stage2_43[55]}
   );
   gpc615_5 gpc5465 (
      {stage1_43[191], stage1_43[192], stage1_43[193], stage1_43[194], stage1_43[195]},
      {stage1_44[8]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[3],stage2_45[33],stage2_44[56],stage2_43[56]}
   );
   gpc615_5 gpc5466 (
      {stage1_43[196], stage1_43[197], stage1_43[198], stage1_43[199], stage1_43[200]},
      {stage1_44[9]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[4],stage2_45[34],stage2_44[57],stage2_43[57]}
   );
   gpc615_5 gpc5467 (
      {stage1_43[201], stage1_43[202], stage1_43[203], stage1_43[204], stage1_43[205]},
      {stage1_44[10]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[5],stage2_45[35],stage2_44[58],stage2_43[58]}
   );
   gpc615_5 gpc5468 (
      {stage1_43[206], stage1_43[207], stage1_43[208], stage1_43[209], stage1_43[210]},
      {stage1_44[11]},
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage2_47[5],stage2_46[6],stage2_45[36],stage2_44[59],stage2_43[59]}
   );
   gpc615_5 gpc5469 (
      {stage1_43[211], stage1_43[212], stage1_43[213], stage1_43[214], stage1_43[215]},
      {stage1_44[12]},
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage2_47[6],stage2_46[7],stage2_45[37],stage2_44[60],stage2_43[60]}
   );
   gpc615_5 gpc5470 (
      {stage1_43[216], stage1_43[217], stage1_43[218], stage1_43[219], stage1_43[220]},
      {stage1_44[13]},
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage2_47[7],stage2_46[8],stage2_45[38],stage2_44[61],stage2_43[61]}
   );
   gpc615_5 gpc5471 (
      {stage1_43[221], stage1_43[222], stage1_43[223], stage1_43[224], stage1_43[225]},
      {stage1_44[14]},
      {stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51], stage1_45[52], stage1_45[53]},
      {stage2_47[8],stage2_46[9],stage2_45[39],stage2_44[62],stage2_43[62]}
   );
   gpc615_5 gpc5472 (
      {stage1_43[226], stage1_43[227], stage1_43[228], stage1_43[229], stage1_43[230]},
      {stage1_44[15]},
      {stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57], stage1_45[58], stage1_45[59]},
      {stage2_47[9],stage2_46[10],stage2_45[40],stage2_44[63],stage2_43[63]}
   );
   gpc615_5 gpc5473 (
      {stage1_43[231], stage1_43[232], stage1_43[233], stage1_43[234], stage1_43[235]},
      {stage1_44[16]},
      {stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63], stage1_45[64], stage1_45[65]},
      {stage2_47[10],stage2_46[11],stage2_45[41],stage2_44[64],stage2_43[64]}
   );
   gpc615_5 gpc5474 (
      {stage1_43[236], stage1_43[237], stage1_43[238], stage1_43[239], stage1_43[240]},
      {stage1_44[17]},
      {stage1_45[66], stage1_45[67], stage1_45[68], stage1_45[69], stage1_45[70], stage1_45[71]},
      {stage2_47[11],stage2_46[12],stage2_45[42],stage2_44[65],stage2_43[65]}
   );
   gpc606_5 gpc5475 (
      {stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[12],stage2_46[13],stage2_45[43],stage2_44[66]}
   );
   gpc606_5 gpc5476 (
      {stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[13],stage2_46[14],stage2_45[44],stage2_44[67]}
   );
   gpc606_5 gpc5477 (
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34], stage1_44[35]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage2_48[2],stage2_47[14],stage2_46[15],stage2_45[45],stage2_44[68]}
   );
   gpc606_5 gpc5478 (
      {stage1_44[36], stage1_44[37], stage1_44[38], stage1_44[39], stage1_44[40], stage1_44[41]},
      {stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21], stage1_46[22], stage1_46[23]},
      {stage2_48[3],stage2_47[15],stage2_46[16],stage2_45[46],stage2_44[69]}
   );
   gpc606_5 gpc5479 (
      {stage1_44[42], stage1_44[43], stage1_44[44], stage1_44[45], stage1_44[46], stage1_44[47]},
      {stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27], stage1_46[28], stage1_46[29]},
      {stage2_48[4],stage2_47[16],stage2_46[17],stage2_45[47],stage2_44[70]}
   );
   gpc606_5 gpc5480 (
      {stage1_44[48], stage1_44[49], stage1_44[50], stage1_44[51], stage1_44[52], stage1_44[53]},
      {stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35]},
      {stage2_48[5],stage2_47[17],stage2_46[18],stage2_45[48],stage2_44[71]}
   );
   gpc606_5 gpc5481 (
      {stage1_44[54], stage1_44[55], stage1_44[56], stage1_44[57], stage1_44[58], stage1_44[59]},
      {stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage2_48[6],stage2_47[18],stage2_46[19],stage2_45[49],stage2_44[72]}
   );
   gpc606_5 gpc5482 (
      {stage1_44[60], stage1_44[61], stage1_44[62], stage1_44[63], stage1_44[64], stage1_44[65]},
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46], stage1_46[47]},
      {stage2_48[7],stage2_47[19],stage2_46[20],stage2_45[50],stage2_44[73]}
   );
   gpc606_5 gpc5483 (
      {stage1_44[66], stage1_44[67], stage1_44[68], stage1_44[69], stage1_44[70], stage1_44[71]},
      {stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51], stage1_46[52], stage1_46[53]},
      {stage2_48[8],stage2_47[20],stage2_46[21],stage2_45[51],stage2_44[74]}
   );
   gpc606_5 gpc5484 (
      {stage1_44[72], stage1_44[73], stage1_44[74], stage1_44[75], stage1_44[76], stage1_44[77]},
      {stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57], stage1_46[58], stage1_46[59]},
      {stage2_48[9],stage2_47[21],stage2_46[22],stage2_45[52],stage2_44[75]}
   );
   gpc606_5 gpc5485 (
      {stage1_44[78], stage1_44[79], stage1_44[80], stage1_44[81], stage1_44[82], stage1_44[83]},
      {stage1_46[60], stage1_46[61], stage1_46[62], stage1_46[63], stage1_46[64], stage1_46[65]},
      {stage2_48[10],stage2_47[22],stage2_46[23],stage2_45[53],stage2_44[76]}
   );
   gpc606_5 gpc5486 (
      {stage1_44[84], stage1_44[85], stage1_44[86], stage1_44[87], stage1_44[88], stage1_44[89]},
      {stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69], stage1_46[70], stage1_46[71]},
      {stage2_48[11],stage2_47[23],stage2_46[24],stage2_45[54],stage2_44[77]}
   );
   gpc606_5 gpc5487 (
      {stage1_44[90], stage1_44[91], stage1_44[92], stage1_44[93], stage1_44[94], stage1_44[95]},
      {stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75], stage1_46[76], stage1_46[77]},
      {stage2_48[12],stage2_47[24],stage2_46[25],stage2_45[55],stage2_44[78]}
   );
   gpc606_5 gpc5488 (
      {stage1_44[96], stage1_44[97], stage1_44[98], stage1_44[99], stage1_44[100], stage1_44[101]},
      {stage1_46[78], stage1_46[79], stage1_46[80], stage1_46[81], stage1_46[82], stage1_46[83]},
      {stage2_48[13],stage2_47[25],stage2_46[26],stage2_45[56],stage2_44[79]}
   );
   gpc606_5 gpc5489 (
      {stage1_44[102], stage1_44[103], stage1_44[104], stage1_44[105], stage1_44[106], stage1_44[107]},
      {stage1_46[84], stage1_46[85], stage1_46[86], stage1_46[87], stage1_46[88], stage1_46[89]},
      {stage2_48[14],stage2_47[26],stage2_46[27],stage2_45[57],stage2_44[80]}
   );
   gpc606_5 gpc5490 (
      {stage1_44[108], stage1_44[109], stage1_44[110], stage1_44[111], stage1_44[112], stage1_44[113]},
      {stage1_46[90], stage1_46[91], stage1_46[92], stage1_46[93], stage1_46[94], stage1_46[95]},
      {stage2_48[15],stage2_47[27],stage2_46[28],stage2_45[58],stage2_44[81]}
   );
   gpc606_5 gpc5491 (
      {stage1_44[114], stage1_44[115], stage1_44[116], stage1_44[117], stage1_44[118], stage1_44[119]},
      {stage1_46[96], stage1_46[97], stage1_46[98], stage1_46[99], stage1_46[100], stage1_46[101]},
      {stage2_48[16],stage2_47[28],stage2_46[29],stage2_45[59],stage2_44[82]}
   );
   gpc606_5 gpc5492 (
      {stage1_44[120], stage1_44[121], stage1_44[122], stage1_44[123], stage1_44[124], stage1_44[125]},
      {stage1_46[102], stage1_46[103], stage1_46[104], stage1_46[105], stage1_46[106], stage1_46[107]},
      {stage2_48[17],stage2_47[29],stage2_46[30],stage2_45[60],stage2_44[83]}
   );
   gpc606_5 gpc5493 (
      {stage1_44[126], stage1_44[127], stage1_44[128], stage1_44[129], stage1_44[130], stage1_44[131]},
      {stage1_46[108], stage1_46[109], stage1_46[110], stage1_46[111], stage1_46[112], stage1_46[113]},
      {stage2_48[18],stage2_47[30],stage2_46[31],stage2_45[61],stage2_44[84]}
   );
   gpc606_5 gpc5494 (
      {stage1_44[132], stage1_44[133], stage1_44[134], stage1_44[135], stage1_44[136], stage1_44[137]},
      {stage1_46[114], stage1_46[115], stage1_46[116], stage1_46[117], stage1_46[118], stage1_46[119]},
      {stage2_48[19],stage2_47[31],stage2_46[32],stage2_45[62],stage2_44[85]}
   );
   gpc606_5 gpc5495 (
      {stage1_44[138], stage1_44[139], stage1_44[140], stage1_44[141], stage1_44[142], stage1_44[143]},
      {stage1_46[120], stage1_46[121], stage1_46[122], stage1_46[123], stage1_46[124], stage1_46[125]},
      {stage2_48[20],stage2_47[32],stage2_46[33],stage2_45[63],stage2_44[86]}
   );
   gpc606_5 gpc5496 (
      {stage1_44[144], stage1_44[145], stage1_44[146], stage1_44[147], stage1_44[148], stage1_44[149]},
      {stage1_46[126], stage1_46[127], stage1_46[128], stage1_46[129], stage1_46[130], stage1_46[131]},
      {stage2_48[21],stage2_47[33],stage2_46[34],stage2_45[64],stage2_44[87]}
   );
   gpc606_5 gpc5497 (
      {stage1_44[150], stage1_44[151], stage1_44[152], stage1_44[153], stage1_44[154], stage1_44[155]},
      {stage1_46[132], stage1_46[133], stage1_46[134], stage1_46[135], stage1_46[136], stage1_46[137]},
      {stage2_48[22],stage2_47[34],stage2_46[35],stage2_45[65],stage2_44[88]}
   );
   gpc606_5 gpc5498 (
      {stage1_44[156], stage1_44[157], stage1_44[158], stage1_44[159], stage1_44[160], stage1_44[161]},
      {stage1_46[138], stage1_46[139], stage1_46[140], stage1_46[141], stage1_46[142], stage1_46[143]},
      {stage2_48[23],stage2_47[35],stage2_46[36],stage2_45[66],stage2_44[89]}
   );
   gpc606_5 gpc5499 (
      {stage1_44[162], stage1_44[163], stage1_44[164], stage1_44[165], stage1_44[166], stage1_44[167]},
      {stage1_46[144], stage1_46[145], stage1_46[146], stage1_46[147], stage1_46[148], stage1_46[149]},
      {stage2_48[24],stage2_47[36],stage2_46[37],stage2_45[67],stage2_44[90]}
   );
   gpc606_5 gpc5500 (
      {stage1_44[168], stage1_44[169], stage1_44[170], stage1_44[171], stage1_44[172], stage1_44[173]},
      {stage1_46[150], stage1_46[151], stage1_46[152], stage1_46[153], stage1_46[154], stage1_46[155]},
      {stage2_48[25],stage2_47[37],stage2_46[38],stage2_45[68],stage2_44[91]}
   );
   gpc606_5 gpc5501 (
      {stage1_44[174], stage1_44[175], stage1_44[176], stage1_44[177], stage1_44[178], stage1_44[179]},
      {stage1_46[156], stage1_46[157], stage1_46[158], stage1_46[159], stage1_46[160], stage1_46[161]},
      {stage2_48[26],stage2_47[38],stage2_46[39],stage2_45[69],stage2_44[92]}
   );
   gpc606_5 gpc5502 (
      {stage1_44[180], stage1_44[181], stage1_44[182], stage1_44[183], stage1_44[184], stage1_44[185]},
      {stage1_46[162], stage1_46[163], stage1_46[164], stage1_46[165], stage1_46[166], stage1_46[167]},
      {stage2_48[27],stage2_47[39],stage2_46[40],stage2_45[70],stage2_44[93]}
   );
   gpc606_5 gpc5503 (
      {stage1_44[186], stage1_44[187], stage1_44[188], stage1_44[189], stage1_44[190], stage1_44[191]},
      {stage1_46[168], stage1_46[169], stage1_46[170], stage1_46[171], stage1_46[172], stage1_46[173]},
      {stage2_48[28],stage2_47[40],stage2_46[41],stage2_45[71],stage2_44[94]}
   );
   gpc606_5 gpc5504 (
      {stage1_44[192], stage1_44[193], stage1_44[194], stage1_44[195], stage1_44[196], stage1_44[197]},
      {stage1_46[174], stage1_46[175], stage1_46[176], stage1_46[177], stage1_46[178], stage1_46[179]},
      {stage2_48[29],stage2_47[41],stage2_46[42],stage2_45[72],stage2_44[95]}
   );
   gpc606_5 gpc5505 (
      {stage1_44[198], stage1_44[199], stage1_44[200], stage1_44[201], stage1_44[202], stage1_44[203]},
      {stage1_46[180], stage1_46[181], stage1_46[182], stage1_46[183], stage1_46[184], stage1_46[185]},
      {stage2_48[30],stage2_47[42],stage2_46[43],stage2_45[73],stage2_44[96]}
   );
   gpc606_5 gpc5506 (
      {stage1_44[204], stage1_44[205], stage1_44[206], stage1_44[207], stage1_44[208], stage1_44[209]},
      {stage1_46[186], stage1_46[187], stage1_46[188], stage1_46[189], stage1_46[190], stage1_46[191]},
      {stage2_48[31],stage2_47[43],stage2_46[44],stage2_45[74],stage2_44[97]}
   );
   gpc606_5 gpc5507 (
      {stage1_44[210], stage1_44[211], stage1_44[212], stage1_44[213], stage1_44[214], stage1_44[215]},
      {stage1_46[192], stage1_46[193], stage1_46[194], stage1_46[195], stage1_46[196], stage1_46[197]},
      {stage2_48[32],stage2_47[44],stage2_46[45],stage2_45[75],stage2_44[98]}
   );
   gpc606_5 gpc5508 (
      {stage1_44[216], stage1_44[217], stage1_44[218], stage1_44[219], stage1_44[220], stage1_44[221]},
      {stage1_46[198], stage1_46[199], stage1_46[200], stage1_46[201], stage1_46[202], stage1_46[203]},
      {stage2_48[33],stage2_47[45],stage2_46[46],stage2_45[76],stage2_44[99]}
   );
   gpc606_5 gpc5509 (
      {stage1_44[222], stage1_44[223], stage1_44[224], stage1_44[225], stage1_44[226], stage1_44[227]},
      {stage1_46[204], stage1_46[205], stage1_46[206], stage1_46[207], stage1_46[208], stage1_46[209]},
      {stage2_48[34],stage2_47[46],stage2_46[47],stage2_45[77],stage2_44[100]}
   );
   gpc606_5 gpc5510 (
      {stage1_44[228], stage1_44[229], stage1_44[230], stage1_44[231], stage1_44[232], stage1_44[233]},
      {stage1_46[210], stage1_46[211], stage1_46[212], stage1_46[213], stage1_46[214], stage1_46[215]},
      {stage2_48[35],stage2_47[47],stage2_46[48],stage2_45[78],stage2_44[101]}
   );
   gpc606_5 gpc5511 (
      {stage1_44[234], stage1_44[235], stage1_44[236], stage1_44[237], stage1_44[238], stage1_44[239]},
      {stage1_46[216], stage1_46[217], stage1_46[218], stage1_46[219], stage1_46[220], stage1_46[221]},
      {stage2_48[36],stage2_47[48],stage2_46[49],stage2_45[79],stage2_44[102]}
   );
   gpc606_5 gpc5512 (
      {stage1_45[72], stage1_45[73], stage1_45[74], stage1_45[75], stage1_45[76], stage1_45[77]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[37],stage2_47[49],stage2_46[50],stage2_45[80]}
   );
   gpc606_5 gpc5513 (
      {stage1_45[78], stage1_45[79], stage1_45[80], stage1_45[81], stage1_45[82], stage1_45[83]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[38],stage2_47[50],stage2_46[51],stage2_45[81]}
   );
   gpc615_5 gpc5514 (
      {stage1_45[84], stage1_45[85], stage1_45[86], stage1_45[87], stage1_45[88]},
      {stage1_46[222]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[39],stage2_47[51],stage2_46[52],stage2_45[82]}
   );
   gpc615_5 gpc5515 (
      {stage1_45[89], stage1_45[90], stage1_45[91], stage1_45[92], stage1_45[93]},
      {stage1_46[223]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[40],stage2_47[52],stage2_46[53],stage2_45[83]}
   );
   gpc615_5 gpc5516 (
      {stage1_45[94], stage1_45[95], stage1_45[96], stage1_45[97], stage1_45[98]},
      {stage1_46[224]},
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage2_49[4],stage2_48[41],stage2_47[53],stage2_46[54],stage2_45[84]}
   );
   gpc615_5 gpc5517 (
      {stage1_45[99], stage1_45[100], stage1_45[101], stage1_45[102], stage1_45[103]},
      {stage1_46[225]},
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage2_49[5],stage2_48[42],stage2_47[54],stage2_46[55],stage2_45[85]}
   );
   gpc615_5 gpc5518 (
      {stage1_45[104], stage1_45[105], stage1_45[106], stage1_45[107], stage1_45[108]},
      {stage1_46[226]},
      {stage1_47[36], stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41]},
      {stage2_49[6],stage2_48[43],stage2_47[55],stage2_46[56],stage2_45[86]}
   );
   gpc615_5 gpc5519 (
      {stage1_45[109], stage1_45[110], stage1_45[111], stage1_45[112], stage1_45[113]},
      {stage1_46[227]},
      {stage1_47[42], stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47]},
      {stage2_49[7],stage2_48[44],stage2_47[56],stage2_46[57],stage2_45[87]}
   );
   gpc615_5 gpc5520 (
      {stage1_45[114], stage1_45[115], stage1_45[116], stage1_45[117], stage1_45[118]},
      {stage1_46[228]},
      {stage1_47[48], stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage2_49[8],stage2_48[45],stage2_47[57],stage2_46[58],stage2_45[88]}
   );
   gpc615_5 gpc5521 (
      {stage1_45[119], stage1_45[120], stage1_45[121], stage1_45[122], stage1_45[123]},
      {stage1_46[229]},
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58], stage1_47[59]},
      {stage2_49[9],stage2_48[46],stage2_47[58],stage2_46[59],stage2_45[89]}
   );
   gpc615_5 gpc5522 (
      {stage1_45[124], stage1_45[125], stage1_45[126], stage1_45[127], stage1_45[128]},
      {stage1_46[230]},
      {stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63], stage1_47[64], stage1_47[65]},
      {stage2_49[10],stage2_48[47],stage2_47[59],stage2_46[60],stage2_45[90]}
   );
   gpc615_5 gpc5523 (
      {stage1_45[129], stage1_45[130], stage1_45[131], stage1_45[132], stage1_45[133]},
      {stage1_46[231]},
      {stage1_47[66], stage1_47[67], stage1_47[68], stage1_47[69], stage1_47[70], stage1_47[71]},
      {stage2_49[11],stage2_48[48],stage2_47[60],stage2_46[61],stage2_45[91]}
   );
   gpc615_5 gpc5524 (
      {stage1_45[134], stage1_45[135], stage1_45[136], stage1_45[137], stage1_45[138]},
      {stage1_46[232]},
      {stage1_47[72], stage1_47[73], stage1_47[74], stage1_47[75], stage1_47[76], stage1_47[77]},
      {stage2_49[12],stage2_48[49],stage2_47[61],stage2_46[62],stage2_45[92]}
   );
   gpc615_5 gpc5525 (
      {stage1_45[139], stage1_45[140], stage1_45[141], stage1_45[142], stage1_45[143]},
      {stage1_46[233]},
      {stage1_47[78], stage1_47[79], stage1_47[80], stage1_47[81], stage1_47[82], stage1_47[83]},
      {stage2_49[13],stage2_48[50],stage2_47[62],stage2_46[63],stage2_45[93]}
   );
   gpc615_5 gpc5526 (
      {stage1_45[144], stage1_45[145], stage1_45[146], stage1_45[147], stage1_45[148]},
      {stage1_46[234]},
      {stage1_47[84], stage1_47[85], stage1_47[86], stage1_47[87], stage1_47[88], stage1_47[89]},
      {stage2_49[14],stage2_48[51],stage2_47[63],stage2_46[64],stage2_45[94]}
   );
   gpc615_5 gpc5527 (
      {stage1_45[149], stage1_45[150], stage1_45[151], stage1_45[152], stage1_45[153]},
      {stage1_46[235]},
      {stage1_47[90], stage1_47[91], stage1_47[92], stage1_47[93], stage1_47[94], stage1_47[95]},
      {stage2_49[15],stage2_48[52],stage2_47[64],stage2_46[65],stage2_45[95]}
   );
   gpc615_5 gpc5528 (
      {stage1_45[154], stage1_45[155], stage1_45[156], stage1_45[157], stage1_45[158]},
      {stage1_46[236]},
      {stage1_47[96], stage1_47[97], stage1_47[98], stage1_47[99], stage1_47[100], stage1_47[101]},
      {stage2_49[16],stage2_48[53],stage2_47[65],stage2_46[66],stage2_45[96]}
   );
   gpc615_5 gpc5529 (
      {stage1_45[159], stage1_45[160], stage1_45[161], stage1_45[162], stage1_45[163]},
      {stage1_46[237]},
      {stage1_47[102], stage1_47[103], stage1_47[104], stage1_47[105], stage1_47[106], stage1_47[107]},
      {stage2_49[17],stage2_48[54],stage2_47[66],stage2_46[67],stage2_45[97]}
   );
   gpc615_5 gpc5530 (
      {stage1_45[164], stage1_45[165], stage1_45[166], stage1_45[167], stage1_45[168]},
      {stage1_46[238]},
      {stage1_47[108], stage1_47[109], stage1_47[110], stage1_47[111], stage1_47[112], stage1_47[113]},
      {stage2_49[18],stage2_48[55],stage2_47[67],stage2_46[68],stage2_45[98]}
   );
   gpc615_5 gpc5531 (
      {stage1_45[169], stage1_45[170], stage1_45[171], stage1_45[172], stage1_45[173]},
      {stage1_46[239]},
      {stage1_47[114], stage1_47[115], stage1_47[116], stage1_47[117], stage1_47[118], stage1_47[119]},
      {stage2_49[19],stage2_48[56],stage2_47[68],stage2_46[69],stage2_45[99]}
   );
   gpc615_5 gpc5532 (
      {stage1_45[174], stage1_45[175], stage1_45[176], stage1_45[177], stage1_45[178]},
      {stage1_46[240]},
      {stage1_47[120], stage1_47[121], stage1_47[122], stage1_47[123], stage1_47[124], stage1_47[125]},
      {stage2_49[20],stage2_48[57],stage2_47[69],stage2_46[70],stage2_45[100]}
   );
   gpc615_5 gpc5533 (
      {stage1_45[179], stage1_45[180], stage1_45[181], stage1_45[182], stage1_45[183]},
      {stage1_46[241]},
      {stage1_47[126], stage1_47[127], stage1_47[128], stage1_47[129], stage1_47[130], stage1_47[131]},
      {stage2_49[21],stage2_48[58],stage2_47[70],stage2_46[71],stage2_45[101]}
   );
   gpc615_5 gpc5534 (
      {stage1_45[184], stage1_45[185], stage1_45[186], stage1_45[187], stage1_45[188]},
      {stage1_46[242]},
      {stage1_47[132], stage1_47[133], stage1_47[134], stage1_47[135], stage1_47[136], stage1_47[137]},
      {stage2_49[22],stage2_48[59],stage2_47[71],stage2_46[72],stage2_45[102]}
   );
   gpc615_5 gpc5535 (
      {stage1_45[189], stage1_45[190], stage1_45[191], stage1_45[192], stage1_45[193]},
      {stage1_46[243]},
      {stage1_47[138], stage1_47[139], stage1_47[140], stage1_47[141], stage1_47[142], stage1_47[143]},
      {stage2_49[23],stage2_48[60],stage2_47[72],stage2_46[73],stage2_45[103]}
   );
   gpc615_5 gpc5536 (
      {stage1_45[194], stage1_45[195], stage1_45[196], stage1_45[197], stage1_45[198]},
      {stage1_46[244]},
      {stage1_47[144], stage1_47[145], stage1_47[146], stage1_47[147], stage1_47[148], stage1_47[149]},
      {stage2_49[24],stage2_48[61],stage2_47[73],stage2_46[74],stage2_45[104]}
   );
   gpc615_5 gpc5537 (
      {stage1_46[245], stage1_46[246], stage1_46[247], stage1_46[248], stage1_46[249]},
      {stage1_47[150]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[25],stage2_48[62],stage2_47[74],stage2_46[75]}
   );
   gpc615_5 gpc5538 (
      {stage1_46[250], stage1_46[251], stage1_46[252], stage1_46[253], stage1_46[254]},
      {stage1_47[151]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[26],stage2_48[63],stage2_47[75],stage2_46[76]}
   );
   gpc615_5 gpc5539 (
      {stage1_46[255], stage1_46[256], stage1_46[257], stage1_46[258], stage1_46[259]},
      {stage1_47[152]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[27],stage2_48[64],stage2_47[76],stage2_46[77]}
   );
   gpc615_5 gpc5540 (
      {stage1_46[260], stage1_46[261], stage1_46[262], stage1_46[263], stage1_46[264]},
      {stage1_47[153]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[28],stage2_48[65],stage2_47[77],stage2_46[78]}
   );
   gpc615_5 gpc5541 (
      {stage1_46[265], stage1_46[266], stage1_46[267], stage1_46[268], stage1_46[269]},
      {stage1_47[154]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[29],stage2_48[66],stage2_47[78],stage2_46[79]}
   );
   gpc615_5 gpc5542 (
      {stage1_46[270], stage1_46[271], stage1_46[272], stage1_46[273], stage1_46[274]},
      {stage1_47[155]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[30],stage2_48[67],stage2_47[79],stage2_46[80]}
   );
   gpc615_5 gpc5543 (
      {stage1_46[275], stage1_46[276], stage1_46[277], stage1_46[278], stage1_46[279]},
      {stage1_47[156]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[31],stage2_48[68],stage2_47[80],stage2_46[81]}
   );
   gpc615_5 gpc5544 (
      {stage1_46[280], stage1_46[281], stage1_46[282], stage1_46[283], stage1_46[284]},
      {stage1_47[157]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[32],stage2_48[69],stage2_47[81],stage2_46[82]}
   );
   gpc615_5 gpc5545 (
      {stage1_46[285], stage1_46[286], stage1_46[287], stage1_46[288], stage1_46[289]},
      {stage1_47[158]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[33],stage2_48[70],stage2_47[82],stage2_46[83]}
   );
   gpc615_5 gpc5546 (
      {stage1_46[290], stage1_46[291], stage1_46[292], stage1_46[293], stage1_46[294]},
      {stage1_47[159]},
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage2_50[9],stage2_49[34],stage2_48[71],stage2_47[83],stage2_46[84]}
   );
   gpc615_5 gpc5547 (
      {stage1_47[160], stage1_47[161], stage1_47[162], stage1_47[163], stage1_47[164]},
      {stage1_48[60]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[10],stage2_49[35],stage2_48[72],stage2_47[84]}
   );
   gpc615_5 gpc5548 (
      {stage1_47[165], stage1_47[166], stage1_47[167], stage1_47[168], stage1_47[169]},
      {stage1_48[61]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[11],stage2_49[36],stage2_48[73],stage2_47[85]}
   );
   gpc615_5 gpc5549 (
      {stage1_47[170], stage1_47[171], stage1_47[172], stage1_47[173], stage1_47[174]},
      {stage1_48[62]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[12],stage2_49[37],stage2_48[74],stage2_47[86]}
   );
   gpc615_5 gpc5550 (
      {stage1_47[175], stage1_47[176], stage1_47[177], stage1_47[178], stage1_47[179]},
      {stage1_48[63]},
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage2_51[3],stage2_50[13],stage2_49[38],stage2_48[75],stage2_47[87]}
   );
   gpc615_5 gpc5551 (
      {stage1_47[180], stage1_47[181], stage1_47[182], stage1_47[183], stage1_47[184]},
      {stage1_48[64]},
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage2_51[4],stage2_50[14],stage2_49[39],stage2_48[76],stage2_47[88]}
   );
   gpc615_5 gpc5552 (
      {stage1_47[185], stage1_47[186], stage1_47[187], stage1_47[188], stage1_47[189]},
      {stage1_48[65]},
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage2_51[5],stage2_50[15],stage2_49[40],stage2_48[77],stage2_47[89]}
   );
   gpc615_5 gpc5553 (
      {stage1_47[190], stage1_47[191], stage1_47[192], stage1_47[193], stage1_47[194]},
      {stage1_48[66]},
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage2_51[6],stage2_50[16],stage2_49[41],stage2_48[78],stage2_47[90]}
   );
   gpc615_5 gpc5554 (
      {stage1_47[195], stage1_47[196], stage1_47[197], stage1_47[198], stage1_47[199]},
      {stage1_48[67]},
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage2_51[7],stage2_50[17],stage2_49[42],stage2_48[79],stage2_47[91]}
   );
   gpc615_5 gpc5555 (
      {stage1_47[200], stage1_47[201], stage1_47[202], stage1_47[203], stage1_47[204]},
      {stage1_48[68]},
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage2_51[8],stage2_50[18],stage2_49[43],stage2_48[80],stage2_47[92]}
   );
   gpc615_5 gpc5556 (
      {stage1_47[205], stage1_47[206], stage1_47[207], stage1_47[208], stage1_47[209]},
      {stage1_48[69]},
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage2_51[9],stage2_50[19],stage2_49[44],stage2_48[81],stage2_47[93]}
   );
   gpc615_5 gpc5557 (
      {stage1_47[210], stage1_47[211], stage1_47[212], stage1_47[213], stage1_47[214]},
      {stage1_48[70]},
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage2_51[10],stage2_50[20],stage2_49[45],stage2_48[82],stage2_47[94]}
   );
   gpc615_5 gpc5558 (
      {stage1_47[215], stage1_47[216], stage1_47[217], stage1_47[218], stage1_47[219]},
      {stage1_48[71]},
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage2_51[11],stage2_50[21],stage2_49[46],stage2_48[83],stage2_47[95]}
   );
   gpc615_5 gpc5559 (
      {stage1_47[220], stage1_47[221], stage1_47[222], stage1_47[223], stage1_47[224]},
      {stage1_48[72]},
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage2_51[12],stage2_50[22],stage2_49[47],stage2_48[84],stage2_47[96]}
   );
   gpc615_5 gpc5560 (
      {stage1_47[225], stage1_47[226], stage1_47[227], stage1_47[228], stage1_47[229]},
      {stage1_48[73]},
      {stage1_49[78], stage1_49[79], stage1_49[80], stage1_49[81], stage1_49[82], stage1_49[83]},
      {stage2_51[13],stage2_50[23],stage2_49[48],stage2_48[85],stage2_47[97]}
   );
   gpc606_5 gpc5561 (
      {stage1_48[74], stage1_48[75], stage1_48[76], stage1_48[77], stage1_48[78], stage1_48[79]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[14],stage2_50[24],stage2_49[49],stage2_48[86]}
   );
   gpc606_5 gpc5562 (
      {stage1_48[80], stage1_48[81], stage1_48[82], stage1_48[83], stage1_48[84], stage1_48[85]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[15],stage2_50[25],stage2_49[50],stage2_48[87]}
   );
   gpc606_5 gpc5563 (
      {stage1_48[86], stage1_48[87], stage1_48[88], stage1_48[89], stage1_48[90], stage1_48[91]},
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17]},
      {stage2_52[2],stage2_51[16],stage2_50[26],stage2_49[51],stage2_48[88]}
   );
   gpc606_5 gpc5564 (
      {stage1_48[92], stage1_48[93], stage1_48[94], stage1_48[95], stage1_48[96], stage1_48[97]},
      {stage1_50[18], stage1_50[19], stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23]},
      {stage2_52[3],stage2_51[17],stage2_50[27],stage2_49[52],stage2_48[89]}
   );
   gpc606_5 gpc5565 (
      {stage1_48[98], stage1_48[99], stage1_48[100], stage1_48[101], stage1_48[102], stage1_48[103]},
      {stage1_50[24], stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage2_52[4],stage2_51[18],stage2_50[28],stage2_49[53],stage2_48[90]}
   );
   gpc606_5 gpc5566 (
      {stage1_48[104], stage1_48[105], stage1_48[106], stage1_48[107], stage1_48[108], stage1_48[109]},
      {stage1_50[30], stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35]},
      {stage2_52[5],stage2_51[19],stage2_50[29],stage2_49[54],stage2_48[91]}
   );
   gpc606_5 gpc5567 (
      {stage1_48[110], stage1_48[111], stage1_48[112], stage1_48[113], stage1_48[114], stage1_48[115]},
      {stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage2_52[6],stage2_51[20],stage2_50[30],stage2_49[55],stage2_48[92]}
   );
   gpc606_5 gpc5568 (
      {stage1_48[116], stage1_48[117], stage1_48[118], stage1_48[119], stage1_48[120], stage1_48[121]},
      {stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45], stage1_50[46], stage1_50[47]},
      {stage2_52[7],stage2_51[21],stage2_50[31],stage2_49[56],stage2_48[93]}
   );
   gpc615_5 gpc5569 (
      {stage1_48[122], stage1_48[123], stage1_48[124], stage1_48[125], stage1_48[126]},
      {stage1_49[84]},
      {stage1_50[48], stage1_50[49], stage1_50[50], stage1_50[51], stage1_50[52], stage1_50[53]},
      {stage2_52[8],stage2_51[22],stage2_50[32],stage2_49[57],stage2_48[94]}
   );
   gpc615_5 gpc5570 (
      {stage1_48[127], stage1_48[128], stage1_48[129], stage1_48[130], stage1_48[131]},
      {stage1_49[85]},
      {stage1_50[54], stage1_50[55], stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59]},
      {stage2_52[9],stage2_51[23],stage2_50[33],stage2_49[58],stage2_48[95]}
   );
   gpc615_5 gpc5571 (
      {stage1_48[132], stage1_48[133], stage1_48[134], stage1_48[135], stage1_48[136]},
      {stage1_49[86]},
      {stage1_50[60], stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64], stage1_50[65]},
      {stage2_52[10],stage2_51[24],stage2_50[34],stage2_49[59],stage2_48[96]}
   );
   gpc615_5 gpc5572 (
      {stage1_48[137], stage1_48[138], stage1_48[139], stage1_48[140], stage1_48[141]},
      {stage1_49[87]},
      {stage1_50[66], stage1_50[67], stage1_50[68], stage1_50[69], stage1_50[70], stage1_50[71]},
      {stage2_52[11],stage2_51[25],stage2_50[35],stage2_49[60],stage2_48[97]}
   );
   gpc615_5 gpc5573 (
      {stage1_48[142], stage1_48[143], stage1_48[144], stage1_48[145], stage1_48[146]},
      {stage1_49[88]},
      {stage1_50[72], stage1_50[73], stage1_50[74], stage1_50[75], stage1_50[76], stage1_50[77]},
      {stage2_52[12],stage2_51[26],stage2_50[36],stage2_49[61],stage2_48[98]}
   );
   gpc615_5 gpc5574 (
      {stage1_48[147], stage1_48[148], stage1_48[149], stage1_48[150], stage1_48[151]},
      {stage1_49[89]},
      {stage1_50[78], stage1_50[79], stage1_50[80], stage1_50[81], stage1_50[82], stage1_50[83]},
      {stage2_52[13],stage2_51[27],stage2_50[37],stage2_49[62],stage2_48[99]}
   );
   gpc615_5 gpc5575 (
      {stage1_48[152], stage1_48[153], stage1_48[154], stage1_48[155], stage1_48[156]},
      {stage1_49[90]},
      {stage1_50[84], stage1_50[85], stage1_50[86], stage1_50[87], stage1_50[88], stage1_50[89]},
      {stage2_52[14],stage2_51[28],stage2_50[38],stage2_49[63],stage2_48[100]}
   );
   gpc615_5 gpc5576 (
      {stage1_48[157], stage1_48[158], stage1_48[159], stage1_48[160], stage1_48[161]},
      {stage1_49[91]},
      {stage1_50[90], stage1_50[91], stage1_50[92], stage1_50[93], stage1_50[94], stage1_50[95]},
      {stage2_52[15],stage2_51[29],stage2_50[39],stage2_49[64],stage2_48[101]}
   );
   gpc615_5 gpc5577 (
      {stage1_48[162], stage1_48[163], stage1_48[164], stage1_48[165], stage1_48[166]},
      {stage1_49[92]},
      {stage1_50[96], stage1_50[97], stage1_50[98], stage1_50[99], stage1_50[100], stage1_50[101]},
      {stage2_52[16],stage2_51[30],stage2_50[40],stage2_49[65],stage2_48[102]}
   );
   gpc615_5 gpc5578 (
      {stage1_48[167], stage1_48[168], stage1_48[169], stage1_48[170], stage1_48[171]},
      {stage1_49[93]},
      {stage1_50[102], stage1_50[103], stage1_50[104], stage1_50[105], stage1_50[106], stage1_50[107]},
      {stage2_52[17],stage2_51[31],stage2_50[41],stage2_49[66],stage2_48[103]}
   );
   gpc606_5 gpc5579 (
      {stage1_49[94], stage1_49[95], stage1_49[96], stage1_49[97], stage1_49[98], stage1_49[99]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[18],stage2_51[32],stage2_50[42],stage2_49[67]}
   );
   gpc606_5 gpc5580 (
      {stage1_49[100], stage1_49[101], stage1_49[102], stage1_49[103], stage1_49[104], stage1_49[105]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[19],stage2_51[33],stage2_50[43],stage2_49[68]}
   );
   gpc606_5 gpc5581 (
      {stage1_49[106], stage1_49[107], stage1_49[108], stage1_49[109], stage1_49[110], stage1_49[111]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[20],stage2_51[34],stage2_50[44],stage2_49[69]}
   );
   gpc606_5 gpc5582 (
      {stage1_49[112], stage1_49[113], stage1_49[114], stage1_49[115], stage1_49[116], stage1_49[117]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage2_53[3],stage2_52[21],stage2_51[35],stage2_50[45],stage2_49[70]}
   );
   gpc606_5 gpc5583 (
      {stage1_49[118], stage1_49[119], stage1_49[120], stage1_49[121], stage1_49[122], stage1_49[123]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage2_53[4],stage2_52[22],stage2_51[36],stage2_50[46],stage2_49[71]}
   );
   gpc606_5 gpc5584 (
      {stage1_49[124], stage1_49[125], stage1_49[126], stage1_49[127], stage1_49[128], stage1_49[129]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage2_53[5],stage2_52[23],stage2_51[37],stage2_50[47],stage2_49[72]}
   );
   gpc606_5 gpc5585 (
      {stage1_49[130], stage1_49[131], stage1_49[132], stage1_49[133], stage1_49[134], stage1_49[135]},
      {stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39], stage1_51[40], stage1_51[41]},
      {stage2_53[6],stage2_52[24],stage2_51[38],stage2_50[48],stage2_49[73]}
   );
   gpc606_5 gpc5586 (
      {stage1_49[136], stage1_49[137], stage1_49[138], stage1_49[139], stage1_49[140], stage1_49[141]},
      {stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45], stage1_51[46], stage1_51[47]},
      {stage2_53[7],stage2_52[25],stage2_51[39],stage2_50[49],stage2_49[74]}
   );
   gpc606_5 gpc5587 (
      {stage1_49[142], stage1_49[143], stage1_49[144], stage1_49[145], stage1_49[146], stage1_49[147]},
      {stage1_51[48], stage1_51[49], stage1_51[50], stage1_51[51], stage1_51[52], stage1_51[53]},
      {stage2_53[8],stage2_52[26],stage2_51[40],stage2_50[50],stage2_49[75]}
   );
   gpc606_5 gpc5588 (
      {stage1_49[148], stage1_49[149], stage1_49[150], stage1_49[151], stage1_49[152], stage1_49[153]},
      {stage1_51[54], stage1_51[55], stage1_51[56], stage1_51[57], stage1_51[58], stage1_51[59]},
      {stage2_53[9],stage2_52[27],stage2_51[41],stage2_50[51],stage2_49[76]}
   );
   gpc2135_5 gpc5589 (
      {stage1_50[108], stage1_50[109], stage1_50[110], stage1_50[111], stage1_50[112]},
      {stage1_51[60], stage1_51[61], stage1_51[62]},
      {stage1_52[0]},
      {stage1_53[0], stage1_53[1]},
      {stage2_54[0],stage2_53[10],stage2_52[28],stage2_51[42],stage2_50[52]}
   );
   gpc1163_5 gpc5590 (
      {stage1_50[113], stage1_50[114], stage1_50[115]},
      {stage1_51[63], stage1_51[64], stage1_51[65], stage1_51[66], stage1_51[67], stage1_51[68]},
      {stage1_52[1]},
      {stage1_53[2]},
      {stage2_54[1],stage2_53[11],stage2_52[29],stage2_51[43],stage2_50[53]}
   );
   gpc1163_5 gpc5591 (
      {stage1_50[116], stage1_50[117], stage1_50[118]},
      {stage1_51[69], stage1_51[70], stage1_51[71], stage1_51[72], stage1_51[73], stage1_51[74]},
      {stage1_52[2]},
      {stage1_53[3]},
      {stage2_54[2],stage2_53[12],stage2_52[30],stage2_51[44],stage2_50[54]}
   );
   gpc1163_5 gpc5592 (
      {stage1_50[119], stage1_50[120], stage1_50[121]},
      {stage1_51[75], stage1_51[76], stage1_51[77], stage1_51[78], stage1_51[79], stage1_51[80]},
      {stage1_52[3]},
      {stage1_53[4]},
      {stage2_54[3],stage2_53[13],stage2_52[31],stage2_51[45],stage2_50[55]}
   );
   gpc1163_5 gpc5593 (
      {stage1_50[122], stage1_50[123], stage1_50[124]},
      {stage1_51[81], stage1_51[82], stage1_51[83], stage1_51[84], stage1_51[85], stage1_51[86]},
      {stage1_52[4]},
      {stage1_53[5]},
      {stage2_54[4],stage2_53[14],stage2_52[32],stage2_51[46],stage2_50[56]}
   );
   gpc1163_5 gpc5594 (
      {stage1_50[125], stage1_50[126], stage1_50[127]},
      {stage1_51[87], stage1_51[88], stage1_51[89], stage1_51[90], stage1_51[91], stage1_51[92]},
      {stage1_52[5]},
      {stage1_53[6]},
      {stage2_54[5],stage2_53[15],stage2_52[33],stage2_51[47],stage2_50[57]}
   );
   gpc1163_5 gpc5595 (
      {stage1_50[128], stage1_50[129], stage1_50[130]},
      {stage1_51[93], stage1_51[94], stage1_51[95], stage1_51[96], stage1_51[97], stage1_51[98]},
      {stage1_52[6]},
      {stage1_53[7]},
      {stage2_54[6],stage2_53[16],stage2_52[34],stage2_51[48],stage2_50[58]}
   );
   gpc1163_5 gpc5596 (
      {stage1_50[131], stage1_50[132], stage1_50[133]},
      {stage1_51[99], stage1_51[100], stage1_51[101], stage1_51[102], stage1_51[103], stage1_51[104]},
      {stage1_52[7]},
      {stage1_53[8]},
      {stage2_54[7],stage2_53[17],stage2_52[35],stage2_51[49],stage2_50[59]}
   );
   gpc1163_5 gpc5597 (
      {stage1_50[134], stage1_50[135], stage1_50[136]},
      {stage1_51[105], stage1_51[106], stage1_51[107], stage1_51[108], stage1_51[109], stage1_51[110]},
      {stage1_52[8]},
      {stage1_53[9]},
      {stage2_54[8],stage2_53[18],stage2_52[36],stage2_51[50],stage2_50[60]}
   );
   gpc1163_5 gpc5598 (
      {stage1_50[137], stage1_50[138], stage1_50[139]},
      {stage1_51[111], stage1_51[112], stage1_51[113], stage1_51[114], stage1_51[115], stage1_51[116]},
      {stage1_52[9]},
      {stage1_53[10]},
      {stage2_54[9],stage2_53[19],stage2_52[37],stage2_51[51],stage2_50[61]}
   );
   gpc1163_5 gpc5599 (
      {stage1_50[140], stage1_50[141], stage1_50[142]},
      {stage1_51[117], stage1_51[118], stage1_51[119], stage1_51[120], stage1_51[121], stage1_51[122]},
      {stage1_52[10]},
      {stage1_53[11]},
      {stage2_54[10],stage2_53[20],stage2_52[38],stage2_51[52],stage2_50[62]}
   );
   gpc1163_5 gpc5600 (
      {stage1_50[143], stage1_50[144], stage1_50[145]},
      {stage1_51[123], stage1_51[124], stage1_51[125], stage1_51[126], stage1_51[127], stage1_51[128]},
      {stage1_52[11]},
      {stage1_53[12]},
      {stage2_54[11],stage2_53[21],stage2_52[39],stage2_51[53],stage2_50[63]}
   );
   gpc1163_5 gpc5601 (
      {stage1_50[146], stage1_50[147], stage1_50[148]},
      {stage1_51[129], stage1_51[130], stage1_51[131], stage1_51[132], stage1_51[133], stage1_51[134]},
      {stage1_52[12]},
      {stage1_53[13]},
      {stage2_54[12],stage2_53[22],stage2_52[40],stage2_51[54],stage2_50[64]}
   );
   gpc1163_5 gpc5602 (
      {stage1_50[149], stage1_50[150], stage1_50[151]},
      {stage1_51[135], stage1_51[136], stage1_51[137], stage1_51[138], stage1_51[139], stage1_51[140]},
      {stage1_52[13]},
      {stage1_53[14]},
      {stage2_54[13],stage2_53[23],stage2_52[41],stage2_51[55],stage2_50[65]}
   );
   gpc1163_5 gpc5603 (
      {stage1_50[152], stage1_50[153], stage1_50[154]},
      {stage1_51[141], stage1_51[142], stage1_51[143], stage1_51[144], stage1_51[145], stage1_51[146]},
      {stage1_52[14]},
      {stage1_53[15]},
      {stage2_54[14],stage2_53[24],stage2_52[42],stage2_51[56],stage2_50[66]}
   );
   gpc1163_5 gpc5604 (
      {stage1_50[155], stage1_50[156], stage1_50[157]},
      {stage1_51[147], stage1_51[148], stage1_51[149], stage1_51[150], stage1_51[151], stage1_51[152]},
      {stage1_52[15]},
      {stage1_53[16]},
      {stage2_54[15],stage2_53[25],stage2_52[43],stage2_51[57],stage2_50[67]}
   );
   gpc1163_5 gpc5605 (
      {stage1_50[158], stage1_50[159], stage1_50[160]},
      {stage1_51[153], stage1_51[154], stage1_51[155], stage1_51[156], stage1_51[157], stage1_51[158]},
      {stage1_52[16]},
      {stage1_53[17]},
      {stage2_54[16],stage2_53[26],stage2_52[44],stage2_51[58],stage2_50[68]}
   );
   gpc1163_5 gpc5606 (
      {stage1_50[161], stage1_50[162], stage1_50[163]},
      {stage1_51[159], stage1_51[160], stage1_51[161], stage1_51[162], stage1_51[163], stage1_51[164]},
      {stage1_52[17]},
      {stage1_53[18]},
      {stage2_54[17],stage2_53[27],stage2_52[45],stage2_51[59],stage2_50[69]}
   );
   gpc1163_5 gpc5607 (
      {stage1_50[164], stage1_50[165], stage1_50[166]},
      {stage1_51[165], stage1_51[166], stage1_51[167], stage1_51[168], stage1_51[169], stage1_51[170]},
      {stage1_52[18]},
      {stage1_53[19]},
      {stage2_54[18],stage2_53[28],stage2_52[46],stage2_51[60],stage2_50[70]}
   );
   gpc1163_5 gpc5608 (
      {stage1_50[167], stage1_50[168], stage1_50[169]},
      {stage1_51[171], stage1_51[172], stage1_51[173], stage1_51[174], stage1_51[175], stage1_51[176]},
      {stage1_52[19]},
      {stage1_53[20]},
      {stage2_54[19],stage2_53[29],stage2_52[47],stage2_51[61],stage2_50[71]}
   );
   gpc1163_5 gpc5609 (
      {stage1_50[170], stage1_50[171], stage1_50[172]},
      {stage1_51[177], stage1_51[178], stage1_51[179], stage1_51[180], stage1_51[181], stage1_51[182]},
      {stage1_52[20]},
      {stage1_53[21]},
      {stage2_54[20],stage2_53[30],stage2_52[48],stage2_51[62],stage2_50[72]}
   );
   gpc1163_5 gpc5610 (
      {stage1_50[173], stage1_50[174], stage1_50[175]},
      {stage1_51[183], stage1_51[184], stage1_51[185], stage1_51[186], stage1_51[187], stage1_51[188]},
      {stage1_52[21]},
      {stage1_53[22]},
      {stage2_54[21],stage2_53[31],stage2_52[49],stage2_51[63],stage2_50[73]}
   );
   gpc1163_5 gpc5611 (
      {stage1_50[176], stage1_50[177], stage1_50[178]},
      {stage1_51[189], stage1_51[190], stage1_51[191], stage1_51[192], stage1_51[193], stage1_51[194]},
      {stage1_52[22]},
      {stage1_53[23]},
      {stage2_54[22],stage2_53[32],stage2_52[50],stage2_51[64],stage2_50[74]}
   );
   gpc606_5 gpc5612 (
      {stage1_51[195], stage1_51[196], stage1_51[197], stage1_51[198], stage1_51[199], stage1_51[200]},
      {stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage2_55[0],stage2_54[23],stage2_53[33],stage2_52[51],stage2_51[65]}
   );
   gpc615_5 gpc5613 (
      {stage1_51[201], stage1_51[202], stage1_51[203], stage1_51[204], stage1_51[205]},
      {stage1_52[23]},
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34], stage1_53[35]},
      {stage2_55[1],stage2_54[24],stage2_53[34],stage2_52[52],stage2_51[66]}
   );
   gpc615_5 gpc5614 (
      {stage1_51[206], stage1_51[207], stage1_51[208], stage1_51[209], stage1_51[210]},
      {stage1_52[24]},
      {stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39], stage1_53[40], stage1_53[41]},
      {stage2_55[2],stage2_54[25],stage2_53[35],stage2_52[53],stage2_51[67]}
   );
   gpc615_5 gpc5615 (
      {stage1_51[211], stage1_51[212], stage1_51[213], stage1_51[214], stage1_51[215]},
      {stage1_52[25]},
      {stage1_53[42], stage1_53[43], stage1_53[44], stage1_53[45], stage1_53[46], stage1_53[47]},
      {stage2_55[3],stage2_54[26],stage2_53[36],stage2_52[54],stage2_51[68]}
   );
   gpc615_5 gpc5616 (
      {stage1_51[216], stage1_51[217], stage1_51[218], stage1_51[219], stage1_51[220]},
      {stage1_52[26]},
      {stage1_53[48], stage1_53[49], stage1_53[50], stage1_53[51], stage1_53[52], stage1_53[53]},
      {stage2_55[4],stage2_54[27],stage2_53[37],stage2_52[55],stage2_51[69]}
   );
   gpc615_5 gpc5617 (
      {stage1_51[221], stage1_51[222], stage1_51[223], stage1_51[224], stage1_51[225]},
      {stage1_52[27]},
      {stage1_53[54], stage1_53[55], stage1_53[56], stage1_53[57], stage1_53[58], stage1_53[59]},
      {stage2_55[5],stage2_54[28],stage2_53[38],stage2_52[56],stage2_51[70]}
   );
   gpc615_5 gpc5618 (
      {stage1_51[226], stage1_51[227], stage1_51[228], stage1_51[229], stage1_51[230]},
      {stage1_52[28]},
      {stage1_53[60], stage1_53[61], stage1_53[62], stage1_53[63], stage1_53[64], stage1_53[65]},
      {stage2_55[6],stage2_54[29],stage2_53[39],stage2_52[57],stage2_51[71]}
   );
   gpc615_5 gpc5619 (
      {stage1_51[231], stage1_51[232], stage1_51[233], stage1_51[234], stage1_51[235]},
      {stage1_52[29]},
      {stage1_53[66], stage1_53[67], stage1_53[68], stage1_53[69], stage1_53[70], stage1_53[71]},
      {stage2_55[7],stage2_54[30],stage2_53[40],stage2_52[58],stage2_51[72]}
   );
   gpc615_5 gpc5620 (
      {stage1_51[236], stage1_51[237], stage1_51[238], stage1_51[239], stage1_51[240]},
      {stage1_52[30]},
      {stage1_53[72], stage1_53[73], stage1_53[74], stage1_53[75], stage1_53[76], stage1_53[77]},
      {stage2_55[8],stage2_54[31],stage2_53[41],stage2_52[59],stage2_51[73]}
   );
   gpc615_5 gpc5621 (
      {stage1_51[241], stage1_51[242], stage1_51[243], stage1_51[244], stage1_51[245]},
      {stage1_52[31]},
      {stage1_53[78], stage1_53[79], stage1_53[80], stage1_53[81], stage1_53[82], stage1_53[83]},
      {stage2_55[9],stage2_54[32],stage2_53[42],stage2_52[60],stage2_51[74]}
   );
   gpc615_5 gpc5622 (
      {stage1_51[246], stage1_51[247], stage1_51[248], stage1_51[249], stage1_51[250]},
      {stage1_52[32]},
      {stage1_53[84], stage1_53[85], stage1_53[86], stage1_53[87], stage1_53[88], stage1_53[89]},
      {stage2_55[10],stage2_54[33],stage2_53[43],stage2_52[61],stage2_51[75]}
   );
   gpc615_5 gpc5623 (
      {stage1_51[251], stage1_51[252], stage1_51[253], stage1_51[254], stage1_51[255]},
      {stage1_52[33]},
      {stage1_53[90], stage1_53[91], stage1_53[92], stage1_53[93], stage1_53[94], stage1_53[95]},
      {stage2_55[11],stage2_54[34],stage2_53[44],stage2_52[62],stage2_51[76]}
   );
   gpc615_5 gpc5624 (
      {stage1_51[256], stage1_51[257], stage1_51[258], stage1_51[259], stage1_51[260]},
      {stage1_52[34]},
      {stage1_53[96], stage1_53[97], stage1_53[98], stage1_53[99], stage1_53[100], stage1_53[101]},
      {stage2_55[12],stage2_54[35],stage2_53[45],stage2_52[63],stage2_51[77]}
   );
   gpc615_5 gpc5625 (
      {stage1_51[261], stage1_51[262], stage1_51[263], stage1_51[264], stage1_51[265]},
      {stage1_52[35]},
      {stage1_53[102], stage1_53[103], stage1_53[104], stage1_53[105], stage1_53[106], stage1_53[107]},
      {stage2_55[13],stage2_54[36],stage2_53[46],stage2_52[64],stage2_51[78]}
   );
   gpc606_5 gpc5626 (
      {stage1_52[36], stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[14],stage2_54[37],stage2_53[47],stage2_52[65]}
   );
   gpc606_5 gpc5627 (
      {stage1_52[42], stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[15],stage2_54[38],stage2_53[48],stage2_52[66]}
   );
   gpc606_5 gpc5628 (
      {stage1_52[48], stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[16],stage2_54[39],stage2_53[49],stage2_52[67]}
   );
   gpc606_5 gpc5629 (
      {stage1_52[54], stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[17],stage2_54[40],stage2_53[50],stage2_52[68]}
   );
   gpc606_5 gpc5630 (
      {stage1_52[60], stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64], stage1_52[65]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[18],stage2_54[41],stage2_53[51],stage2_52[69]}
   );
   gpc606_5 gpc5631 (
      {stage1_52[66], stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70], stage1_52[71]},
      {stage1_54[30], stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage2_56[5],stage2_55[19],stage2_54[42],stage2_53[52],stage2_52[70]}
   );
   gpc606_5 gpc5632 (
      {stage1_52[72], stage1_52[73], stage1_52[74], stage1_52[75], stage1_52[76], stage1_52[77]},
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40], stage1_54[41]},
      {stage2_56[6],stage2_55[20],stage2_54[43],stage2_53[53],stage2_52[71]}
   );
   gpc606_5 gpc5633 (
      {stage1_52[78], stage1_52[79], stage1_52[80], stage1_52[81], stage1_52[82], stage1_52[83]},
      {stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46], stage1_54[47]},
      {stage2_56[7],stage2_55[21],stage2_54[44],stage2_53[54],stage2_52[72]}
   );
   gpc606_5 gpc5634 (
      {stage1_52[84], stage1_52[85], stage1_52[86], stage1_52[87], stage1_52[88], stage1_52[89]},
      {stage1_54[48], stage1_54[49], stage1_54[50], stage1_54[51], stage1_54[52], stage1_54[53]},
      {stage2_56[8],stage2_55[22],stage2_54[45],stage2_53[55],stage2_52[73]}
   );
   gpc606_5 gpc5635 (
      {stage1_52[90], stage1_52[91], stage1_52[92], stage1_52[93], stage1_52[94], stage1_52[95]},
      {stage1_54[54], stage1_54[55], stage1_54[56], stage1_54[57], stage1_54[58], stage1_54[59]},
      {stage2_56[9],stage2_55[23],stage2_54[46],stage2_53[56],stage2_52[74]}
   );
   gpc606_5 gpc5636 (
      {stage1_52[96], stage1_52[97], stage1_52[98], stage1_52[99], stage1_52[100], stage1_52[101]},
      {stage1_54[60], stage1_54[61], stage1_54[62], stage1_54[63], stage1_54[64], stage1_54[65]},
      {stage2_56[10],stage2_55[24],stage2_54[47],stage2_53[57],stage2_52[75]}
   );
   gpc615_5 gpc5637 (
      {stage1_52[102], stage1_52[103], stage1_52[104], stage1_52[105], stage1_52[106]},
      {stage1_53[108]},
      {stage1_54[66], stage1_54[67], stage1_54[68], stage1_54[69], stage1_54[70], stage1_54[71]},
      {stage2_56[11],stage2_55[25],stage2_54[48],stage2_53[58],stage2_52[76]}
   );
   gpc615_5 gpc5638 (
      {stage1_52[107], stage1_52[108], stage1_52[109], stage1_52[110], stage1_52[111]},
      {stage1_53[109]},
      {stage1_54[72], stage1_54[73], stage1_54[74], stage1_54[75], stage1_54[76], stage1_54[77]},
      {stage2_56[12],stage2_55[26],stage2_54[49],stage2_53[59],stage2_52[77]}
   );
   gpc615_5 gpc5639 (
      {stage1_52[112], stage1_52[113], stage1_52[114], stage1_52[115], stage1_52[116]},
      {stage1_53[110]},
      {stage1_54[78], stage1_54[79], stage1_54[80], stage1_54[81], stage1_54[82], stage1_54[83]},
      {stage2_56[13],stage2_55[27],stage2_54[50],stage2_53[60],stage2_52[78]}
   );
   gpc615_5 gpc5640 (
      {stage1_52[117], stage1_52[118], stage1_52[119], stage1_52[120], stage1_52[121]},
      {stage1_53[111]},
      {stage1_54[84], stage1_54[85], stage1_54[86], stage1_54[87], stage1_54[88], stage1_54[89]},
      {stage2_56[14],stage2_55[28],stage2_54[51],stage2_53[61],stage2_52[79]}
   );
   gpc615_5 gpc5641 (
      {stage1_52[122], stage1_52[123], stage1_52[124], stage1_52[125], stage1_52[126]},
      {stage1_53[112]},
      {stage1_54[90], stage1_54[91], stage1_54[92], stage1_54[93], stage1_54[94], stage1_54[95]},
      {stage2_56[15],stage2_55[29],stage2_54[52],stage2_53[62],stage2_52[80]}
   );
   gpc615_5 gpc5642 (
      {stage1_52[127], stage1_52[128], stage1_52[129], stage1_52[130], stage1_52[131]},
      {stage1_53[113]},
      {stage1_54[96], stage1_54[97], stage1_54[98], stage1_54[99], stage1_54[100], stage1_54[101]},
      {stage2_56[16],stage2_55[30],stage2_54[53],stage2_53[63],stage2_52[81]}
   );
   gpc615_5 gpc5643 (
      {stage1_52[132], stage1_52[133], stage1_52[134], stage1_52[135], stage1_52[136]},
      {stage1_53[114]},
      {stage1_54[102], stage1_54[103], stage1_54[104], stage1_54[105], stage1_54[106], stage1_54[107]},
      {stage2_56[17],stage2_55[31],stage2_54[54],stage2_53[64],stage2_52[82]}
   );
   gpc615_5 gpc5644 (
      {stage1_52[137], stage1_52[138], stage1_52[139], stage1_52[140], stage1_52[141]},
      {stage1_53[115]},
      {stage1_54[108], stage1_54[109], stage1_54[110], stage1_54[111], stage1_54[112], stage1_54[113]},
      {stage2_56[18],stage2_55[32],stage2_54[55],stage2_53[65],stage2_52[83]}
   );
   gpc615_5 gpc5645 (
      {stage1_52[142], stage1_52[143], stage1_52[144], stage1_52[145], stage1_52[146]},
      {stage1_53[116]},
      {stage1_54[114], stage1_54[115], stage1_54[116], stage1_54[117], stage1_54[118], stage1_54[119]},
      {stage2_56[19],stage2_55[33],stage2_54[56],stage2_53[66],stage2_52[84]}
   );
   gpc615_5 gpc5646 (
      {stage1_52[147], stage1_52[148], stage1_52[149], stage1_52[150], stage1_52[151]},
      {stage1_53[117]},
      {stage1_54[120], stage1_54[121], stage1_54[122], stage1_54[123], stage1_54[124], stage1_54[125]},
      {stage2_56[20],stage2_55[34],stage2_54[57],stage2_53[67],stage2_52[85]}
   );
   gpc615_5 gpc5647 (
      {stage1_52[152], stage1_52[153], stage1_52[154], stage1_52[155], stage1_52[156]},
      {stage1_53[118]},
      {stage1_54[126], stage1_54[127], stage1_54[128], stage1_54[129], stage1_54[130], stage1_54[131]},
      {stage2_56[21],stage2_55[35],stage2_54[58],stage2_53[68],stage2_52[86]}
   );
   gpc615_5 gpc5648 (
      {stage1_52[157], stage1_52[158], stage1_52[159], stage1_52[160], stage1_52[161]},
      {stage1_53[119]},
      {stage1_54[132], stage1_54[133], stage1_54[134], stage1_54[135], stage1_54[136], stage1_54[137]},
      {stage2_56[22],stage2_55[36],stage2_54[59],stage2_53[69],stage2_52[87]}
   );
   gpc615_5 gpc5649 (
      {stage1_52[162], stage1_52[163], stage1_52[164], stage1_52[165], stage1_52[166]},
      {stage1_53[120]},
      {stage1_54[138], stage1_54[139], stage1_54[140], stage1_54[141], stage1_54[142], stage1_54[143]},
      {stage2_56[23],stage2_55[37],stage2_54[60],stage2_53[70],stage2_52[88]}
   );
   gpc615_5 gpc5650 (
      {stage1_52[167], stage1_52[168], stage1_52[169], stage1_52[170], stage1_52[171]},
      {stage1_53[121]},
      {stage1_54[144], stage1_54[145], stage1_54[146], stage1_54[147], stage1_54[148], stage1_54[149]},
      {stage2_56[24],stage2_55[38],stage2_54[61],stage2_53[71],stage2_52[89]}
   );
   gpc615_5 gpc5651 (
      {stage1_52[172], stage1_52[173], stage1_52[174], stage1_52[175], stage1_52[176]},
      {stage1_53[122]},
      {stage1_54[150], stage1_54[151], stage1_54[152], stage1_54[153], stage1_54[154], stage1_54[155]},
      {stage2_56[25],stage2_55[39],stage2_54[62],stage2_53[72],stage2_52[90]}
   );
   gpc615_5 gpc5652 (
      {stage1_52[177], stage1_52[178], stage1_52[179], stage1_52[180], stage1_52[181]},
      {stage1_53[123]},
      {stage1_54[156], stage1_54[157], stage1_54[158], stage1_54[159], stage1_54[160], stage1_54[161]},
      {stage2_56[26],stage2_55[40],stage2_54[63],stage2_53[73],stage2_52[91]}
   );
   gpc615_5 gpc5653 (
      {stage1_52[182], stage1_52[183], stage1_52[184], stage1_52[185], stage1_52[186]},
      {stage1_53[124]},
      {stage1_54[162], stage1_54[163], stage1_54[164], stage1_54[165], stage1_54[166], stage1_54[167]},
      {stage2_56[27],stage2_55[41],stage2_54[64],stage2_53[74],stage2_52[92]}
   );
   gpc615_5 gpc5654 (
      {stage1_53[125], stage1_53[126], stage1_53[127], stage1_53[128], stage1_53[129]},
      {stage1_54[168]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[28],stage2_55[42],stage2_54[65],stage2_53[75]}
   );
   gpc606_5 gpc5655 (
      {stage1_54[169], stage1_54[170], stage1_54[171], stage1_54[172], stage1_54[173], stage1_54[174]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[1],stage2_56[29],stage2_55[43],stage2_54[66]}
   );
   gpc606_5 gpc5656 (
      {stage1_54[175], stage1_54[176], stage1_54[177], stage1_54[178], stage1_54[179], stage1_54[180]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[2],stage2_56[30],stage2_55[44],stage2_54[67]}
   );
   gpc606_5 gpc5657 (
      {stage1_54[181], stage1_54[182], stage1_54[183], stage1_54[184], stage1_54[185], stage1_54[186]},
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage2_58[2],stage2_57[3],stage2_56[31],stage2_55[45],stage2_54[68]}
   );
   gpc606_5 gpc5658 (
      {stage1_54[187], stage1_54[188], stage1_54[189], stage1_54[190], stage1_54[191], stage1_54[192]},
      {stage1_56[18], stage1_56[19], stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage2_58[3],stage2_57[4],stage2_56[32],stage2_55[46],stage2_54[69]}
   );
   gpc615_5 gpc5659 (
      {stage1_54[193], stage1_54[194], stage1_54[195], stage1_54[196], stage1_54[197]},
      {stage1_55[6]},
      {stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage2_58[4],stage2_57[5],stage2_56[33],stage2_55[47],stage2_54[70]}
   );
   gpc615_5 gpc5660 (
      {stage1_54[198], stage1_54[199], stage1_54[200], stage1_54[201], stage1_54[202]},
      {stage1_55[7]},
      {stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage2_58[5],stage2_57[6],stage2_56[34],stage2_55[48],stage2_54[71]}
   );
   gpc2135_5 gpc5661 (
      {stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11], stage1_55[12]},
      {stage1_56[36], stage1_56[37], stage1_56[38]},
      {stage1_57[0]},
      {stage1_58[0], stage1_58[1]},
      {stage2_59[0],stage2_58[6],stage2_57[7],stage2_56[35],stage2_55[49]}
   );
   gpc2135_5 gpc5662 (
      {stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage1_56[39], stage1_56[40], stage1_56[41]},
      {stage1_57[1]},
      {stage1_58[2], stage1_58[3]},
      {stage2_59[1],stage2_58[7],stage2_57[8],stage2_56[36],stage2_55[50]}
   );
   gpc2135_5 gpc5663 (
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22]},
      {stage1_56[42], stage1_56[43], stage1_56[44]},
      {stage1_57[2]},
      {stage1_58[4], stage1_58[5]},
      {stage2_59[2],stage2_58[8],stage2_57[9],stage2_56[37],stage2_55[51]}
   );
   gpc2135_5 gpc5664 (
      {stage1_55[23], stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27]},
      {stage1_56[45], stage1_56[46], stage1_56[47]},
      {stage1_57[3]},
      {stage1_58[6], stage1_58[7]},
      {stage2_59[3],stage2_58[9],stage2_57[10],stage2_56[38],stage2_55[52]}
   );
   gpc2135_5 gpc5665 (
      {stage1_55[28], stage1_55[29], stage1_55[30], stage1_55[31], stage1_55[32]},
      {stage1_56[48], stage1_56[49], stage1_56[50]},
      {stage1_57[4]},
      {stage1_58[8], stage1_58[9]},
      {stage2_59[4],stage2_58[10],stage2_57[11],stage2_56[39],stage2_55[53]}
   );
   gpc2135_5 gpc5666 (
      {stage1_55[33], stage1_55[34], stage1_55[35], stage1_55[36], stage1_55[37]},
      {stage1_56[51], stage1_56[52], stage1_56[53]},
      {stage1_57[5]},
      {stage1_58[10], stage1_58[11]},
      {stage2_59[5],stage2_58[11],stage2_57[12],stage2_56[40],stage2_55[54]}
   );
   gpc2135_5 gpc5667 (
      {stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41], stage1_55[42]},
      {stage1_56[54], stage1_56[55], stage1_56[56]},
      {stage1_57[6]},
      {stage1_58[12], stage1_58[13]},
      {stage2_59[6],stage2_58[12],stage2_57[13],stage2_56[41],stage2_55[55]}
   );
   gpc2135_5 gpc5668 (
      {stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage1_56[57], stage1_56[58], stage1_56[59]},
      {stage1_57[7]},
      {stage1_58[14], stage1_58[15]},
      {stage2_59[7],stage2_58[13],stage2_57[14],stage2_56[42],stage2_55[56]}
   );
   gpc2135_5 gpc5669 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[60], stage1_56[61], stage1_56[62]},
      {stage1_57[8]},
      {stage1_58[16], stage1_58[17]},
      {stage2_59[8],stage2_58[14],stage2_57[15],stage2_56[43],stage2_55[57]}
   );
   gpc2135_5 gpc5670 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[63], stage1_56[64], stage1_56[65]},
      {stage1_57[9]},
      {stage1_58[18], stage1_58[19]},
      {stage2_59[9],stage2_58[15],stage2_57[16],stage2_56[44],stage2_55[58]}
   );
   gpc2135_5 gpc5671 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[66], stage1_56[67], stage1_56[68]},
      {stage1_57[10]},
      {stage1_58[20], stage1_58[21]},
      {stage2_59[10],stage2_58[16],stage2_57[17],stage2_56[45],stage2_55[59]}
   );
   gpc2135_5 gpc5672 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[69], stage1_56[70], stage1_56[71]},
      {stage1_57[11]},
      {stage1_58[22], stage1_58[23]},
      {stage2_59[11],stage2_58[17],stage2_57[18],stage2_56[46],stage2_55[60]}
   );
   gpc2135_5 gpc5673 (
      {stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71], stage1_55[72]},
      {stage1_56[72], stage1_56[73], stage1_56[74]},
      {stage1_57[12]},
      {stage1_58[24], stage1_58[25]},
      {stage2_59[12],stage2_58[18],stage2_57[19],stage2_56[47],stage2_55[61]}
   );
   gpc2135_5 gpc5674 (
      {stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage1_56[75], stage1_56[76], stage1_56[77]},
      {stage1_57[13]},
      {stage1_58[26], stage1_58[27]},
      {stage2_59[13],stage2_58[19],stage2_57[20],stage2_56[48],stage2_55[62]}
   );
   gpc2135_5 gpc5675 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82]},
      {stage1_56[78], stage1_56[79], stage1_56[80]},
      {stage1_57[14]},
      {stage1_58[28], stage1_58[29]},
      {stage2_59[14],stage2_58[20],stage2_57[21],stage2_56[49],stage2_55[63]}
   );
   gpc2135_5 gpc5676 (
      {stage1_55[83], stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87]},
      {stage1_56[81], stage1_56[82], stage1_56[83]},
      {stage1_57[15]},
      {stage1_58[30], stage1_58[31]},
      {stage2_59[15],stage2_58[21],stage2_57[22],stage2_56[50],stage2_55[64]}
   );
   gpc2135_5 gpc5677 (
      {stage1_55[88], stage1_55[89], stage1_55[90], stage1_55[91], stage1_55[92]},
      {stage1_56[84], stage1_56[85], stage1_56[86]},
      {stage1_57[16]},
      {stage1_58[32], stage1_58[33]},
      {stage2_59[16],stage2_58[22],stage2_57[23],stage2_56[51],stage2_55[65]}
   );
   gpc2135_5 gpc5678 (
      {stage1_55[93], stage1_55[94], stage1_55[95], stage1_55[96], stage1_55[97]},
      {stage1_56[87], stage1_56[88], stage1_56[89]},
      {stage1_57[17]},
      {stage1_58[34], stage1_58[35]},
      {stage2_59[17],stage2_58[23],stage2_57[24],stage2_56[52],stage2_55[66]}
   );
   gpc606_5 gpc5679 (
      {stage1_55[98], stage1_55[99], stage1_55[100], stage1_55[101], stage1_55[102], stage1_55[103]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[18],stage2_58[24],stage2_57[25],stage2_56[53],stage2_55[67]}
   );
   gpc606_5 gpc5680 (
      {stage1_55[104], stage1_55[105], stage1_55[106], stage1_55[107], stage1_55[108], stage1_55[109]},
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage2_59[19],stage2_58[25],stage2_57[26],stage2_56[54],stage2_55[68]}
   );
   gpc606_5 gpc5681 (
      {stage1_55[110], stage1_55[111], stage1_55[112], stage1_55[113], stage1_55[114], stage1_55[115]},
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage2_59[20],stage2_58[26],stage2_57[27],stage2_56[55],stage2_55[69]}
   );
   gpc606_5 gpc5682 (
      {stage1_55[116], stage1_55[117], stage1_55[118], stage1_55[119], stage1_55[120], stage1_55[121]},
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage2_59[21],stage2_58[27],stage2_57[28],stage2_56[56],stage2_55[70]}
   );
   gpc606_5 gpc5683 (
      {stage1_55[122], stage1_55[123], stage1_55[124], stage1_55[125], stage1_55[126], stage1_55[127]},
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage2_59[22],stage2_58[28],stage2_57[29],stage2_56[57],stage2_55[71]}
   );
   gpc606_5 gpc5684 (
      {stage1_55[128], stage1_55[129], stage1_55[130], stage1_55[131], stage1_55[132], stage1_55[133]},
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage2_59[23],stage2_58[29],stage2_57[30],stage2_56[58],stage2_55[72]}
   );
   gpc606_5 gpc5685 (
      {stage1_55[134], stage1_55[135], stage1_55[136], stage1_55[137], stage1_55[138], stage1_55[139]},
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage2_59[24],stage2_58[30],stage2_57[31],stage2_56[59],stage2_55[73]}
   );
   gpc606_5 gpc5686 (
      {stage1_55[140], stage1_55[141], stage1_55[142], stage1_55[143], stage1_55[144], stage1_55[145]},
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage2_59[25],stage2_58[31],stage2_57[32],stage2_56[60],stage2_55[74]}
   );
   gpc606_5 gpc5687 (
      {stage1_55[146], stage1_55[147], stage1_55[148], stage1_55[149], stage1_55[150], stage1_55[151]},
      {stage1_57[66], stage1_57[67], stage1_57[68], stage1_57[69], stage1_57[70], stage1_57[71]},
      {stage2_59[26],stage2_58[32],stage2_57[33],stage2_56[61],stage2_55[75]}
   );
   gpc606_5 gpc5688 (
      {stage1_55[152], stage1_55[153], stage1_55[154], stage1_55[155], stage1_55[156], stage1_55[157]},
      {stage1_57[72], stage1_57[73], stage1_57[74], stage1_57[75], stage1_57[76], stage1_57[77]},
      {stage2_59[27],stage2_58[33],stage2_57[34],stage2_56[62],stage2_55[76]}
   );
   gpc606_5 gpc5689 (
      {stage1_55[158], stage1_55[159], stage1_55[160], stage1_55[161], stage1_55[162], stage1_55[163]},
      {stage1_57[78], stage1_57[79], stage1_57[80], stage1_57[81], stage1_57[82], stage1_57[83]},
      {stage2_59[28],stage2_58[34],stage2_57[35],stage2_56[63],stage2_55[77]}
   );
   gpc606_5 gpc5690 (
      {stage1_55[164], stage1_55[165], stage1_55[166], stage1_55[167], stage1_55[168], stage1_55[169]},
      {stage1_57[84], stage1_57[85], stage1_57[86], stage1_57[87], stage1_57[88], stage1_57[89]},
      {stage2_59[29],stage2_58[35],stage2_57[36],stage2_56[64],stage2_55[78]}
   );
   gpc606_5 gpc5691 (
      {stage1_55[170], stage1_55[171], stage1_55[172], stage1_55[173], stage1_55[174], stage1_55[175]},
      {stage1_57[90], stage1_57[91], stage1_57[92], stage1_57[93], stage1_57[94], stage1_57[95]},
      {stage2_59[30],stage2_58[36],stage2_57[37],stage2_56[65],stage2_55[79]}
   );
   gpc606_5 gpc5692 (
      {stage1_55[176], stage1_55[177], stage1_55[178], stage1_55[179], stage1_55[180], stage1_55[181]},
      {stage1_57[96], stage1_57[97], stage1_57[98], stage1_57[99], stage1_57[100], stage1_57[101]},
      {stage2_59[31],stage2_58[37],stage2_57[38],stage2_56[66],stage2_55[80]}
   );
   gpc606_5 gpc5693 (
      {stage1_55[182], stage1_55[183], stage1_55[184], stage1_55[185], stage1_55[186], stage1_55[187]},
      {stage1_57[102], stage1_57[103], stage1_57[104], stage1_57[105], stage1_57[106], stage1_57[107]},
      {stage2_59[32],stage2_58[38],stage2_57[39],stage2_56[67],stage2_55[81]}
   );
   gpc606_5 gpc5694 (
      {stage1_55[188], stage1_55[189], stage1_55[190], stage1_55[191], stage1_55[192], stage1_55[193]},
      {stage1_57[108], stage1_57[109], stage1_57[110], stage1_57[111], stage1_57[112], stage1_57[113]},
      {stage2_59[33],stage2_58[39],stage2_57[40],stage2_56[68],stage2_55[82]}
   );
   gpc606_5 gpc5695 (
      {stage1_55[194], stage1_55[195], stage1_55[196], stage1_55[197], stage1_55[198], stage1_55[199]},
      {stage1_57[114], stage1_57[115], stage1_57[116], stage1_57[117], stage1_57[118], stage1_57[119]},
      {stage2_59[34],stage2_58[40],stage2_57[41],stage2_56[69],stage2_55[83]}
   );
   gpc606_5 gpc5696 (
      {stage1_55[200], stage1_55[201], stage1_55[202], stage1_55[203], stage1_55[204], stage1_55[205]},
      {stage1_57[120], stage1_57[121], stage1_57[122], stage1_57[123], stage1_57[124], stage1_57[125]},
      {stage2_59[35],stage2_58[41],stage2_57[42],stage2_56[70],stage2_55[84]}
   );
   gpc606_5 gpc5697 (
      {stage1_55[206], stage1_55[207], stage1_55[208], stage1_55[209], stage1_55[210], stage1_55[211]},
      {stage1_57[126], stage1_57[127], stage1_57[128], stage1_57[129], stage1_57[130], stage1_57[131]},
      {stage2_59[36],stage2_58[42],stage2_57[43],stage2_56[71],stage2_55[85]}
   );
   gpc606_5 gpc5698 (
      {stage1_55[212], stage1_55[213], stage1_55[214], stage1_55[215], stage1_55[216], stage1_55[217]},
      {stage1_57[132], stage1_57[133], stage1_57[134], stage1_57[135], stage1_57[136], stage1_57[137]},
      {stage2_59[37],stage2_58[43],stage2_57[44],stage2_56[72],stage2_55[86]}
   );
   gpc606_5 gpc5699 (
      {stage1_55[218], stage1_55[219], stage1_55[220], stage1_55[221], stage1_55[222], stage1_55[223]},
      {stage1_57[138], stage1_57[139], stage1_57[140], stage1_57[141], stage1_57[142], stage1_57[143]},
      {stage2_59[38],stage2_58[44],stage2_57[45],stage2_56[73],stage2_55[87]}
   );
   gpc606_5 gpc5700 (
      {stage1_55[224], stage1_55[225], stage1_55[226], stage1_55[227], stage1_55[228], stage1_55[229]},
      {stage1_57[144], stage1_57[145], stage1_57[146], stage1_57[147], stage1_57[148], stage1_57[149]},
      {stage2_59[39],stage2_58[45],stage2_57[46],stage2_56[74],stage2_55[88]}
   );
   gpc606_5 gpc5701 (
      {stage1_55[230], stage1_55[231], stage1_55[232], stage1_55[233], stage1_55[234], stage1_55[235]},
      {stage1_57[150], stage1_57[151], stage1_57[152], stage1_57[153], stage1_57[154], stage1_57[155]},
      {stage2_59[40],stage2_58[46],stage2_57[47],stage2_56[75],stage2_55[89]}
   );
   gpc606_5 gpc5702 (
      {stage1_55[236], stage1_55[237], stage1_55[238], stage1_55[239], stage1_55[240], stage1_55[241]},
      {stage1_57[156], stage1_57[157], stage1_57[158], stage1_57[159], stage1_57[160], stage1_57[161]},
      {stage2_59[41],stage2_58[47],stage2_57[48],stage2_56[76],stage2_55[90]}
   );
   gpc606_5 gpc5703 (
      {stage1_55[242], stage1_55[243], stage1_55[244], stage1_55[245], stage1_55[246], stage1_55[247]},
      {stage1_57[162], stage1_57[163], stage1_57[164], stage1_57[165], stage1_57[166], stage1_57[167]},
      {stage2_59[42],stage2_58[48],stage2_57[49],stage2_56[77],stage2_55[91]}
   );
   gpc606_5 gpc5704 (
      {stage1_55[248], stage1_55[249], stage1_55[250], stage1_55[251], stage1_55[252], stage1_55[253]},
      {stage1_57[168], stage1_57[169], stage1_57[170], stage1_57[171], stage1_57[172], stage1_57[173]},
      {stage2_59[43],stage2_58[49],stage2_57[50],stage2_56[78],stage2_55[92]}
   );
   gpc606_5 gpc5705 (
      {stage1_56[90], stage1_56[91], stage1_56[92], stage1_56[93], stage1_56[94], stage1_56[95]},
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage2_60[0],stage2_59[44],stage2_58[50],stage2_57[51],stage2_56[79]}
   );
   gpc606_5 gpc5706 (
      {stage1_56[96], stage1_56[97], stage1_56[98], stage1_56[99], stage1_56[100], stage1_56[101]},
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage2_60[1],stage2_59[45],stage2_58[51],stage2_57[52],stage2_56[80]}
   );
   gpc606_5 gpc5707 (
      {stage1_56[102], stage1_56[103], stage1_56[104], stage1_56[105], stage1_56[106], stage1_56[107]},
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage2_60[2],stage2_59[46],stage2_58[52],stage2_57[53],stage2_56[81]}
   );
   gpc606_5 gpc5708 (
      {stage1_56[108], stage1_56[109], stage1_56[110], stage1_56[111], stage1_56[112], stage1_56[113]},
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage2_60[3],stage2_59[47],stage2_58[53],stage2_57[54],stage2_56[82]}
   );
   gpc606_5 gpc5709 (
      {stage1_56[114], stage1_56[115], stage1_56[116], stage1_56[117], stage1_56[118], stage1_56[119]},
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64], stage1_58[65]},
      {stage2_60[4],stage2_59[48],stage2_58[54],stage2_57[55],stage2_56[83]}
   );
   gpc606_5 gpc5710 (
      {stage1_56[120], stage1_56[121], stage1_56[122], stage1_56[123], stage1_56[124], stage1_56[125]},
      {stage1_58[66], stage1_58[67], stage1_58[68], stage1_58[69], stage1_58[70], stage1_58[71]},
      {stage2_60[5],stage2_59[49],stage2_58[55],stage2_57[56],stage2_56[84]}
   );
   gpc606_5 gpc5711 (
      {stage1_56[126], stage1_56[127], stage1_56[128], stage1_56[129], stage1_56[130], stage1_56[131]},
      {stage1_58[72], stage1_58[73], stage1_58[74], stage1_58[75], stage1_58[76], stage1_58[77]},
      {stage2_60[6],stage2_59[50],stage2_58[56],stage2_57[57],stage2_56[85]}
   );
   gpc606_5 gpc5712 (
      {stage1_56[132], stage1_56[133], stage1_56[134], stage1_56[135], stage1_56[136], stage1_56[137]},
      {stage1_58[78], stage1_58[79], stage1_58[80], stage1_58[81], stage1_58[82], stage1_58[83]},
      {stage2_60[7],stage2_59[51],stage2_58[57],stage2_57[58],stage2_56[86]}
   );
   gpc606_5 gpc5713 (
      {stage1_56[138], stage1_56[139], stage1_56[140], stage1_56[141], stage1_56[142], stage1_56[143]},
      {stage1_58[84], stage1_58[85], stage1_58[86], stage1_58[87], stage1_58[88], stage1_58[89]},
      {stage2_60[8],stage2_59[52],stage2_58[58],stage2_57[59],stage2_56[87]}
   );
   gpc615_5 gpc5714 (
      {stage1_56[144], stage1_56[145], stage1_56[146], stage1_56[147], stage1_56[148]},
      {stage1_57[174]},
      {stage1_58[90], stage1_58[91], stage1_58[92], stage1_58[93], stage1_58[94], stage1_58[95]},
      {stage2_60[9],stage2_59[53],stage2_58[59],stage2_57[60],stage2_56[88]}
   );
   gpc615_5 gpc5715 (
      {stage1_56[149], stage1_56[150], stage1_56[151], stage1_56[152], stage1_56[153]},
      {stage1_57[175]},
      {stage1_58[96], stage1_58[97], stage1_58[98], stage1_58[99], stage1_58[100], stage1_58[101]},
      {stage2_60[10],stage2_59[54],stage2_58[60],stage2_57[61],stage2_56[89]}
   );
   gpc615_5 gpc5716 (
      {stage1_56[154], stage1_56[155], stage1_56[156], stage1_56[157], stage1_56[158]},
      {stage1_57[176]},
      {stage1_58[102], stage1_58[103], stage1_58[104], stage1_58[105], stage1_58[106], stage1_58[107]},
      {stage2_60[11],stage2_59[55],stage2_58[61],stage2_57[62],stage2_56[90]}
   );
   gpc615_5 gpc5717 (
      {stage1_56[159], stage1_56[160], stage1_56[161], stage1_56[162], stage1_56[163]},
      {stage1_57[177]},
      {stage1_58[108], stage1_58[109], stage1_58[110], stage1_58[111], stage1_58[112], stage1_58[113]},
      {stage2_60[12],stage2_59[56],stage2_58[62],stage2_57[63],stage2_56[91]}
   );
   gpc606_5 gpc5718 (
      {stage1_57[178], stage1_57[179], stage1_57[180], stage1_57[181], stage1_57[182], stage1_57[183]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[13],stage2_59[57],stage2_58[63],stage2_57[64]}
   );
   gpc615_5 gpc5719 (
      {stage1_57[184], stage1_57[185], stage1_57[186], stage1_57[187], stage1_57[188]},
      {stage1_58[114]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[14],stage2_59[58],stage2_58[64],stage2_57[65]}
   );
   gpc615_5 gpc5720 (
      {stage1_58[115], stage1_58[116], stage1_58[117], stage1_58[118], stage1_58[119]},
      {stage1_59[12]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[2],stage2_60[15],stage2_59[59],stage2_58[65]}
   );
   gpc615_5 gpc5721 (
      {stage1_58[120], stage1_58[121], stage1_58[122], stage1_58[123], stage1_58[124]},
      {stage1_59[13]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[3],stage2_60[16],stage2_59[60],stage2_58[66]}
   );
   gpc615_5 gpc5722 (
      {stage1_58[125], stage1_58[126], stage1_58[127], stage1_58[128], stage1_58[129]},
      {stage1_59[14]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[4],stage2_60[17],stage2_59[61],stage2_58[67]}
   );
   gpc615_5 gpc5723 (
      {stage1_58[130], stage1_58[131], stage1_58[132], stage1_58[133], stage1_58[134]},
      {stage1_59[15]},
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage2_62[3],stage2_61[5],stage2_60[18],stage2_59[62],stage2_58[68]}
   );
   gpc615_5 gpc5724 (
      {stage1_58[135], stage1_58[136], stage1_58[137], stage1_58[138], stage1_58[139]},
      {stage1_59[16]},
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage2_62[4],stage2_61[6],stage2_60[19],stage2_59[63],stage2_58[69]}
   );
   gpc615_5 gpc5725 (
      {stage1_58[140], stage1_58[141], stage1_58[142], stage1_58[143], stage1_58[144]},
      {stage1_59[17]},
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage2_62[5],stage2_61[7],stage2_60[20],stage2_59[64],stage2_58[70]}
   );
   gpc615_5 gpc5726 (
      {stage1_58[145], stage1_58[146], stage1_58[147], stage1_58[148], stage1_58[149]},
      {stage1_59[18]},
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage2_62[6],stage2_61[8],stage2_60[21],stage2_59[65],stage2_58[71]}
   );
   gpc615_5 gpc5727 (
      {stage1_58[150], stage1_58[151], stage1_58[152], stage1_58[153], stage1_58[154]},
      {stage1_59[19]},
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage2_62[7],stage2_61[9],stage2_60[22],stage2_59[66],stage2_58[72]}
   );
   gpc615_5 gpc5728 (
      {stage1_58[155], stage1_58[156], stage1_58[157], stage1_58[158], stage1_58[159]},
      {stage1_59[20]},
      {stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51], stage1_60[52], stage1_60[53]},
      {stage2_62[8],stage2_61[10],stage2_60[23],stage2_59[67],stage2_58[73]}
   );
   gpc615_5 gpc5729 (
      {stage1_58[160], stage1_58[161], stage1_58[162], stage1_58[163], stage1_58[164]},
      {stage1_59[21]},
      {stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57], stage1_60[58], stage1_60[59]},
      {stage2_62[9],stage2_61[11],stage2_60[24],stage2_59[68],stage2_58[74]}
   );
   gpc615_5 gpc5730 (
      {stage1_58[165], stage1_58[166], stage1_58[167], stage1_58[168], stage1_58[169]},
      {stage1_59[22]},
      {stage1_60[60], stage1_60[61], stage1_60[62], stage1_60[63], stage1_60[64], stage1_60[65]},
      {stage2_62[10],stage2_61[12],stage2_60[25],stage2_59[69],stage2_58[75]}
   );
   gpc615_5 gpc5731 (
      {stage1_58[170], stage1_58[171], stage1_58[172], stage1_58[173], stage1_58[174]},
      {stage1_59[23]},
      {stage1_60[66], stage1_60[67], stage1_60[68], stage1_60[69], stage1_60[70], stage1_60[71]},
      {stage2_62[11],stage2_61[13],stage2_60[26],stage2_59[70],stage2_58[76]}
   );
   gpc615_5 gpc5732 (
      {stage1_58[175], stage1_58[176], stage1_58[177], stage1_58[178], stage1_58[179]},
      {stage1_59[24]},
      {stage1_60[72], stage1_60[73], stage1_60[74], stage1_60[75], stage1_60[76], stage1_60[77]},
      {stage2_62[12],stage2_61[14],stage2_60[27],stage2_59[71],stage2_58[77]}
   );
   gpc615_5 gpc5733 (
      {stage1_58[180], stage1_58[181], stage1_58[182], stage1_58[183], stage1_58[184]},
      {stage1_59[25]},
      {stage1_60[78], stage1_60[79], stage1_60[80], stage1_60[81], stage1_60[82], stage1_60[83]},
      {stage2_62[13],stage2_61[15],stage2_60[28],stage2_59[72],stage2_58[78]}
   );
   gpc615_5 gpc5734 (
      {stage1_58[185], stage1_58[186], stage1_58[187], stage1_58[188], stage1_58[189]},
      {stage1_59[26]},
      {stage1_60[84], stage1_60[85], stage1_60[86], stage1_60[87], stage1_60[88], stage1_60[89]},
      {stage2_62[14],stage2_61[16],stage2_60[29],stage2_59[73],stage2_58[79]}
   );
   gpc615_5 gpc5735 (
      {stage1_58[190], stage1_58[191], stage1_58[192], stage1_58[193], stage1_58[194]},
      {stage1_59[27]},
      {stage1_60[90], stage1_60[91], stage1_60[92], stage1_60[93], stage1_60[94], stage1_60[95]},
      {stage2_62[15],stage2_61[17],stage2_60[30],stage2_59[74],stage2_58[80]}
   );
   gpc615_5 gpc5736 (
      {stage1_58[195], stage1_58[196], stage1_58[197], stage1_58[198], stage1_58[199]},
      {stage1_59[28]},
      {stage1_60[96], stage1_60[97], stage1_60[98], stage1_60[99], stage1_60[100], stage1_60[101]},
      {stage2_62[16],stage2_61[18],stage2_60[31],stage2_59[75],stage2_58[81]}
   );
   gpc615_5 gpc5737 (
      {stage1_58[200], stage1_58[201], stage1_58[202], stage1_58[203], stage1_58[204]},
      {stage1_59[29]},
      {stage1_60[102], stage1_60[103], stage1_60[104], stage1_60[105], stage1_60[106], stage1_60[107]},
      {stage2_62[17],stage2_61[19],stage2_60[32],stage2_59[76],stage2_58[82]}
   );
   gpc615_5 gpc5738 (
      {stage1_58[205], stage1_58[206], stage1_58[207], stage1_58[208], stage1_58[209]},
      {stage1_59[30]},
      {stage1_60[108], stage1_60[109], stage1_60[110], stage1_60[111], stage1_60[112], stage1_60[113]},
      {stage2_62[18],stage2_61[20],stage2_60[33],stage2_59[77],stage2_58[83]}
   );
   gpc615_5 gpc5739 (
      {stage1_58[210], stage1_58[211], stage1_58[212], stage1_58[213], stage1_58[214]},
      {stage1_59[31]},
      {stage1_60[114], stage1_60[115], stage1_60[116], stage1_60[117], stage1_60[118], stage1_60[119]},
      {stage2_62[19],stage2_61[21],stage2_60[34],stage2_59[78],stage2_58[84]}
   );
   gpc615_5 gpc5740 (
      {stage1_58[215], stage1_58[216], stage1_58[217], stage1_58[218], stage1_58[219]},
      {stage1_59[32]},
      {stage1_60[120], stage1_60[121], stage1_60[122], stage1_60[123], stage1_60[124], stage1_60[125]},
      {stage2_62[20],stage2_61[22],stage2_60[35],stage2_59[79],stage2_58[85]}
   );
   gpc2135_5 gpc5741 (
      {stage1_59[33], stage1_59[34], stage1_59[35], stage1_59[36], stage1_59[37]},
      {stage1_60[126], stage1_60[127], stage1_60[128]},
      {stage1_61[0]},
      {stage1_62[0], stage1_62[1]},
      {stage2_63[0],stage2_62[21],stage2_61[23],stage2_60[36],stage2_59[80]}
   );
   gpc606_5 gpc5742 (
      {stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41], stage1_59[42], stage1_59[43]},
      {stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5], stage1_61[6]},
      {stage2_63[1],stage2_62[22],stage2_61[24],stage2_60[37],stage2_59[81]}
   );
   gpc606_5 gpc5743 (
      {stage1_59[44], stage1_59[45], stage1_59[46], stage1_59[47], stage1_59[48], stage1_59[49]},
      {stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11], stage1_61[12]},
      {stage2_63[2],stage2_62[23],stage2_61[25],stage2_60[38],stage2_59[82]}
   );
   gpc606_5 gpc5744 (
      {stage1_59[50], stage1_59[51], stage1_59[52], stage1_59[53], stage1_59[54], stage1_59[55]},
      {stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17], stage1_61[18]},
      {stage2_63[3],stage2_62[24],stage2_61[26],stage2_60[39],stage2_59[83]}
   );
   gpc606_5 gpc5745 (
      {stage1_59[56], stage1_59[57], stage1_59[58], stage1_59[59], stage1_59[60], stage1_59[61]},
      {stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23], stage1_61[24]},
      {stage2_63[4],stage2_62[25],stage2_61[27],stage2_60[40],stage2_59[84]}
   );
   gpc606_5 gpc5746 (
      {stage1_59[62], stage1_59[63], stage1_59[64], stage1_59[65], stage1_59[66], stage1_59[67]},
      {stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29], stage1_61[30]},
      {stage2_63[5],stage2_62[26],stage2_61[28],stage2_60[41],stage2_59[85]}
   );
   gpc606_5 gpc5747 (
      {stage1_59[68], stage1_59[69], stage1_59[70], stage1_59[71], stage1_59[72], stage1_59[73]},
      {stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35], stage1_61[36]},
      {stage2_63[6],stage2_62[27],stage2_61[29],stage2_60[42],stage2_59[86]}
   );
   gpc606_5 gpc5748 (
      {stage1_59[74], stage1_59[75], stage1_59[76], stage1_59[77], stage1_59[78], stage1_59[79]},
      {stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41], stage1_61[42]},
      {stage2_63[7],stage2_62[28],stage2_61[30],stage2_60[43],stage2_59[87]}
   );
   gpc606_5 gpc5749 (
      {stage1_59[80], stage1_59[81], stage1_59[82], stage1_59[83], stage1_59[84], stage1_59[85]},
      {stage1_61[43], stage1_61[44], stage1_61[45], stage1_61[46], stage1_61[47], stage1_61[48]},
      {stage2_63[8],stage2_62[29],stage2_61[31],stage2_60[44],stage2_59[88]}
   );
   gpc606_5 gpc5750 (
      {stage1_59[86], stage1_59[87], stage1_59[88], stage1_59[89], stage1_59[90], stage1_59[91]},
      {stage1_61[49], stage1_61[50], stage1_61[51], stage1_61[52], stage1_61[53], stage1_61[54]},
      {stage2_63[9],stage2_62[30],stage2_61[32],stage2_60[45],stage2_59[89]}
   );
   gpc606_5 gpc5751 (
      {stage1_59[92], stage1_59[93], stage1_59[94], stage1_59[95], stage1_59[96], stage1_59[97]},
      {stage1_61[55], stage1_61[56], stage1_61[57], stage1_61[58], stage1_61[59], stage1_61[60]},
      {stage2_63[10],stage2_62[31],stage2_61[33],stage2_60[46],stage2_59[90]}
   );
   gpc606_5 gpc5752 (
      {stage1_59[98], stage1_59[99], stage1_59[100], stage1_59[101], stage1_59[102], stage1_59[103]},
      {stage1_61[61], stage1_61[62], stage1_61[63], stage1_61[64], stage1_61[65], stage1_61[66]},
      {stage2_63[11],stage2_62[32],stage2_61[34],stage2_60[47],stage2_59[91]}
   );
   gpc606_5 gpc5753 (
      {stage1_59[104], stage1_59[105], stage1_59[106], stage1_59[107], stage1_59[108], stage1_59[109]},
      {stage1_61[67], stage1_61[68], stage1_61[69], stage1_61[70], stage1_61[71], stage1_61[72]},
      {stage2_63[12],stage2_62[33],stage2_61[35],stage2_60[48],stage2_59[92]}
   );
   gpc606_5 gpc5754 (
      {stage1_59[110], stage1_59[111], stage1_59[112], stage1_59[113], stage1_59[114], stage1_59[115]},
      {stage1_61[73], stage1_61[74], stage1_61[75], stage1_61[76], stage1_61[77], stage1_61[78]},
      {stage2_63[13],stage2_62[34],stage2_61[36],stage2_60[49],stage2_59[93]}
   );
   gpc606_5 gpc5755 (
      {stage1_59[116], stage1_59[117], stage1_59[118], stage1_59[119], stage1_59[120], stage1_59[121]},
      {stage1_61[79], stage1_61[80], stage1_61[81], stage1_61[82], stage1_61[83], stage1_61[84]},
      {stage2_63[14],stage2_62[35],stage2_61[37],stage2_60[50],stage2_59[94]}
   );
   gpc606_5 gpc5756 (
      {stage1_59[122], stage1_59[123], stage1_59[124], stage1_59[125], stage1_59[126], stage1_59[127]},
      {stage1_61[85], stage1_61[86], stage1_61[87], stage1_61[88], stage1_61[89], stage1_61[90]},
      {stage2_63[15],stage2_62[36],stage2_61[38],stage2_60[51],stage2_59[95]}
   );
   gpc606_5 gpc5757 (
      {stage1_59[128], stage1_59[129], stage1_59[130], stage1_59[131], stage1_59[132], stage1_59[133]},
      {stage1_61[91], stage1_61[92], stage1_61[93], stage1_61[94], stage1_61[95], stage1_61[96]},
      {stage2_63[16],stage2_62[37],stage2_61[39],stage2_60[52],stage2_59[96]}
   );
   gpc606_5 gpc5758 (
      {stage1_59[134], stage1_59[135], stage1_59[136], stage1_59[137], stage1_59[138], stage1_59[139]},
      {stage1_61[97], stage1_61[98], stage1_61[99], stage1_61[100], stage1_61[101], stage1_61[102]},
      {stage2_63[17],stage2_62[38],stage2_61[40],stage2_60[53],stage2_59[97]}
   );
   gpc606_5 gpc5759 (
      {stage1_59[140], stage1_59[141], stage1_59[142], stage1_59[143], stage1_59[144], stage1_59[145]},
      {stage1_61[103], stage1_61[104], stage1_61[105], stage1_61[106], stage1_61[107], stage1_61[108]},
      {stage2_63[18],stage2_62[39],stage2_61[41],stage2_60[54],stage2_59[98]}
   );
   gpc606_5 gpc5760 (
      {stage1_59[146], stage1_59[147], stage1_59[148], stage1_59[149], stage1_59[150], stage1_59[151]},
      {stage1_61[109], stage1_61[110], stage1_61[111], stage1_61[112], stage1_61[113], stage1_61[114]},
      {stage2_63[19],stage2_62[40],stage2_61[42],stage2_60[55],stage2_59[99]}
   );
   gpc606_5 gpc5761 (
      {stage1_59[152], stage1_59[153], stage1_59[154], stage1_59[155], stage1_59[156], stage1_59[157]},
      {stage1_61[115], stage1_61[116], stage1_61[117], stage1_61[118], stage1_61[119], stage1_61[120]},
      {stage2_63[20],stage2_62[41],stage2_61[43],stage2_60[56],stage2_59[100]}
   );
   gpc606_5 gpc5762 (
      {stage1_59[158], stage1_59[159], stage1_59[160], stage1_59[161], stage1_59[162], stage1_59[163]},
      {stage1_61[121], stage1_61[122], stage1_61[123], stage1_61[124], stage1_61[125], stage1_61[126]},
      {stage2_63[21],stage2_62[42],stage2_61[44],stage2_60[57],stage2_59[101]}
   );
   gpc606_5 gpc5763 (
      {stage1_59[164], stage1_59[165], stage1_59[166], stage1_59[167], stage1_59[168], stage1_59[169]},
      {stage1_61[127], stage1_61[128], stage1_61[129], stage1_61[130], stage1_61[131], stage1_61[132]},
      {stage2_63[22],stage2_62[43],stage2_61[45],stage2_60[58],stage2_59[102]}
   );
   gpc606_5 gpc5764 (
      {stage1_59[170], stage1_59[171], stage1_59[172], stage1_59[173], stage1_59[174], stage1_59[175]},
      {stage1_61[133], stage1_61[134], stage1_61[135], stage1_61[136], stage1_61[137], stage1_61[138]},
      {stage2_63[23],stage2_62[44],stage2_61[46],stage2_60[59],stage2_59[103]}
   );
   gpc606_5 gpc5765 (
      {stage1_59[176], stage1_59[177], stage1_59[178], stage1_59[179], stage1_59[180], stage1_59[181]},
      {stage1_61[139], stage1_61[140], stage1_61[141], stage1_61[142], stage1_61[143], stage1_61[144]},
      {stage2_63[24],stage2_62[45],stage2_61[47],stage2_60[60],stage2_59[104]}
   );
   gpc606_5 gpc5766 (
      {stage1_59[182], stage1_59[183], stage1_59[184], stage1_59[185], stage1_59[186], stage1_59[187]},
      {stage1_61[145], stage1_61[146], stage1_61[147], stage1_61[148], stage1_61[149], stage1_61[150]},
      {stage2_63[25],stage2_62[46],stage2_61[48],stage2_60[61],stage2_59[105]}
   );
   gpc606_5 gpc5767 (
      {stage1_59[188], stage1_59[189], stage1_59[190], stage1_59[191], stage1_59[192], stage1_59[193]},
      {stage1_61[151], stage1_61[152], stage1_61[153], stage1_61[154], stage1_61[155], stage1_61[156]},
      {stage2_63[26],stage2_62[47],stage2_61[49],stage2_60[62],stage2_59[106]}
   );
   gpc606_5 gpc5768 (
      {stage1_59[194], stage1_59[195], stage1_59[196], stage1_59[197], stage1_59[198], stage1_59[199]},
      {stage1_61[157], stage1_61[158], stage1_61[159], stage1_61[160], stage1_61[161], stage1_61[162]},
      {stage2_63[27],stage2_62[48],stage2_61[50],stage2_60[63],stage2_59[107]}
   );
   gpc615_5 gpc5769 (
      {stage1_59[200], stage1_59[201], stage1_59[202], stage1_59[203], stage1_59[204]},
      {stage1_60[129]},
      {stage1_61[163], stage1_61[164], stage1_61[165], stage1_61[166], stage1_61[167], stage1_61[168]},
      {stage2_63[28],stage2_62[49],stage2_61[51],stage2_60[64],stage2_59[108]}
   );
   gpc606_5 gpc5770 (
      {stage1_60[130], stage1_60[131], stage1_60[132], stage1_60[133], stage1_60[134], stage1_60[135]},
      {stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5], stage1_62[6], stage1_62[7]},
      {stage2_64[0],stage2_63[29],stage2_62[50],stage2_61[52],stage2_60[65]}
   );
   gpc606_5 gpc5771 (
      {stage1_60[136], stage1_60[137], stage1_60[138], stage1_60[139], stage1_60[140], stage1_60[141]},
      {stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11], stage1_62[12], stage1_62[13]},
      {stage2_64[1],stage2_63[30],stage2_62[51],stage2_61[53],stage2_60[66]}
   );
   gpc606_5 gpc5772 (
      {stage1_60[142], stage1_60[143], stage1_60[144], stage1_60[145], stage1_60[146], stage1_60[147]},
      {stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17], stage1_62[18], stage1_62[19]},
      {stage2_64[2],stage2_63[31],stage2_62[52],stage2_61[54],stage2_60[67]}
   );
   gpc606_5 gpc5773 (
      {stage1_60[148], stage1_60[149], stage1_60[150], stage1_60[151], stage1_60[152], stage1_60[153]},
      {stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23], stage1_62[24], stage1_62[25]},
      {stage2_64[3],stage2_63[32],stage2_62[53],stage2_61[55],stage2_60[68]}
   );
   gpc606_5 gpc5774 (
      {stage1_60[154], stage1_60[155], stage1_60[156], stage1_60[157], stage1_60[158], stage1_60[159]},
      {stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29], stage1_62[30], stage1_62[31]},
      {stage2_64[4],stage2_63[33],stage2_62[54],stage2_61[56],stage2_60[69]}
   );
   gpc606_5 gpc5775 (
      {stage1_60[160], stage1_60[161], stage1_60[162], stage1_60[163], stage1_60[164], stage1_60[165]},
      {stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35], stage1_62[36], stage1_62[37]},
      {stage2_64[5],stage2_63[34],stage2_62[55],stage2_61[57],stage2_60[70]}
   );
   gpc606_5 gpc5776 (
      {stage1_60[166], stage1_60[167], stage1_60[168], stage1_60[169], stage1_60[170], stage1_60[171]},
      {stage1_62[38], stage1_62[39], stage1_62[40], stage1_62[41], stage1_62[42], stage1_62[43]},
      {stage2_64[6],stage2_63[35],stage2_62[56],stage2_61[58],stage2_60[71]}
   );
   gpc606_5 gpc5777 (
      {stage1_60[172], stage1_60[173], stage1_60[174], stage1_60[175], stage1_60[176], stage1_60[177]},
      {stage1_62[44], stage1_62[45], stage1_62[46], stage1_62[47], stage1_62[48], stage1_62[49]},
      {stage2_64[7],stage2_63[36],stage2_62[57],stage2_61[59],stage2_60[72]}
   );
   gpc606_5 gpc5778 (
      {stage1_60[178], stage1_60[179], stage1_60[180], stage1_60[181], stage1_60[182], stage1_60[183]},
      {stage1_62[50], stage1_62[51], stage1_62[52], stage1_62[53], stage1_62[54], stage1_62[55]},
      {stage2_64[8],stage2_63[37],stage2_62[58],stage2_61[60],stage2_60[73]}
   );
   gpc615_5 gpc5779 (
      {stage1_60[184], stage1_60[185], stage1_60[186], stage1_60[187], stage1_60[188]},
      {stage1_61[169]},
      {stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59], stage1_62[60], stage1_62[61]},
      {stage2_64[9],stage2_63[38],stage2_62[59],stage2_61[61],stage2_60[74]}
   );
   gpc615_5 gpc5780 (
      {stage1_60[189], stage1_60[190], stage1_60[191], stage1_60[192], stage1_60[193]},
      {stage1_61[170]},
      {stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65], stage1_62[66], stage1_62[67]},
      {stage2_64[10],stage2_63[39],stage2_62[60],stage2_61[62],stage2_60[75]}
   );
   gpc615_5 gpc5781 (
      {stage1_60[194], stage1_60[195], stage1_60[196], stage1_60[197], stage1_60[198]},
      {stage1_61[171]},
      {stage1_62[68], stage1_62[69], stage1_62[70], stage1_62[71], stage1_62[72], stage1_62[73]},
      {stage2_64[11],stage2_63[40],stage2_62[61],stage2_61[63],stage2_60[76]}
   );
   gpc615_5 gpc5782 (
      {stage1_60[199], stage1_60[200], stage1_60[201], stage1_60[202], stage1_60[203]},
      {stage1_61[172]},
      {stage1_62[74], stage1_62[75], stage1_62[76], stage1_62[77], stage1_62[78], stage1_62[79]},
      {stage2_64[12],stage2_63[41],stage2_62[62],stage2_61[64],stage2_60[77]}
   );
   gpc615_5 gpc5783 (
      {stage1_60[204], stage1_60[205], stage1_60[206], stage1_60[207], stage1_60[208]},
      {stage1_61[173]},
      {stage1_62[80], stage1_62[81], stage1_62[82], stage1_62[83], stage1_62[84], stage1_62[85]},
      {stage2_64[13],stage2_63[42],stage2_62[63],stage2_61[65],stage2_60[78]}
   );
   gpc615_5 gpc5784 (
      {stage1_61[174], stage1_61[175], stage1_61[176], stage1_61[177], stage1_61[178]},
      {stage1_62[86]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[14],stage2_63[43],stage2_62[64],stage2_61[66]}
   );
   gpc615_5 gpc5785 (
      {stage1_61[179], stage1_61[180], stage1_61[181], stage1_61[182], stage1_61[183]},
      {stage1_62[87]},
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage2_65[1],stage2_64[15],stage2_63[44],stage2_62[65],stage2_61[67]}
   );
   gpc615_5 gpc5786 (
      {stage1_61[184], stage1_61[185], stage1_61[186], stage1_61[187], stage1_61[188]},
      {stage1_62[88]},
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage2_65[2],stage2_64[16],stage2_63[45],stage2_62[66],stage2_61[68]}
   );
   gpc615_5 gpc5787 (
      {stage1_61[189], stage1_61[190], stage1_61[191], stage1_61[192], stage1_61[193]},
      {stage1_62[89]},
      {stage1_63[18], stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage2_65[3],stage2_64[17],stage2_63[46],stage2_62[67],stage2_61[69]}
   );
   gpc615_5 gpc5788 (
      {stage1_61[194], stage1_61[195], stage1_61[196], stage1_61[197], stage1_61[198]},
      {stage1_62[90]},
      {stage1_63[24], stage1_63[25], stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29]},
      {stage2_65[4],stage2_64[18],stage2_63[47],stage2_62[68],stage2_61[70]}
   );
   gpc615_5 gpc5789 (
      {stage1_61[199], stage1_61[200], stage1_61[201], stage1_61[202], stage1_61[203]},
      {stage1_62[91]},
      {stage1_63[30], stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage2_65[5],stage2_64[19],stage2_63[48],stage2_62[69],stage2_61[71]}
   );
   gpc615_5 gpc5790 (
      {stage1_61[204], stage1_61[205], stage1_61[206], stage1_61[207], stage1_61[208]},
      {stage1_62[92]},
      {stage1_63[36], stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41]},
      {stage2_65[6],stage2_64[20],stage2_63[49],stage2_62[70],stage2_61[72]}
   );
   gpc615_5 gpc5791 (
      {stage1_61[209], stage1_61[210], stage1_61[211], stage1_61[212], stage1_61[213]},
      {stage1_62[93]},
      {stage1_63[42], stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47]},
      {stage2_65[7],stage2_64[21],stage2_63[50],stage2_62[71],stage2_61[73]}
   );
   gpc615_5 gpc5792 (
      {stage1_61[214], stage1_61[215], stage1_61[216], stage1_61[217], stage1_61[218]},
      {stage1_62[94]},
      {stage1_63[48], stage1_63[49], stage1_63[50], stage1_63[51], stage1_63[52], stage1_63[53]},
      {stage2_65[8],stage2_64[22],stage2_63[51],stage2_62[72],stage2_61[74]}
   );
   gpc1163_5 gpc5793 (
      {stage1_62[95], stage1_62[96], stage1_62[97]},
      {stage1_63[54], stage1_63[55], stage1_63[56], stage1_63[57], stage1_63[58], stage1_63[59]},
      {stage1_64[0]},
      {stage1_65[0]},
      {stage2_66[0],stage2_65[9],stage2_64[23],stage2_63[52],stage2_62[73]}
   );
   gpc1163_5 gpc5794 (
      {stage1_62[98], stage1_62[99], stage1_62[100]},
      {stage1_63[60], stage1_63[61], stage1_63[62], stage1_63[63], stage1_63[64], stage1_63[65]},
      {stage1_64[1]},
      {stage1_65[1]},
      {stage2_66[1],stage2_65[10],stage2_64[24],stage2_63[53],stage2_62[74]}
   );
   gpc1163_5 gpc5795 (
      {stage1_62[101], stage1_62[102], stage1_62[103]},
      {stage1_63[66], stage1_63[67], stage1_63[68], stage1_63[69], stage1_63[70], stage1_63[71]},
      {stage1_64[2]},
      {stage1_65[2]},
      {stage2_66[2],stage2_65[11],stage2_64[25],stage2_63[54],stage2_62[75]}
   );
   gpc1163_5 gpc5796 (
      {stage1_62[104], stage1_62[105], stage1_62[106]},
      {stage1_63[72], stage1_63[73], stage1_63[74], stage1_63[75], stage1_63[76], stage1_63[77]},
      {stage1_64[3]},
      {stage1_65[3]},
      {stage2_66[3],stage2_65[12],stage2_64[26],stage2_63[55],stage2_62[76]}
   );
   gpc1163_5 gpc5797 (
      {stage1_62[107], stage1_62[108], stage1_62[109]},
      {stage1_63[78], stage1_63[79], stage1_63[80], stage1_63[81], stage1_63[82], stage1_63[83]},
      {stage1_64[4]},
      {stage1_65[4]},
      {stage2_66[4],stage2_65[13],stage2_64[27],stage2_63[56],stage2_62[77]}
   );
   gpc1163_5 gpc5798 (
      {stage1_62[110], stage1_62[111], stage1_62[112]},
      {stage1_63[84], stage1_63[85], stage1_63[86], stage1_63[87], stage1_63[88], stage1_63[89]},
      {stage1_64[5]},
      {stage1_65[5]},
      {stage2_66[5],stage2_65[14],stage2_64[28],stage2_63[57],stage2_62[78]}
   );
   gpc1163_5 gpc5799 (
      {stage1_62[113], stage1_62[114], stage1_62[115]},
      {stage1_63[90], stage1_63[91], stage1_63[92], stage1_63[93], stage1_63[94], stage1_63[95]},
      {stage1_64[6]},
      {stage1_65[6]},
      {stage2_66[6],stage2_65[15],stage2_64[29],stage2_63[58],stage2_62[79]}
   );
   gpc1163_5 gpc5800 (
      {stage1_62[116], stage1_62[117], stage1_62[118]},
      {stage1_63[96], stage1_63[97], stage1_63[98], stage1_63[99], stage1_63[100], stage1_63[101]},
      {stage1_64[7]},
      {stage1_65[7]},
      {stage2_66[7],stage2_65[16],stage2_64[30],stage2_63[59],stage2_62[80]}
   );
   gpc1163_5 gpc5801 (
      {stage1_62[119], stage1_62[120], stage1_62[121]},
      {stage1_63[102], stage1_63[103], stage1_63[104], stage1_63[105], stage1_63[106], stage1_63[107]},
      {stage1_64[8]},
      {stage1_65[8]},
      {stage2_66[8],stage2_65[17],stage2_64[31],stage2_63[60],stage2_62[81]}
   );
   gpc1163_5 gpc5802 (
      {stage1_62[122], stage1_62[123], stage1_62[124]},
      {stage1_63[108], stage1_63[109], stage1_63[110], stage1_63[111], stage1_63[112], stage1_63[113]},
      {stage1_64[9]},
      {stage1_65[9]},
      {stage2_66[9],stage2_65[18],stage2_64[32],stage2_63[61],stage2_62[82]}
   );
   gpc1163_5 gpc5803 (
      {stage1_62[125], stage1_62[126], stage1_62[127]},
      {stage1_63[114], stage1_63[115], stage1_63[116], stage1_63[117], stage1_63[118], stage1_63[119]},
      {stage1_64[10]},
      {stage1_65[10]},
      {stage2_66[10],stage2_65[19],stage2_64[33],stage2_63[62],stage2_62[83]}
   );
   gpc1163_5 gpc5804 (
      {stage1_62[128], stage1_62[129], stage1_62[130]},
      {stage1_63[120], stage1_63[121], stage1_63[122], stage1_63[123], stage1_63[124], stage1_63[125]},
      {stage1_64[11]},
      {stage1_65[11]},
      {stage2_66[11],stage2_65[20],stage2_64[34],stage2_63[63],stage2_62[84]}
   );
   gpc1163_5 gpc5805 (
      {stage1_62[131], stage1_62[132], stage1_62[133]},
      {stage1_63[126], stage1_63[127], stage1_63[128], stage1_63[129], stage1_63[130], stage1_63[131]},
      {stage1_64[12]},
      {stage1_65[12]},
      {stage2_66[12],stage2_65[21],stage2_64[35],stage2_63[64],stage2_62[85]}
   );
   gpc1163_5 gpc5806 (
      {stage1_62[134], stage1_62[135], stage1_62[136]},
      {stage1_63[132], stage1_63[133], stage1_63[134], stage1_63[135], stage1_63[136], stage1_63[137]},
      {stage1_64[13]},
      {stage1_65[13]},
      {stage2_66[13],stage2_65[22],stage2_64[36],stage2_63[65],stage2_62[86]}
   );
   gpc1163_5 gpc5807 (
      {stage1_62[137], stage1_62[138], stage1_62[139]},
      {stage1_63[138], stage1_63[139], stage1_63[140], stage1_63[141], stage1_63[142], stage1_63[143]},
      {stage1_64[14]},
      {stage1_65[14]},
      {stage2_66[14],stage2_65[23],stage2_64[37],stage2_63[66],stage2_62[87]}
   );
   gpc1163_5 gpc5808 (
      {stage1_62[140], stage1_62[141], stage1_62[142]},
      {stage1_63[144], stage1_63[145], stage1_63[146], stage1_63[147], stage1_63[148], stage1_63[149]},
      {stage1_64[15]},
      {stage1_65[15]},
      {stage2_66[15],stage2_65[24],stage2_64[38],stage2_63[67],stage2_62[88]}
   );
   gpc1163_5 gpc5809 (
      {stage1_62[143], stage1_62[144], stage1_62[145]},
      {stage1_63[150], stage1_63[151], stage1_63[152], stage1_63[153], stage1_63[154], stage1_63[155]},
      {stage1_64[16]},
      {stage1_65[16]},
      {stage2_66[16],stage2_65[25],stage2_64[39],stage2_63[68],stage2_62[89]}
   );
   gpc1163_5 gpc5810 (
      {stage1_62[146], stage1_62[147], stage1_62[148]},
      {stage1_63[156], stage1_63[157], stage1_63[158], stage1_63[159], stage1_63[160], stage1_63[161]},
      {stage1_64[17]},
      {stage1_65[17]},
      {stage2_66[17],stage2_65[26],stage2_64[40],stage2_63[69],stage2_62[90]}
   );
   gpc1163_5 gpc5811 (
      {stage1_62[149], stage1_62[150], stage1_62[151]},
      {stage1_63[162], stage1_63[163], stage1_63[164], stage1_63[165], stage1_63[166], stage1_63[167]},
      {stage1_64[18]},
      {stage1_65[18]},
      {stage2_66[18],stage2_65[27],stage2_64[41],stage2_63[70],stage2_62[91]}
   );
   gpc1163_5 gpc5812 (
      {stage1_62[152], stage1_62[153], stage1_62[154]},
      {stage1_63[168], stage1_63[169], stage1_63[170], stage1_63[171], stage1_63[172], stage1_63[173]},
      {stage1_64[19]},
      {stage1_65[19]},
      {stage2_66[19],stage2_65[28],stage2_64[42],stage2_63[71],stage2_62[92]}
   );
   gpc1163_5 gpc5813 (
      {stage1_62[155], stage1_62[156], stage1_62[157]},
      {stage1_63[174], stage1_63[175], stage1_63[176], stage1_63[177], stage1_63[178], stage1_63[179]},
      {stage1_64[20]},
      {stage1_65[20]},
      {stage2_66[20],stage2_65[29],stage2_64[43],stage2_63[72],stage2_62[93]}
   );
   gpc1163_5 gpc5814 (
      {stage1_62[158], stage1_62[159], stage1_62[160]},
      {stage1_63[180], stage1_63[181], stage1_63[182], stage1_63[183], stage1_63[184], stage1_63[185]},
      {stage1_64[21]},
      {stage1_65[21]},
      {stage2_66[21],stage2_65[30],stage2_64[44],stage2_63[73],stage2_62[94]}
   );
   gpc1163_5 gpc5815 (
      {stage1_62[161], stage1_62[162], stage1_62[163]},
      {stage1_63[186], stage1_63[187], stage1_63[188], stage1_63[189], stage1_63[190], stage1_63[191]},
      {stage1_64[22]},
      {stage1_65[22]},
      {stage2_66[22],stage2_65[31],stage2_64[45],stage2_63[74],stage2_62[95]}
   );
   gpc1163_5 gpc5816 (
      {stage1_62[164], stage1_62[165], stage1_62[166]},
      {stage1_63[192], stage1_63[193], stage1_63[194], stage1_63[195], stage1_63[196], stage1_63[197]},
      {stage1_64[23]},
      {stage1_65[23]},
      {stage2_66[23],stage2_65[32],stage2_64[46],stage2_63[75],stage2_62[96]}
   );
   gpc1163_5 gpc5817 (
      {stage1_62[167], stage1_62[168], stage1_62[169]},
      {stage1_63[198], stage1_63[199], stage1_63[200], stage1_63[201], stage1_63[202], stage1_63[203]},
      {stage1_64[24]},
      {stage1_65[24]},
      {stage2_66[24],stage2_65[33],stage2_64[47],stage2_63[76],stage2_62[97]}
   );
   gpc1163_5 gpc5818 (
      {stage1_62[170], stage1_62[171], stage1_62[172]},
      {stage1_63[204], stage1_63[205], stage1_63[206], stage1_63[207], stage1_63[208], stage1_63[209]},
      {stage1_64[25]},
      {stage1_65[25]},
      {stage2_66[25],stage2_65[34],stage2_64[48],stage2_63[77],stage2_62[98]}
   );
   gpc1163_5 gpc5819 (
      {stage1_62[173], stage1_62[174], stage1_62[175]},
      {stage1_63[210], stage1_63[211], stage1_63[212], stage1_63[213], stage1_63[214], stage1_63[215]},
      {stage1_64[26]},
      {stage1_65[26]},
      {stage2_66[26],stage2_65[35],stage2_64[49],stage2_63[78],stage2_62[99]}
   );
   gpc1163_5 gpc5820 (
      {stage1_62[176], stage1_62[177], stage1_62[178]},
      {stage1_63[216], stage1_63[217], stage1_63[218], stage1_63[219], stage1_63[220], stage1_63[221]},
      {stage1_64[27]},
      {stage1_65[27]},
      {stage2_66[27],stage2_65[36],stage2_64[50],stage2_63[79],stage2_62[100]}
   );
   gpc1163_5 gpc5821 (
      {stage1_62[179], stage1_62[180], stage1_62[181]},
      {stage1_63[222], stage1_63[223], stage1_63[224], stage1_63[225], stage1_63[226], stage1_63[227]},
      {stage1_64[28]},
      {stage1_65[28]},
      {stage2_66[28],stage2_65[37],stage2_64[51],stage2_63[80],stage2_62[101]}
   );
   gpc615_5 gpc5822 (
      {stage1_62[182], stage1_62[183], stage1_62[184], stage1_62[185], stage1_62[186]},
      {stage1_63[228]},
      {stage1_64[29], stage1_64[30], stage1_64[31], stage1_64[32], stage1_64[33], stage1_64[34]},
      {stage2_66[29],stage2_65[38],stage2_64[52],stage2_63[81],stage2_62[102]}
   );
   gpc615_5 gpc5823 (
      {stage1_62[187], stage1_62[188], stage1_62[189], stage1_62[190], stage1_62[191]},
      {stage1_63[229]},
      {stage1_64[35], stage1_64[36], stage1_64[37], stage1_64[38], stage1_64[39], stage1_64[40]},
      {stage2_66[30],stage2_65[39],stage2_64[53],stage2_63[82],stage2_62[103]}
   );
   gpc135_4 gpc5824 (
      {stage1_63[230], stage1_63[231], stage1_63[232], stage1_63[233], stage1_63[234]},
      {stage1_64[41], stage1_64[42], stage1_64[43]},
      {stage1_65[29]},
      {stage2_66[31],stage2_65[40],stage2_64[54],stage2_63[83]}
   );
   gpc135_4 gpc5825 (
      {stage1_63[235], stage1_63[236], stage1_63[237], stage1_63[238], stage1_63[239]},
      {stage1_64[44], stage1_64[45], stage1_64[46]},
      {stage1_65[30]},
      {stage2_66[32],stage2_65[41],stage2_64[55],stage2_63[84]}
   );
   gpc207_4 gpc5826 (
      {stage1_63[240], stage1_63[241], stage1_63[242], stage1_63[243], stage1_63[244], stage1_63[245], stage1_63[246]},
      {stage1_65[31], stage1_65[32]},
      {stage2_66[33],stage2_65[42],stage2_64[56],stage2_63[85]}
   );
   gpc207_4 gpc5827 (
      {stage1_63[247], stage1_63[248], stage1_63[249], stage1_63[250], stage1_63[251], stage1_63[252], stage1_63[253]},
      {stage1_65[33], stage1_65[34]},
      {stage2_66[34],stage2_65[43],stage2_64[57],stage2_63[86]}
   );
   gpc207_4 gpc5828 (
      {stage1_63[254], stage1_63[255], stage1_63[256], stage1_63[257], stage1_63[258], stage1_63[259], stage1_63[260]},
      {stage1_65[35], stage1_65[36]},
      {stage2_66[35],stage2_65[44],stage2_64[58],stage2_63[87]}
   );
   gpc207_4 gpc5829 (
      {stage1_63[261], stage1_63[262], stage1_63[263], stage1_63[264], stage1_63[265], stage1_63[266], stage1_63[267]},
      {stage1_65[37], stage1_65[38]},
      {stage2_66[36],stage2_65[45],stage2_64[59],stage2_63[88]}
   );
   gpc207_4 gpc5830 (
      {stage1_63[268], stage1_63[269], stage1_63[270], stage1_63[271], stage1_63[272], stage1_63[273], stage1_63[274]},
      {stage1_65[39], stage1_65[40]},
      {stage2_66[37],stage2_65[46],stage2_64[60],stage2_63[89]}
   );
   gpc207_4 gpc5831 (
      {stage1_63[275], stage1_63[276], stage1_63[277], stage1_63[278], stage1_63[279], stage1_63[280], stage1_63[281]},
      {stage1_65[41], stage1_65[42]},
      {stage2_66[38],stage2_65[47],stage2_64[61],stage2_63[90]}
   );
   gpc207_4 gpc5832 (
      {stage1_63[282], stage1_63[283], stage1_63[284], stage1_63[285], stage1_63[286], stage1_63[287], stage1_63[288]},
      {stage1_65[43], stage1_65[44]},
      {stage2_66[39],stage2_65[48],stage2_64[62],stage2_63[91]}
   );
   gpc207_4 gpc5833 (
      {stage1_63[289], stage1_63[290], stage1_63[291], stage1_63[292], stage1_63[293], stage1_63[294], stage1_63[295]},
      {stage1_65[45], stage1_65[46]},
      {stage2_66[40],stage2_65[49],stage2_64[63],stage2_63[92]}
   );
   gpc207_4 gpc5834 (
      {stage1_63[296], stage1_63[297], stage1_63[298], stage1_63[299], stage1_63[300], stage1_63[301], stage1_63[302]},
      {stage1_65[47], stage1_65[48]},
      {stage2_66[41],stage2_65[50],stage2_64[64],stage2_63[93]}
   );
   gpc1_1 gpc5835 (
      {stage1_0[108]},
      {stage2_0[21]}
   );
   gpc1_1 gpc5836 (
      {stage1_0[109]},
      {stage2_0[22]}
   );
   gpc1_1 gpc5837 (
      {stage1_0[110]},
      {stage2_0[23]}
   );
   gpc1_1 gpc5838 (
      {stage1_0[111]},
      {stage2_0[24]}
   );
   gpc1_1 gpc5839 (
      {stage1_0[112]},
      {stage2_0[25]}
   );
   gpc1_1 gpc5840 (
      {stage1_0[113]},
      {stage2_0[26]}
   );
   gpc1_1 gpc5841 (
      {stage1_0[114]},
      {stage2_0[27]}
   );
   gpc1_1 gpc5842 (
      {stage1_0[115]},
      {stage2_0[28]}
   );
   gpc1_1 gpc5843 (
      {stage1_0[116]},
      {stage2_0[29]}
   );
   gpc1_1 gpc5844 (
      {stage1_0[117]},
      {stage2_0[30]}
   );
   gpc1_1 gpc5845 (
      {stage1_0[118]},
      {stage2_0[31]}
   );
   gpc1_1 gpc5846 (
      {stage1_0[119]},
      {stage2_0[32]}
   );
   gpc1_1 gpc5847 (
      {stage1_0[120]},
      {stage2_0[33]}
   );
   gpc1_1 gpc5848 (
      {stage1_0[121]},
      {stage2_0[34]}
   );
   gpc1_1 gpc5849 (
      {stage1_0[122]},
      {stage2_0[35]}
   );
   gpc1_1 gpc5850 (
      {stage1_0[123]},
      {stage2_0[36]}
   );
   gpc1_1 gpc5851 (
      {stage1_0[124]},
      {stage2_0[37]}
   );
   gpc1_1 gpc5852 (
      {stage1_1[168]},
      {stage2_1[46]}
   );
   gpc1_1 gpc5853 (
      {stage1_1[169]},
      {stage2_1[47]}
   );
   gpc1_1 gpc5854 (
      {stage1_1[170]},
      {stage2_1[48]}
   );
   gpc1_1 gpc5855 (
      {stage1_1[171]},
      {stage2_1[49]}
   );
   gpc1_1 gpc5856 (
      {stage1_1[172]},
      {stage2_1[50]}
   );
   gpc1_1 gpc5857 (
      {stage1_1[173]},
      {stage2_1[51]}
   );
   gpc1_1 gpc5858 (
      {stage1_1[174]},
      {stage2_1[52]}
   );
   gpc1_1 gpc5859 (
      {stage1_1[175]},
      {stage2_1[53]}
   );
   gpc1_1 gpc5860 (
      {stage1_2[144]},
      {stage2_2[49]}
   );
   gpc1_1 gpc5861 (
      {stage1_2[145]},
      {stage2_2[50]}
   );
   gpc1_1 gpc5862 (
      {stage1_2[146]},
      {stage2_2[51]}
   );
   gpc1_1 gpc5863 (
      {stage1_2[147]},
      {stage2_2[52]}
   );
   gpc1_1 gpc5864 (
      {stage1_2[148]},
      {stage2_2[53]}
   );
   gpc1_1 gpc5865 (
      {stage1_2[149]},
      {stage2_2[54]}
   );
   gpc1_1 gpc5866 (
      {stage1_2[150]},
      {stage2_2[55]}
   );
   gpc1_1 gpc5867 (
      {stage1_2[151]},
      {stage2_2[56]}
   );
   gpc1_1 gpc5868 (
      {stage1_2[152]},
      {stage2_2[57]}
   );
   gpc1_1 gpc5869 (
      {stage1_2[153]},
      {stage2_2[58]}
   );
   gpc1_1 gpc5870 (
      {stage1_2[154]},
      {stage2_2[59]}
   );
   gpc1_1 gpc5871 (
      {stage1_2[155]},
      {stage2_2[60]}
   );
   gpc1_1 gpc5872 (
      {stage1_2[156]},
      {stage2_2[61]}
   );
   gpc1_1 gpc5873 (
      {stage1_2[157]},
      {stage2_2[62]}
   );
   gpc1_1 gpc5874 (
      {stage1_3[150]},
      {stage2_3[49]}
   );
   gpc1_1 gpc5875 (
      {stage1_3[151]},
      {stage2_3[50]}
   );
   gpc1_1 gpc5876 (
      {stage1_3[152]},
      {stage2_3[51]}
   );
   gpc1_1 gpc5877 (
      {stage1_3[153]},
      {stage2_3[52]}
   );
   gpc1_1 gpc5878 (
      {stage1_3[154]},
      {stage2_3[53]}
   );
   gpc1_1 gpc5879 (
      {stage1_3[155]},
      {stage2_3[54]}
   );
   gpc1_1 gpc5880 (
      {stage1_3[156]},
      {stage2_3[55]}
   );
   gpc1_1 gpc5881 (
      {stage1_3[157]},
      {stage2_3[56]}
   );
   gpc1_1 gpc5882 (
      {stage1_3[158]},
      {stage2_3[57]}
   );
   gpc1_1 gpc5883 (
      {stage1_3[159]},
      {stage2_3[58]}
   );
   gpc1_1 gpc5884 (
      {stage1_3[160]},
      {stage2_3[59]}
   );
   gpc1_1 gpc5885 (
      {stage1_3[161]},
      {stage2_3[60]}
   );
   gpc1_1 gpc5886 (
      {stage1_3[162]},
      {stage2_3[61]}
   );
   gpc1_1 gpc5887 (
      {stage1_3[163]},
      {stage2_3[62]}
   );
   gpc1_1 gpc5888 (
      {stage1_3[164]},
      {stage2_3[63]}
   );
   gpc1_1 gpc5889 (
      {stage1_3[165]},
      {stage2_3[64]}
   );
   gpc1_1 gpc5890 (
      {stage1_3[166]},
      {stage2_3[65]}
   );
   gpc1_1 gpc5891 (
      {stage1_3[167]},
      {stage2_3[66]}
   );
   gpc1_1 gpc5892 (
      {stage1_3[168]},
      {stage2_3[67]}
   );
   gpc1_1 gpc5893 (
      {stage1_3[169]},
      {stage2_3[68]}
   );
   gpc1_1 gpc5894 (
      {stage1_3[170]},
      {stage2_3[69]}
   );
   gpc1_1 gpc5895 (
      {stage1_3[171]},
      {stage2_3[70]}
   );
   gpc1_1 gpc5896 (
      {stage1_3[172]},
      {stage2_3[71]}
   );
   gpc1_1 gpc5897 (
      {stage1_3[173]},
      {stage2_3[72]}
   );
   gpc1_1 gpc5898 (
      {stage1_3[174]},
      {stage2_3[73]}
   );
   gpc1_1 gpc5899 (
      {stage1_3[175]},
      {stage2_3[74]}
   );
   gpc1_1 gpc5900 (
      {stage1_3[176]},
      {stage2_3[75]}
   );
   gpc1_1 gpc5901 (
      {stage1_3[177]},
      {stage2_3[76]}
   );
   gpc1_1 gpc5902 (
      {stage1_3[178]},
      {stage2_3[77]}
   );
   gpc1_1 gpc5903 (
      {stage1_3[179]},
      {stage2_3[78]}
   );
   gpc1_1 gpc5904 (
      {stage1_3[180]},
      {stage2_3[79]}
   );
   gpc1_1 gpc5905 (
      {stage1_3[181]},
      {stage2_3[80]}
   );
   gpc1_1 gpc5906 (
      {stage1_3[182]},
      {stage2_3[81]}
   );
   gpc1_1 gpc5907 (
      {stage1_3[183]},
      {stage2_3[82]}
   );
   gpc1_1 gpc5908 (
      {stage1_3[184]},
      {stage2_3[83]}
   );
   gpc1_1 gpc5909 (
      {stage1_3[185]},
      {stage2_3[84]}
   );
   gpc1_1 gpc5910 (
      {stage1_3[186]},
      {stage2_3[85]}
   );
   gpc1_1 gpc5911 (
      {stage1_3[187]},
      {stage2_3[86]}
   );
   gpc1_1 gpc5912 (
      {stage1_3[188]},
      {stage2_3[87]}
   );
   gpc1_1 gpc5913 (
      {stage1_3[189]},
      {stage2_3[88]}
   );
   gpc1_1 gpc5914 (
      {stage1_3[190]},
      {stage2_3[89]}
   );
   gpc1_1 gpc5915 (
      {stage1_3[191]},
      {stage2_3[90]}
   );
   gpc1_1 gpc5916 (
      {stage1_3[192]},
      {stage2_3[91]}
   );
   gpc1_1 gpc5917 (
      {stage1_3[193]},
      {stage2_3[92]}
   );
   gpc1_1 gpc5918 (
      {stage1_3[194]},
      {stage2_3[93]}
   );
   gpc1_1 gpc5919 (
      {stage1_3[195]},
      {stage2_3[94]}
   );
   gpc1_1 gpc5920 (
      {stage1_3[196]},
      {stage2_3[95]}
   );
   gpc1_1 gpc5921 (
      {stage1_3[197]},
      {stage2_3[96]}
   );
   gpc1_1 gpc5922 (
      {stage1_3[198]},
      {stage2_3[97]}
   );
   gpc1_1 gpc5923 (
      {stage1_3[199]},
      {stage2_3[98]}
   );
   gpc1_1 gpc5924 (
      {stage1_3[200]},
      {stage2_3[99]}
   );
   gpc1_1 gpc5925 (
      {stage1_3[201]},
      {stage2_3[100]}
   );
   gpc1_1 gpc5926 (
      {stage1_3[202]},
      {stage2_3[101]}
   );
   gpc1_1 gpc5927 (
      {stage1_3[203]},
      {stage2_3[102]}
   );
   gpc1_1 gpc5928 (
      {stage1_3[204]},
      {stage2_3[103]}
   );
   gpc1_1 gpc5929 (
      {stage1_3[205]},
      {stage2_3[104]}
   );
   gpc1_1 gpc5930 (
      {stage1_3[206]},
      {stage2_3[105]}
   );
   gpc1_1 gpc5931 (
      {stage1_3[207]},
      {stage2_3[106]}
   );
   gpc1_1 gpc5932 (
      {stage1_3[208]},
      {stage2_3[107]}
   );
   gpc1_1 gpc5933 (
      {stage1_3[209]},
      {stage2_3[108]}
   );
   gpc1_1 gpc5934 (
      {stage1_3[210]},
      {stage2_3[109]}
   );
   gpc1_1 gpc5935 (
      {stage1_3[211]},
      {stage2_3[110]}
   );
   gpc1_1 gpc5936 (
      {stage1_3[212]},
      {stage2_3[111]}
   );
   gpc1_1 gpc5937 (
      {stage1_3[213]},
      {stage2_3[112]}
   );
   gpc1_1 gpc5938 (
      {stage1_3[214]},
      {stage2_3[113]}
   );
   gpc1_1 gpc5939 (
      {stage1_4[195]},
      {stage2_4[79]}
   );
   gpc1_1 gpc5940 (
      {stage1_4[196]},
      {stage2_4[80]}
   );
   gpc1_1 gpc5941 (
      {stage1_4[197]},
      {stage2_4[81]}
   );
   gpc1_1 gpc5942 (
      {stage1_4[198]},
      {stage2_4[82]}
   );
   gpc1_1 gpc5943 (
      {stage1_4[199]},
      {stage2_4[83]}
   );
   gpc1_1 gpc5944 (
      {stage1_4[200]},
      {stage2_4[84]}
   );
   gpc1_1 gpc5945 (
      {stage1_4[201]},
      {stage2_4[85]}
   );
   gpc1_1 gpc5946 (
      {stage1_4[202]},
      {stage2_4[86]}
   );
   gpc1_1 gpc5947 (
      {stage1_4[203]},
      {stage2_4[87]}
   );
   gpc1_1 gpc5948 (
      {stage1_4[204]},
      {stage2_4[88]}
   );
   gpc1_1 gpc5949 (
      {stage1_4[205]},
      {stage2_4[89]}
   );
   gpc1_1 gpc5950 (
      {stage1_4[206]},
      {stage2_4[90]}
   );
   gpc1_1 gpc5951 (
      {stage1_4[207]},
      {stage2_4[91]}
   );
   gpc1_1 gpc5952 (
      {stage1_4[208]},
      {stage2_4[92]}
   );
   gpc1_1 gpc5953 (
      {stage1_4[209]},
      {stage2_4[93]}
   );
   gpc1_1 gpc5954 (
      {stage1_4[210]},
      {stage2_4[94]}
   );
   gpc1_1 gpc5955 (
      {stage1_4[211]},
      {stage2_4[95]}
   );
   gpc1_1 gpc5956 (
      {stage1_4[212]},
      {stage2_4[96]}
   );
   gpc1_1 gpc5957 (
      {stage1_4[213]},
      {stage2_4[97]}
   );
   gpc1_1 gpc5958 (
      {stage1_4[214]},
      {stage2_4[98]}
   );
   gpc1_1 gpc5959 (
      {stage1_4[215]},
      {stage2_4[99]}
   );
   gpc1_1 gpc5960 (
      {stage1_4[216]},
      {stage2_4[100]}
   );
   gpc1_1 gpc5961 (
      {stage1_4[217]},
      {stage2_4[101]}
   );
   gpc1_1 gpc5962 (
      {stage1_4[218]},
      {stage2_4[102]}
   );
   gpc1_1 gpc5963 (
      {stage1_4[219]},
      {stage2_4[103]}
   );
   gpc1_1 gpc5964 (
      {stage1_4[220]},
      {stage2_4[104]}
   );
   gpc1_1 gpc5965 (
      {stage1_4[221]},
      {stage2_4[105]}
   );
   gpc1_1 gpc5966 (
      {stage1_4[222]},
      {stage2_4[106]}
   );
   gpc1_1 gpc5967 (
      {stage1_4[223]},
      {stage2_4[107]}
   );
   gpc1_1 gpc5968 (
      {stage1_4[224]},
      {stage2_4[108]}
   );
   gpc1_1 gpc5969 (
      {stage1_4[225]},
      {stage2_4[109]}
   );
   gpc1_1 gpc5970 (
      {stage1_4[226]},
      {stage2_4[110]}
   );
   gpc1_1 gpc5971 (
      {stage1_4[227]},
      {stage2_4[111]}
   );
   gpc1_1 gpc5972 (
      {stage1_5[124]},
      {stage2_5[78]}
   );
   gpc1_1 gpc5973 (
      {stage1_5[125]},
      {stage2_5[79]}
   );
   gpc1_1 gpc5974 (
      {stage1_5[126]},
      {stage2_5[80]}
   );
   gpc1_1 gpc5975 (
      {stage1_5[127]},
      {stage2_5[81]}
   );
   gpc1_1 gpc5976 (
      {stage1_5[128]},
      {stage2_5[82]}
   );
   gpc1_1 gpc5977 (
      {stage1_5[129]},
      {stage2_5[83]}
   );
   gpc1_1 gpc5978 (
      {stage1_5[130]},
      {stage2_5[84]}
   );
   gpc1_1 gpc5979 (
      {stage1_5[131]},
      {stage2_5[85]}
   );
   gpc1_1 gpc5980 (
      {stage1_5[132]},
      {stage2_5[86]}
   );
   gpc1_1 gpc5981 (
      {stage1_5[133]},
      {stage2_5[87]}
   );
   gpc1_1 gpc5982 (
      {stage1_5[134]},
      {stage2_5[88]}
   );
   gpc1_1 gpc5983 (
      {stage1_5[135]},
      {stage2_5[89]}
   );
   gpc1_1 gpc5984 (
      {stage1_5[136]},
      {stage2_5[90]}
   );
   gpc1_1 gpc5985 (
      {stage1_5[137]},
      {stage2_5[91]}
   );
   gpc1_1 gpc5986 (
      {stage1_5[138]},
      {stage2_5[92]}
   );
   gpc1_1 gpc5987 (
      {stage1_5[139]},
      {stage2_5[93]}
   );
   gpc1_1 gpc5988 (
      {stage1_5[140]},
      {stage2_5[94]}
   );
   gpc1_1 gpc5989 (
      {stage1_5[141]},
      {stage2_5[95]}
   );
   gpc1_1 gpc5990 (
      {stage1_5[142]},
      {stage2_5[96]}
   );
   gpc1_1 gpc5991 (
      {stage1_5[143]},
      {stage2_5[97]}
   );
   gpc1_1 gpc5992 (
      {stage1_5[144]},
      {stage2_5[98]}
   );
   gpc1_1 gpc5993 (
      {stage1_5[145]},
      {stage2_5[99]}
   );
   gpc1_1 gpc5994 (
      {stage1_5[146]},
      {stage2_5[100]}
   );
   gpc1_1 gpc5995 (
      {stage1_5[147]},
      {stage2_5[101]}
   );
   gpc1_1 gpc5996 (
      {stage1_5[148]},
      {stage2_5[102]}
   );
   gpc1_1 gpc5997 (
      {stage1_5[149]},
      {stage2_5[103]}
   );
   gpc1_1 gpc5998 (
      {stage1_5[150]},
      {stage2_5[104]}
   );
   gpc1_1 gpc5999 (
      {stage1_5[151]},
      {stage2_5[105]}
   );
   gpc1_1 gpc6000 (
      {stage1_5[152]},
      {stage2_5[106]}
   );
   gpc1_1 gpc6001 (
      {stage1_5[153]},
      {stage2_5[107]}
   );
   gpc1_1 gpc6002 (
      {stage1_5[154]},
      {stage2_5[108]}
   );
   gpc1_1 gpc6003 (
      {stage1_5[155]},
      {stage2_5[109]}
   );
   gpc1_1 gpc6004 (
      {stage1_5[156]},
      {stage2_5[110]}
   );
   gpc1_1 gpc6005 (
      {stage1_5[157]},
      {stage2_5[111]}
   );
   gpc1_1 gpc6006 (
      {stage1_5[158]},
      {stage2_5[112]}
   );
   gpc1_1 gpc6007 (
      {stage1_5[159]},
      {stage2_5[113]}
   );
   gpc1_1 gpc6008 (
      {stage1_5[160]},
      {stage2_5[114]}
   );
   gpc1_1 gpc6009 (
      {stage1_5[161]},
      {stage2_5[115]}
   );
   gpc1_1 gpc6010 (
      {stage1_5[162]},
      {stage2_5[116]}
   );
   gpc1_1 gpc6011 (
      {stage1_5[163]},
      {stage2_5[117]}
   );
   gpc1_1 gpc6012 (
      {stage1_5[164]},
      {stage2_5[118]}
   );
   gpc1_1 gpc6013 (
      {stage1_5[165]},
      {stage2_5[119]}
   );
   gpc1_1 gpc6014 (
      {stage1_5[166]},
      {stage2_5[120]}
   );
   gpc1_1 gpc6015 (
      {stage1_5[167]},
      {stage2_5[121]}
   );
   gpc1_1 gpc6016 (
      {stage1_5[168]},
      {stage2_5[122]}
   );
   gpc1_1 gpc6017 (
      {stage1_5[169]},
      {stage2_5[123]}
   );
   gpc1_1 gpc6018 (
      {stage1_5[170]},
      {stage2_5[124]}
   );
   gpc1_1 gpc6019 (
      {stage1_5[171]},
      {stage2_5[125]}
   );
   gpc1_1 gpc6020 (
      {stage1_5[172]},
      {stage2_5[126]}
   );
   gpc1_1 gpc6021 (
      {stage1_5[173]},
      {stage2_5[127]}
   );
   gpc1_1 gpc6022 (
      {stage1_5[174]},
      {stage2_5[128]}
   );
   gpc1_1 gpc6023 (
      {stage1_5[175]},
      {stage2_5[129]}
   );
   gpc1_1 gpc6024 (
      {stage1_5[176]},
      {stage2_5[130]}
   );
   gpc1_1 gpc6025 (
      {stage1_5[177]},
      {stage2_5[131]}
   );
   gpc1_1 gpc6026 (
      {stage1_5[178]},
      {stage2_5[132]}
   );
   gpc1_1 gpc6027 (
      {stage1_5[179]},
      {stage2_5[133]}
   );
   gpc1_1 gpc6028 (
      {stage1_5[180]},
      {stage2_5[134]}
   );
   gpc1_1 gpc6029 (
      {stage1_5[181]},
      {stage2_5[135]}
   );
   gpc1_1 gpc6030 (
      {stage1_5[182]},
      {stage2_5[136]}
   );
   gpc1_1 gpc6031 (
      {stage1_5[183]},
      {stage2_5[137]}
   );
   gpc1_1 gpc6032 (
      {stage1_5[184]},
      {stage2_5[138]}
   );
   gpc1_1 gpc6033 (
      {stage1_5[185]},
      {stage2_5[139]}
   );
   gpc1_1 gpc6034 (
      {stage1_5[186]},
      {stage2_5[140]}
   );
   gpc1_1 gpc6035 (
      {stage1_5[187]},
      {stage2_5[141]}
   );
   gpc1_1 gpc6036 (
      {stage1_5[188]},
      {stage2_5[142]}
   );
   gpc1_1 gpc6037 (
      {stage1_5[189]},
      {stage2_5[143]}
   );
   gpc1_1 gpc6038 (
      {stage1_5[190]},
      {stage2_5[144]}
   );
   gpc1_1 gpc6039 (
      {stage1_5[191]},
      {stage2_5[145]}
   );
   gpc1_1 gpc6040 (
      {stage1_5[192]},
      {stage2_5[146]}
   );
   gpc1_1 gpc6041 (
      {stage1_5[193]},
      {stage2_5[147]}
   );
   gpc1_1 gpc6042 (
      {stage1_5[194]},
      {stage2_5[148]}
   );
   gpc1_1 gpc6043 (
      {stage1_5[195]},
      {stage2_5[149]}
   );
   gpc1_1 gpc6044 (
      {stage1_5[196]},
      {stage2_5[150]}
   );
   gpc1_1 gpc6045 (
      {stage1_5[197]},
      {stage2_5[151]}
   );
   gpc1_1 gpc6046 (
      {stage1_6[175]},
      {stage2_6[53]}
   );
   gpc1_1 gpc6047 (
      {stage1_6[176]},
      {stage2_6[54]}
   );
   gpc1_1 gpc6048 (
      {stage1_6[177]},
      {stage2_6[55]}
   );
   gpc1_1 gpc6049 (
      {stage1_6[178]},
      {stage2_6[56]}
   );
   gpc1_1 gpc6050 (
      {stage1_6[179]},
      {stage2_6[57]}
   );
   gpc1_1 gpc6051 (
      {stage1_6[180]},
      {stage2_6[58]}
   );
   gpc1_1 gpc6052 (
      {stage1_6[181]},
      {stage2_6[59]}
   );
   gpc1_1 gpc6053 (
      {stage1_6[182]},
      {stage2_6[60]}
   );
   gpc1_1 gpc6054 (
      {stage1_6[183]},
      {stage2_6[61]}
   );
   gpc1_1 gpc6055 (
      {stage1_6[184]},
      {stage2_6[62]}
   );
   gpc1_1 gpc6056 (
      {stage1_6[185]},
      {stage2_6[63]}
   );
   gpc1_1 gpc6057 (
      {stage1_6[186]},
      {stage2_6[64]}
   );
   gpc1_1 gpc6058 (
      {stage1_6[187]},
      {stage2_6[65]}
   );
   gpc1_1 gpc6059 (
      {stage1_6[188]},
      {stage2_6[66]}
   );
   gpc1_1 gpc6060 (
      {stage1_6[189]},
      {stage2_6[67]}
   );
   gpc1_1 gpc6061 (
      {stage1_6[190]},
      {stage2_6[68]}
   );
   gpc1_1 gpc6062 (
      {stage1_6[191]},
      {stage2_6[69]}
   );
   gpc1_1 gpc6063 (
      {stage1_6[192]},
      {stage2_6[70]}
   );
   gpc1_1 gpc6064 (
      {stage1_6[193]},
      {stage2_6[71]}
   );
   gpc1_1 gpc6065 (
      {stage1_6[194]},
      {stage2_6[72]}
   );
   gpc1_1 gpc6066 (
      {stage1_6[195]},
      {stage2_6[73]}
   );
   gpc1_1 gpc6067 (
      {stage1_6[196]},
      {stage2_6[74]}
   );
   gpc1_1 gpc6068 (
      {stage1_6[197]},
      {stage2_6[75]}
   );
   gpc1_1 gpc6069 (
      {stage1_6[198]},
      {stage2_6[76]}
   );
   gpc1_1 gpc6070 (
      {stage1_6[199]},
      {stage2_6[77]}
   );
   gpc1_1 gpc6071 (
      {stage1_6[200]},
      {stage2_6[78]}
   );
   gpc1_1 gpc6072 (
      {stage1_6[201]},
      {stage2_6[79]}
   );
   gpc1_1 gpc6073 (
      {stage1_6[202]},
      {stage2_6[80]}
   );
   gpc1_1 gpc6074 (
      {stage1_6[203]},
      {stage2_6[81]}
   );
   gpc1_1 gpc6075 (
      {stage1_6[204]},
      {stage2_6[82]}
   );
   gpc1_1 gpc6076 (
      {stage1_6[205]},
      {stage2_6[83]}
   );
   gpc1_1 gpc6077 (
      {stage1_6[206]},
      {stage2_6[84]}
   );
   gpc1_1 gpc6078 (
      {stage1_6[207]},
      {stage2_6[85]}
   );
   gpc1_1 gpc6079 (
      {stage1_6[208]},
      {stage2_6[86]}
   );
   gpc1_1 gpc6080 (
      {stage1_6[209]},
      {stage2_6[87]}
   );
   gpc1_1 gpc6081 (
      {stage1_6[210]},
      {stage2_6[88]}
   );
   gpc1_1 gpc6082 (
      {stage1_6[211]},
      {stage2_6[89]}
   );
   gpc1_1 gpc6083 (
      {stage1_6[212]},
      {stage2_6[90]}
   );
   gpc1_1 gpc6084 (
      {stage1_6[213]},
      {stage2_6[91]}
   );
   gpc1_1 gpc6085 (
      {stage1_7[217]},
      {stage2_7[69]}
   );
   gpc1_1 gpc6086 (
      {stage1_7[218]},
      {stage2_7[70]}
   );
   gpc1_1 gpc6087 (
      {stage1_7[219]},
      {stage2_7[71]}
   );
   gpc1_1 gpc6088 (
      {stage1_7[220]},
      {stage2_7[72]}
   );
   gpc1_1 gpc6089 (
      {stage1_8[134]},
      {stage2_8[88]}
   );
   gpc1_1 gpc6090 (
      {stage1_8[135]},
      {stage2_8[89]}
   );
   gpc1_1 gpc6091 (
      {stage1_8[136]},
      {stage2_8[90]}
   );
   gpc1_1 gpc6092 (
      {stage1_8[137]},
      {stage2_8[91]}
   );
   gpc1_1 gpc6093 (
      {stage1_8[138]},
      {stage2_8[92]}
   );
   gpc1_1 gpc6094 (
      {stage1_8[139]},
      {stage2_8[93]}
   );
   gpc1_1 gpc6095 (
      {stage1_8[140]},
      {stage2_8[94]}
   );
   gpc1_1 gpc6096 (
      {stage1_8[141]},
      {stage2_8[95]}
   );
   gpc1_1 gpc6097 (
      {stage1_8[142]},
      {stage2_8[96]}
   );
   gpc1_1 gpc6098 (
      {stage1_8[143]},
      {stage2_8[97]}
   );
   gpc1_1 gpc6099 (
      {stage1_8[144]},
      {stage2_8[98]}
   );
   gpc1_1 gpc6100 (
      {stage1_8[145]},
      {stage2_8[99]}
   );
   gpc1_1 gpc6101 (
      {stage1_8[146]},
      {stage2_8[100]}
   );
   gpc1_1 gpc6102 (
      {stage1_8[147]},
      {stage2_8[101]}
   );
   gpc1_1 gpc6103 (
      {stage1_8[148]},
      {stage2_8[102]}
   );
   gpc1_1 gpc6104 (
      {stage1_8[149]},
      {stage2_8[103]}
   );
   gpc1_1 gpc6105 (
      {stage1_8[150]},
      {stage2_8[104]}
   );
   gpc1_1 gpc6106 (
      {stage1_8[151]},
      {stage2_8[105]}
   );
   gpc1_1 gpc6107 (
      {stage1_8[152]},
      {stage2_8[106]}
   );
   gpc1_1 gpc6108 (
      {stage1_8[153]},
      {stage2_8[107]}
   );
   gpc1_1 gpc6109 (
      {stage1_8[154]},
      {stage2_8[108]}
   );
   gpc1_1 gpc6110 (
      {stage1_8[155]},
      {stage2_8[109]}
   );
   gpc1_1 gpc6111 (
      {stage1_8[156]},
      {stage2_8[110]}
   );
   gpc1_1 gpc6112 (
      {stage1_8[157]},
      {stage2_8[111]}
   );
   gpc1_1 gpc6113 (
      {stage1_8[158]},
      {stage2_8[112]}
   );
   gpc1_1 gpc6114 (
      {stage1_8[159]},
      {stage2_8[113]}
   );
   gpc1_1 gpc6115 (
      {stage1_8[160]},
      {stage2_8[114]}
   );
   gpc1_1 gpc6116 (
      {stage1_8[161]},
      {stage2_8[115]}
   );
   gpc1_1 gpc6117 (
      {stage1_8[162]},
      {stage2_8[116]}
   );
   gpc1_1 gpc6118 (
      {stage1_8[163]},
      {stage2_8[117]}
   );
   gpc1_1 gpc6119 (
      {stage1_8[164]},
      {stage2_8[118]}
   );
   gpc1_1 gpc6120 (
      {stage1_8[165]},
      {stage2_8[119]}
   );
   gpc1_1 gpc6121 (
      {stage1_8[166]},
      {stage2_8[120]}
   );
   gpc1_1 gpc6122 (
      {stage1_8[167]},
      {stage2_8[121]}
   );
   gpc1_1 gpc6123 (
      {stage1_8[168]},
      {stage2_8[122]}
   );
   gpc1_1 gpc6124 (
      {stage1_8[169]},
      {stage2_8[123]}
   );
   gpc1_1 gpc6125 (
      {stage1_8[170]},
      {stage2_8[124]}
   );
   gpc1_1 gpc6126 (
      {stage1_8[171]},
      {stage2_8[125]}
   );
   gpc1_1 gpc6127 (
      {stage1_8[172]},
      {stage2_8[126]}
   );
   gpc1_1 gpc6128 (
      {stage1_8[173]},
      {stage2_8[127]}
   );
   gpc1_1 gpc6129 (
      {stage1_8[174]},
      {stage2_8[128]}
   );
   gpc1_1 gpc6130 (
      {stage1_8[175]},
      {stage2_8[129]}
   );
   gpc1_1 gpc6131 (
      {stage1_8[176]},
      {stage2_8[130]}
   );
   gpc1_1 gpc6132 (
      {stage1_8[177]},
      {stage2_8[131]}
   );
   gpc1_1 gpc6133 (
      {stage1_8[178]},
      {stage2_8[132]}
   );
   gpc1_1 gpc6134 (
      {stage1_8[179]},
      {stage2_8[133]}
   );
   gpc1_1 gpc6135 (
      {stage1_8[180]},
      {stage2_8[134]}
   );
   gpc1_1 gpc6136 (
      {stage1_8[181]},
      {stage2_8[135]}
   );
   gpc1_1 gpc6137 (
      {stage1_8[182]},
      {stage2_8[136]}
   );
   gpc1_1 gpc6138 (
      {stage1_8[183]},
      {stage2_8[137]}
   );
   gpc1_1 gpc6139 (
      {stage1_8[184]},
      {stage2_8[138]}
   );
   gpc1_1 gpc6140 (
      {stage1_8[185]},
      {stage2_8[139]}
   );
   gpc1_1 gpc6141 (
      {stage1_8[186]},
      {stage2_8[140]}
   );
   gpc1_1 gpc6142 (
      {stage1_8[187]},
      {stage2_8[141]}
   );
   gpc1_1 gpc6143 (
      {stage1_8[188]},
      {stage2_8[142]}
   );
   gpc1_1 gpc6144 (
      {stage1_8[189]},
      {stage2_8[143]}
   );
   gpc1_1 gpc6145 (
      {stage1_8[190]},
      {stage2_8[144]}
   );
   gpc1_1 gpc6146 (
      {stage1_8[191]},
      {stage2_8[145]}
   );
   gpc1_1 gpc6147 (
      {stage1_8[192]},
      {stage2_8[146]}
   );
   gpc1_1 gpc6148 (
      {stage1_8[193]},
      {stage2_8[147]}
   );
   gpc1_1 gpc6149 (
      {stage1_8[194]},
      {stage2_8[148]}
   );
   gpc1_1 gpc6150 (
      {stage1_8[195]},
      {stage2_8[149]}
   );
   gpc1_1 gpc6151 (
      {stage1_8[196]},
      {stage2_8[150]}
   );
   gpc1_1 gpc6152 (
      {stage1_8[197]},
      {stage2_8[151]}
   );
   gpc1_1 gpc6153 (
      {stage1_8[198]},
      {stage2_8[152]}
   );
   gpc1_1 gpc6154 (
      {stage1_8[199]},
      {stage2_8[153]}
   );
   gpc1_1 gpc6155 (
      {stage1_8[200]},
      {stage2_8[154]}
   );
   gpc1_1 gpc6156 (
      {stage1_8[201]},
      {stage2_8[155]}
   );
   gpc1_1 gpc6157 (
      {stage1_8[202]},
      {stage2_8[156]}
   );
   gpc1_1 gpc6158 (
      {stage1_8[203]},
      {stage2_8[157]}
   );
   gpc1_1 gpc6159 (
      {stage1_8[204]},
      {stage2_8[158]}
   );
   gpc1_1 gpc6160 (
      {stage1_8[205]},
      {stage2_8[159]}
   );
   gpc1_1 gpc6161 (
      {stage1_9[132]},
      {stage2_9[61]}
   );
   gpc1_1 gpc6162 (
      {stage1_9[133]},
      {stage2_9[62]}
   );
   gpc1_1 gpc6163 (
      {stage1_9[134]},
      {stage2_9[63]}
   );
   gpc1_1 gpc6164 (
      {stage1_9[135]},
      {stage2_9[64]}
   );
   gpc1_1 gpc6165 (
      {stage1_9[136]},
      {stage2_9[65]}
   );
   gpc1_1 gpc6166 (
      {stage1_9[137]},
      {stage2_9[66]}
   );
   gpc1_1 gpc6167 (
      {stage1_9[138]},
      {stage2_9[67]}
   );
   gpc1_1 gpc6168 (
      {stage1_9[139]},
      {stage2_9[68]}
   );
   gpc1_1 gpc6169 (
      {stage1_9[140]},
      {stage2_9[69]}
   );
   gpc1_1 gpc6170 (
      {stage1_9[141]},
      {stage2_9[70]}
   );
   gpc1_1 gpc6171 (
      {stage1_9[142]},
      {stage2_9[71]}
   );
   gpc1_1 gpc6172 (
      {stage1_9[143]},
      {stage2_9[72]}
   );
   gpc1_1 gpc6173 (
      {stage1_9[144]},
      {stage2_9[73]}
   );
   gpc1_1 gpc6174 (
      {stage1_9[145]},
      {stage2_9[74]}
   );
   gpc1_1 gpc6175 (
      {stage1_9[146]},
      {stage2_9[75]}
   );
   gpc1_1 gpc6176 (
      {stage1_9[147]},
      {stage2_9[76]}
   );
   gpc1_1 gpc6177 (
      {stage1_9[148]},
      {stage2_9[77]}
   );
   gpc1_1 gpc6178 (
      {stage1_9[149]},
      {stage2_9[78]}
   );
   gpc1_1 gpc6179 (
      {stage1_9[150]},
      {stage2_9[79]}
   );
   gpc1_1 gpc6180 (
      {stage1_9[151]},
      {stage2_9[80]}
   );
   gpc1_1 gpc6181 (
      {stage1_9[152]},
      {stage2_9[81]}
   );
   gpc1_1 gpc6182 (
      {stage1_9[153]},
      {stage2_9[82]}
   );
   gpc1_1 gpc6183 (
      {stage1_9[154]},
      {stage2_9[83]}
   );
   gpc1_1 gpc6184 (
      {stage1_9[155]},
      {stage2_9[84]}
   );
   gpc1_1 gpc6185 (
      {stage1_9[156]},
      {stage2_9[85]}
   );
   gpc1_1 gpc6186 (
      {stage1_9[157]},
      {stage2_9[86]}
   );
   gpc1_1 gpc6187 (
      {stage1_9[158]},
      {stage2_9[87]}
   );
   gpc1_1 gpc6188 (
      {stage1_9[159]},
      {stage2_9[88]}
   );
   gpc1_1 gpc6189 (
      {stage1_9[160]},
      {stage2_9[89]}
   );
   gpc1_1 gpc6190 (
      {stage1_9[161]},
      {stage2_9[90]}
   );
   gpc1_1 gpc6191 (
      {stage1_9[162]},
      {stage2_9[91]}
   );
   gpc1_1 gpc6192 (
      {stage1_9[163]},
      {stage2_9[92]}
   );
   gpc1_1 gpc6193 (
      {stage1_9[164]},
      {stage2_9[93]}
   );
   gpc1_1 gpc6194 (
      {stage1_9[165]},
      {stage2_9[94]}
   );
   gpc1_1 gpc6195 (
      {stage1_9[166]},
      {stage2_9[95]}
   );
   gpc1_1 gpc6196 (
      {stage1_9[167]},
      {stage2_9[96]}
   );
   gpc1_1 gpc6197 (
      {stage1_9[168]},
      {stage2_9[97]}
   );
   gpc1_1 gpc6198 (
      {stage1_9[169]},
      {stage2_9[98]}
   );
   gpc1_1 gpc6199 (
      {stage1_9[170]},
      {stage2_9[99]}
   );
   gpc1_1 gpc6200 (
      {stage1_9[171]},
      {stage2_9[100]}
   );
   gpc1_1 gpc6201 (
      {stage1_9[172]},
      {stage2_9[101]}
   );
   gpc1_1 gpc6202 (
      {stage1_9[173]},
      {stage2_9[102]}
   );
   gpc1_1 gpc6203 (
      {stage1_9[174]},
      {stage2_9[103]}
   );
   gpc1_1 gpc6204 (
      {stage1_9[175]},
      {stage2_9[104]}
   );
   gpc1_1 gpc6205 (
      {stage1_9[176]},
      {stage2_9[105]}
   );
   gpc1_1 gpc6206 (
      {stage1_9[177]},
      {stage2_9[106]}
   );
   gpc1_1 gpc6207 (
      {stage1_9[178]},
      {stage2_9[107]}
   );
   gpc1_1 gpc6208 (
      {stage1_9[179]},
      {stage2_9[108]}
   );
   gpc1_1 gpc6209 (
      {stage1_9[180]},
      {stage2_9[109]}
   );
   gpc1_1 gpc6210 (
      {stage1_9[181]},
      {stage2_9[110]}
   );
   gpc1_1 gpc6211 (
      {stage1_9[182]},
      {stage2_9[111]}
   );
   gpc1_1 gpc6212 (
      {stage1_9[183]},
      {stage2_9[112]}
   );
   gpc1_1 gpc6213 (
      {stage1_9[184]},
      {stage2_9[113]}
   );
   gpc1_1 gpc6214 (
      {stage1_9[185]},
      {stage2_9[114]}
   );
   gpc1_1 gpc6215 (
      {stage1_9[186]},
      {stage2_9[115]}
   );
   gpc1_1 gpc6216 (
      {stage1_9[187]},
      {stage2_9[116]}
   );
   gpc1_1 gpc6217 (
      {stage1_9[188]},
      {stage2_9[117]}
   );
   gpc1_1 gpc6218 (
      {stage1_9[189]},
      {stage2_9[118]}
   );
   gpc1_1 gpc6219 (
      {stage1_9[190]},
      {stage2_9[119]}
   );
   gpc1_1 gpc6220 (
      {stage1_9[191]},
      {stage2_9[120]}
   );
   gpc1_1 gpc6221 (
      {stage1_9[192]},
      {stage2_9[121]}
   );
   gpc1_1 gpc6222 (
      {stage1_9[193]},
      {stage2_9[122]}
   );
   gpc1_1 gpc6223 (
      {stage1_9[194]},
      {stage2_9[123]}
   );
   gpc1_1 gpc6224 (
      {stage1_9[195]},
      {stage2_9[124]}
   );
   gpc1_1 gpc6225 (
      {stage1_9[196]},
      {stage2_9[125]}
   );
   gpc1_1 gpc6226 (
      {stage1_9[197]},
      {stage2_9[126]}
   );
   gpc1_1 gpc6227 (
      {stage1_9[198]},
      {stage2_9[127]}
   );
   gpc1_1 gpc6228 (
      {stage1_9[199]},
      {stage2_9[128]}
   );
   gpc1_1 gpc6229 (
      {stage1_9[200]},
      {stage2_9[129]}
   );
   gpc1_1 gpc6230 (
      {stage1_9[201]},
      {stage2_9[130]}
   );
   gpc1_1 gpc6231 (
      {stage1_9[202]},
      {stage2_9[131]}
   );
   gpc1_1 gpc6232 (
      {stage1_9[203]},
      {stage2_9[132]}
   );
   gpc1_1 gpc6233 (
      {stage1_9[204]},
      {stage2_9[133]}
   );
   gpc1_1 gpc6234 (
      {stage1_9[205]},
      {stage2_9[134]}
   );
   gpc1_1 gpc6235 (
      {stage1_9[206]},
      {stage2_9[135]}
   );
   gpc1_1 gpc6236 (
      {stage1_9[207]},
      {stage2_9[136]}
   );
   gpc1_1 gpc6237 (
      {stage1_9[208]},
      {stage2_9[137]}
   );
   gpc1_1 gpc6238 (
      {stage1_9[209]},
      {stage2_9[138]}
   );
   gpc1_1 gpc6239 (
      {stage1_9[210]},
      {stage2_9[139]}
   );
   gpc1_1 gpc6240 (
      {stage1_9[211]},
      {stage2_9[140]}
   );
   gpc1_1 gpc6241 (
      {stage1_9[212]},
      {stage2_9[141]}
   );
   gpc1_1 gpc6242 (
      {stage1_9[213]},
      {stage2_9[142]}
   );
   gpc1_1 gpc6243 (
      {stage1_10[175]},
      {stage2_10[54]}
   );
   gpc1_1 gpc6244 (
      {stage1_10[176]},
      {stage2_10[55]}
   );
   gpc1_1 gpc6245 (
      {stage1_10[177]},
      {stage2_10[56]}
   );
   gpc1_1 gpc6246 (
      {stage1_10[178]},
      {stage2_10[57]}
   );
   gpc1_1 gpc6247 (
      {stage1_10[179]},
      {stage2_10[58]}
   );
   gpc1_1 gpc6248 (
      {stage1_10[180]},
      {stage2_10[59]}
   );
   gpc1_1 gpc6249 (
      {stage1_10[181]},
      {stage2_10[60]}
   );
   gpc1_1 gpc6250 (
      {stage1_10[182]},
      {stage2_10[61]}
   );
   gpc1_1 gpc6251 (
      {stage1_10[183]},
      {stage2_10[62]}
   );
   gpc1_1 gpc6252 (
      {stage1_10[184]},
      {stage2_10[63]}
   );
   gpc1_1 gpc6253 (
      {stage1_10[185]},
      {stage2_10[64]}
   );
   gpc1_1 gpc6254 (
      {stage1_10[186]},
      {stage2_10[65]}
   );
   gpc1_1 gpc6255 (
      {stage1_10[187]},
      {stage2_10[66]}
   );
   gpc1_1 gpc6256 (
      {stage1_10[188]},
      {stage2_10[67]}
   );
   gpc1_1 gpc6257 (
      {stage1_10[189]},
      {stage2_10[68]}
   );
   gpc1_1 gpc6258 (
      {stage1_10[190]},
      {stage2_10[69]}
   );
   gpc1_1 gpc6259 (
      {stage1_10[191]},
      {stage2_10[70]}
   );
   gpc1_1 gpc6260 (
      {stage1_10[192]},
      {stage2_10[71]}
   );
   gpc1_1 gpc6261 (
      {stage1_10[193]},
      {stage2_10[72]}
   );
   gpc1_1 gpc6262 (
      {stage1_10[194]},
      {stage2_10[73]}
   );
   gpc1_1 gpc6263 (
      {stage1_10[195]},
      {stage2_10[74]}
   );
   gpc1_1 gpc6264 (
      {stage1_10[196]},
      {stage2_10[75]}
   );
   gpc1_1 gpc6265 (
      {stage1_10[197]},
      {stage2_10[76]}
   );
   gpc1_1 gpc6266 (
      {stage1_10[198]},
      {stage2_10[77]}
   );
   gpc1_1 gpc6267 (
      {stage1_10[199]},
      {stage2_10[78]}
   );
   gpc1_1 gpc6268 (
      {stage1_10[200]},
      {stage2_10[79]}
   );
   gpc1_1 gpc6269 (
      {stage1_10[201]},
      {stage2_10[80]}
   );
   gpc1_1 gpc6270 (
      {stage1_10[202]},
      {stage2_10[81]}
   );
   gpc1_1 gpc6271 (
      {stage1_10[203]},
      {stage2_10[82]}
   );
   gpc1_1 gpc6272 (
      {stage1_10[204]},
      {stage2_10[83]}
   );
   gpc1_1 gpc6273 (
      {stage1_10[205]},
      {stage2_10[84]}
   );
   gpc1_1 gpc6274 (
      {stage1_10[206]},
      {stage2_10[85]}
   );
   gpc1_1 gpc6275 (
      {stage1_10[207]},
      {stage2_10[86]}
   );
   gpc1_1 gpc6276 (
      {stage1_10[208]},
      {stage2_10[87]}
   );
   gpc1_1 gpc6277 (
      {stage1_10[209]},
      {stage2_10[88]}
   );
   gpc1_1 gpc6278 (
      {stage1_10[210]},
      {stage2_10[89]}
   );
   gpc1_1 gpc6279 (
      {stage1_10[211]},
      {stage2_10[90]}
   );
   gpc1_1 gpc6280 (
      {stage1_10[212]},
      {stage2_10[91]}
   );
   gpc1_1 gpc6281 (
      {stage1_10[213]},
      {stage2_10[92]}
   );
   gpc1_1 gpc6282 (
      {stage1_10[214]},
      {stage2_10[93]}
   );
   gpc1_1 gpc6283 (
      {stage1_10[215]},
      {stage2_10[94]}
   );
   gpc1_1 gpc6284 (
      {stage1_10[216]},
      {stage2_10[95]}
   );
   gpc1_1 gpc6285 (
      {stage1_10[217]},
      {stage2_10[96]}
   );
   gpc1_1 gpc6286 (
      {stage1_10[218]},
      {stage2_10[97]}
   );
   gpc1_1 gpc6287 (
      {stage1_10[219]},
      {stage2_10[98]}
   );
   gpc1_1 gpc6288 (
      {stage1_10[220]},
      {stage2_10[99]}
   );
   gpc1_1 gpc6289 (
      {stage1_10[221]},
      {stage2_10[100]}
   );
   gpc1_1 gpc6290 (
      {stage1_10[222]},
      {stage2_10[101]}
   );
   gpc1_1 gpc6291 (
      {stage1_10[223]},
      {stage2_10[102]}
   );
   gpc1_1 gpc6292 (
      {stage1_10[224]},
      {stage2_10[103]}
   );
   gpc1_1 gpc6293 (
      {stage1_10[225]},
      {stage2_10[104]}
   );
   gpc1_1 gpc6294 (
      {stage1_10[226]},
      {stage2_10[105]}
   );
   gpc1_1 gpc6295 (
      {stage1_10[227]},
      {stage2_10[106]}
   );
   gpc1_1 gpc6296 (
      {stage1_10[228]},
      {stage2_10[107]}
   );
   gpc1_1 gpc6297 (
      {stage1_10[229]},
      {stage2_10[108]}
   );
   gpc1_1 gpc6298 (
      {stage1_10[230]},
      {stage2_10[109]}
   );
   gpc1_1 gpc6299 (
      {stage1_10[231]},
      {stage2_10[110]}
   );
   gpc1_1 gpc6300 (
      {stage1_10[232]},
      {stage2_10[111]}
   );
   gpc1_1 gpc6301 (
      {stage1_10[233]},
      {stage2_10[112]}
   );
   gpc1_1 gpc6302 (
      {stage1_10[234]},
      {stage2_10[113]}
   );
   gpc1_1 gpc6303 (
      {stage1_10[235]},
      {stage2_10[114]}
   );
   gpc1_1 gpc6304 (
      {stage1_10[236]},
      {stage2_10[115]}
   );
   gpc1_1 gpc6305 (
      {stage1_10[237]},
      {stage2_10[116]}
   );
   gpc1_1 gpc6306 (
      {stage1_10[238]},
      {stage2_10[117]}
   );
   gpc1_1 gpc6307 (
      {stage1_10[239]},
      {stage2_10[118]}
   );
   gpc1_1 gpc6308 (
      {stage1_10[240]},
      {stage2_10[119]}
   );
   gpc1_1 gpc6309 (
      {stage1_10[241]},
      {stage2_10[120]}
   );
   gpc1_1 gpc6310 (
      {stage1_10[242]},
      {stage2_10[121]}
   );
   gpc1_1 gpc6311 (
      {stage1_10[243]},
      {stage2_10[122]}
   );
   gpc1_1 gpc6312 (
      {stage1_10[244]},
      {stage2_10[123]}
   );
   gpc1_1 gpc6313 (
      {stage1_10[245]},
      {stage2_10[124]}
   );
   gpc1_1 gpc6314 (
      {stage1_10[246]},
      {stage2_10[125]}
   );
   gpc1_1 gpc6315 (
      {stage1_10[247]},
      {stage2_10[126]}
   );
   gpc1_1 gpc6316 (
      {stage1_10[248]},
      {stage2_10[127]}
   );
   gpc1_1 gpc6317 (
      {stage1_10[249]},
      {stage2_10[128]}
   );
   gpc1_1 gpc6318 (
      {stage1_10[250]},
      {stage2_10[129]}
   );
   gpc1_1 gpc6319 (
      {stage1_10[251]},
      {stage2_10[130]}
   );
   gpc1_1 gpc6320 (
      {stage1_10[252]},
      {stage2_10[131]}
   );
   gpc1_1 gpc6321 (
      {stage1_10[253]},
      {stage2_10[132]}
   );
   gpc1_1 gpc6322 (
      {stage1_10[254]},
      {stage2_10[133]}
   );
   gpc1_1 gpc6323 (
      {stage1_10[255]},
      {stage2_10[134]}
   );
   gpc1_1 gpc6324 (
      {stage1_10[256]},
      {stage2_10[135]}
   );
   gpc1_1 gpc6325 (
      {stage1_10[257]},
      {stage2_10[136]}
   );
   gpc1_1 gpc6326 (
      {stage1_10[258]},
      {stage2_10[137]}
   );
   gpc1_1 gpc6327 (
      {stage1_10[259]},
      {stage2_10[138]}
   );
   gpc1_1 gpc6328 (
      {stage1_10[260]},
      {stage2_10[139]}
   );
   gpc1_1 gpc6329 (
      {stage1_10[261]},
      {stage2_10[140]}
   );
   gpc1_1 gpc6330 (
      {stage1_10[262]},
      {stage2_10[141]}
   );
   gpc1_1 gpc6331 (
      {stage1_10[263]},
      {stage2_10[142]}
   );
   gpc1_1 gpc6332 (
      {stage1_10[264]},
      {stage2_10[143]}
   );
   gpc1_1 gpc6333 (
      {stage1_10[265]},
      {stage2_10[144]}
   );
   gpc1_1 gpc6334 (
      {stage1_10[266]},
      {stage2_10[145]}
   );
   gpc1_1 gpc6335 (
      {stage1_10[267]},
      {stage2_10[146]}
   );
   gpc1_1 gpc6336 (
      {stage1_10[268]},
      {stage2_10[147]}
   );
   gpc1_1 gpc6337 (
      {stage1_10[269]},
      {stage2_10[148]}
   );
   gpc1_1 gpc6338 (
      {stage1_10[270]},
      {stage2_10[149]}
   );
   gpc1_1 gpc6339 (
      {stage1_10[271]},
      {stage2_10[150]}
   );
   gpc1_1 gpc6340 (
      {stage1_10[272]},
      {stage2_10[151]}
   );
   gpc1_1 gpc6341 (
      {stage1_10[273]},
      {stage2_10[152]}
   );
   gpc1_1 gpc6342 (
      {stage1_10[274]},
      {stage2_10[153]}
   );
   gpc1_1 gpc6343 (
      {stage1_10[275]},
      {stage2_10[154]}
   );
   gpc1_1 gpc6344 (
      {stage1_10[276]},
      {stage2_10[155]}
   );
   gpc1_1 gpc6345 (
      {stage1_10[277]},
      {stage2_10[156]}
   );
   gpc1_1 gpc6346 (
      {stage1_10[278]},
      {stage2_10[157]}
   );
   gpc1_1 gpc6347 (
      {stage1_10[279]},
      {stage2_10[158]}
   );
   gpc1_1 gpc6348 (
      {stage1_10[280]},
      {stage2_10[159]}
   );
   gpc1_1 gpc6349 (
      {stage1_10[281]},
      {stage2_10[160]}
   );
   gpc1_1 gpc6350 (
      {stage1_10[282]},
      {stage2_10[161]}
   );
   gpc1_1 gpc6351 (
      {stage1_10[283]},
      {stage2_10[162]}
   );
   gpc1_1 gpc6352 (
      {stage1_10[284]},
      {stage2_10[163]}
   );
   gpc1_1 gpc6353 (
      {stage1_11[228]},
      {stage2_11[90]}
   );
   gpc1_1 gpc6354 (
      {stage1_11[229]},
      {stage2_11[91]}
   );
   gpc1_1 gpc6355 (
      {stage1_11[230]},
      {stage2_11[92]}
   );
   gpc1_1 gpc6356 (
      {stage1_11[231]},
      {stage2_11[93]}
   );
   gpc1_1 gpc6357 (
      {stage1_11[232]},
      {stage2_11[94]}
   );
   gpc1_1 gpc6358 (
      {stage1_11[233]},
      {stage2_11[95]}
   );
   gpc1_1 gpc6359 (
      {stage1_11[234]},
      {stage2_11[96]}
   );
   gpc1_1 gpc6360 (
      {stage1_11[235]},
      {stage2_11[97]}
   );
   gpc1_1 gpc6361 (
      {stage1_11[236]},
      {stage2_11[98]}
   );
   gpc1_1 gpc6362 (
      {stage1_11[237]},
      {stage2_11[99]}
   );
   gpc1_1 gpc6363 (
      {stage1_11[238]},
      {stage2_11[100]}
   );
   gpc1_1 gpc6364 (
      {stage1_11[239]},
      {stage2_11[101]}
   );
   gpc1_1 gpc6365 (
      {stage1_11[240]},
      {stage2_11[102]}
   );
   gpc1_1 gpc6366 (
      {stage1_11[241]},
      {stage2_11[103]}
   );
   gpc1_1 gpc6367 (
      {stage1_11[242]},
      {stage2_11[104]}
   );
   gpc1_1 gpc6368 (
      {stage1_11[243]},
      {stage2_11[105]}
   );
   gpc1_1 gpc6369 (
      {stage1_11[244]},
      {stage2_11[106]}
   );
   gpc1_1 gpc6370 (
      {stage1_11[245]},
      {stage2_11[107]}
   );
   gpc1_1 gpc6371 (
      {stage1_11[246]},
      {stage2_11[108]}
   );
   gpc1_1 gpc6372 (
      {stage1_11[247]},
      {stage2_11[109]}
   );
   gpc1_1 gpc6373 (
      {stage1_11[248]},
      {stage2_11[110]}
   );
   gpc1_1 gpc6374 (
      {stage1_11[249]},
      {stage2_11[111]}
   );
   gpc1_1 gpc6375 (
      {stage1_11[250]},
      {stage2_11[112]}
   );
   gpc1_1 gpc6376 (
      {stage1_11[251]},
      {stage2_11[113]}
   );
   gpc1_1 gpc6377 (
      {stage1_11[252]},
      {stage2_11[114]}
   );
   gpc1_1 gpc6378 (
      {stage1_11[253]},
      {stage2_11[115]}
   );
   gpc1_1 gpc6379 (
      {stage1_11[254]},
      {stage2_11[116]}
   );
   gpc1_1 gpc6380 (
      {stage1_11[255]},
      {stage2_11[117]}
   );
   gpc1_1 gpc6381 (
      {stage1_11[256]},
      {stage2_11[118]}
   );
   gpc1_1 gpc6382 (
      {stage1_11[257]},
      {stage2_11[119]}
   );
   gpc1_1 gpc6383 (
      {stage1_11[258]},
      {stage2_11[120]}
   );
   gpc1_1 gpc6384 (
      {stage1_11[259]},
      {stage2_11[121]}
   );
   gpc1_1 gpc6385 (
      {stage1_11[260]},
      {stage2_11[122]}
   );
   gpc1_1 gpc6386 (
      {stage1_11[261]},
      {stage2_11[123]}
   );
   gpc1_1 gpc6387 (
      {stage1_11[262]},
      {stage2_11[124]}
   );
   gpc1_1 gpc6388 (
      {stage1_11[263]},
      {stage2_11[125]}
   );
   gpc1_1 gpc6389 (
      {stage1_11[264]},
      {stage2_11[126]}
   );
   gpc1_1 gpc6390 (
      {stage1_11[265]},
      {stage2_11[127]}
   );
   gpc1_1 gpc6391 (
      {stage1_11[266]},
      {stage2_11[128]}
   );
   gpc1_1 gpc6392 (
      {stage1_11[267]},
      {stage2_11[129]}
   );
   gpc1_1 gpc6393 (
      {stage1_11[268]},
      {stage2_11[130]}
   );
   gpc1_1 gpc6394 (
      {stage1_11[269]},
      {stage2_11[131]}
   );
   gpc1_1 gpc6395 (
      {stage1_11[270]},
      {stage2_11[132]}
   );
   gpc1_1 gpc6396 (
      {stage1_11[271]},
      {stage2_11[133]}
   );
   gpc1_1 gpc6397 (
      {stage1_11[272]},
      {stage2_11[134]}
   );
   gpc1_1 gpc6398 (
      {stage1_11[273]},
      {stage2_11[135]}
   );
   gpc1_1 gpc6399 (
      {stage1_11[274]},
      {stage2_11[136]}
   );
   gpc1_1 gpc6400 (
      {stage1_11[275]},
      {stage2_11[137]}
   );
   gpc1_1 gpc6401 (
      {stage1_11[276]},
      {stage2_11[138]}
   );
   gpc1_1 gpc6402 (
      {stage1_12[163]},
      {stage2_12[81]}
   );
   gpc1_1 gpc6403 (
      {stage1_12[164]},
      {stage2_12[82]}
   );
   gpc1_1 gpc6404 (
      {stage1_12[165]},
      {stage2_12[83]}
   );
   gpc1_1 gpc6405 (
      {stage1_12[166]},
      {stage2_12[84]}
   );
   gpc1_1 gpc6406 (
      {stage1_12[167]},
      {stage2_12[85]}
   );
   gpc1_1 gpc6407 (
      {stage1_12[168]},
      {stage2_12[86]}
   );
   gpc1_1 gpc6408 (
      {stage1_12[169]},
      {stage2_12[87]}
   );
   gpc1_1 gpc6409 (
      {stage1_12[170]},
      {stage2_12[88]}
   );
   gpc1_1 gpc6410 (
      {stage1_12[171]},
      {stage2_12[89]}
   );
   gpc1_1 gpc6411 (
      {stage1_12[172]},
      {stage2_12[90]}
   );
   gpc1_1 gpc6412 (
      {stage1_12[173]},
      {stage2_12[91]}
   );
   gpc1_1 gpc6413 (
      {stage1_12[174]},
      {stage2_12[92]}
   );
   gpc1_1 gpc6414 (
      {stage1_12[175]},
      {stage2_12[93]}
   );
   gpc1_1 gpc6415 (
      {stage1_12[176]},
      {stage2_12[94]}
   );
   gpc1_1 gpc6416 (
      {stage1_12[177]},
      {stage2_12[95]}
   );
   gpc1_1 gpc6417 (
      {stage1_12[178]},
      {stage2_12[96]}
   );
   gpc1_1 gpc6418 (
      {stage1_12[179]},
      {stage2_12[97]}
   );
   gpc1_1 gpc6419 (
      {stage1_12[180]},
      {stage2_12[98]}
   );
   gpc1_1 gpc6420 (
      {stage1_12[181]},
      {stage2_12[99]}
   );
   gpc1_1 gpc6421 (
      {stage1_12[182]},
      {stage2_12[100]}
   );
   gpc1_1 gpc6422 (
      {stage1_12[183]},
      {stage2_12[101]}
   );
   gpc1_1 gpc6423 (
      {stage1_12[184]},
      {stage2_12[102]}
   );
   gpc1_1 gpc6424 (
      {stage1_12[185]},
      {stage2_12[103]}
   );
   gpc1_1 gpc6425 (
      {stage1_12[186]},
      {stage2_12[104]}
   );
   gpc1_1 gpc6426 (
      {stage1_12[187]},
      {stage2_12[105]}
   );
   gpc1_1 gpc6427 (
      {stage1_12[188]},
      {stage2_12[106]}
   );
   gpc1_1 gpc6428 (
      {stage1_14[217]},
      {stage2_14[106]}
   );
   gpc1_1 gpc6429 (
      {stage1_14[218]},
      {stage2_14[107]}
   );
   gpc1_1 gpc6430 (
      {stage1_15[123]},
      {stage2_15[93]}
   );
   gpc1_1 gpc6431 (
      {stage1_15[124]},
      {stage2_15[94]}
   );
   gpc1_1 gpc6432 (
      {stage1_15[125]},
      {stage2_15[95]}
   );
   gpc1_1 gpc6433 (
      {stage1_15[126]},
      {stage2_15[96]}
   );
   gpc1_1 gpc6434 (
      {stage1_15[127]},
      {stage2_15[97]}
   );
   gpc1_1 gpc6435 (
      {stage1_15[128]},
      {stage2_15[98]}
   );
   gpc1_1 gpc6436 (
      {stage1_15[129]},
      {stage2_15[99]}
   );
   gpc1_1 gpc6437 (
      {stage1_15[130]},
      {stage2_15[100]}
   );
   gpc1_1 gpc6438 (
      {stage1_15[131]},
      {stage2_15[101]}
   );
   gpc1_1 gpc6439 (
      {stage1_15[132]},
      {stage2_15[102]}
   );
   gpc1_1 gpc6440 (
      {stage1_15[133]},
      {stage2_15[103]}
   );
   gpc1_1 gpc6441 (
      {stage1_15[134]},
      {stage2_15[104]}
   );
   gpc1_1 gpc6442 (
      {stage1_15[135]},
      {stage2_15[105]}
   );
   gpc1_1 gpc6443 (
      {stage1_15[136]},
      {stage2_15[106]}
   );
   gpc1_1 gpc6444 (
      {stage1_15[137]},
      {stage2_15[107]}
   );
   gpc1_1 gpc6445 (
      {stage1_15[138]},
      {stage2_15[108]}
   );
   gpc1_1 gpc6446 (
      {stage1_15[139]},
      {stage2_15[109]}
   );
   gpc1_1 gpc6447 (
      {stage1_15[140]},
      {stage2_15[110]}
   );
   gpc1_1 gpc6448 (
      {stage1_15[141]},
      {stage2_15[111]}
   );
   gpc1_1 gpc6449 (
      {stage1_15[142]},
      {stage2_15[112]}
   );
   gpc1_1 gpc6450 (
      {stage1_15[143]},
      {stage2_15[113]}
   );
   gpc1_1 gpc6451 (
      {stage1_15[144]},
      {stage2_15[114]}
   );
   gpc1_1 gpc6452 (
      {stage1_15[145]},
      {stage2_15[115]}
   );
   gpc1_1 gpc6453 (
      {stage1_15[146]},
      {stage2_15[116]}
   );
   gpc1_1 gpc6454 (
      {stage1_15[147]},
      {stage2_15[117]}
   );
   gpc1_1 gpc6455 (
      {stage1_15[148]},
      {stage2_15[118]}
   );
   gpc1_1 gpc6456 (
      {stage1_15[149]},
      {stage2_15[119]}
   );
   gpc1_1 gpc6457 (
      {stage1_15[150]},
      {stage2_15[120]}
   );
   gpc1_1 gpc6458 (
      {stage1_15[151]},
      {stage2_15[121]}
   );
   gpc1_1 gpc6459 (
      {stage1_15[152]},
      {stage2_15[122]}
   );
   gpc1_1 gpc6460 (
      {stage1_15[153]},
      {stage2_15[123]}
   );
   gpc1_1 gpc6461 (
      {stage1_15[154]},
      {stage2_15[124]}
   );
   gpc1_1 gpc6462 (
      {stage1_15[155]},
      {stage2_15[125]}
   );
   gpc1_1 gpc6463 (
      {stage1_15[156]},
      {stage2_15[126]}
   );
   gpc1_1 gpc6464 (
      {stage1_15[157]},
      {stage2_15[127]}
   );
   gpc1_1 gpc6465 (
      {stage1_15[158]},
      {stage2_15[128]}
   );
   gpc1_1 gpc6466 (
      {stage1_15[159]},
      {stage2_15[129]}
   );
   gpc1_1 gpc6467 (
      {stage1_15[160]},
      {stage2_15[130]}
   );
   gpc1_1 gpc6468 (
      {stage1_15[161]},
      {stage2_15[131]}
   );
   gpc1_1 gpc6469 (
      {stage1_15[162]},
      {stage2_15[132]}
   );
   gpc1_1 gpc6470 (
      {stage1_15[163]},
      {stage2_15[133]}
   );
   gpc1_1 gpc6471 (
      {stage1_15[164]},
      {stage2_15[134]}
   );
   gpc1_1 gpc6472 (
      {stage1_15[165]},
      {stage2_15[135]}
   );
   gpc1_1 gpc6473 (
      {stage1_15[166]},
      {stage2_15[136]}
   );
   gpc1_1 gpc6474 (
      {stage1_15[167]},
      {stage2_15[137]}
   );
   gpc1_1 gpc6475 (
      {stage1_15[168]},
      {stage2_15[138]}
   );
   gpc1_1 gpc6476 (
      {stage1_15[169]},
      {stage2_15[139]}
   );
   gpc1_1 gpc6477 (
      {stage1_15[170]},
      {stage2_15[140]}
   );
   gpc1_1 gpc6478 (
      {stage1_16[198]},
      {stage2_16[59]}
   );
   gpc1_1 gpc6479 (
      {stage1_16[199]},
      {stage2_16[60]}
   );
   gpc1_1 gpc6480 (
      {stage1_16[200]},
      {stage2_16[61]}
   );
   gpc1_1 gpc6481 (
      {stage1_16[201]},
      {stage2_16[62]}
   );
   gpc1_1 gpc6482 (
      {stage1_16[202]},
      {stage2_16[63]}
   );
   gpc1_1 gpc6483 (
      {stage1_16[203]},
      {stage2_16[64]}
   );
   gpc1_1 gpc6484 (
      {stage1_16[204]},
      {stage2_16[65]}
   );
   gpc1_1 gpc6485 (
      {stage1_16[205]},
      {stage2_16[66]}
   );
   gpc1_1 gpc6486 (
      {stage1_16[206]},
      {stage2_16[67]}
   );
   gpc1_1 gpc6487 (
      {stage1_16[207]},
      {stage2_16[68]}
   );
   gpc1_1 gpc6488 (
      {stage1_16[208]},
      {stage2_16[69]}
   );
   gpc1_1 gpc6489 (
      {stage1_16[209]},
      {stage2_16[70]}
   );
   gpc1_1 gpc6490 (
      {stage1_16[210]},
      {stage2_16[71]}
   );
   gpc1_1 gpc6491 (
      {stage1_16[211]},
      {stage2_16[72]}
   );
   gpc1_1 gpc6492 (
      {stage1_16[212]},
      {stage2_16[73]}
   );
   gpc1_1 gpc6493 (
      {stage1_16[213]},
      {stage2_16[74]}
   );
   gpc1_1 gpc6494 (
      {stage1_16[214]},
      {stage2_16[75]}
   );
   gpc1_1 gpc6495 (
      {stage1_16[215]},
      {stage2_16[76]}
   );
   gpc1_1 gpc6496 (
      {stage1_16[216]},
      {stage2_16[77]}
   );
   gpc1_1 gpc6497 (
      {stage1_16[217]},
      {stage2_16[78]}
   );
   gpc1_1 gpc6498 (
      {stage1_16[218]},
      {stage2_16[79]}
   );
   gpc1_1 gpc6499 (
      {stage1_16[219]},
      {stage2_16[80]}
   );
   gpc1_1 gpc6500 (
      {stage1_16[220]},
      {stage2_16[81]}
   );
   gpc1_1 gpc6501 (
      {stage1_16[221]},
      {stage2_16[82]}
   );
   gpc1_1 gpc6502 (
      {stage1_17[228]},
      {stage2_17[86]}
   );
   gpc1_1 gpc6503 (
      {stage1_18[191]},
      {stage2_18[101]}
   );
   gpc1_1 gpc6504 (
      {stage1_18[192]},
      {stage2_18[102]}
   );
   gpc1_1 gpc6505 (
      {stage1_18[193]},
      {stage2_18[103]}
   );
   gpc1_1 gpc6506 (
      {stage1_18[194]},
      {stage2_18[104]}
   );
   gpc1_1 gpc6507 (
      {stage1_18[195]},
      {stage2_18[105]}
   );
   gpc1_1 gpc6508 (
      {stage1_18[196]},
      {stage2_18[106]}
   );
   gpc1_1 gpc6509 (
      {stage1_18[197]},
      {stage2_18[107]}
   );
   gpc1_1 gpc6510 (
      {stage1_18[198]},
      {stage2_18[108]}
   );
   gpc1_1 gpc6511 (
      {stage1_18[199]},
      {stage2_18[109]}
   );
   gpc1_1 gpc6512 (
      {stage1_18[200]},
      {stage2_18[110]}
   );
   gpc1_1 gpc6513 (
      {stage1_18[201]},
      {stage2_18[111]}
   );
   gpc1_1 gpc6514 (
      {stage1_18[202]},
      {stage2_18[112]}
   );
   gpc1_1 gpc6515 (
      {stage1_18[203]},
      {stage2_18[113]}
   );
   gpc1_1 gpc6516 (
      {stage1_18[204]},
      {stage2_18[114]}
   );
   gpc1_1 gpc6517 (
      {stage1_18[205]},
      {stage2_18[115]}
   );
   gpc1_1 gpc6518 (
      {stage1_18[206]},
      {stage2_18[116]}
   );
   gpc1_1 gpc6519 (
      {stage1_18[207]},
      {stage2_18[117]}
   );
   gpc1_1 gpc6520 (
      {stage1_18[208]},
      {stage2_18[118]}
   );
   gpc1_1 gpc6521 (
      {stage1_19[234]},
      {stage2_19[71]}
   );
   gpc1_1 gpc6522 (
      {stage1_19[235]},
      {stage2_19[72]}
   );
   gpc1_1 gpc6523 (
      {stage1_19[236]},
      {stage2_19[73]}
   );
   gpc1_1 gpc6524 (
      {stage1_19[237]},
      {stage2_19[74]}
   );
   gpc1_1 gpc6525 (
      {stage1_19[238]},
      {stage2_19[75]}
   );
   gpc1_1 gpc6526 (
      {stage1_19[239]},
      {stage2_19[76]}
   );
   gpc1_1 gpc6527 (
      {stage1_19[240]},
      {stage2_19[77]}
   );
   gpc1_1 gpc6528 (
      {stage1_19[241]},
      {stage2_19[78]}
   );
   gpc1_1 gpc6529 (
      {stage1_19[242]},
      {stage2_19[79]}
   );
   gpc1_1 gpc6530 (
      {stage1_19[243]},
      {stage2_19[80]}
   );
   gpc1_1 gpc6531 (
      {stage1_19[244]},
      {stage2_19[81]}
   );
   gpc1_1 gpc6532 (
      {stage1_19[245]},
      {stage2_19[82]}
   );
   gpc1_1 gpc6533 (
      {stage1_19[246]},
      {stage2_19[83]}
   );
   gpc1_1 gpc6534 (
      {stage1_19[247]},
      {stage2_19[84]}
   );
   gpc1_1 gpc6535 (
      {stage1_19[248]},
      {stage2_19[85]}
   );
   gpc1_1 gpc6536 (
      {stage1_19[249]},
      {stage2_19[86]}
   );
   gpc1_1 gpc6537 (
      {stage1_19[250]},
      {stage2_19[87]}
   );
   gpc1_1 gpc6538 (
      {stage1_19[251]},
      {stage2_19[88]}
   );
   gpc1_1 gpc6539 (
      {stage1_19[252]},
      {stage2_19[89]}
   );
   gpc1_1 gpc6540 (
      {stage1_19[253]},
      {stage2_19[90]}
   );
   gpc1_1 gpc6541 (
      {stage1_19[254]},
      {stage2_19[91]}
   );
   gpc1_1 gpc6542 (
      {stage1_19[255]},
      {stage2_19[92]}
   );
   gpc1_1 gpc6543 (
      {stage1_19[256]},
      {stage2_19[93]}
   );
   gpc1_1 gpc6544 (
      {stage1_19[257]},
      {stage2_19[94]}
   );
   gpc1_1 gpc6545 (
      {stage1_19[258]},
      {stage2_19[95]}
   );
   gpc1_1 gpc6546 (
      {stage1_19[259]},
      {stage2_19[96]}
   );
   gpc1_1 gpc6547 (
      {stage1_19[260]},
      {stage2_19[97]}
   );
   gpc1_1 gpc6548 (
      {stage1_19[261]},
      {stage2_19[98]}
   );
   gpc1_1 gpc6549 (
      {stage1_19[262]},
      {stage2_19[99]}
   );
   gpc1_1 gpc6550 (
      {stage1_19[263]},
      {stage2_19[100]}
   );
   gpc1_1 gpc6551 (
      {stage1_19[264]},
      {stage2_19[101]}
   );
   gpc1_1 gpc6552 (
      {stage1_19[265]},
      {stage2_19[102]}
   );
   gpc1_1 gpc6553 (
      {stage1_19[266]},
      {stage2_19[103]}
   );
   gpc1_1 gpc6554 (
      {stage1_19[267]},
      {stage2_19[104]}
   );
   gpc1_1 gpc6555 (
      {stage1_19[268]},
      {stage2_19[105]}
   );
   gpc1_1 gpc6556 (
      {stage1_19[269]},
      {stage2_19[106]}
   );
   gpc1_1 gpc6557 (
      {stage1_19[270]},
      {stage2_19[107]}
   );
   gpc1_1 gpc6558 (
      {stage1_19[271]},
      {stage2_19[108]}
   );
   gpc1_1 gpc6559 (
      {stage1_19[272]},
      {stage2_19[109]}
   );
   gpc1_1 gpc6560 (
      {stage1_19[273]},
      {stage2_19[110]}
   );
   gpc1_1 gpc6561 (
      {stage1_19[274]},
      {stage2_19[111]}
   );
   gpc1_1 gpc6562 (
      {stage1_19[275]},
      {stage2_19[112]}
   );
   gpc1_1 gpc6563 (
      {stage1_20[262]},
      {stage2_20[87]}
   );
   gpc1_1 gpc6564 (
      {stage1_20[263]},
      {stage2_20[88]}
   );
   gpc1_1 gpc6565 (
      {stage1_20[264]},
      {stage2_20[89]}
   );
   gpc1_1 gpc6566 (
      {stage1_20[265]},
      {stage2_20[90]}
   );
   gpc1_1 gpc6567 (
      {stage1_20[266]},
      {stage2_20[91]}
   );
   gpc1_1 gpc6568 (
      {stage1_20[267]},
      {stage2_20[92]}
   );
   gpc1_1 gpc6569 (
      {stage1_21[174]},
      {stage2_21[112]}
   );
   gpc1_1 gpc6570 (
      {stage1_21[175]},
      {stage2_21[113]}
   );
   gpc1_1 gpc6571 (
      {stage1_21[176]},
      {stage2_21[114]}
   );
   gpc1_1 gpc6572 (
      {stage1_21[177]},
      {stage2_21[115]}
   );
   gpc1_1 gpc6573 (
      {stage1_21[178]},
      {stage2_21[116]}
   );
   gpc1_1 gpc6574 (
      {stage1_21[179]},
      {stage2_21[117]}
   );
   gpc1_1 gpc6575 (
      {stage1_21[180]},
      {stage2_21[118]}
   );
   gpc1_1 gpc6576 (
      {stage1_21[181]},
      {stage2_21[119]}
   );
   gpc1_1 gpc6577 (
      {stage1_21[182]},
      {stage2_21[120]}
   );
   gpc1_1 gpc6578 (
      {stage1_21[183]},
      {stage2_21[121]}
   );
   gpc1_1 gpc6579 (
      {stage1_21[184]},
      {stage2_21[122]}
   );
   gpc1_1 gpc6580 (
      {stage1_21[185]},
      {stage2_21[123]}
   );
   gpc1_1 gpc6581 (
      {stage1_21[186]},
      {stage2_21[124]}
   );
   gpc1_1 gpc6582 (
      {stage1_21[187]},
      {stage2_21[125]}
   );
   gpc1_1 gpc6583 (
      {stage1_21[188]},
      {stage2_21[126]}
   );
   gpc1_1 gpc6584 (
      {stage1_21[189]},
      {stage2_21[127]}
   );
   gpc1_1 gpc6585 (
      {stage1_22[145]},
      {stage2_22[82]}
   );
   gpc1_1 gpc6586 (
      {stage1_22[146]},
      {stage2_22[83]}
   );
   gpc1_1 gpc6587 (
      {stage1_22[147]},
      {stage2_22[84]}
   );
   gpc1_1 gpc6588 (
      {stage1_22[148]},
      {stage2_22[85]}
   );
   gpc1_1 gpc6589 (
      {stage1_22[149]},
      {stage2_22[86]}
   );
   gpc1_1 gpc6590 (
      {stage1_22[150]},
      {stage2_22[87]}
   );
   gpc1_1 gpc6591 (
      {stage1_22[151]},
      {stage2_22[88]}
   );
   gpc1_1 gpc6592 (
      {stage1_22[152]},
      {stage2_22[89]}
   );
   gpc1_1 gpc6593 (
      {stage1_22[153]},
      {stage2_22[90]}
   );
   gpc1_1 gpc6594 (
      {stage1_22[154]},
      {stage2_22[91]}
   );
   gpc1_1 gpc6595 (
      {stage1_22[155]},
      {stage2_22[92]}
   );
   gpc1_1 gpc6596 (
      {stage1_22[156]},
      {stage2_22[93]}
   );
   gpc1_1 gpc6597 (
      {stage1_22[157]},
      {stage2_22[94]}
   );
   gpc1_1 gpc6598 (
      {stage1_22[158]},
      {stage2_22[95]}
   );
   gpc1_1 gpc6599 (
      {stage1_22[159]},
      {stage2_22[96]}
   );
   gpc1_1 gpc6600 (
      {stage1_22[160]},
      {stage2_22[97]}
   );
   gpc1_1 gpc6601 (
      {stage1_22[161]},
      {stage2_22[98]}
   );
   gpc1_1 gpc6602 (
      {stage1_22[162]},
      {stage2_22[99]}
   );
   gpc1_1 gpc6603 (
      {stage1_22[163]},
      {stage2_22[100]}
   );
   gpc1_1 gpc6604 (
      {stage1_22[164]},
      {stage2_22[101]}
   );
   gpc1_1 gpc6605 (
      {stage1_22[165]},
      {stage2_22[102]}
   );
   gpc1_1 gpc6606 (
      {stage1_22[166]},
      {stage2_22[103]}
   );
   gpc1_1 gpc6607 (
      {stage1_22[167]},
      {stage2_22[104]}
   );
   gpc1_1 gpc6608 (
      {stage1_22[168]},
      {stage2_22[105]}
   );
   gpc1_1 gpc6609 (
      {stage1_22[169]},
      {stage2_22[106]}
   );
   gpc1_1 gpc6610 (
      {stage1_22[170]},
      {stage2_22[107]}
   );
   gpc1_1 gpc6611 (
      {stage1_24[210]},
      {stage2_24[98]}
   );
   gpc1_1 gpc6612 (
      {stage1_24[211]},
      {stage2_24[99]}
   );
   gpc1_1 gpc6613 (
      {stage1_24[212]},
      {stage2_24[100]}
   );
   gpc1_1 gpc6614 (
      {stage1_24[213]},
      {stage2_24[101]}
   );
   gpc1_1 gpc6615 (
      {stage1_25[175]},
      {stage2_25[87]}
   );
   gpc1_1 gpc6616 (
      {stage1_25[176]},
      {stage2_25[88]}
   );
   gpc1_1 gpc6617 (
      {stage1_25[177]},
      {stage2_25[89]}
   );
   gpc1_1 gpc6618 (
      {stage1_25[178]},
      {stage2_25[90]}
   );
   gpc1_1 gpc6619 (
      {stage1_25[179]},
      {stage2_25[91]}
   );
   gpc1_1 gpc6620 (
      {stage1_25[180]},
      {stage2_25[92]}
   );
   gpc1_1 gpc6621 (
      {stage1_25[181]},
      {stage2_25[93]}
   );
   gpc1_1 gpc6622 (
      {stage1_25[182]},
      {stage2_25[94]}
   );
   gpc1_1 gpc6623 (
      {stage1_25[183]},
      {stage2_25[95]}
   );
   gpc1_1 gpc6624 (
      {stage1_26[248]},
      {stage2_26[82]}
   );
   gpc1_1 gpc6625 (
      {stage1_26[249]},
      {stage2_26[83]}
   );
   gpc1_1 gpc6626 (
      {stage1_26[250]},
      {stage2_26[84]}
   );
   gpc1_1 gpc6627 (
      {stage1_29[216]},
      {stage2_29[74]}
   );
   gpc1_1 gpc6628 (
      {stage1_29[217]},
      {stage2_29[75]}
   );
   gpc1_1 gpc6629 (
      {stage1_29[218]},
      {stage2_29[76]}
   );
   gpc1_1 gpc6630 (
      {stage1_29[219]},
      {stage2_29[77]}
   );
   gpc1_1 gpc6631 (
      {stage1_29[220]},
      {stage2_29[78]}
   );
   gpc1_1 gpc6632 (
      {stage1_29[221]},
      {stage2_29[79]}
   );
   gpc1_1 gpc6633 (
      {stage1_29[222]},
      {stage2_29[80]}
   );
   gpc1_1 gpc6634 (
      {stage1_29[223]},
      {stage2_29[81]}
   );
   gpc1_1 gpc6635 (
      {stage1_29[224]},
      {stage2_29[82]}
   );
   gpc1_1 gpc6636 (
      {stage1_29[225]},
      {stage2_29[83]}
   );
   gpc1_1 gpc6637 (
      {stage1_29[226]},
      {stage2_29[84]}
   );
   gpc1_1 gpc6638 (
      {stage1_29[227]},
      {stage2_29[85]}
   );
   gpc1_1 gpc6639 (
      {stage1_29[228]},
      {stage2_29[86]}
   );
   gpc1_1 gpc6640 (
      {stage1_30[160]},
      {stage2_30[85]}
   );
   gpc1_1 gpc6641 (
      {stage1_30[161]},
      {stage2_30[86]}
   );
   gpc1_1 gpc6642 (
      {stage1_30[162]},
      {stage2_30[87]}
   );
   gpc1_1 gpc6643 (
      {stage1_30[163]},
      {stage2_30[88]}
   );
   gpc1_1 gpc6644 (
      {stage1_30[164]},
      {stage2_30[89]}
   );
   gpc1_1 gpc6645 (
      {stage1_30[165]},
      {stage2_30[90]}
   );
   gpc1_1 gpc6646 (
      {stage1_30[166]},
      {stage2_30[91]}
   );
   gpc1_1 gpc6647 (
      {stage1_30[167]},
      {stage2_30[92]}
   );
   gpc1_1 gpc6648 (
      {stage1_30[168]},
      {stage2_30[93]}
   );
   gpc1_1 gpc6649 (
      {stage1_30[169]},
      {stage2_30[94]}
   );
   gpc1_1 gpc6650 (
      {stage1_30[170]},
      {stage2_30[95]}
   );
   gpc1_1 gpc6651 (
      {stage1_30[171]},
      {stage2_30[96]}
   );
   gpc1_1 gpc6652 (
      {stage1_30[172]},
      {stage2_30[97]}
   );
   gpc1_1 gpc6653 (
      {stage1_30[173]},
      {stage2_30[98]}
   );
   gpc1_1 gpc6654 (
      {stage1_30[174]},
      {stage2_30[99]}
   );
   gpc1_1 gpc6655 (
      {stage1_30[175]},
      {stage2_30[100]}
   );
   gpc1_1 gpc6656 (
      {stage1_30[176]},
      {stage2_30[101]}
   );
   gpc1_1 gpc6657 (
      {stage1_30[177]},
      {stage2_30[102]}
   );
   gpc1_1 gpc6658 (
      {stage1_30[178]},
      {stage2_30[103]}
   );
   gpc1_1 gpc6659 (
      {stage1_30[179]},
      {stage2_30[104]}
   );
   gpc1_1 gpc6660 (
      {stage1_30[180]},
      {stage2_30[105]}
   );
   gpc1_1 gpc6661 (
      {stage1_30[181]},
      {stage2_30[106]}
   );
   gpc1_1 gpc6662 (
      {stage1_30[182]},
      {stage2_30[107]}
   );
   gpc1_1 gpc6663 (
      {stage1_30[183]},
      {stage2_30[108]}
   );
   gpc1_1 gpc6664 (
      {stage1_30[184]},
      {stage2_30[109]}
   );
   gpc1_1 gpc6665 (
      {stage1_30[185]},
      {stage2_30[110]}
   );
   gpc1_1 gpc6666 (
      {stage1_30[186]},
      {stage2_30[111]}
   );
   gpc1_1 gpc6667 (
      {stage1_30[187]},
      {stage2_30[112]}
   );
   gpc1_1 gpc6668 (
      {stage1_30[188]},
      {stage2_30[113]}
   );
   gpc1_1 gpc6669 (
      {stage1_30[189]},
      {stage2_30[114]}
   );
   gpc1_1 gpc6670 (
      {stage1_30[190]},
      {stage2_30[115]}
   );
   gpc1_1 gpc6671 (
      {stage1_30[191]},
      {stage2_30[116]}
   );
   gpc1_1 gpc6672 (
      {stage1_32[189]},
      {stage2_32[78]}
   );
   gpc1_1 gpc6673 (
      {stage1_32[190]},
      {stage2_32[79]}
   );
   gpc1_1 gpc6674 (
      {stage1_32[191]},
      {stage2_32[80]}
   );
   gpc1_1 gpc6675 (
      {stage1_32[192]},
      {stage2_32[81]}
   );
   gpc1_1 gpc6676 (
      {stage1_32[193]},
      {stage2_32[82]}
   );
   gpc1_1 gpc6677 (
      {stage1_32[194]},
      {stage2_32[83]}
   );
   gpc1_1 gpc6678 (
      {stage1_32[195]},
      {stage2_32[84]}
   );
   gpc1_1 gpc6679 (
      {stage1_32[196]},
      {stage2_32[85]}
   );
   gpc1_1 gpc6680 (
      {stage1_32[197]},
      {stage2_32[86]}
   );
   gpc1_1 gpc6681 (
      {stage1_32[198]},
      {stage2_32[87]}
   );
   gpc1_1 gpc6682 (
      {stage1_32[199]},
      {stage2_32[88]}
   );
   gpc1_1 gpc6683 (
      {stage1_32[200]},
      {stage2_32[89]}
   );
   gpc1_1 gpc6684 (
      {stage1_32[201]},
      {stage2_32[90]}
   );
   gpc1_1 gpc6685 (
      {stage1_32[202]},
      {stage2_32[91]}
   );
   gpc1_1 gpc6686 (
      {stage1_32[203]},
      {stage2_32[92]}
   );
   gpc1_1 gpc6687 (
      {stage1_32[204]},
      {stage2_32[93]}
   );
   gpc1_1 gpc6688 (
      {stage1_32[205]},
      {stage2_32[94]}
   );
   gpc1_1 gpc6689 (
      {stage1_32[206]},
      {stage2_32[95]}
   );
   gpc1_1 gpc6690 (
      {stage1_32[207]},
      {stage2_32[96]}
   );
   gpc1_1 gpc6691 (
      {stage1_32[208]},
      {stage2_32[97]}
   );
   gpc1_1 gpc6692 (
      {stage1_32[209]},
      {stage2_32[98]}
   );
   gpc1_1 gpc6693 (
      {stage1_32[210]},
      {stage2_32[99]}
   );
   gpc1_1 gpc6694 (
      {stage1_32[211]},
      {stage2_32[100]}
   );
   gpc1_1 gpc6695 (
      {stage1_32[212]},
      {stage2_32[101]}
   );
   gpc1_1 gpc6696 (
      {stage1_32[213]},
      {stage2_32[102]}
   );
   gpc1_1 gpc6697 (
      {stage1_32[214]},
      {stage2_32[103]}
   );
   gpc1_1 gpc6698 (
      {stage1_32[215]},
      {stage2_32[104]}
   );
   gpc1_1 gpc6699 (
      {stage1_32[216]},
      {stage2_32[105]}
   );
   gpc1_1 gpc6700 (
      {stage1_34[140]},
      {stage2_34[82]}
   );
   gpc1_1 gpc6701 (
      {stage1_34[141]},
      {stage2_34[83]}
   );
   gpc1_1 gpc6702 (
      {stage1_34[142]},
      {stage2_34[84]}
   );
   gpc1_1 gpc6703 (
      {stage1_34[143]},
      {stage2_34[85]}
   );
   gpc1_1 gpc6704 (
      {stage1_34[144]},
      {stage2_34[86]}
   );
   gpc1_1 gpc6705 (
      {stage1_34[145]},
      {stage2_34[87]}
   );
   gpc1_1 gpc6706 (
      {stage1_34[146]},
      {stage2_34[88]}
   );
   gpc1_1 gpc6707 (
      {stage1_34[147]},
      {stage2_34[89]}
   );
   gpc1_1 gpc6708 (
      {stage1_34[148]},
      {stage2_34[90]}
   );
   gpc1_1 gpc6709 (
      {stage1_34[149]},
      {stage2_34[91]}
   );
   gpc1_1 gpc6710 (
      {stage1_34[150]},
      {stage2_34[92]}
   );
   gpc1_1 gpc6711 (
      {stage1_34[151]},
      {stage2_34[93]}
   );
   gpc1_1 gpc6712 (
      {stage1_34[152]},
      {stage2_34[94]}
   );
   gpc1_1 gpc6713 (
      {stage1_34[153]},
      {stage2_34[95]}
   );
   gpc1_1 gpc6714 (
      {stage1_34[154]},
      {stage2_34[96]}
   );
   gpc1_1 gpc6715 (
      {stage1_34[155]},
      {stage2_34[97]}
   );
   gpc1_1 gpc6716 (
      {stage1_34[156]},
      {stage2_34[98]}
   );
   gpc1_1 gpc6717 (
      {stage1_34[157]},
      {stage2_34[99]}
   );
   gpc1_1 gpc6718 (
      {stage1_34[158]},
      {stage2_34[100]}
   );
   gpc1_1 gpc6719 (
      {stage1_34[159]},
      {stage2_34[101]}
   );
   gpc1_1 gpc6720 (
      {stage1_34[160]},
      {stage2_34[102]}
   );
   gpc1_1 gpc6721 (
      {stage1_34[161]},
      {stage2_34[103]}
   );
   gpc1_1 gpc6722 (
      {stage1_34[162]},
      {stage2_34[104]}
   );
   gpc1_1 gpc6723 (
      {stage1_34[163]},
      {stage2_34[105]}
   );
   gpc1_1 gpc6724 (
      {stage1_34[164]},
      {stage2_34[106]}
   );
   gpc1_1 gpc6725 (
      {stage1_34[165]},
      {stage2_34[107]}
   );
   gpc1_1 gpc6726 (
      {stage1_34[166]},
      {stage2_34[108]}
   );
   gpc1_1 gpc6727 (
      {stage1_34[167]},
      {stage2_34[109]}
   );
   gpc1_1 gpc6728 (
      {stage1_34[168]},
      {stage2_34[110]}
   );
   gpc1_1 gpc6729 (
      {stage1_34[169]},
      {stage2_34[111]}
   );
   gpc1_1 gpc6730 (
      {stage1_34[170]},
      {stage2_34[112]}
   );
   gpc1_1 gpc6731 (
      {stage1_34[171]},
      {stage2_34[113]}
   );
   gpc1_1 gpc6732 (
      {stage1_34[172]},
      {stage2_34[114]}
   );
   gpc1_1 gpc6733 (
      {stage1_34[173]},
      {stage2_34[115]}
   );
   gpc1_1 gpc6734 (
      {stage1_34[174]},
      {stage2_34[116]}
   );
   gpc1_1 gpc6735 (
      {stage1_34[175]},
      {stage2_34[117]}
   );
   gpc1_1 gpc6736 (
      {stage1_34[176]},
      {stage2_34[118]}
   );
   gpc1_1 gpc6737 (
      {stage1_34[177]},
      {stage2_34[119]}
   );
   gpc1_1 gpc6738 (
      {stage1_34[178]},
      {stage2_34[120]}
   );
   gpc1_1 gpc6739 (
      {stage1_34[179]},
      {stage2_34[121]}
   );
   gpc1_1 gpc6740 (
      {stage1_34[180]},
      {stage2_34[122]}
   );
   gpc1_1 gpc6741 (
      {stage1_34[181]},
      {stage2_34[123]}
   );
   gpc1_1 gpc6742 (
      {stage1_34[182]},
      {stage2_34[124]}
   );
   gpc1_1 gpc6743 (
      {stage1_34[183]},
      {stage2_34[125]}
   );
   gpc1_1 gpc6744 (
      {stage1_34[184]},
      {stage2_34[126]}
   );
   gpc1_1 gpc6745 (
      {stage1_34[185]},
      {stage2_34[127]}
   );
   gpc1_1 gpc6746 (
      {stage1_34[186]},
      {stage2_34[128]}
   );
   gpc1_1 gpc6747 (
      {stage1_34[187]},
      {stage2_34[129]}
   );
   gpc1_1 gpc6748 (
      {stage1_34[188]},
      {stage2_34[130]}
   );
   gpc1_1 gpc6749 (
      {stage1_34[189]},
      {stage2_34[131]}
   );
   gpc1_1 gpc6750 (
      {stage1_35[178]},
      {stage2_35[94]}
   );
   gpc1_1 gpc6751 (
      {stage1_35[179]},
      {stage2_35[95]}
   );
   gpc1_1 gpc6752 (
      {stage1_35[180]},
      {stage2_35[96]}
   );
   gpc1_1 gpc6753 (
      {stage1_35[181]},
      {stage2_35[97]}
   );
   gpc1_1 gpc6754 (
      {stage1_35[182]},
      {stage2_35[98]}
   );
   gpc1_1 gpc6755 (
      {stage1_35[183]},
      {stage2_35[99]}
   );
   gpc1_1 gpc6756 (
      {stage1_35[184]},
      {stage2_35[100]}
   );
   gpc1_1 gpc6757 (
      {stage1_35[185]},
      {stage2_35[101]}
   );
   gpc1_1 gpc6758 (
      {stage1_35[186]},
      {stage2_35[102]}
   );
   gpc1_1 gpc6759 (
      {stage1_35[187]},
      {stage2_35[103]}
   );
   gpc1_1 gpc6760 (
      {stage1_35[188]},
      {stage2_35[104]}
   );
   gpc1_1 gpc6761 (
      {stage1_35[189]},
      {stage2_35[105]}
   );
   gpc1_1 gpc6762 (
      {stage1_35[190]},
      {stage2_35[106]}
   );
   gpc1_1 gpc6763 (
      {stage1_35[191]},
      {stage2_35[107]}
   );
   gpc1_1 gpc6764 (
      {stage1_35[192]},
      {stage2_35[108]}
   );
   gpc1_1 gpc6765 (
      {stage1_35[193]},
      {stage2_35[109]}
   );
   gpc1_1 gpc6766 (
      {stage1_35[194]},
      {stage2_35[110]}
   );
   gpc1_1 gpc6767 (
      {stage1_35[195]},
      {stage2_35[111]}
   );
   gpc1_1 gpc6768 (
      {stage1_35[196]},
      {stage2_35[112]}
   );
   gpc1_1 gpc6769 (
      {stage1_35[197]},
      {stage2_35[113]}
   );
   gpc1_1 gpc6770 (
      {stage1_35[198]},
      {stage2_35[114]}
   );
   gpc1_1 gpc6771 (
      {stage1_35[199]},
      {stage2_35[115]}
   );
   gpc1_1 gpc6772 (
      {stage1_35[200]},
      {stage2_35[116]}
   );
   gpc1_1 gpc6773 (
      {stage1_35[201]},
      {stage2_35[117]}
   );
   gpc1_1 gpc6774 (
      {stage1_35[202]},
      {stage2_35[118]}
   );
   gpc1_1 gpc6775 (
      {stage1_35[203]},
      {stage2_35[119]}
   );
   gpc1_1 gpc6776 (
      {stage1_35[204]},
      {stage2_35[120]}
   );
   gpc1_1 gpc6777 (
      {stage1_35[205]},
      {stage2_35[121]}
   );
   gpc1_1 gpc6778 (
      {stage1_35[206]},
      {stage2_35[122]}
   );
   gpc1_1 gpc6779 (
      {stage1_35[207]},
      {stage2_35[123]}
   );
   gpc1_1 gpc6780 (
      {stage1_35[208]},
      {stage2_35[124]}
   );
   gpc1_1 gpc6781 (
      {stage1_35[209]},
      {stage2_35[125]}
   );
   gpc1_1 gpc6782 (
      {stage1_35[210]},
      {stage2_35[126]}
   );
   gpc1_1 gpc6783 (
      {stage1_35[211]},
      {stage2_35[127]}
   );
   gpc1_1 gpc6784 (
      {stage1_35[212]},
      {stage2_35[128]}
   );
   gpc1_1 gpc6785 (
      {stage1_35[213]},
      {stage2_35[129]}
   );
   gpc1_1 gpc6786 (
      {stage1_35[214]},
      {stage2_35[130]}
   );
   gpc1_1 gpc6787 (
      {stage1_35[215]},
      {stage2_35[131]}
   );
   gpc1_1 gpc6788 (
      {stage1_35[216]},
      {stage2_35[132]}
   );
   gpc1_1 gpc6789 (
      {stage1_37[306]},
      {stage2_37[88]}
   );
   gpc1_1 gpc6790 (
      {stage1_37[307]},
      {stage2_37[89]}
   );
   gpc1_1 gpc6791 (
      {stage1_38[231]},
      {stage2_38[106]}
   );
   gpc1_1 gpc6792 (
      {stage1_38[232]},
      {stage2_38[107]}
   );
   gpc1_1 gpc6793 (
      {stage1_38[233]},
      {stage2_38[108]}
   );
   gpc1_1 gpc6794 (
      {stage1_38[234]},
      {stage2_38[109]}
   );
   gpc1_1 gpc6795 (
      {stage1_38[235]},
      {stage2_38[110]}
   );
   gpc1_1 gpc6796 (
      {stage1_38[236]},
      {stage2_38[111]}
   );
   gpc1_1 gpc6797 (
      {stage1_38[237]},
      {stage2_38[112]}
   );
   gpc1_1 gpc6798 (
      {stage1_38[238]},
      {stage2_38[113]}
   );
   gpc1_1 gpc6799 (
      {stage1_38[239]},
      {stage2_38[114]}
   );
   gpc1_1 gpc6800 (
      {stage1_38[240]},
      {stage2_38[115]}
   );
   gpc1_1 gpc6801 (
      {stage1_38[241]},
      {stage2_38[116]}
   );
   gpc1_1 gpc6802 (
      {stage1_38[242]},
      {stage2_38[117]}
   );
   gpc1_1 gpc6803 (
      {stage1_38[243]},
      {stage2_38[118]}
   );
   gpc1_1 gpc6804 (
      {stage1_38[244]},
      {stage2_38[119]}
   );
   gpc1_1 gpc6805 (
      {stage1_38[245]},
      {stage2_38[120]}
   );
   gpc1_1 gpc6806 (
      {stage1_38[246]},
      {stage2_38[121]}
   );
   gpc1_1 gpc6807 (
      {stage1_38[247]},
      {stage2_38[122]}
   );
   gpc1_1 gpc6808 (
      {stage1_38[248]},
      {stage2_38[123]}
   );
   gpc1_1 gpc6809 (
      {stage1_38[249]},
      {stage2_38[124]}
   );
   gpc1_1 gpc6810 (
      {stage1_38[250]},
      {stage2_38[125]}
   );
   gpc1_1 gpc6811 (
      {stage1_38[251]},
      {stage2_38[126]}
   );
   gpc1_1 gpc6812 (
      {stage1_38[252]},
      {stage2_38[127]}
   );
   gpc1_1 gpc6813 (
      {stage1_38[253]},
      {stage2_38[128]}
   );
   gpc1_1 gpc6814 (
      {stage1_38[254]},
      {stage2_38[129]}
   );
   gpc1_1 gpc6815 (
      {stage1_38[255]},
      {stage2_38[130]}
   );
   gpc1_1 gpc6816 (
      {stage1_38[256]},
      {stage2_38[131]}
   );
   gpc1_1 gpc6817 (
      {stage1_38[257]},
      {stage2_38[132]}
   );
   gpc1_1 gpc6818 (
      {stage1_38[258]},
      {stage2_38[133]}
   );
   gpc1_1 gpc6819 (
      {stage1_38[259]},
      {stage2_38[134]}
   );
   gpc1_1 gpc6820 (
      {stage1_38[260]},
      {stage2_38[135]}
   );
   gpc1_1 gpc6821 (
      {stage1_38[261]},
      {stage2_38[136]}
   );
   gpc1_1 gpc6822 (
      {stage1_38[262]},
      {stage2_38[137]}
   );
   gpc1_1 gpc6823 (
      {stage1_38[263]},
      {stage2_38[138]}
   );
   gpc1_1 gpc6824 (
      {stage1_38[264]},
      {stage2_38[139]}
   );
   gpc1_1 gpc6825 (
      {stage1_39[170]},
      {stage2_39[94]}
   );
   gpc1_1 gpc6826 (
      {stage1_39[171]},
      {stage2_39[95]}
   );
   gpc1_1 gpc6827 (
      {stage1_39[172]},
      {stage2_39[96]}
   );
   gpc1_1 gpc6828 (
      {stage1_39[173]},
      {stage2_39[97]}
   );
   gpc1_1 gpc6829 (
      {stage1_39[174]},
      {stage2_39[98]}
   );
   gpc1_1 gpc6830 (
      {stage1_39[175]},
      {stage2_39[99]}
   );
   gpc1_1 gpc6831 (
      {stage1_39[176]},
      {stage2_39[100]}
   );
   gpc1_1 gpc6832 (
      {stage1_39[177]},
      {stage2_39[101]}
   );
   gpc1_1 gpc6833 (
      {stage1_39[178]},
      {stage2_39[102]}
   );
   gpc1_1 gpc6834 (
      {stage1_39[179]},
      {stage2_39[103]}
   );
   gpc1_1 gpc6835 (
      {stage1_39[180]},
      {stage2_39[104]}
   );
   gpc1_1 gpc6836 (
      {stage1_39[181]},
      {stage2_39[105]}
   );
   gpc1_1 gpc6837 (
      {stage1_39[182]},
      {stage2_39[106]}
   );
   gpc1_1 gpc6838 (
      {stage1_39[183]},
      {stage2_39[107]}
   );
   gpc1_1 gpc6839 (
      {stage1_39[184]},
      {stage2_39[108]}
   );
   gpc1_1 gpc6840 (
      {stage1_39[185]},
      {stage2_39[109]}
   );
   gpc1_1 gpc6841 (
      {stage1_39[186]},
      {stage2_39[110]}
   );
   gpc1_1 gpc6842 (
      {stage1_39[187]},
      {stage2_39[111]}
   );
   gpc1_1 gpc6843 (
      {stage1_39[188]},
      {stage2_39[112]}
   );
   gpc1_1 gpc6844 (
      {stage1_39[189]},
      {stage2_39[113]}
   );
   gpc1_1 gpc6845 (
      {stage1_39[190]},
      {stage2_39[114]}
   );
   gpc1_1 gpc6846 (
      {stage1_39[191]},
      {stage2_39[115]}
   );
   gpc1_1 gpc6847 (
      {stage1_39[192]},
      {stage2_39[116]}
   );
   gpc1_1 gpc6848 (
      {stage1_39[193]},
      {stage2_39[117]}
   );
   gpc1_1 gpc6849 (
      {stage1_39[194]},
      {stage2_39[118]}
   );
   gpc1_1 gpc6850 (
      {stage1_39[195]},
      {stage2_39[119]}
   );
   gpc1_1 gpc6851 (
      {stage1_39[196]},
      {stage2_39[120]}
   );
   gpc1_1 gpc6852 (
      {stage1_39[197]},
      {stage2_39[121]}
   );
   gpc1_1 gpc6853 (
      {stage1_39[198]},
      {stage2_39[122]}
   );
   gpc1_1 gpc6854 (
      {stage1_39[199]},
      {stage2_39[123]}
   );
   gpc1_1 gpc6855 (
      {stage1_39[200]},
      {stage2_39[124]}
   );
   gpc1_1 gpc6856 (
      {stage1_39[201]},
      {stage2_39[125]}
   );
   gpc1_1 gpc6857 (
      {stage1_39[202]},
      {stage2_39[126]}
   );
   gpc1_1 gpc6858 (
      {stage1_39[203]},
      {stage2_39[127]}
   );
   gpc1_1 gpc6859 (
      {stage1_39[204]},
      {stage2_39[128]}
   );
   gpc1_1 gpc6860 (
      {stage1_39[205]},
      {stage2_39[129]}
   );
   gpc1_1 gpc6861 (
      {stage1_39[206]},
      {stage2_39[130]}
   );
   gpc1_1 gpc6862 (
      {stage1_39[207]},
      {stage2_39[131]}
   );
   gpc1_1 gpc6863 (
      {stage1_39[208]},
      {stage2_39[132]}
   );
   gpc1_1 gpc6864 (
      {stage1_39[209]},
      {stage2_39[133]}
   );
   gpc1_1 gpc6865 (
      {stage1_39[210]},
      {stage2_39[134]}
   );
   gpc1_1 gpc6866 (
      {stage1_39[211]},
      {stage2_39[135]}
   );
   gpc1_1 gpc6867 (
      {stage1_39[212]},
      {stage2_39[136]}
   );
   gpc1_1 gpc6868 (
      {stage1_40[281]},
      {stage2_40[90]}
   );
   gpc1_1 gpc6869 (
      {stage1_40[282]},
      {stage2_40[91]}
   );
   gpc1_1 gpc6870 (
      {stage1_40[283]},
      {stage2_40[92]}
   );
   gpc1_1 gpc6871 (
      {stage1_40[284]},
      {stage2_40[93]}
   );
   gpc1_1 gpc6872 (
      {stage1_40[285]},
      {stage2_40[94]}
   );
   gpc1_1 gpc6873 (
      {stage1_40[286]},
      {stage2_40[95]}
   );
   gpc1_1 gpc6874 (
      {stage1_40[287]},
      {stage2_40[96]}
   );
   gpc1_1 gpc6875 (
      {stage1_40[288]},
      {stage2_40[97]}
   );
   gpc1_1 gpc6876 (
      {stage1_40[289]},
      {stage2_40[98]}
   );
   gpc1_1 gpc6877 (
      {stage1_40[290]},
      {stage2_40[99]}
   );
   gpc1_1 gpc6878 (
      {stage1_40[291]},
      {stage2_40[100]}
   );
   gpc1_1 gpc6879 (
      {stage1_40[292]},
      {stage2_40[101]}
   );
   gpc1_1 gpc6880 (
      {stage1_40[293]},
      {stage2_40[102]}
   );
   gpc1_1 gpc6881 (
      {stage1_40[294]},
      {stage2_40[103]}
   );
   gpc1_1 gpc6882 (
      {stage1_40[295]},
      {stage2_40[104]}
   );
   gpc1_1 gpc6883 (
      {stage1_40[296]},
      {stage2_40[105]}
   );
   gpc1_1 gpc6884 (
      {stage1_40[297]},
      {stage2_40[106]}
   );
   gpc1_1 gpc6885 (
      {stage1_40[298]},
      {stage2_40[107]}
   );
   gpc1_1 gpc6886 (
      {stage1_40[299]},
      {stage2_40[108]}
   );
   gpc1_1 gpc6887 (
      {stage1_40[300]},
      {stage2_40[109]}
   );
   gpc1_1 gpc6888 (
      {stage1_40[301]},
      {stage2_40[110]}
   );
   gpc1_1 gpc6889 (
      {stage1_40[302]},
      {stage2_40[111]}
   );
   gpc1_1 gpc6890 (
      {stage1_40[303]},
      {stage2_40[112]}
   );
   gpc1_1 gpc6891 (
      {stage1_41[168]},
      {stage2_41[103]}
   );
   gpc1_1 gpc6892 (
      {stage1_41[169]},
      {stage2_41[104]}
   );
   gpc1_1 gpc6893 (
      {stage1_41[170]},
      {stage2_41[105]}
   );
   gpc1_1 gpc6894 (
      {stage1_42[168]},
      {stage2_42[80]}
   );
   gpc1_1 gpc6895 (
      {stage1_42[169]},
      {stage2_42[81]}
   );
   gpc1_1 gpc6896 (
      {stage1_42[170]},
      {stage2_42[82]}
   );
   gpc1_1 gpc6897 (
      {stage1_42[171]},
      {stage2_42[83]}
   );
   gpc1_1 gpc6898 (
      {stage1_42[172]},
      {stage2_42[84]}
   );
   gpc1_1 gpc6899 (
      {stage1_42[173]},
      {stage2_42[85]}
   );
   gpc1_1 gpc6900 (
      {stage1_43[241]},
      {stage2_43[66]}
   );
   gpc1_1 gpc6901 (
      {stage1_43[242]},
      {stage2_43[67]}
   );
   gpc1_1 gpc6902 (
      {stage1_43[243]},
      {stage2_43[68]}
   );
   gpc1_1 gpc6903 (
      {stage1_43[244]},
      {stage2_43[69]}
   );
   gpc1_1 gpc6904 (
      {stage1_43[245]},
      {stage2_43[70]}
   );
   gpc1_1 gpc6905 (
      {stage1_43[246]},
      {stage2_43[71]}
   );
   gpc1_1 gpc6906 (
      {stage1_43[247]},
      {stage2_43[72]}
   );
   gpc1_1 gpc6907 (
      {stage1_43[248]},
      {stage2_43[73]}
   );
   gpc1_1 gpc6908 (
      {stage1_43[249]},
      {stage2_43[74]}
   );
   gpc1_1 gpc6909 (
      {stage1_43[250]},
      {stage2_43[75]}
   );
   gpc1_1 gpc6910 (
      {stage1_43[251]},
      {stage2_43[76]}
   );
   gpc1_1 gpc6911 (
      {stage1_43[252]},
      {stage2_43[77]}
   );
   gpc1_1 gpc6912 (
      {stage1_43[253]},
      {stage2_43[78]}
   );
   gpc1_1 gpc6913 (
      {stage1_44[240]},
      {stage2_44[103]}
   );
   gpc1_1 gpc6914 (
      {stage1_44[241]},
      {stage2_44[104]}
   );
   gpc1_1 gpc6915 (
      {stage1_44[242]},
      {stage2_44[105]}
   );
   gpc1_1 gpc6916 (
      {stage1_44[243]},
      {stage2_44[106]}
   );
   gpc1_1 gpc6917 (
      {stage1_44[244]},
      {stage2_44[107]}
   );
   gpc1_1 gpc6918 (
      {stage1_44[245]},
      {stage2_44[108]}
   );
   gpc1_1 gpc6919 (
      {stage1_44[246]},
      {stage2_44[109]}
   );
   gpc1_1 gpc6920 (
      {stage1_44[247]},
      {stage2_44[110]}
   );
   gpc1_1 gpc6921 (
      {stage1_44[248]},
      {stage2_44[111]}
   );
   gpc1_1 gpc6922 (
      {stage1_44[249]},
      {stage2_44[112]}
   );
   gpc1_1 gpc6923 (
      {stage1_44[250]},
      {stage2_44[113]}
   );
   gpc1_1 gpc6924 (
      {stage1_44[251]},
      {stage2_44[114]}
   );
   gpc1_1 gpc6925 (
      {stage1_44[252]},
      {stage2_44[115]}
   );
   gpc1_1 gpc6926 (
      {stage1_44[253]},
      {stage2_44[116]}
   );
   gpc1_1 gpc6927 (
      {stage1_44[254]},
      {stage2_44[117]}
   );
   gpc1_1 gpc6928 (
      {stage1_44[255]},
      {stage2_44[118]}
   );
   gpc1_1 gpc6929 (
      {stage1_45[199]},
      {stage2_45[105]}
   );
   gpc1_1 gpc6930 (
      {stage1_45[200]},
      {stage2_45[106]}
   );
   gpc1_1 gpc6931 (
      {stage1_45[201]},
      {stage2_45[107]}
   );
   gpc1_1 gpc6932 (
      {stage1_45[202]},
      {stage2_45[108]}
   );
   gpc1_1 gpc6933 (
      {stage1_45[203]},
      {stage2_45[109]}
   );
   gpc1_1 gpc6934 (
      {stage1_45[204]},
      {stage2_45[110]}
   );
   gpc1_1 gpc6935 (
      {stage1_45[205]},
      {stage2_45[111]}
   );
   gpc1_1 gpc6936 (
      {stage1_45[206]},
      {stage2_45[112]}
   );
   gpc1_1 gpc6937 (
      {stage1_45[207]},
      {stage2_45[113]}
   );
   gpc1_1 gpc6938 (
      {stage1_45[208]},
      {stage2_45[114]}
   );
   gpc1_1 gpc6939 (
      {stage1_45[209]},
      {stage2_45[115]}
   );
   gpc1_1 gpc6940 (
      {stage1_45[210]},
      {stage2_45[116]}
   );
   gpc1_1 gpc6941 (
      {stage1_45[211]},
      {stage2_45[117]}
   );
   gpc1_1 gpc6942 (
      {stage1_46[295]},
      {stage2_46[85]}
   );
   gpc1_1 gpc6943 (
      {stage1_46[296]},
      {stage2_46[86]}
   );
   gpc1_1 gpc6944 (
      {stage1_46[297]},
      {stage2_46[87]}
   );
   gpc1_1 gpc6945 (
      {stage1_47[230]},
      {stage2_47[98]}
   );
   gpc1_1 gpc6946 (
      {stage1_47[231]},
      {stage2_47[99]}
   );
   gpc1_1 gpc6947 (
      {stage1_47[232]},
      {stage2_47[100]}
   );
   gpc1_1 gpc6948 (
      {stage1_47[233]},
      {stage2_47[101]}
   );
   gpc1_1 gpc6949 (
      {stage1_47[234]},
      {stage2_47[102]}
   );
   gpc1_1 gpc6950 (
      {stage1_47[235]},
      {stage2_47[103]}
   );
   gpc1_1 gpc6951 (
      {stage1_48[172]},
      {stage2_48[104]}
   );
   gpc1_1 gpc6952 (
      {stage1_48[173]},
      {stage2_48[105]}
   );
   gpc1_1 gpc6953 (
      {stage1_48[174]},
      {stage2_48[106]}
   );
   gpc1_1 gpc6954 (
      {stage1_48[175]},
      {stage2_48[107]}
   );
   gpc1_1 gpc6955 (
      {stage1_48[176]},
      {stage2_48[108]}
   );
   gpc1_1 gpc6956 (
      {stage1_48[177]},
      {stage2_48[109]}
   );
   gpc1_1 gpc6957 (
      {stage1_48[178]},
      {stage2_48[110]}
   );
   gpc1_1 gpc6958 (
      {stage1_48[179]},
      {stage2_48[111]}
   );
   gpc1_1 gpc6959 (
      {stage1_48[180]},
      {stage2_48[112]}
   );
   gpc1_1 gpc6960 (
      {stage1_48[181]},
      {stage2_48[113]}
   );
   gpc1_1 gpc6961 (
      {stage1_48[182]},
      {stage2_48[114]}
   );
   gpc1_1 gpc6962 (
      {stage1_48[183]},
      {stage2_48[115]}
   );
   gpc1_1 gpc6963 (
      {stage1_48[184]},
      {stage2_48[116]}
   );
   gpc1_1 gpc6964 (
      {stage1_48[185]},
      {stage2_48[117]}
   );
   gpc1_1 gpc6965 (
      {stage1_48[186]},
      {stage2_48[118]}
   );
   gpc1_1 gpc6966 (
      {stage1_48[187]},
      {stage2_48[119]}
   );
   gpc1_1 gpc6967 (
      {stage1_48[188]},
      {stage2_48[120]}
   );
   gpc1_1 gpc6968 (
      {stage1_48[189]},
      {stage2_48[121]}
   );
   gpc1_1 gpc6969 (
      {stage1_48[190]},
      {stage2_48[122]}
   );
   gpc1_1 gpc6970 (
      {stage1_48[191]},
      {stage2_48[123]}
   );
   gpc1_1 gpc6971 (
      {stage1_48[192]},
      {stage2_48[124]}
   );
   gpc1_1 gpc6972 (
      {stage1_48[193]},
      {stage2_48[125]}
   );
   gpc1_1 gpc6973 (
      {stage1_48[194]},
      {stage2_48[126]}
   );
   gpc1_1 gpc6974 (
      {stage1_48[195]},
      {stage2_48[127]}
   );
   gpc1_1 gpc6975 (
      {stage1_48[196]},
      {stage2_48[128]}
   );
   gpc1_1 gpc6976 (
      {stage1_48[197]},
      {stage2_48[129]}
   );
   gpc1_1 gpc6977 (
      {stage1_49[154]},
      {stage2_49[77]}
   );
   gpc1_1 gpc6978 (
      {stage1_49[155]},
      {stage2_49[78]}
   );
   gpc1_1 gpc6979 (
      {stage1_49[156]},
      {stage2_49[79]}
   );
   gpc1_1 gpc6980 (
      {stage1_49[157]},
      {stage2_49[80]}
   );
   gpc1_1 gpc6981 (
      {stage1_49[158]},
      {stage2_49[81]}
   );
   gpc1_1 gpc6982 (
      {stage1_49[159]},
      {stage2_49[82]}
   );
   gpc1_1 gpc6983 (
      {stage1_49[160]},
      {stage2_49[83]}
   );
   gpc1_1 gpc6984 (
      {stage1_49[161]},
      {stage2_49[84]}
   );
   gpc1_1 gpc6985 (
      {stage1_49[162]},
      {stage2_49[85]}
   );
   gpc1_1 gpc6986 (
      {stage1_49[163]},
      {stage2_49[86]}
   );
   gpc1_1 gpc6987 (
      {stage1_49[164]},
      {stage2_49[87]}
   );
   gpc1_1 gpc6988 (
      {stage1_49[165]},
      {stage2_49[88]}
   );
   gpc1_1 gpc6989 (
      {stage1_49[166]},
      {stage2_49[89]}
   );
   gpc1_1 gpc6990 (
      {stage1_49[167]},
      {stage2_49[90]}
   );
   gpc1_1 gpc6991 (
      {stage1_49[168]},
      {stage2_49[91]}
   );
   gpc1_1 gpc6992 (
      {stage1_49[169]},
      {stage2_49[92]}
   );
   gpc1_1 gpc6993 (
      {stage1_49[170]},
      {stage2_49[93]}
   );
   gpc1_1 gpc6994 (
      {stage1_49[171]},
      {stage2_49[94]}
   );
   gpc1_1 gpc6995 (
      {stage1_49[172]},
      {stage2_49[95]}
   );
   gpc1_1 gpc6996 (
      {stage1_50[179]},
      {stage2_50[75]}
   );
   gpc1_1 gpc6997 (
      {stage1_50[180]},
      {stage2_50[76]}
   );
   gpc1_1 gpc6998 (
      {stage1_50[181]},
      {stage2_50[77]}
   );
   gpc1_1 gpc6999 (
      {stage1_50[182]},
      {stage2_50[78]}
   );
   gpc1_1 gpc7000 (
      {stage1_50[183]},
      {stage2_50[79]}
   );
   gpc1_1 gpc7001 (
      {stage1_50[184]},
      {stage2_50[80]}
   );
   gpc1_1 gpc7002 (
      {stage1_50[185]},
      {stage2_50[81]}
   );
   gpc1_1 gpc7003 (
      {stage1_50[186]},
      {stage2_50[82]}
   );
   gpc1_1 gpc7004 (
      {stage1_50[187]},
      {stage2_50[83]}
   );
   gpc1_1 gpc7005 (
      {stage1_50[188]},
      {stage2_50[84]}
   );
   gpc1_1 gpc7006 (
      {stage1_50[189]},
      {stage2_50[85]}
   );
   gpc1_1 gpc7007 (
      {stage1_51[266]},
      {stage2_51[79]}
   );
   gpc1_1 gpc7008 (
      {stage1_51[267]},
      {stage2_51[80]}
   );
   gpc1_1 gpc7009 (
      {stage1_51[268]},
      {stage2_51[81]}
   );
   gpc1_1 gpc7010 (
      {stage1_51[269]},
      {stage2_51[82]}
   );
   gpc1_1 gpc7011 (
      {stage1_51[270]},
      {stage2_51[83]}
   );
   gpc1_1 gpc7012 (
      {stage1_51[271]},
      {stage2_51[84]}
   );
   gpc1_1 gpc7013 (
      {stage1_51[272]},
      {stage2_51[85]}
   );
   gpc1_1 gpc7014 (
      {stage1_51[273]},
      {stage2_51[86]}
   );
   gpc1_1 gpc7015 (
      {stage1_51[274]},
      {stage2_51[87]}
   );
   gpc1_1 gpc7016 (
      {stage1_52[187]},
      {stage2_52[93]}
   );
   gpc1_1 gpc7017 (
      {stage1_52[188]},
      {stage2_52[94]}
   );
   gpc1_1 gpc7018 (
      {stage1_52[189]},
      {stage2_52[95]}
   );
   gpc1_1 gpc7019 (
      {stage1_52[190]},
      {stage2_52[96]}
   );
   gpc1_1 gpc7020 (
      {stage1_52[191]},
      {stage2_52[97]}
   );
   gpc1_1 gpc7021 (
      {stage1_52[192]},
      {stage2_52[98]}
   );
   gpc1_1 gpc7022 (
      {stage1_52[193]},
      {stage2_52[99]}
   );
   gpc1_1 gpc7023 (
      {stage1_52[194]},
      {stage2_52[100]}
   );
   gpc1_1 gpc7024 (
      {stage1_52[195]},
      {stage2_52[101]}
   );
   gpc1_1 gpc7025 (
      {stage1_52[196]},
      {stage2_52[102]}
   );
   gpc1_1 gpc7026 (
      {stage1_52[197]},
      {stage2_52[103]}
   );
   gpc1_1 gpc7027 (
      {stage1_52[198]},
      {stage2_52[104]}
   );
   gpc1_1 gpc7028 (
      {stage1_53[130]},
      {stage2_53[76]}
   );
   gpc1_1 gpc7029 (
      {stage1_53[131]},
      {stage2_53[77]}
   );
   gpc1_1 gpc7030 (
      {stage1_53[132]},
      {stage2_53[78]}
   );
   gpc1_1 gpc7031 (
      {stage1_53[133]},
      {stage2_53[79]}
   );
   gpc1_1 gpc7032 (
      {stage1_53[134]},
      {stage2_53[80]}
   );
   gpc1_1 gpc7033 (
      {stage1_53[135]},
      {stage2_53[81]}
   );
   gpc1_1 gpc7034 (
      {stage1_53[136]},
      {stage2_53[82]}
   );
   gpc1_1 gpc7035 (
      {stage1_53[137]},
      {stage2_53[83]}
   );
   gpc1_1 gpc7036 (
      {stage1_53[138]},
      {stage2_53[84]}
   );
   gpc1_1 gpc7037 (
      {stage1_53[139]},
      {stage2_53[85]}
   );
   gpc1_1 gpc7038 (
      {stage1_53[140]},
      {stage2_53[86]}
   );
   gpc1_1 gpc7039 (
      {stage1_53[141]},
      {stage2_53[87]}
   );
   gpc1_1 gpc7040 (
      {stage1_53[142]},
      {stage2_53[88]}
   );
   gpc1_1 gpc7041 (
      {stage1_53[143]},
      {stage2_53[89]}
   );
   gpc1_1 gpc7042 (
      {stage1_53[144]},
      {stage2_53[90]}
   );
   gpc1_1 gpc7043 (
      {stage1_53[145]},
      {stage2_53[91]}
   );
   gpc1_1 gpc7044 (
      {stage1_53[146]},
      {stage2_53[92]}
   );
   gpc1_1 gpc7045 (
      {stage1_53[147]},
      {stage2_53[93]}
   );
   gpc1_1 gpc7046 (
      {stage1_53[148]},
      {stage2_53[94]}
   );
   gpc1_1 gpc7047 (
      {stage1_53[149]},
      {stage2_53[95]}
   );
   gpc1_1 gpc7048 (
      {stage1_53[150]},
      {stage2_53[96]}
   );
   gpc1_1 gpc7049 (
      {stage1_53[151]},
      {stage2_53[97]}
   );
   gpc1_1 gpc7050 (
      {stage1_53[152]},
      {stage2_53[98]}
   );
   gpc1_1 gpc7051 (
      {stage1_53[153]},
      {stage2_53[99]}
   );
   gpc1_1 gpc7052 (
      {stage1_53[154]},
      {stage2_53[100]}
   );
   gpc1_1 gpc7053 (
      {stage1_53[155]},
      {stage2_53[101]}
   );
   gpc1_1 gpc7054 (
      {stage1_53[156]},
      {stage2_53[102]}
   );
   gpc1_1 gpc7055 (
      {stage1_53[157]},
      {stage2_53[103]}
   );
   gpc1_1 gpc7056 (
      {stage1_53[158]},
      {stage2_53[104]}
   );
   gpc1_1 gpc7057 (
      {stage1_53[159]},
      {stage2_53[105]}
   );
   gpc1_1 gpc7058 (
      {stage1_53[160]},
      {stage2_53[106]}
   );
   gpc1_1 gpc7059 (
      {stage1_53[161]},
      {stage2_53[107]}
   );
   gpc1_1 gpc7060 (
      {stage1_53[162]},
      {stage2_53[108]}
   );
   gpc1_1 gpc7061 (
      {stage1_53[163]},
      {stage2_53[109]}
   );
   gpc1_1 gpc7062 (
      {stage1_53[164]},
      {stage2_53[110]}
   );
   gpc1_1 gpc7063 (
      {stage1_53[165]},
      {stage2_53[111]}
   );
   gpc1_1 gpc7064 (
      {stage1_53[166]},
      {stage2_53[112]}
   );
   gpc1_1 gpc7065 (
      {stage1_53[167]},
      {stage2_53[113]}
   );
   gpc1_1 gpc7066 (
      {stage1_53[168]},
      {stage2_53[114]}
   );
   gpc1_1 gpc7067 (
      {stage1_54[203]},
      {stage2_54[72]}
   );
   gpc1_1 gpc7068 (
      {stage1_54[204]},
      {stage2_54[73]}
   );
   gpc1_1 gpc7069 (
      {stage1_54[205]},
      {stage2_54[74]}
   );
   gpc1_1 gpc7070 (
      {stage1_54[206]},
      {stage2_54[75]}
   );
   gpc1_1 gpc7071 (
      {stage1_54[207]},
      {stage2_54[76]}
   );
   gpc1_1 gpc7072 (
      {stage1_54[208]},
      {stage2_54[77]}
   );
   gpc1_1 gpc7073 (
      {stage1_54[209]},
      {stage2_54[78]}
   );
   gpc1_1 gpc7074 (
      {stage1_54[210]},
      {stage2_54[79]}
   );
   gpc1_1 gpc7075 (
      {stage1_54[211]},
      {stage2_54[80]}
   );
   gpc1_1 gpc7076 (
      {stage1_54[212]},
      {stage2_54[81]}
   );
   gpc1_1 gpc7077 (
      {stage1_54[213]},
      {stage2_54[82]}
   );
   gpc1_1 gpc7078 (
      {stage1_54[214]},
      {stage2_54[83]}
   );
   gpc1_1 gpc7079 (
      {stage1_54[215]},
      {stage2_54[84]}
   );
   gpc1_1 gpc7080 (
      {stage1_54[216]},
      {stage2_54[85]}
   );
   gpc1_1 gpc7081 (
      {stage1_54[217]},
      {stage2_54[86]}
   );
   gpc1_1 gpc7082 (
      {stage1_54[218]},
      {stage2_54[87]}
   );
   gpc1_1 gpc7083 (
      {stage1_54[219]},
      {stage2_54[88]}
   );
   gpc1_1 gpc7084 (
      {stage1_54[220]},
      {stage2_54[89]}
   );
   gpc1_1 gpc7085 (
      {stage1_54[221]},
      {stage2_54[90]}
   );
   gpc1_1 gpc7086 (
      {stage1_54[222]},
      {stage2_54[91]}
   );
   gpc1_1 gpc7087 (
      {stage1_54[223]},
      {stage2_54[92]}
   );
   gpc1_1 gpc7088 (
      {stage1_54[224]},
      {stage2_54[93]}
   );
   gpc1_1 gpc7089 (
      {stage1_54[225]},
      {stage2_54[94]}
   );
   gpc1_1 gpc7090 (
      {stage1_54[226]},
      {stage2_54[95]}
   );
   gpc1_1 gpc7091 (
      {stage1_54[227]},
      {stage2_54[96]}
   );
   gpc1_1 gpc7092 (
      {stage1_54[228]},
      {stage2_54[97]}
   );
   gpc1_1 gpc7093 (
      {stage1_54[229]},
      {stage2_54[98]}
   );
   gpc1_1 gpc7094 (
      {stage1_54[230]},
      {stage2_54[99]}
   );
   gpc1_1 gpc7095 (
      {stage1_55[254]},
      {stage2_55[93]}
   );
   gpc1_1 gpc7096 (
      {stage1_55[255]},
      {stage2_55[94]}
   );
   gpc1_1 gpc7097 (
      {stage1_55[256]},
      {stage2_55[95]}
   );
   gpc1_1 gpc7098 (
      {stage1_55[257]},
      {stage2_55[96]}
   );
   gpc1_1 gpc7099 (
      {stage1_55[258]},
      {stage2_55[97]}
   );
   gpc1_1 gpc7100 (
      {stage1_55[259]},
      {stage2_55[98]}
   );
   gpc1_1 gpc7101 (
      {stage1_55[260]},
      {stage2_55[99]}
   );
   gpc1_1 gpc7102 (
      {stage1_55[261]},
      {stage2_55[100]}
   );
   gpc1_1 gpc7103 (
      {stage1_55[262]},
      {stage2_55[101]}
   );
   gpc1_1 gpc7104 (
      {stage1_55[263]},
      {stage2_55[102]}
   );
   gpc1_1 gpc7105 (
      {stage1_55[264]},
      {stage2_55[103]}
   );
   gpc1_1 gpc7106 (
      {stage1_55[265]},
      {stage2_55[104]}
   );
   gpc1_1 gpc7107 (
      {stage1_55[266]},
      {stage2_55[105]}
   );
   gpc1_1 gpc7108 (
      {stage1_56[164]},
      {stage2_56[92]}
   );
   gpc1_1 gpc7109 (
      {stage1_56[165]},
      {stage2_56[93]}
   );
   gpc1_1 gpc7110 (
      {stage1_56[166]},
      {stage2_56[94]}
   );
   gpc1_1 gpc7111 (
      {stage1_56[167]},
      {stage2_56[95]}
   );
   gpc1_1 gpc7112 (
      {stage1_56[168]},
      {stage2_56[96]}
   );
   gpc1_1 gpc7113 (
      {stage1_56[169]},
      {stage2_56[97]}
   );
   gpc1_1 gpc7114 (
      {stage1_56[170]},
      {stage2_56[98]}
   );
   gpc1_1 gpc7115 (
      {stage1_56[171]},
      {stage2_56[99]}
   );
   gpc1_1 gpc7116 (
      {stage1_56[172]},
      {stage2_56[100]}
   );
   gpc1_1 gpc7117 (
      {stage1_56[173]},
      {stage2_56[101]}
   );
   gpc1_1 gpc7118 (
      {stage1_56[174]},
      {stage2_56[102]}
   );
   gpc1_1 gpc7119 (
      {stage1_56[175]},
      {stage2_56[103]}
   );
   gpc1_1 gpc7120 (
      {stage1_56[176]},
      {stage2_56[104]}
   );
   gpc1_1 gpc7121 (
      {stage1_56[177]},
      {stage2_56[105]}
   );
   gpc1_1 gpc7122 (
      {stage1_56[178]},
      {stage2_56[106]}
   );
   gpc1_1 gpc7123 (
      {stage1_56[179]},
      {stage2_56[107]}
   );
   gpc1_1 gpc7124 (
      {stage1_56[180]},
      {stage2_56[108]}
   );
   gpc1_1 gpc7125 (
      {stage1_56[181]},
      {stage2_56[109]}
   );
   gpc1_1 gpc7126 (
      {stage1_56[182]},
      {stage2_56[110]}
   );
   gpc1_1 gpc7127 (
      {stage1_56[183]},
      {stage2_56[111]}
   );
   gpc1_1 gpc7128 (
      {stage1_56[184]},
      {stage2_56[112]}
   );
   gpc1_1 gpc7129 (
      {stage1_56[185]},
      {stage2_56[113]}
   );
   gpc1_1 gpc7130 (
      {stage1_56[186]},
      {stage2_56[114]}
   );
   gpc1_1 gpc7131 (
      {stage1_59[205]},
      {stage2_59[109]}
   );
   gpc1_1 gpc7132 (
      {stage1_60[209]},
      {stage2_60[79]}
   );
   gpc1_1 gpc7133 (
      {stage1_60[210]},
      {stage2_60[80]}
   );
   gpc1_1 gpc7134 (
      {stage1_60[211]},
      {stage2_60[81]}
   );
   gpc1_1 gpc7135 (
      {stage1_60[212]},
      {stage2_60[82]}
   );
   gpc1_1 gpc7136 (
      {stage1_60[213]},
      {stage2_60[83]}
   );
   gpc1_1 gpc7137 (
      {stage1_60[214]},
      {stage2_60[84]}
   );
   gpc1_1 gpc7138 (
      {stage1_62[192]},
      {stage2_62[104]}
   );
   gpc1_1 gpc7139 (
      {stage1_63[303]},
      {stage2_63[94]}
   );
   gpc1_1 gpc7140 (
      {stage1_63[304]},
      {stage2_63[95]}
   );
   gpc1_1 gpc7141 (
      {stage1_63[305]},
      {stage2_63[96]}
   );
   gpc1_1 gpc7142 (
      {stage1_63[306]},
      {stage2_63[97]}
   );
   gpc1_1 gpc7143 (
      {stage1_63[307]},
      {stage2_63[98]}
   );
   gpc1_1 gpc7144 (
      {stage1_64[47]},
      {stage2_64[65]}
   );
   gpc1_1 gpc7145 (
      {stage1_64[48]},
      {stage2_64[66]}
   );
   gpc1_1 gpc7146 (
      {stage1_64[49]},
      {stage2_64[67]}
   );
   gpc1_1 gpc7147 (
      {stage1_64[50]},
      {stage2_64[68]}
   );
   gpc1_1 gpc7148 (
      {stage1_64[51]},
      {stage2_64[69]}
   );
   gpc1_1 gpc7149 (
      {stage1_64[52]},
      {stage2_64[70]}
   );
   gpc1_1 gpc7150 (
      {stage1_64[53]},
      {stage2_64[71]}
   );
   gpc1_1 gpc7151 (
      {stage1_64[54]},
      {stage2_64[72]}
   );
   gpc1_1 gpc7152 (
      {stage1_64[55]},
      {stage2_64[73]}
   );
   gpc1_1 gpc7153 (
      {stage1_64[56]},
      {stage2_64[74]}
   );
   gpc1_1 gpc7154 (
      {stage1_64[57]},
      {stage2_64[75]}
   );
   gpc1_1 gpc7155 (
      {stage1_64[58]},
      {stage2_64[76]}
   );
   gpc1_1 gpc7156 (
      {stage1_64[59]},
      {stage2_64[77]}
   );
   gpc1_1 gpc7157 (
      {stage1_64[60]},
      {stage2_64[78]}
   );
   gpc1_1 gpc7158 (
      {stage1_64[61]},
      {stage2_64[79]}
   );
   gpc1_1 gpc7159 (
      {stage1_64[62]},
      {stage2_64[80]}
   );
   gpc1_1 gpc7160 (
      {stage1_64[63]},
      {stage2_64[81]}
   );
   gpc1_1 gpc7161 (
      {stage1_64[64]},
      {stage2_64[82]}
   );
   gpc1_1 gpc7162 (
      {stage1_64[65]},
      {stage2_64[83]}
   );
   gpc1_1 gpc7163 (
      {stage1_64[66]},
      {stage2_64[84]}
   );
   gpc1_1 gpc7164 (
      {stage1_64[67]},
      {stage2_64[85]}
   );
   gpc1_1 gpc7165 (
      {stage1_64[68]},
      {stage2_64[86]}
   );
   gpc1_1 gpc7166 (
      {stage1_64[69]},
      {stage2_64[87]}
   );
   gpc1_1 gpc7167 (
      {stage1_64[70]},
      {stage2_64[88]}
   );
   gpc1_1 gpc7168 (
      {stage1_64[71]},
      {stage2_64[89]}
   );
   gpc1_1 gpc7169 (
      {stage1_64[72]},
      {stage2_64[90]}
   );
   gpc1_1 gpc7170 (
      {stage1_64[73]},
      {stage2_64[91]}
   );
   gpc1_1 gpc7171 (
      {stage1_64[74]},
      {stage2_64[92]}
   );
   gpc1_1 gpc7172 (
      {stage1_64[75]},
      {stage2_64[93]}
   );
   gpc1_1 gpc7173 (
      {stage1_64[76]},
      {stage2_64[94]}
   );
   gpc1_1 gpc7174 (
      {stage1_64[77]},
      {stage2_64[95]}
   );
   gpc1_1 gpc7175 (
      {stage1_64[78]},
      {stage2_64[96]}
   );
   gpc1_1 gpc7176 (
      {stage1_64[79]},
      {stage2_64[97]}
   );
   gpc1_1 gpc7177 (
      {stage1_64[80]},
      {stage2_64[98]}
   );
   gpc1_1 gpc7178 (
      {stage1_64[81]},
      {stage2_64[99]}
   );
   gpc1_1 gpc7179 (
      {stage1_64[82]},
      {stage2_64[100]}
   );
   gpc1_1 gpc7180 (
      {stage1_64[83]},
      {stage2_64[101]}
   );
   gpc1_1 gpc7181 (
      {stage1_64[84]},
      {stage2_64[102]}
   );
   gpc1_1 gpc7182 (
      {stage1_64[85]},
      {stage2_64[103]}
   );
   gpc1_1 gpc7183 (
      {stage1_64[86]},
      {stage2_64[104]}
   );
   gpc1_1 gpc7184 (
      {stage1_64[87]},
      {stage2_64[105]}
   );
   gpc1_1 gpc7185 (
      {stage1_64[88]},
      {stage2_64[106]}
   );
   gpc1_1 gpc7186 (
      {stage1_64[89]},
      {stage2_64[107]}
   );
   gpc1_1 gpc7187 (
      {stage1_64[90]},
      {stage2_64[108]}
   );
   gpc1_1 gpc7188 (
      {stage1_64[91]},
      {stage2_64[109]}
   );
   gpc1_1 gpc7189 (
      {stage1_64[92]},
      {stage2_64[110]}
   );
   gpc1_1 gpc7190 (
      {stage1_64[93]},
      {stage2_64[111]}
   );
   gpc1_1 gpc7191 (
      {stage1_64[94]},
      {stage2_64[112]}
   );
   gpc1_1 gpc7192 (
      {stage1_64[95]},
      {stage2_64[113]}
   );
   gpc1_1 gpc7193 (
      {stage1_64[96]},
      {stage2_64[114]}
   );
   gpc1_1 gpc7194 (
      {stage1_64[97]},
      {stage2_64[115]}
   );
   gpc1_1 gpc7195 (
      {stage1_64[98]},
      {stage2_64[116]}
   );
   gpc1_1 gpc7196 (
      {stage1_64[99]},
      {stage2_64[117]}
   );
   gpc1_1 gpc7197 (
      {stage1_64[100]},
      {stage2_64[118]}
   );
   gpc1_1 gpc7198 (
      {stage1_64[101]},
      {stage2_64[119]}
   );
   gpc1_1 gpc7199 (
      {stage1_64[102]},
      {stage2_64[120]}
   );
   gpc1_1 gpc7200 (
      {stage1_64[103]},
      {stage2_64[121]}
   );
   gpc1_1 gpc7201 (
      {stage1_64[104]},
      {stage2_64[122]}
   );
   gpc1_1 gpc7202 (
      {stage1_64[105]},
      {stage2_64[123]}
   );
   gpc1_1 gpc7203 (
      {stage1_64[106]},
      {stage2_64[124]}
   );
   gpc1_1 gpc7204 (
      {stage1_64[107]},
      {stage2_64[125]}
   );
   gpc1_1 gpc7205 (
      {stage1_64[108]},
      {stage2_64[126]}
   );
   gpc1_1 gpc7206 (
      {stage1_64[109]},
      {stage2_64[127]}
   );
   gpc1_1 gpc7207 (
      {stage1_64[110]},
      {stage2_64[128]}
   );
   gpc1_1 gpc7208 (
      {stage1_64[111]},
      {stage2_64[129]}
   );
   gpc1_1 gpc7209 (
      {stage1_64[112]},
      {stage2_64[130]}
   );
   gpc1_1 gpc7210 (
      {stage1_64[113]},
      {stage2_64[131]}
   );
   gpc1_1 gpc7211 (
      {stage1_64[114]},
      {stage2_64[132]}
   );
   gpc1_1 gpc7212 (
      {stage1_64[115]},
      {stage2_64[133]}
   );
   gpc1_1 gpc7213 (
      {stage1_64[116]},
      {stage2_64[134]}
   );
   gpc1_1 gpc7214 (
      {stage1_64[117]},
      {stage2_64[135]}
   );
   gpc1_1 gpc7215 (
      {stage1_64[118]},
      {stage2_64[136]}
   );
   gpc1_1 gpc7216 (
      {stage1_64[119]},
      {stage2_64[137]}
   );
   gpc1_1 gpc7217 (
      {stage1_64[120]},
      {stage2_64[138]}
   );
   gpc1_1 gpc7218 (
      {stage1_64[121]},
      {stage2_64[139]}
   );
   gpc1_1 gpc7219 (
      {stage1_64[122]},
      {stage2_64[140]}
   );
   gpc1_1 gpc7220 (
      {stage1_64[123]},
      {stage2_64[141]}
   );
   gpc1_1 gpc7221 (
      {stage1_65[49]},
      {stage2_65[51]}
   );
   gpc1_1 gpc7222 (
      {stage1_65[50]},
      {stage2_65[52]}
   );
   gpc1_1 gpc7223 (
      {stage1_65[51]},
      {stage2_65[53]}
   );
   gpc1_1 gpc7224 (
      {stage1_65[52]},
      {stage2_65[54]}
   );
   gpc1_1 gpc7225 (
      {stage1_65[53]},
      {stage2_65[55]}
   );
   gpc1343_5 gpc7226 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3]},
      {stage2_2[0], stage2_2[1], stage2_2[2]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1343_5 gpc7227 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7]},
      {stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1343_5 gpc7228 (
      {stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[6], stage2_2[7], stage2_2[8]},
      {stage2_3[2]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc1343_5 gpc7229 (
      {stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15]},
      {stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_3[3]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc2135_5 gpc7230 (
      {stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15], stage2_0[16]},
      {stage2_1[16], stage2_1[17], stage2_1[18]},
      {stage2_2[12]},
      {stage2_3[4], stage2_3[5]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc606_5 gpc7231 (
      {stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20], stage2_0[21], stage2_0[22]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc606_5 gpc7232 (
      {stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23], stage2_1[24]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[0],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc7233 (
      {stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29], stage2_1[30]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[1],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc7234 (
      {stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35], stage2_1[36]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[2],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc615_5 gpc7235 (
      {stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_2[19]},
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage3_5[3],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc7236 (
      {stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24], stage2_2[25]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[4],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc606_5 gpc7237 (
      {stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30], stage2_2[31]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[5],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc7238 (
      {stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34]},
      {stage2_4[12]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[2],stage3_5[6],stage3_4[12],stage3_3[12]}
   );
   gpc615_5 gpc7239 (
      {stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39]},
      {stage2_4[13]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[3],stage3_5[7],stage3_4[13],stage3_3[13]}
   );
   gpc615_5 gpc7240 (
      {stage2_3[40], stage2_3[41], stage2_3[42], stage2_3[43], stage2_3[44]},
      {stage2_4[14]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[4],stage3_5[8],stage3_4[14],stage3_3[14]}
   );
   gpc615_5 gpc7241 (
      {stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48], stage2_3[49]},
      {stage2_4[15]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[5],stage3_5[9],stage3_4[15],stage3_3[15]}
   );
   gpc615_5 gpc7242 (
      {stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53], stage2_3[54]},
      {stage2_4[16]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[6],stage3_5[10],stage3_4[16],stage3_3[16]}
   );
   gpc615_5 gpc7243 (
      {stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58], stage2_3[59]},
      {stage2_4[17]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[7],stage3_5[11],stage3_4[17],stage3_3[17]}
   );
   gpc615_5 gpc7244 (
      {stage2_3[60], stage2_3[61], stage2_3[62], stage2_3[63], stage2_3[64]},
      {stage2_4[18]},
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage3_7[6],stage3_6[8],stage3_5[12],stage3_4[18],stage3_3[18]}
   );
   gpc615_5 gpc7245 (
      {stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68], stage2_3[69]},
      {stage2_4[19]},
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage3_7[7],stage3_6[9],stage3_5[13],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc7246 (
      {stage2_3[70], stage2_3[71], stage2_3[72], stage2_3[73], stage2_3[74]},
      {stage2_4[20]},
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage3_7[8],stage3_6[10],stage3_5[14],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc7247 (
      {stage2_3[75], stage2_3[76], stage2_3[77], stage2_3[78], stage2_3[79]},
      {stage2_4[21]},
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage3_7[9],stage3_6[11],stage3_5[15],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc7248 (
      {stage2_3[80], stage2_3[81], stage2_3[82], stage2_3[83], stage2_3[84]},
      {stage2_4[22]},
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage3_7[10],stage3_6[12],stage3_5[16],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc7249 (
      {stage2_3[85], stage2_3[86], stage2_3[87], stage2_3[88], stage2_3[89]},
      {stage2_4[23]},
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage3_7[11],stage3_6[13],stage3_5[17],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc7250 (
      {stage2_3[90], stage2_3[91], stage2_3[92], stage2_3[93], stage2_3[94]},
      {stage2_4[24]},
      {stage2_5[72], stage2_5[73], stage2_5[74], stage2_5[75], stage2_5[76], stage2_5[77]},
      {stage3_7[12],stage3_6[14],stage3_5[18],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc7251 (
      {stage2_3[95], stage2_3[96], stage2_3[97], stage2_3[98], stage2_3[99]},
      {stage2_4[25]},
      {stage2_5[78], stage2_5[79], stage2_5[80], stage2_5[81], stage2_5[82], stage2_5[83]},
      {stage3_7[13],stage3_6[15],stage3_5[19],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc7252 (
      {stage2_3[100], stage2_3[101], stage2_3[102], stage2_3[103], stage2_3[104]},
      {stage2_4[26]},
      {stage2_5[84], stage2_5[85], stage2_5[86], stage2_5[87], stage2_5[88], stage2_5[89]},
      {stage3_7[14],stage3_6[16],stage3_5[20],stage3_4[26],stage3_3[26]}
   );
   gpc615_5 gpc7253 (
      {stage2_3[105], stage2_3[106], stage2_3[107], stage2_3[108], stage2_3[109]},
      {stage2_4[27]},
      {stage2_5[90], stage2_5[91], stage2_5[92], stage2_5[93], stage2_5[94], stage2_5[95]},
      {stage3_7[15],stage3_6[17],stage3_5[21],stage3_4[27],stage3_3[27]}
   );
   gpc615_5 gpc7254 (
      {stage2_3[110], stage2_3[111], stage2_3[112], stage2_3[113], 1'b0},
      {stage2_4[28]},
      {stage2_5[96], stage2_5[97], stage2_5[98], stage2_5[99], stage2_5[100], stage2_5[101]},
      {stage3_7[16],stage3_6[18],stage3_5[22],stage3_4[28],stage3_3[28]}
   );
   gpc606_5 gpc7255 (
      {stage2_5[102], stage2_5[103], stage2_5[104], stage2_5[105], stage2_5[106], stage2_5[107]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[17],stage3_6[19],stage3_5[23]}
   );
   gpc606_5 gpc7256 (
      {stage2_5[108], stage2_5[109], stage2_5[110], stage2_5[111], stage2_5[112], stage2_5[113]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[1],stage3_7[18],stage3_6[20],stage3_5[24]}
   );
   gpc606_5 gpc7257 (
      {stage2_5[114], stage2_5[115], stage2_5[116], stage2_5[117], stage2_5[118], stage2_5[119]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[2],stage3_7[19],stage3_6[21],stage3_5[25]}
   );
   gpc606_5 gpc7258 (
      {stage2_5[120], stage2_5[121], stage2_5[122], stage2_5[123], stage2_5[124], stage2_5[125]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[3],stage3_7[20],stage3_6[22],stage3_5[26]}
   );
   gpc606_5 gpc7259 (
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[4],stage3_8[4],stage3_7[21],stage3_6[23]}
   );
   gpc615_5 gpc7260 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10]},
      {stage2_7[24]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[5],stage3_8[5],stage3_7[22],stage3_6[24]}
   );
   gpc615_5 gpc7261 (
      {stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15]},
      {stage2_7[25]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[6],stage3_8[6],stage3_7[23],stage3_6[25]}
   );
   gpc615_5 gpc7262 (
      {stage2_6[16], stage2_6[17], stage2_6[18], stage2_6[19], stage2_6[20]},
      {stage2_7[26]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[7],stage3_8[7],stage3_7[24],stage3_6[26]}
   );
   gpc615_5 gpc7263 (
      {stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24], stage2_6[25]},
      {stage2_7[27]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[8],stage3_8[8],stage3_7[25],stage3_6[27]}
   );
   gpc615_5 gpc7264 (
      {stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29], stage2_6[30]},
      {stage2_7[28]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[9],stage3_8[9],stage3_7[26],stage3_6[28]}
   );
   gpc615_5 gpc7265 (
      {stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_7[29]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[10],stage3_8[10],stage3_7[27],stage3_6[29]}
   );
   gpc615_5 gpc7266 (
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40]},
      {stage2_7[30]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[11],stage3_8[11],stage3_7[28],stage3_6[30]}
   );
   gpc615_5 gpc7267 (
      {stage2_6[41], stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45]},
      {stage2_7[31]},
      {stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage3_10[8],stage3_9[12],stage3_8[12],stage3_7[29],stage3_6[31]}
   );
   gpc615_5 gpc7268 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[54]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[9],stage3_9[13],stage3_8[13],stage3_7[30]}
   );
   gpc615_5 gpc7269 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[55]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[10],stage3_9[14],stage3_8[14],stage3_7[31]}
   );
   gpc615_5 gpc7270 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[56]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[11],stage3_9[15],stage3_8[15],stage3_7[32]}
   );
   gpc615_5 gpc7271 (
      {stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_8[57]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[12],stage3_9[16],stage3_8[16],stage3_7[33]}
   );
   gpc615_5 gpc7272 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[58]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[13],stage3_9[17],stage3_8[17],stage3_7[34]}
   );
   gpc606_5 gpc7273 (
      {stage2_8[59], stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[5],stage3_10[14],stage3_9[18],stage3_8[18]}
   );
   gpc606_5 gpc7274 (
      {stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[6],stage3_10[15],stage3_9[19],stage3_8[19]}
   );
   gpc606_5 gpc7275 (
      {stage2_8[71], stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[7],stage3_10[16],stage3_9[20],stage3_8[20]}
   );
   gpc606_5 gpc7276 (
      {stage2_8[77], stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81], stage2_8[82]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[8],stage3_10[17],stage3_9[21],stage3_8[21]}
   );
   gpc606_5 gpc7277 (
      {stage2_8[83], stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87], stage2_8[88]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[9],stage3_10[18],stage3_9[22],stage3_8[22]}
   );
   gpc606_5 gpc7278 (
      {stage2_8[89], stage2_8[90], stage2_8[91], stage2_8[92], stage2_8[93], stage2_8[94]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[10],stage3_10[19],stage3_9[23],stage3_8[23]}
   );
   gpc606_5 gpc7279 (
      {stage2_8[95], stage2_8[96], stage2_8[97], stage2_8[98], stage2_8[99], stage2_8[100]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[11],stage3_10[20],stage3_9[24],stage3_8[24]}
   );
   gpc606_5 gpc7280 (
      {stage2_8[101], stage2_8[102], stage2_8[103], stage2_8[104], stage2_8[105], stage2_8[106]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[7],stage3_11[12],stage3_10[21],stage3_9[25],stage3_8[25]}
   );
   gpc606_5 gpc7281 (
      {stage2_8[107], stage2_8[108], stage2_8[109], stage2_8[110], stage2_8[111], stage2_8[112]},
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage3_12[8],stage3_11[13],stage3_10[22],stage3_9[26],stage3_8[26]}
   );
   gpc606_5 gpc7282 (
      {stage2_8[113], stage2_8[114], stage2_8[115], stage2_8[116], stage2_8[117], stage2_8[118]},
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage3_12[9],stage3_11[14],stage3_10[23],stage3_9[27],stage3_8[27]}
   );
   gpc606_5 gpc7283 (
      {stage2_8[119], stage2_8[120], stage2_8[121], stage2_8[122], stage2_8[123], stage2_8[124]},
      {stage2_10[60], stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65]},
      {stage3_12[10],stage3_11[15],stage3_10[24],stage3_9[28],stage3_8[28]}
   );
   gpc606_5 gpc7284 (
      {stage2_8[125], stage2_8[126], stage2_8[127], stage2_8[128], stage2_8[129], stage2_8[130]},
      {stage2_10[66], stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage3_12[11],stage3_11[16],stage3_10[25],stage3_9[29],stage3_8[29]}
   );
   gpc606_5 gpc7285 (
      {stage2_8[131], stage2_8[132], stage2_8[133], stage2_8[134], stage2_8[135], stage2_8[136]},
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76], stage2_10[77]},
      {stage3_12[12],stage3_11[17],stage3_10[26],stage3_9[30],stage3_8[30]}
   );
   gpc606_5 gpc7286 (
      {stage2_8[137], stage2_8[138], stage2_8[139], stage2_8[140], stage2_8[141], stage2_8[142]},
      {stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81], stage2_10[82], stage2_10[83]},
      {stage3_12[13],stage3_11[18],stage3_10[27],stage3_9[31],stage3_8[31]}
   );
   gpc606_5 gpc7287 (
      {stage2_8[143], stage2_8[144], stage2_8[145], stage2_8[146], stage2_8[147], stage2_8[148]},
      {stage2_10[84], stage2_10[85], stage2_10[86], stage2_10[87], stage2_10[88], stage2_10[89]},
      {stage3_12[14],stage3_11[19],stage3_10[28],stage3_9[32],stage3_8[32]}
   );
   gpc606_5 gpc7288 (
      {stage2_8[149], stage2_8[150], stage2_8[151], stage2_8[152], stage2_8[153], stage2_8[154]},
      {stage2_10[90], stage2_10[91], stage2_10[92], stage2_10[93], stage2_10[94], stage2_10[95]},
      {stage3_12[15],stage3_11[20],stage3_10[29],stage3_9[33],stage3_8[33]}
   );
   gpc606_5 gpc7289 (
      {stage2_8[155], stage2_8[156], stage2_8[157], stage2_8[158], stage2_8[159], 1'b0},
      {stage2_10[96], stage2_10[97], stage2_10[98], stage2_10[99], stage2_10[100], stage2_10[101]},
      {stage3_12[16],stage3_11[21],stage3_10[30],stage3_9[34],stage3_8[34]}
   );
   gpc606_5 gpc7290 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[17],stage3_11[22],stage3_10[31],stage3_9[35]}
   );
   gpc606_5 gpc7291 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[18],stage3_11[23],stage3_10[32],stage3_9[36]}
   );
   gpc606_5 gpc7292 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[19],stage3_11[24],stage3_10[33],stage3_9[37]}
   );
   gpc606_5 gpc7293 (
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[20],stage3_11[25],stage3_10[34],stage3_9[38]}
   );
   gpc606_5 gpc7294 (
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage3_13[4],stage3_12[21],stage3_11[26],stage3_10[35],stage3_9[39]}
   );
   gpc606_5 gpc7295 (
      {stage2_9[60], stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage3_13[5],stage3_12[22],stage3_11[27],stage3_10[36],stage3_9[40]}
   );
   gpc606_5 gpc7296 (
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71]},
      {stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41]},
      {stage3_13[6],stage3_12[23],stage3_11[28],stage3_10[37],stage3_9[41]}
   );
   gpc606_5 gpc7297 (
      {stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77]},
      {stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47]},
      {stage3_13[7],stage3_12[24],stage3_11[29],stage3_10[38],stage3_9[42]}
   );
   gpc606_5 gpc7298 (
      {stage2_9[78], stage2_9[79], stage2_9[80], stage2_9[81], stage2_9[82], stage2_9[83]},
      {stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53]},
      {stage3_13[8],stage3_12[25],stage3_11[30],stage3_10[39],stage3_9[43]}
   );
   gpc606_5 gpc7299 (
      {stage2_9[84], stage2_9[85], stage2_9[86], stage2_9[87], stage2_9[88], stage2_9[89]},
      {stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59]},
      {stage3_13[9],stage3_12[26],stage3_11[31],stage3_10[40],stage3_9[44]}
   );
   gpc606_5 gpc7300 (
      {stage2_9[90], stage2_9[91], stage2_9[92], stage2_9[93], stage2_9[94], stage2_9[95]},
      {stage2_11[60], stage2_11[61], stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65]},
      {stage3_13[10],stage3_12[27],stage3_11[32],stage3_10[41],stage3_9[45]}
   );
   gpc606_5 gpc7301 (
      {stage2_9[96], stage2_9[97], stage2_9[98], stage2_9[99], stage2_9[100], stage2_9[101]},
      {stage2_11[66], stage2_11[67], stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71]},
      {stage3_13[11],stage3_12[28],stage3_11[33],stage3_10[42],stage3_9[46]}
   );
   gpc606_5 gpc7302 (
      {stage2_9[102], stage2_9[103], stage2_9[104], stage2_9[105], stage2_9[106], stage2_9[107]},
      {stage2_11[72], stage2_11[73], stage2_11[74], stage2_11[75], stage2_11[76], stage2_11[77]},
      {stage3_13[12],stage3_12[29],stage3_11[34],stage3_10[43],stage3_9[47]}
   );
   gpc606_5 gpc7303 (
      {stage2_9[108], stage2_9[109], stage2_9[110], stage2_9[111], stage2_9[112], stage2_9[113]},
      {stage2_11[78], stage2_11[79], stage2_11[80], stage2_11[81], stage2_11[82], stage2_11[83]},
      {stage3_13[13],stage3_12[30],stage3_11[35],stage3_10[44],stage3_9[48]}
   );
   gpc606_5 gpc7304 (
      {stage2_9[114], stage2_9[115], stage2_9[116], stage2_9[117], stage2_9[118], stage2_9[119]},
      {stage2_11[84], stage2_11[85], stage2_11[86], stage2_11[87], stage2_11[88], stage2_11[89]},
      {stage3_13[14],stage3_12[31],stage3_11[36],stage3_10[45],stage3_9[49]}
   );
   gpc606_5 gpc7305 (
      {stage2_9[120], stage2_9[121], stage2_9[122], stage2_9[123], stage2_9[124], stage2_9[125]},
      {stage2_11[90], stage2_11[91], stage2_11[92], stage2_11[93], stage2_11[94], stage2_11[95]},
      {stage3_13[15],stage3_12[32],stage3_11[37],stage3_10[46],stage3_9[50]}
   );
   gpc606_5 gpc7306 (
      {stage2_9[126], stage2_9[127], stage2_9[128], stage2_9[129], stage2_9[130], stage2_9[131]},
      {stage2_11[96], stage2_11[97], stage2_11[98], stage2_11[99], stage2_11[100], stage2_11[101]},
      {stage3_13[16],stage3_12[33],stage3_11[38],stage3_10[47],stage3_9[51]}
   );
   gpc606_5 gpc7307 (
      {stage2_9[132], stage2_9[133], stage2_9[134], stage2_9[135], stage2_9[136], stage2_9[137]},
      {stage2_11[102], stage2_11[103], stage2_11[104], stage2_11[105], stage2_11[106], stage2_11[107]},
      {stage3_13[17],stage3_12[34],stage3_11[39],stage3_10[48],stage3_9[52]}
   );
   gpc606_5 gpc7308 (
      {stage2_9[138], stage2_9[139], stage2_9[140], stage2_9[141], stage2_9[142], 1'b0},
      {stage2_11[108], stage2_11[109], stage2_11[110], stage2_11[111], stage2_11[112], stage2_11[113]},
      {stage3_13[18],stage3_12[35],stage3_11[40],stage3_10[49],stage3_9[53]}
   );
   gpc615_5 gpc7309 (
      {stage2_10[102], stage2_10[103], stage2_10[104], stage2_10[105], stage2_10[106]},
      {stage2_11[114]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[19],stage3_12[36],stage3_11[41],stage3_10[50]}
   );
   gpc615_5 gpc7310 (
      {stage2_10[107], stage2_10[108], stage2_10[109], stage2_10[110], stage2_10[111]},
      {stage2_11[115]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[20],stage3_12[37],stage3_11[42],stage3_10[51]}
   );
   gpc615_5 gpc7311 (
      {stage2_10[112], stage2_10[113], stage2_10[114], stage2_10[115], stage2_10[116]},
      {stage2_11[116]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[21],stage3_12[38],stage3_11[43],stage3_10[52]}
   );
   gpc615_5 gpc7312 (
      {stage2_11[117], stage2_11[118], stage2_11[119], stage2_11[120], stage2_11[121]},
      {stage2_12[18]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[22],stage3_12[39],stage3_11[44]}
   );
   gpc615_5 gpc7313 (
      {stage2_11[122], stage2_11[123], stage2_11[124], stage2_11[125], stage2_11[126]},
      {stage2_12[19]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[23],stage3_12[40],stage3_11[45]}
   );
   gpc606_5 gpc7314 (
      {stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[5],stage3_13[24],stage3_12[41]}
   );
   gpc606_5 gpc7315 (
      {stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30], stage2_12[31]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[3],stage3_14[6],stage3_13[25],stage3_12[42]}
   );
   gpc606_5 gpc7316 (
      {stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[4],stage3_14[7],stage3_13[26],stage3_12[43]}
   );
   gpc606_5 gpc7317 (
      {stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[5],stage3_14[8],stage3_13[27],stage3_12[44]}
   );
   gpc606_5 gpc7318 (
      {stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47], stage2_12[48], stage2_12[49]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[6],stage3_14[9],stage3_13[28],stage3_12[45]}
   );
   gpc606_5 gpc7319 (
      {stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53], stage2_12[54], stage2_12[55]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[7],stage3_14[10],stage3_13[29],stage3_12[46]}
   );
   gpc606_5 gpc7320 (
      {stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59], stage2_12[60], stage2_12[61]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[8],stage3_14[11],stage3_13[30],stage3_12[47]}
   );
   gpc606_5 gpc7321 (
      {stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[9],stage3_14[12],stage3_13[31],stage3_12[48]}
   );
   gpc606_5 gpc7322 (
      {stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72], stage2_12[73]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[10],stage3_14[13],stage3_13[32],stage3_12[49]}
   );
   gpc606_5 gpc7323 (
      {stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77], stage2_12[78], stage2_12[79]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[11],stage3_14[14],stage3_13[33],stage3_12[50]}
   );
   gpc606_5 gpc7324 (
      {stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83], stage2_12[84], stage2_12[85]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[12],stage3_14[15],stage3_13[34],stage3_12[51]}
   );
   gpc606_5 gpc7325 (
      {stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89], stage2_12[90], stage2_12[91]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[13],stage3_14[16],stage3_13[35],stage3_12[52]}
   );
   gpc606_5 gpc7326 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[12],stage3_15[14],stage3_14[17],stage3_13[36]}
   );
   gpc606_5 gpc7327 (
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[13],stage3_15[15],stage3_14[18],stage3_13[37]}
   );
   gpc606_5 gpc7328 (
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[14],stage3_15[16],stage3_14[19],stage3_13[38]}
   );
   gpc606_5 gpc7329 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[15],stage3_15[17],stage3_14[20],stage3_13[39]}
   );
   gpc606_5 gpc7330 (
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[16],stage3_15[18],stage3_14[21],stage3_13[40]}
   );
   gpc606_5 gpc7331 (
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34], stage2_15[35]},
      {stage3_17[5],stage3_16[17],stage3_15[19],stage3_14[22],stage3_13[41]}
   );
   gpc606_5 gpc7332 (
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41]},
      {stage3_17[6],stage3_16[18],stage3_15[20],stage3_14[23],stage3_13[42]}
   );
   gpc606_5 gpc7333 (
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage3_17[7],stage3_16[19],stage3_15[21],stage3_14[24],stage3_13[43]}
   );
   gpc606_5 gpc7334 (
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53]},
      {stage3_17[8],stage3_16[20],stage3_15[22],stage3_14[25],stage3_13[44]}
   );
   gpc606_5 gpc7335 (
      {stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[9],stage3_16[21],stage3_15[23],stage3_14[26]}
   );
   gpc606_5 gpc7336 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82], stage2_14[83]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[10],stage3_16[22],stage3_15[24],stage3_14[27]}
   );
   gpc606_5 gpc7337 (
      {stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87], stage2_14[88], stage2_14[89]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[11],stage3_16[23],stage3_15[25],stage3_14[28]}
   );
   gpc606_5 gpc7338 (
      {stage2_14[90], stage2_14[91], stage2_14[92], stage2_14[93], stage2_14[94], stage2_14[95]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[12],stage3_16[24],stage3_15[26],stage3_14[29]}
   );
   gpc606_5 gpc7339 (
      {stage2_14[96], stage2_14[97], stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[13],stage3_16[25],stage3_15[27],stage3_14[30]}
   );
   gpc606_5 gpc7340 (
      {stage2_14[102], stage2_14[103], stage2_14[104], stage2_14[105], stage2_14[106], stage2_14[107]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[14],stage3_16[26],stage3_15[28],stage3_14[31]}
   );
   gpc207_4 gpc7341 (
      {stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58], stage2_15[59], stage2_15[60]},
      {stage2_17[0], stage2_17[1]},
      {stage3_18[6],stage3_17[15],stage3_16[27],stage3_15[29]}
   );
   gpc207_4 gpc7342 (
      {stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64], stage2_15[65], stage2_15[66], stage2_15[67]},
      {stage2_17[2], stage2_17[3]},
      {stage3_18[7],stage3_17[16],stage3_16[28],stage3_15[30]}
   );
   gpc615_5 gpc7343 (
      {stage2_15[68], stage2_15[69], stage2_15[70], stage2_15[71], stage2_15[72]},
      {stage2_16[36]},
      {stage2_17[4], stage2_17[5], stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9]},
      {stage3_19[0],stage3_18[8],stage3_17[17],stage3_16[29],stage3_15[31]}
   );
   gpc615_5 gpc7344 (
      {stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76], stage2_15[77]},
      {stage2_16[37]},
      {stage2_17[10], stage2_17[11], stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15]},
      {stage3_19[1],stage3_18[9],stage3_17[18],stage3_16[30],stage3_15[32]}
   );
   gpc615_5 gpc7345 (
      {stage2_15[78], stage2_15[79], stage2_15[80], stage2_15[81], stage2_15[82]},
      {stage2_16[38]},
      {stage2_17[16], stage2_17[17], stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21]},
      {stage3_19[2],stage3_18[10],stage3_17[19],stage3_16[31],stage3_15[33]}
   );
   gpc615_5 gpc7346 (
      {stage2_15[83], stage2_15[84], stage2_15[85], stage2_15[86], stage2_15[87]},
      {stage2_16[39]},
      {stage2_17[22], stage2_17[23], stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27]},
      {stage3_19[3],stage3_18[11],stage3_17[20],stage3_16[32],stage3_15[34]}
   );
   gpc615_5 gpc7347 (
      {stage2_15[88], stage2_15[89], stage2_15[90], stage2_15[91], stage2_15[92]},
      {stage2_16[40]},
      {stage2_17[28], stage2_17[29], stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33]},
      {stage3_19[4],stage3_18[12],stage3_17[21],stage3_16[33],stage3_15[35]}
   );
   gpc615_5 gpc7348 (
      {stage2_15[93], stage2_15[94], stage2_15[95], stage2_15[96], stage2_15[97]},
      {stage2_16[41]},
      {stage2_17[34], stage2_17[35], stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39]},
      {stage3_19[5],stage3_18[13],stage3_17[22],stage3_16[34],stage3_15[36]}
   );
   gpc615_5 gpc7349 (
      {stage2_15[98], stage2_15[99], stage2_15[100], stage2_15[101], stage2_15[102]},
      {stage2_16[42]},
      {stage2_17[40], stage2_17[41], stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45]},
      {stage3_19[6],stage3_18[14],stage3_17[23],stage3_16[35],stage3_15[37]}
   );
   gpc615_5 gpc7350 (
      {stage2_15[103], stage2_15[104], stage2_15[105], stage2_15[106], stage2_15[107]},
      {stage2_16[43]},
      {stage2_17[46], stage2_17[47], stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51]},
      {stage3_19[7],stage3_18[15],stage3_17[24],stage3_16[36],stage3_15[38]}
   );
   gpc615_5 gpc7351 (
      {stage2_15[108], stage2_15[109], stage2_15[110], stage2_15[111], stage2_15[112]},
      {stage2_16[44]},
      {stage2_17[52], stage2_17[53], stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57]},
      {stage3_19[8],stage3_18[16],stage3_17[25],stage3_16[37],stage3_15[39]}
   );
   gpc615_5 gpc7352 (
      {stage2_15[113], stage2_15[114], stage2_15[115], stage2_15[116], stage2_15[117]},
      {stage2_16[45]},
      {stage2_17[58], stage2_17[59], stage2_17[60], stage2_17[61], stage2_17[62], stage2_17[63]},
      {stage3_19[9],stage3_18[17],stage3_17[26],stage3_16[38],stage3_15[40]}
   );
   gpc615_5 gpc7353 (
      {stage2_15[118], stage2_15[119], stage2_15[120], stage2_15[121], stage2_15[122]},
      {stage2_16[46]},
      {stage2_17[64], stage2_17[65], stage2_17[66], stage2_17[67], stage2_17[68], stage2_17[69]},
      {stage3_19[10],stage3_18[18],stage3_17[27],stage3_16[39],stage3_15[41]}
   );
   gpc615_5 gpc7354 (
      {stage2_15[123], stage2_15[124], stage2_15[125], stage2_15[126], stage2_15[127]},
      {stage2_16[47]},
      {stage2_17[70], stage2_17[71], stage2_17[72], stage2_17[73], stage2_17[74], stage2_17[75]},
      {stage3_19[11],stage3_18[19],stage3_17[28],stage3_16[40],stage3_15[42]}
   );
   gpc615_5 gpc7355 (
      {stage2_15[128], stage2_15[129], stage2_15[130], stage2_15[131], stage2_15[132]},
      {stage2_16[48]},
      {stage2_17[76], stage2_17[77], stage2_17[78], stage2_17[79], stage2_17[80], stage2_17[81]},
      {stage3_19[12],stage3_18[20],stage3_17[29],stage3_16[41],stage3_15[43]}
   );
   gpc615_5 gpc7356 (
      {stage2_15[133], stage2_15[134], stage2_15[135], stage2_15[136], stage2_15[137]},
      {stage2_16[49]},
      {stage2_17[82], stage2_17[83], stage2_17[84], stage2_17[85], stage2_17[86], 1'b0},
      {stage3_19[13],stage3_18[21],stage3_17[30],stage3_16[42],stage3_15[44]}
   );
   gpc606_5 gpc7357 (
      {stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53], stage2_16[54], stage2_16[55]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[14],stage3_18[22],stage3_17[31],stage3_16[43]}
   );
   gpc606_5 gpc7358 (
      {stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59], stage2_16[60], stage2_16[61]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[15],stage3_18[23],stage3_17[32],stage3_16[44]}
   );
   gpc606_5 gpc7359 (
      {stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65], stage2_16[66], stage2_16[67]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[16],stage3_18[24],stage3_17[33],stage3_16[45]}
   );
   gpc606_5 gpc7360 (
      {stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71], stage2_16[72], stage2_16[73]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[17],stage3_18[25],stage3_17[34],stage3_16[46]}
   );
   gpc606_5 gpc7361 (
      {stage2_16[74], stage2_16[75], stage2_16[76], stage2_16[77], stage2_16[78], stage2_16[79]},
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage3_20[4],stage3_19[18],stage3_18[26],stage3_17[35],stage3_16[47]}
   );
   gpc2135_5 gpc7362 (
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34]},
      {stage2_19[0], stage2_19[1], stage2_19[2]},
      {stage2_20[0]},
      {stage2_21[0], stage2_21[1]},
      {stage3_22[0],stage3_21[0],stage3_20[5],stage3_19[19],stage3_18[27]}
   );
   gpc2135_5 gpc7363 (
      {stage2_18[35], stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39]},
      {stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage2_20[1]},
      {stage2_21[2], stage2_21[3]},
      {stage3_22[1],stage3_21[1],stage3_20[6],stage3_19[20],stage3_18[28]}
   );
   gpc2135_5 gpc7364 (
      {stage2_18[40], stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44]},
      {stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage2_20[2]},
      {stage2_21[4], stage2_21[5]},
      {stage3_22[2],stage3_21[2],stage3_20[7],stage3_19[21],stage3_18[29]}
   );
   gpc2135_5 gpc7365 (
      {stage2_18[45], stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49]},
      {stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage2_20[3]},
      {stage2_21[6], stage2_21[7]},
      {stage3_22[3],stage3_21[3],stage3_20[8],stage3_19[22],stage3_18[30]}
   );
   gpc2135_5 gpc7366 (
      {stage2_18[50], stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54]},
      {stage2_19[12], stage2_19[13], stage2_19[14]},
      {stage2_20[4]},
      {stage2_21[8], stage2_21[9]},
      {stage3_22[4],stage3_21[4],stage3_20[9],stage3_19[23],stage3_18[31]}
   );
   gpc2135_5 gpc7367 (
      {stage2_18[55], stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59]},
      {stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_20[5]},
      {stage2_21[10], stage2_21[11]},
      {stage3_22[5],stage3_21[5],stage3_20[10],stage3_19[24],stage3_18[32]}
   );
   gpc2135_5 gpc7368 (
      {stage2_18[60], stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64]},
      {stage2_19[18], stage2_19[19], stage2_19[20]},
      {stage2_20[6]},
      {stage2_21[12], stage2_21[13]},
      {stage3_22[6],stage3_21[6],stage3_20[11],stage3_19[25],stage3_18[33]}
   );
   gpc2135_5 gpc7369 (
      {stage2_18[65], stage2_18[66], stage2_18[67], stage2_18[68], stage2_18[69]},
      {stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage2_20[7]},
      {stage2_21[14], stage2_21[15]},
      {stage3_22[7],stage3_21[7],stage3_20[12],stage3_19[26],stage3_18[34]}
   );
   gpc2135_5 gpc7370 (
      {stage2_18[70], stage2_18[71], stage2_18[72], stage2_18[73], stage2_18[74]},
      {stage2_19[24], stage2_19[25], stage2_19[26]},
      {stage2_20[8]},
      {stage2_21[16], stage2_21[17]},
      {stage3_22[8],stage3_21[8],stage3_20[13],stage3_19[27],stage3_18[35]}
   );
   gpc2135_5 gpc7371 (
      {stage2_18[75], stage2_18[76], stage2_18[77], stage2_18[78], stage2_18[79]},
      {stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_20[9]},
      {stage2_21[18], stage2_21[19]},
      {stage3_22[9],stage3_21[9],stage3_20[14],stage3_19[28],stage3_18[36]}
   );
   gpc2135_5 gpc7372 (
      {stage2_18[80], stage2_18[81], stage2_18[82], stage2_18[83], stage2_18[84]},
      {stage2_19[30], stage2_19[31], stage2_19[32]},
      {stage2_20[10]},
      {stage2_21[20], stage2_21[21]},
      {stage3_22[10],stage3_21[10],stage3_20[15],stage3_19[29],stage3_18[37]}
   );
   gpc2135_5 gpc7373 (
      {stage2_18[85], stage2_18[86], stage2_18[87], stage2_18[88], stage2_18[89]},
      {stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage2_20[11]},
      {stage2_21[22], stage2_21[23]},
      {stage3_22[11],stage3_21[11],stage3_20[16],stage3_19[30],stage3_18[38]}
   );
   gpc615_5 gpc7374 (
      {stage2_18[90], stage2_18[91], stage2_18[92], stage2_18[93], stage2_18[94]},
      {stage2_19[36]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[12],stage3_21[12],stage3_20[17],stage3_19[31],stage3_18[39]}
   );
   gpc615_5 gpc7375 (
      {stage2_18[95], stage2_18[96], stage2_18[97], stage2_18[98], stage2_18[99]},
      {stage2_19[37]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[13],stage3_21[13],stage3_20[18],stage3_19[32],stage3_18[40]}
   );
   gpc615_5 gpc7376 (
      {stage2_19[38], stage2_19[39], stage2_19[40], stage2_19[41], stage2_19[42]},
      {stage2_20[24]},
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage3_23[0],stage3_22[14],stage3_21[14],stage3_20[19],stage3_19[33]}
   );
   gpc615_5 gpc7377 (
      {stage2_19[43], stage2_19[44], stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage2_20[25]},
      {stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33], stage2_21[34], stage2_21[35]},
      {stage3_23[1],stage3_22[15],stage3_21[15],stage3_20[20],stage3_19[34]}
   );
   gpc615_5 gpc7378 (
      {stage2_19[48], stage2_19[49], stage2_19[50], stage2_19[51], stage2_19[52]},
      {stage2_20[26]},
      {stage2_21[36], stage2_21[37], stage2_21[38], stage2_21[39], stage2_21[40], stage2_21[41]},
      {stage3_23[2],stage3_22[16],stage3_21[16],stage3_20[21],stage3_19[35]}
   );
   gpc615_5 gpc7379 (
      {stage2_19[53], stage2_19[54], stage2_19[55], stage2_19[56], stage2_19[57]},
      {stage2_20[27]},
      {stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47]},
      {stage3_23[3],stage3_22[17],stage3_21[17],stage3_20[22],stage3_19[36]}
   );
   gpc615_5 gpc7380 (
      {stage2_19[58], stage2_19[59], stage2_19[60], stage2_19[61], stage2_19[62]},
      {stage2_20[28]},
      {stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage3_23[4],stage3_22[18],stage3_21[18],stage3_20[23],stage3_19[37]}
   );
   gpc615_5 gpc7381 (
      {stage2_19[63], stage2_19[64], stage2_19[65], stage2_19[66], stage2_19[67]},
      {stage2_20[29]},
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58], stage2_21[59]},
      {stage3_23[5],stage3_22[19],stage3_21[19],stage3_20[24],stage3_19[38]}
   );
   gpc615_5 gpc7382 (
      {stage2_19[68], stage2_19[69], stage2_19[70], stage2_19[71], stage2_19[72]},
      {stage2_20[30]},
      {stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63], stage2_21[64], stage2_21[65]},
      {stage3_23[6],stage3_22[20],stage3_21[20],stage3_20[25],stage3_19[39]}
   );
   gpc615_5 gpc7383 (
      {stage2_19[73], stage2_19[74], stage2_19[75], stage2_19[76], stage2_19[77]},
      {stage2_20[31]},
      {stage2_21[66], stage2_21[67], stage2_21[68], stage2_21[69], stage2_21[70], stage2_21[71]},
      {stage3_23[7],stage3_22[21],stage3_21[21],stage3_20[26],stage3_19[40]}
   );
   gpc615_5 gpc7384 (
      {stage2_19[78], stage2_19[79], stage2_19[80], stage2_19[81], stage2_19[82]},
      {stage2_20[32]},
      {stage2_21[72], stage2_21[73], stage2_21[74], stage2_21[75], stage2_21[76], stage2_21[77]},
      {stage3_23[8],stage3_22[22],stage3_21[22],stage3_20[27],stage3_19[41]}
   );
   gpc615_5 gpc7385 (
      {stage2_19[83], stage2_19[84], stage2_19[85], stage2_19[86], stage2_19[87]},
      {stage2_20[33]},
      {stage2_21[78], stage2_21[79], stage2_21[80], stage2_21[81], stage2_21[82], stage2_21[83]},
      {stage3_23[9],stage3_22[23],stage3_21[23],stage3_20[28],stage3_19[42]}
   );
   gpc615_5 gpc7386 (
      {stage2_19[88], stage2_19[89], stage2_19[90], stage2_19[91], stage2_19[92]},
      {stage2_20[34]},
      {stage2_21[84], stage2_21[85], stage2_21[86], stage2_21[87], stage2_21[88], stage2_21[89]},
      {stage3_23[10],stage3_22[24],stage3_21[24],stage3_20[29],stage3_19[43]}
   );
   gpc615_5 gpc7387 (
      {stage2_19[93], stage2_19[94], stage2_19[95], stage2_19[96], stage2_19[97]},
      {stage2_20[35]},
      {stage2_21[90], stage2_21[91], stage2_21[92], stage2_21[93], stage2_21[94], stage2_21[95]},
      {stage3_23[11],stage3_22[25],stage3_21[25],stage3_20[30],stage3_19[44]}
   );
   gpc615_5 gpc7388 (
      {stage2_19[98], stage2_19[99], stage2_19[100], stage2_19[101], stage2_19[102]},
      {stage2_20[36]},
      {stage2_21[96], stage2_21[97], stage2_21[98], stage2_21[99], stage2_21[100], stage2_21[101]},
      {stage3_23[12],stage3_22[26],stage3_21[26],stage3_20[31],stage3_19[45]}
   );
   gpc615_5 gpc7389 (
      {stage2_19[103], stage2_19[104], stage2_19[105], stage2_19[106], stage2_19[107]},
      {stage2_20[37]},
      {stage2_21[102], stage2_21[103], stage2_21[104], stage2_21[105], stage2_21[106], stage2_21[107]},
      {stage3_23[13],stage3_22[27],stage3_21[27],stage3_20[32],stage3_19[46]}
   );
   gpc615_5 gpc7390 (
      {stage2_19[108], stage2_19[109], stage2_19[110], stage2_19[111], stage2_19[112]},
      {stage2_20[38]},
      {stage2_21[108], stage2_21[109], stage2_21[110], stage2_21[111], stage2_21[112], stage2_21[113]},
      {stage3_23[14],stage3_22[28],stage3_21[28],stage3_20[33],stage3_19[47]}
   );
   gpc606_5 gpc7391 (
      {stage2_20[39], stage2_20[40], stage2_20[41], stage2_20[42], stage2_20[43], stage2_20[44]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[15],stage3_22[29],stage3_21[29],stage3_20[34]}
   );
   gpc606_5 gpc7392 (
      {stage2_21[114], stage2_21[115], stage2_21[116], stage2_21[117], stage2_21[118], stage2_21[119]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[16],stage3_22[30],stage3_21[30]}
   );
   gpc606_5 gpc7393 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[1],stage3_24[2],stage3_23[17],stage3_22[31]}
   );
   gpc606_5 gpc7394 (
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[2],stage3_24[3],stage3_23[18],stage3_22[32]}
   );
   gpc606_5 gpc7395 (
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[3],stage3_24[4],stage3_23[19],stage3_22[33]}
   );
   gpc606_5 gpc7396 (
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[4],stage3_24[5],stage3_23[20],stage3_22[34]}
   );
   gpc615_5 gpc7397 (
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34]},
      {stage2_23[6]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[5],stage3_24[6],stage3_23[21],stage3_22[35]}
   );
   gpc615_5 gpc7398 (
      {stage2_22[35], stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39]},
      {stage2_23[7]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[6],stage3_24[7],stage3_23[22],stage3_22[36]}
   );
   gpc615_5 gpc7399 (
      {stage2_22[40], stage2_22[41], stage2_22[42], stage2_22[43], stage2_22[44]},
      {stage2_23[8]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[7],stage3_24[8],stage3_23[23],stage3_22[37]}
   );
   gpc615_5 gpc7400 (
      {stage2_22[45], stage2_22[46], stage2_22[47], stage2_22[48], stage2_22[49]},
      {stage2_23[9]},
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage3_26[7],stage3_25[8],stage3_24[9],stage3_23[24],stage3_22[38]}
   );
   gpc615_5 gpc7401 (
      {stage2_22[50], stage2_22[51], stage2_22[52], stage2_22[53], stage2_22[54]},
      {stage2_23[10]},
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage3_26[8],stage3_25[9],stage3_24[10],stage3_23[25],stage3_22[39]}
   );
   gpc615_5 gpc7402 (
      {stage2_22[55], stage2_22[56], stage2_22[57], stage2_22[58], stage2_22[59]},
      {stage2_23[11]},
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage3_26[9],stage3_25[10],stage3_24[11],stage3_23[26],stage3_22[40]}
   );
   gpc615_5 gpc7403 (
      {stage2_22[60], stage2_22[61], stage2_22[62], stage2_22[63], stage2_22[64]},
      {stage2_23[12]},
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage3_26[10],stage3_25[11],stage3_24[12],stage3_23[27],stage3_22[41]}
   );
   gpc615_5 gpc7404 (
      {stage2_22[65], stage2_22[66], stage2_22[67], stage2_22[68], stage2_22[69]},
      {stage2_23[13]},
      {stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70], stage2_24[71]},
      {stage3_26[11],stage3_25[12],stage3_24[13],stage3_23[28],stage3_22[42]}
   );
   gpc615_5 gpc7405 (
      {stage2_22[70], stage2_22[71], stage2_22[72], stage2_22[73], stage2_22[74]},
      {stage2_23[14]},
      {stage2_24[72], stage2_24[73], stage2_24[74], stage2_24[75], stage2_24[76], stage2_24[77]},
      {stage3_26[12],stage3_25[13],stage3_24[14],stage3_23[29],stage3_22[43]}
   );
   gpc615_5 gpc7406 (
      {stage2_22[75], stage2_22[76], stage2_22[77], stage2_22[78], stage2_22[79]},
      {stage2_23[15]},
      {stage2_24[78], stage2_24[79], stage2_24[80], stage2_24[81], stage2_24[82], stage2_24[83]},
      {stage3_26[13],stage3_25[14],stage3_24[15],stage3_23[30],stage3_22[44]}
   );
   gpc2116_5 gpc7407 (
      {stage2_23[16], stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21]},
      {stage2_24[84]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1]},
      {stage3_27[0],stage3_26[14],stage3_25[15],stage3_24[16],stage3_23[31]}
   );
   gpc615_5 gpc7408 (
      {stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26]},
      {stage2_24[85]},
      {stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6]},
      {stage3_27[1],stage3_26[15],stage3_25[16],stage3_24[17],stage3_23[32]}
   );
   gpc615_5 gpc7409 (
      {stage2_23[27], stage2_23[28], stage2_23[29], stage2_23[30], stage2_23[31]},
      {stage2_24[86]},
      {stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12]},
      {stage3_27[2],stage3_26[16],stage3_25[17],stage3_24[18],stage3_23[33]}
   );
   gpc615_5 gpc7410 (
      {stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35], stage2_23[36]},
      {stage2_24[87]},
      {stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17], stage2_25[18]},
      {stage3_27[3],stage3_26[17],stage3_25[18],stage3_24[19],stage3_23[34]}
   );
   gpc615_5 gpc7411 (
      {stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage2_24[88]},
      {stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23], stage2_25[24]},
      {stage3_27[4],stage3_26[18],stage3_25[19],stage3_24[20],stage3_23[35]}
   );
   gpc615_5 gpc7412 (
      {stage2_23[42], stage2_23[43], stage2_23[44], stage2_23[45], stage2_23[46]},
      {stage2_24[89]},
      {stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29], stage2_25[30]},
      {stage3_27[5],stage3_26[19],stage3_25[20],stage3_24[21],stage3_23[36]}
   );
   gpc615_5 gpc7413 (
      {stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50], stage2_23[51]},
      {stage2_24[90]},
      {stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35], stage2_25[36]},
      {stage3_27[6],stage3_26[20],stage3_25[21],stage3_24[22],stage3_23[37]}
   );
   gpc615_5 gpc7414 (
      {stage2_23[52], stage2_23[53], stage2_23[54], stage2_23[55], stage2_23[56]},
      {stage2_24[91]},
      {stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41], stage2_25[42]},
      {stage3_27[7],stage3_26[21],stage3_25[22],stage3_24[23],stage3_23[38]}
   );
   gpc615_5 gpc7415 (
      {stage2_23[57], stage2_23[58], stage2_23[59], stage2_23[60], stage2_23[61]},
      {stage2_24[92]},
      {stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47], stage2_25[48]},
      {stage3_27[8],stage3_26[22],stage3_25[23],stage3_24[24],stage3_23[39]}
   );
   gpc615_5 gpc7416 (
      {stage2_23[62], stage2_23[63], stage2_23[64], stage2_23[65], stage2_23[66]},
      {stage2_24[93]},
      {stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53], stage2_25[54]},
      {stage3_27[9],stage3_26[23],stage3_25[24],stage3_24[25],stage3_23[40]}
   );
   gpc615_5 gpc7417 (
      {stage2_23[67], stage2_23[68], stage2_23[69], stage2_23[70], stage2_23[71]},
      {stage2_24[94]},
      {stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59], stage2_25[60]},
      {stage3_27[10],stage3_26[24],stage3_25[25],stage3_24[26],stage3_23[41]}
   );
   gpc615_5 gpc7418 (
      {stage2_23[72], stage2_23[73], stage2_23[74], stage2_23[75], 1'b0},
      {stage2_24[95]},
      {stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65], stage2_25[66]},
      {stage3_27[11],stage3_26[25],stage3_25[26],stage3_24[27],stage3_23[42]}
   );
   gpc606_5 gpc7419 (
      {stage2_24[96], stage2_24[97], stage2_24[98], stage2_24[99], stage2_24[100], stage2_24[101]},
      {stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6], stage2_26[7]},
      {stage3_28[0],stage3_27[12],stage3_26[26],stage3_25[27],stage3_24[28]}
   );
   gpc606_5 gpc7420 (
      {stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71], stage2_25[72]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[1],stage3_27[13],stage3_26[27],stage3_25[28]}
   );
   gpc606_5 gpc7421 (
      {stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77], stage2_25[78]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[2],stage3_27[14],stage3_26[28],stage3_25[29]}
   );
   gpc606_5 gpc7422 (
      {stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83], stage2_25[84]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[3],stage3_27[15],stage3_26[29],stage3_25[30]}
   );
   gpc606_5 gpc7423 (
      {stage2_25[85], stage2_25[86], stage2_25[87], stage2_25[88], stage2_25[89], stage2_25[90]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[4],stage3_27[16],stage3_26[30],stage3_25[31]}
   );
   gpc606_5 gpc7424 (
      {stage2_25[91], stage2_25[92], stage2_25[93], stage2_25[94], stage2_25[95], 1'b0},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[5],stage3_27[17],stage3_26[31],stage3_25[32]}
   );
   gpc135_4 gpc7425 (
      {stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12]},
      {stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_28[0]},
      {stage3_29[5],stage3_28[6],stage3_27[18],stage3_26[32]}
   );
   gpc135_4 gpc7426 (
      {stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage2_27[33], stage2_27[34], stage2_27[35]},
      {stage2_28[1]},
      {stage3_29[6],stage3_28[7],stage3_27[19],stage3_26[33]}
   );
   gpc135_4 gpc7427 (
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22]},
      {stage2_27[36], stage2_27[37], stage2_27[38]},
      {stage2_28[2]},
      {stage3_29[7],stage3_28[8],stage3_27[20],stage3_26[34]}
   );
   gpc135_4 gpc7428 (
      {stage2_26[23], stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27]},
      {stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage2_28[3]},
      {stage3_29[8],stage3_28[9],stage3_27[21],stage3_26[35]}
   );
   gpc135_4 gpc7429 (
      {stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31], stage2_26[32]},
      {stage2_27[42], stage2_27[43], stage2_27[44]},
      {stage2_28[4]},
      {stage3_29[9],stage3_28[10],stage3_27[22],stage3_26[36]}
   );
   gpc135_4 gpc7430 (
      {stage2_26[33], stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37]},
      {stage2_27[45], stage2_27[46], stage2_27[47]},
      {stage2_28[5]},
      {stage3_29[10],stage3_28[11],stage3_27[23],stage3_26[37]}
   );
   gpc135_4 gpc7431 (
      {stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42]},
      {stage2_27[48], stage2_27[49], stage2_27[50]},
      {stage2_28[6]},
      {stage3_29[11],stage3_28[12],stage3_27[24],stage3_26[38]}
   );
   gpc135_4 gpc7432 (
      {stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47]},
      {stage2_27[51], stage2_27[52], stage2_27[53]},
      {stage2_28[7]},
      {stage3_29[12],stage3_28[13],stage3_27[25],stage3_26[39]}
   );
   gpc135_4 gpc7433 (
      {stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52]},
      {stage2_27[54], stage2_27[55], stage2_27[56]},
      {stage2_28[8]},
      {stage3_29[13],stage3_28[14],stage3_27[26],stage3_26[40]}
   );
   gpc135_4 gpc7434 (
      {stage2_26[53], stage2_26[54], stage2_26[55], stage2_26[56], stage2_26[57]},
      {stage2_27[57], stage2_27[58], stage2_27[59]},
      {stage2_28[9]},
      {stage3_29[14],stage3_28[15],stage3_27[27],stage3_26[41]}
   );
   gpc135_4 gpc7435 (
      {stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_27[60], stage2_27[61], stage2_27[62]},
      {stage2_28[10]},
      {stage3_29[15],stage3_28[16],stage3_27[28],stage3_26[42]}
   );
   gpc135_4 gpc7436 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67]},
      {stage2_27[63], stage2_27[64], stage2_27[65]},
      {stage2_28[11]},
      {stage3_29[16],stage3_28[17],stage3_27[29],stage3_26[43]}
   );
   gpc135_4 gpc7437 (
      {stage2_26[68], stage2_26[69], stage2_26[70], stage2_26[71], stage2_26[72]},
      {stage2_27[66], stage2_27[67], stage2_27[68]},
      {stage2_28[12]},
      {stage3_29[17],stage3_28[18],stage3_27[30],stage3_26[44]}
   );
   gpc1343_5 gpc7438 (
      {stage2_26[73], stage2_26[74], stage2_26[75]},
      {stage2_27[69], stage2_27[70], stage2_27[71], stage2_27[72]},
      {stage2_28[13], stage2_28[14], stage2_28[15]},
      {stage2_29[0]},
      {stage3_30[0],stage3_29[18],stage3_28[19],stage3_27[31],stage3_26[45]}
   );
   gpc117_4 gpc7439 (
      {stage2_26[76], stage2_26[77], stage2_26[78], stage2_26[79], stage2_26[80], stage2_26[81], stage2_26[82]},
      {stage2_27[73]},
      {stage2_28[16]},
      {stage3_29[19],stage3_28[20],stage3_27[32],stage3_26[46]}
   );
   gpc7_3 gpc7440 (
      {stage2_27[74], stage2_27[75], stage2_27[76], stage2_27[77], stage2_27[78], stage2_27[79], stage2_27[80]},
      {stage3_29[20],stage3_28[21],stage3_27[33]}
   );
   gpc7_3 gpc7441 (
      {stage2_27[81], stage2_27[82], stage2_27[83], stage2_27[84], stage2_27[85], stage2_27[86], stage2_27[87]},
      {stage3_29[21],stage3_28[22],stage3_27[34]}
   );
   gpc615_5 gpc7442 (
      {stage2_27[88], stage2_27[89], stage2_27[90], stage2_27[91], stage2_27[92]},
      {stage2_28[17]},
      {stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5], stage2_29[6]},
      {stage3_31[0],stage3_30[1],stage3_29[22],stage3_28[23],stage3_27[35]}
   );
   gpc606_5 gpc7443 (
      {stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[1],stage3_30[2],stage3_29[23],stage3_28[24]}
   );
   gpc615_5 gpc7444 (
      {stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_29[7]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[2],stage3_30[3],stage3_29[24],stage3_28[25]}
   );
   gpc615_5 gpc7445 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33]},
      {stage2_29[8]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[3],stage3_30[4],stage3_29[25],stage3_28[26]}
   );
   gpc615_5 gpc7446 (
      {stage2_28[34], stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38]},
      {stage2_29[9]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[4],stage3_30[5],stage3_29[26],stage3_28[27]}
   );
   gpc615_5 gpc7447 (
      {stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42], stage2_28[43]},
      {stage2_29[10]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[5],stage3_30[6],stage3_29[27],stage3_28[28]}
   );
   gpc615_5 gpc7448 (
      {stage2_28[44], stage2_28[45], stage2_28[46], stage2_28[47], stage2_28[48]},
      {stage2_29[11]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[6],stage3_30[7],stage3_29[28],stage3_28[29]}
   );
   gpc615_5 gpc7449 (
      {stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52], stage2_28[53]},
      {stage2_29[12]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[7],stage3_30[8],stage3_29[29],stage3_28[30]}
   );
   gpc615_5 gpc7450 (
      {stage2_28[54], stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58]},
      {stage2_29[13]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage3_32[7],stage3_31[8],stage3_30[9],stage3_29[30],stage3_28[31]}
   );
   gpc615_5 gpc7451 (
      {stage2_28[59], stage2_28[60], stage2_28[61], stage2_28[62], stage2_28[63]},
      {stage2_29[14]},
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage3_32[8],stage3_31[9],stage3_30[10],stage3_29[31],stage3_28[32]}
   );
   gpc615_5 gpc7452 (
      {stage2_28[64], stage2_28[65], stage2_28[66], stage2_28[67], stage2_28[68]},
      {stage2_29[15]},
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage3_32[9],stage3_31[10],stage3_30[11],stage3_29[32],stage3_28[33]}
   );
   gpc1163_5 gpc7453 (
      {stage2_29[16], stage2_29[17], stage2_29[18]},
      {stage2_30[60], stage2_30[61], stage2_30[62], stage2_30[63], stage2_30[64], stage2_30[65]},
      {stage2_31[0]},
      {stage2_32[0]},
      {stage3_33[0],stage3_32[10],stage3_31[11],stage3_30[12],stage3_29[33]}
   );
   gpc1163_5 gpc7454 (
      {stage2_29[19], stage2_29[20], stage2_29[21]},
      {stage2_30[66], stage2_30[67], stage2_30[68], stage2_30[69], stage2_30[70], stage2_30[71]},
      {stage2_31[1]},
      {stage2_32[1]},
      {stage3_33[1],stage3_32[11],stage3_31[12],stage3_30[13],stage3_29[34]}
   );
   gpc1163_5 gpc7455 (
      {stage2_29[22], stage2_29[23], stage2_29[24]},
      {stage2_30[72], stage2_30[73], stage2_30[74], stage2_30[75], stage2_30[76], stage2_30[77]},
      {stage2_31[2]},
      {stage2_32[2]},
      {stage3_33[2],stage3_32[12],stage3_31[13],stage3_30[14],stage3_29[35]}
   );
   gpc1163_5 gpc7456 (
      {stage2_29[25], stage2_29[26], stage2_29[27]},
      {stage2_30[78], stage2_30[79], stage2_30[80], stage2_30[81], stage2_30[82], stage2_30[83]},
      {stage2_31[3]},
      {stage2_32[3]},
      {stage3_33[3],stage3_32[13],stage3_31[14],stage3_30[15],stage3_29[36]}
   );
   gpc1163_5 gpc7457 (
      {stage2_29[28], stage2_29[29], stage2_29[30]},
      {stage2_30[84], stage2_30[85], stage2_30[86], stage2_30[87], stage2_30[88], stage2_30[89]},
      {stage2_31[4]},
      {stage2_32[4]},
      {stage3_33[4],stage3_32[14],stage3_31[15],stage3_30[16],stage3_29[37]}
   );
   gpc1163_5 gpc7458 (
      {stage2_29[31], stage2_29[32], stage2_29[33]},
      {stage2_30[90], stage2_30[91], stage2_30[92], stage2_30[93], stage2_30[94], stage2_30[95]},
      {stage2_31[5]},
      {stage2_32[5]},
      {stage3_33[5],stage3_32[15],stage3_31[16],stage3_30[17],stage3_29[38]}
   );
   gpc606_5 gpc7459 (
      {stage2_29[34], stage2_29[35], stage2_29[36], stage2_29[37], stage2_29[38], stage2_29[39]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[6],stage3_32[16],stage3_31[17],stage3_30[18],stage3_29[39]}
   );
   gpc606_5 gpc7460 (
      {stage2_29[40], stage2_29[41], stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[7],stage3_32[17],stage3_31[18],stage3_30[19],stage3_29[40]}
   );
   gpc606_5 gpc7461 (
      {stage2_29[46], stage2_29[47], stage2_29[48], stage2_29[49], stage2_29[50], stage2_29[51]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[8],stage3_32[18],stage3_31[19],stage3_30[20],stage3_29[41]}
   );
   gpc606_5 gpc7462 (
      {stage2_29[52], stage2_29[53], stage2_29[54], stage2_29[55], stage2_29[56], stage2_29[57]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[9],stage3_32[19],stage3_31[20],stage3_30[21],stage3_29[42]}
   );
   gpc606_5 gpc7463 (
      {stage2_29[58], stage2_29[59], stage2_29[60], stage2_29[61], stage2_29[62], stage2_29[63]},
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34], stage2_31[35]},
      {stage3_33[10],stage3_32[20],stage3_31[21],stage3_30[22],stage3_29[43]}
   );
   gpc606_5 gpc7464 (
      {stage2_29[64], stage2_29[65], stage2_29[66], stage2_29[67], stage2_29[68], stage2_29[69]},
      {stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40], stage2_31[41]},
      {stage3_33[11],stage3_32[21],stage3_31[22],stage3_30[23],stage3_29[44]}
   );
   gpc606_5 gpc7465 (
      {stage2_29[70], stage2_29[71], stage2_29[72], stage2_29[73], stage2_29[74], stage2_29[75]},
      {stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46], stage2_31[47]},
      {stage3_33[12],stage3_32[22],stage3_31[23],stage3_30[24],stage3_29[45]}
   );
   gpc606_5 gpc7466 (
      {stage2_29[76], stage2_29[77], stage2_29[78], stage2_29[79], stage2_29[80], stage2_29[81]},
      {stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52], stage2_31[53]},
      {stage3_33[13],stage3_32[23],stage3_31[24],stage3_30[25],stage3_29[46]}
   );
   gpc606_5 gpc7467 (
      {stage2_29[82], stage2_29[83], stage2_29[84], stage2_29[85], stage2_29[86], 1'b0},
      {stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57], stage2_31[58], stage2_31[59]},
      {stage3_33[14],stage3_32[24],stage3_31[25],stage3_30[26],stage3_29[47]}
   );
   gpc207_4 gpc7468 (
      {stage2_30[96], stage2_30[97], stage2_30[98], stage2_30[99], stage2_30[100], stage2_30[101], stage2_30[102]},
      {stage2_32[6], stage2_32[7]},
      {stage3_33[15],stage3_32[25],stage3_31[26],stage3_30[27]}
   );
   gpc615_5 gpc7469 (
      {stage2_31[60], stage2_31[61], stage2_31[62], stage2_31[63], stage2_31[64]},
      {stage2_32[8]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[0],stage3_33[16],stage3_32[26],stage3_31[27]}
   );
   gpc615_5 gpc7470 (
      {stage2_31[65], stage2_31[66], stage2_31[67], stage2_31[68], stage2_31[69]},
      {stage2_32[9]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[1],stage3_33[17],stage3_32[27],stage3_31[28]}
   );
   gpc615_5 gpc7471 (
      {stage2_31[70], stage2_31[71], stage2_31[72], stage2_31[73], stage2_31[74]},
      {stage2_32[10]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[2],stage3_33[18],stage3_32[28],stage3_31[29]}
   );
   gpc615_5 gpc7472 (
      {stage2_31[75], stage2_31[76], stage2_31[77], stage2_31[78], stage2_31[79]},
      {stage2_32[11]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[3],stage3_33[19],stage3_32[29],stage3_31[30]}
   );
   gpc615_5 gpc7473 (
      {stage2_31[80], stage2_31[81], stage2_31[82], stage2_31[83], stage2_31[84]},
      {stage2_32[12]},
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage3_35[4],stage3_34[4],stage3_33[20],stage3_32[30],stage3_31[31]}
   );
   gpc615_5 gpc7474 (
      {stage2_31[85], stage2_31[86], stage2_31[87], stage2_31[88], stage2_31[89]},
      {stage2_32[13]},
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage3_35[5],stage3_34[5],stage3_33[21],stage3_32[31],stage3_31[32]}
   );
   gpc615_5 gpc7475 (
      {stage2_31[90], stage2_31[91], stage2_31[92], stage2_31[93], stage2_31[94]},
      {stage2_32[14]},
      {stage2_33[36], stage2_33[37], stage2_33[38], stage2_33[39], stage2_33[40], stage2_33[41]},
      {stage3_35[6],stage3_34[6],stage3_33[22],stage3_32[32],stage3_31[33]}
   );
   gpc606_5 gpc7476 (
      {stage2_32[15], stage2_32[16], stage2_32[17], stage2_32[18], stage2_32[19], stage2_32[20]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[7],stage3_34[7],stage3_33[23],stage3_32[33]}
   );
   gpc606_5 gpc7477 (
      {stage2_32[21], stage2_32[22], stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[8],stage3_34[8],stage3_33[24],stage3_32[34]}
   );
   gpc606_5 gpc7478 (
      {stage2_32[27], stage2_32[28], stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[9],stage3_34[9],stage3_33[25],stage3_32[35]}
   );
   gpc606_5 gpc7479 (
      {stage2_32[33], stage2_32[34], stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38]},
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage3_36[3],stage3_35[10],stage3_34[10],stage3_33[26],stage3_32[36]}
   );
   gpc606_5 gpc7480 (
      {stage2_32[39], stage2_32[40], stage2_32[41], stage2_32[42], stage2_32[43], stage2_32[44]},
      {stage2_34[24], stage2_34[25], stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29]},
      {stage3_36[4],stage3_35[11],stage3_34[11],stage3_33[27],stage3_32[37]}
   );
   gpc606_5 gpc7481 (
      {stage2_32[45], stage2_32[46], stage2_32[47], stage2_32[48], stage2_32[49], stage2_32[50]},
      {stage2_34[30], stage2_34[31], stage2_34[32], stage2_34[33], stage2_34[34], stage2_34[35]},
      {stage3_36[5],stage3_35[12],stage3_34[12],stage3_33[28],stage3_32[38]}
   );
   gpc606_5 gpc7482 (
      {stage2_32[51], stage2_32[52], stage2_32[53], stage2_32[54], stage2_32[55], stage2_32[56]},
      {stage2_34[36], stage2_34[37], stage2_34[38], stage2_34[39], stage2_34[40], stage2_34[41]},
      {stage3_36[6],stage3_35[13],stage3_34[13],stage3_33[29],stage3_32[39]}
   );
   gpc606_5 gpc7483 (
      {stage2_32[57], stage2_32[58], stage2_32[59], stage2_32[60], stage2_32[61], stage2_32[62]},
      {stage2_34[42], stage2_34[43], stage2_34[44], stage2_34[45], stage2_34[46], stage2_34[47]},
      {stage3_36[7],stage3_35[14],stage3_34[14],stage3_33[30],stage3_32[40]}
   );
   gpc606_5 gpc7484 (
      {stage2_32[63], stage2_32[64], stage2_32[65], stage2_32[66], stage2_32[67], stage2_32[68]},
      {stage2_34[48], stage2_34[49], stage2_34[50], stage2_34[51], stage2_34[52], stage2_34[53]},
      {stage3_36[8],stage3_35[15],stage3_34[15],stage3_33[31],stage3_32[41]}
   );
   gpc606_5 gpc7485 (
      {stage2_32[69], stage2_32[70], stage2_32[71], stage2_32[72], stage2_32[73], stage2_32[74]},
      {stage2_34[54], stage2_34[55], stage2_34[56], stage2_34[57], stage2_34[58], stage2_34[59]},
      {stage3_36[9],stage3_35[16],stage3_34[16],stage3_33[32],stage3_32[42]}
   );
   gpc606_5 gpc7486 (
      {stage2_32[75], stage2_32[76], stage2_32[77], stage2_32[78], stage2_32[79], stage2_32[80]},
      {stage2_34[60], stage2_34[61], stage2_34[62], stage2_34[63], stage2_34[64], stage2_34[65]},
      {stage3_36[10],stage3_35[17],stage3_34[17],stage3_33[33],stage3_32[43]}
   );
   gpc606_5 gpc7487 (
      {stage2_32[81], stage2_32[82], stage2_32[83], stage2_32[84], stage2_32[85], stage2_32[86]},
      {stage2_34[66], stage2_34[67], stage2_34[68], stage2_34[69], stage2_34[70], stage2_34[71]},
      {stage3_36[11],stage3_35[18],stage3_34[18],stage3_33[34],stage3_32[44]}
   );
   gpc606_5 gpc7488 (
      {stage2_32[87], stage2_32[88], stage2_32[89], stage2_32[90], stage2_32[91], stage2_32[92]},
      {stage2_34[72], stage2_34[73], stage2_34[74], stage2_34[75], stage2_34[76], stage2_34[77]},
      {stage3_36[12],stage3_35[19],stage3_34[19],stage3_33[35],stage3_32[45]}
   );
   gpc606_5 gpc7489 (
      {stage2_32[93], stage2_32[94], stage2_32[95], stage2_32[96], stage2_32[97], stage2_32[98]},
      {stage2_34[78], stage2_34[79], stage2_34[80], stage2_34[81], stage2_34[82], stage2_34[83]},
      {stage3_36[13],stage3_35[20],stage3_34[20],stage3_33[36],stage3_32[46]}
   );
   gpc606_5 gpc7490 (
      {stage2_33[42], stage2_33[43], stage2_33[44], stage2_33[45], stage2_33[46], stage2_33[47]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[14],stage3_35[21],stage3_34[21],stage3_33[37]}
   );
   gpc606_5 gpc7491 (
      {stage2_33[48], stage2_33[49], stage2_33[50], stage2_33[51], stage2_33[52], stage2_33[53]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[15],stage3_35[22],stage3_34[22],stage3_33[38]}
   );
   gpc606_5 gpc7492 (
      {stage2_33[54], stage2_33[55], stage2_33[56], stage2_33[57], stage2_33[58], stage2_33[59]},
      {stage2_35[12], stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16], stage2_35[17]},
      {stage3_37[2],stage3_36[16],stage3_35[23],stage3_34[23],stage3_33[39]}
   );
   gpc606_5 gpc7493 (
      {stage2_33[60], stage2_33[61], stage2_33[62], stage2_33[63], stage2_33[64], stage2_33[65]},
      {stage2_35[18], stage2_35[19], stage2_35[20], stage2_35[21], stage2_35[22], stage2_35[23]},
      {stage3_37[3],stage3_36[17],stage3_35[24],stage3_34[24],stage3_33[40]}
   );
   gpc606_5 gpc7494 (
      {stage2_33[66], stage2_33[67], stage2_33[68], stage2_33[69], stage2_33[70], stage2_33[71]},
      {stage2_35[24], stage2_35[25], stage2_35[26], stage2_35[27], stage2_35[28], stage2_35[29]},
      {stage3_37[4],stage3_36[18],stage3_35[25],stage3_34[25],stage3_33[41]}
   );
   gpc1163_5 gpc7495 (
      {stage2_34[84], stage2_34[85], stage2_34[86]},
      {stage2_35[30], stage2_35[31], stage2_35[32], stage2_35[33], stage2_35[34], stage2_35[35]},
      {stage2_36[0]},
      {stage2_37[0]},
      {stage3_38[0],stage3_37[5],stage3_36[19],stage3_35[26],stage3_34[26]}
   );
   gpc1163_5 gpc7496 (
      {stage2_34[87], stage2_34[88], stage2_34[89]},
      {stage2_35[36], stage2_35[37], stage2_35[38], stage2_35[39], stage2_35[40], stage2_35[41]},
      {stage2_36[1]},
      {stage2_37[1]},
      {stage3_38[1],stage3_37[6],stage3_36[20],stage3_35[27],stage3_34[27]}
   );
   gpc1163_5 gpc7497 (
      {stage2_34[90], stage2_34[91], stage2_34[92]},
      {stage2_35[42], stage2_35[43], stage2_35[44], stage2_35[45], stage2_35[46], stage2_35[47]},
      {stage2_36[2]},
      {stage2_37[2]},
      {stage3_38[2],stage3_37[7],stage3_36[21],stage3_35[28],stage3_34[28]}
   );
   gpc1163_5 gpc7498 (
      {stage2_34[93], stage2_34[94], stage2_34[95]},
      {stage2_35[48], stage2_35[49], stage2_35[50], stage2_35[51], stage2_35[52], stage2_35[53]},
      {stage2_36[3]},
      {stage2_37[3]},
      {stage3_38[3],stage3_37[8],stage3_36[22],stage3_35[29],stage3_34[29]}
   );
   gpc1163_5 gpc7499 (
      {stage2_34[96], stage2_34[97], stage2_34[98]},
      {stage2_35[54], stage2_35[55], stage2_35[56], stage2_35[57], stage2_35[58], stage2_35[59]},
      {stage2_36[4]},
      {stage2_37[4]},
      {stage3_38[4],stage3_37[9],stage3_36[23],stage3_35[30],stage3_34[30]}
   );
   gpc1163_5 gpc7500 (
      {stage2_34[99], stage2_34[100], stage2_34[101]},
      {stage2_35[60], stage2_35[61], stage2_35[62], stage2_35[63], stage2_35[64], stage2_35[65]},
      {stage2_36[5]},
      {stage2_37[5]},
      {stage3_38[5],stage3_37[10],stage3_36[24],stage3_35[31],stage3_34[31]}
   );
   gpc1163_5 gpc7501 (
      {stage2_34[102], stage2_34[103], stage2_34[104]},
      {stage2_35[66], stage2_35[67], stage2_35[68], stage2_35[69], stage2_35[70], stage2_35[71]},
      {stage2_36[6]},
      {stage2_37[6]},
      {stage3_38[6],stage3_37[11],stage3_36[25],stage3_35[32],stage3_34[32]}
   );
   gpc1163_5 gpc7502 (
      {stage2_34[105], stage2_34[106], stage2_34[107]},
      {stage2_35[72], stage2_35[73], stage2_35[74], stage2_35[75], stage2_35[76], stage2_35[77]},
      {stage2_36[7]},
      {stage2_37[7]},
      {stage3_38[7],stage3_37[12],stage3_36[26],stage3_35[33],stage3_34[33]}
   );
   gpc1163_5 gpc7503 (
      {stage2_34[108], stage2_34[109], stage2_34[110]},
      {stage2_35[78], stage2_35[79], stage2_35[80], stage2_35[81], stage2_35[82], stage2_35[83]},
      {stage2_36[8]},
      {stage2_37[8]},
      {stage3_38[8],stage3_37[13],stage3_36[27],stage3_35[34],stage3_34[34]}
   );
   gpc1163_5 gpc7504 (
      {stage2_34[111], stage2_34[112], stage2_34[113]},
      {stage2_35[84], stage2_35[85], stage2_35[86], stage2_35[87], stage2_35[88], stage2_35[89]},
      {stage2_36[9]},
      {stage2_37[9]},
      {stage3_38[9],stage3_37[14],stage3_36[28],stage3_35[35],stage3_34[35]}
   );
   gpc615_5 gpc7505 (
      {stage2_34[114], stage2_34[115], stage2_34[116], stage2_34[117], stage2_34[118]},
      {stage2_35[90]},
      {stage2_36[10], stage2_36[11], stage2_36[12], stage2_36[13], stage2_36[14], stage2_36[15]},
      {stage3_38[10],stage3_37[15],stage3_36[29],stage3_35[36],stage3_34[36]}
   );
   gpc615_5 gpc7506 (
      {stage2_34[119], stage2_34[120], stage2_34[121], stage2_34[122], stage2_34[123]},
      {stage2_35[91]},
      {stage2_36[16], stage2_36[17], stage2_36[18], stage2_36[19], stage2_36[20], stage2_36[21]},
      {stage3_38[11],stage3_37[16],stage3_36[30],stage3_35[37],stage3_34[37]}
   );
   gpc615_5 gpc7507 (
      {stage2_34[124], stage2_34[125], stage2_34[126], stage2_34[127], stage2_34[128]},
      {stage2_35[92]},
      {stage2_36[22], stage2_36[23], stage2_36[24], stage2_36[25], stage2_36[26], stage2_36[27]},
      {stage3_38[12],stage3_37[17],stage3_36[31],stage3_35[38],stage3_34[38]}
   );
   gpc1406_5 gpc7508 (
      {stage2_35[93], stage2_35[94], stage2_35[95], stage2_35[96], stage2_35[97], stage2_35[98]},
      {stage2_37[10], stage2_37[11], stage2_37[12], stage2_37[13]},
      {stage2_38[0]},
      {stage3_39[0],stage3_38[13],stage3_37[18],stage3_36[32],stage3_35[39]}
   );
   gpc1406_5 gpc7509 (
      {stage2_35[99], stage2_35[100], stage2_35[101], stage2_35[102], stage2_35[103], stage2_35[104]},
      {stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage2_38[1]},
      {stage3_39[1],stage3_38[14],stage3_37[19],stage3_36[33],stage3_35[40]}
   );
   gpc615_5 gpc7510 (
      {stage2_35[105], stage2_35[106], stage2_35[107], stage2_35[108], stage2_35[109]},
      {stage2_36[28]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[2],stage3_38[15],stage3_37[20],stage3_36[34],stage3_35[41]}
   );
   gpc615_5 gpc7511 (
      {stage2_35[110], stage2_35[111], stage2_35[112], stage2_35[113], stage2_35[114]},
      {stage2_36[29]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[3],stage3_38[16],stage3_37[21],stage3_36[35],stage3_35[42]}
   );
   gpc615_5 gpc7512 (
      {stage2_35[115], stage2_35[116], stage2_35[117], stage2_35[118], stage2_35[119]},
      {stage2_36[30]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[4],stage3_38[17],stage3_37[22],stage3_36[36],stage3_35[43]}
   );
   gpc606_5 gpc7513 (
      {stage2_36[31], stage2_36[32], stage2_36[33], stage2_36[34], stage2_36[35], stage2_36[36]},
      {stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5], stage2_38[6], stage2_38[7]},
      {stage3_40[0],stage3_39[5],stage3_38[18],stage3_37[23],stage3_36[37]}
   );
   gpc606_5 gpc7514 (
      {stage2_36[37], stage2_36[38], stage2_36[39], stage2_36[40], stage2_36[41], stage2_36[42]},
      {stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11], stage2_38[12], stage2_38[13]},
      {stage3_40[1],stage3_39[6],stage3_38[19],stage3_37[24],stage3_36[38]}
   );
   gpc606_5 gpc7515 (
      {stage2_36[43], stage2_36[44], stage2_36[45], stage2_36[46], stage2_36[47], stage2_36[48]},
      {stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17], stage2_38[18], stage2_38[19]},
      {stage3_40[2],stage3_39[7],stage3_38[20],stage3_37[25],stage3_36[39]}
   );
   gpc606_5 gpc7516 (
      {stage2_36[49], stage2_36[50], stage2_36[51], stage2_36[52], stage2_36[53], stage2_36[54]},
      {stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23], stage2_38[24], stage2_38[25]},
      {stage3_40[3],stage3_39[8],stage3_38[21],stage3_37[26],stage3_36[40]}
   );
   gpc606_5 gpc7517 (
      {stage2_36[55], stage2_36[56], stage2_36[57], stage2_36[58], stage2_36[59], stage2_36[60]},
      {stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29], stage2_38[30], stage2_38[31]},
      {stage3_40[4],stage3_39[9],stage3_38[22],stage3_37[27],stage3_36[41]}
   );
   gpc606_5 gpc7518 (
      {stage2_36[61], stage2_36[62], stage2_36[63], stage2_36[64], stage2_36[65], stage2_36[66]},
      {stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35], stage2_38[36], stage2_38[37]},
      {stage3_40[5],stage3_39[10],stage3_38[23],stage3_37[28],stage3_36[42]}
   );
   gpc606_5 gpc7519 (
      {stage2_36[67], stage2_36[68], stage2_36[69], stage2_36[70], stage2_36[71], stage2_36[72]},
      {stage2_38[38], stage2_38[39], stage2_38[40], stage2_38[41], stage2_38[42], stage2_38[43]},
      {stage3_40[6],stage3_39[11],stage3_38[24],stage3_37[29],stage3_36[43]}
   );
   gpc606_5 gpc7520 (
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[7],stage3_39[12],stage3_38[25],stage3_37[30]}
   );
   gpc606_5 gpc7521 (
      {stage2_37[42], stage2_37[43], stage2_37[44], stage2_37[45], stage2_37[46], stage2_37[47]},
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage3_41[1],stage3_40[8],stage3_39[13],stage3_38[26],stage3_37[31]}
   );
   gpc606_5 gpc7522 (
      {stage2_37[48], stage2_37[49], stage2_37[50], stage2_37[51], stage2_37[52], stage2_37[53]},
      {stage2_39[12], stage2_39[13], stage2_39[14], stage2_39[15], stage2_39[16], stage2_39[17]},
      {stage3_41[2],stage3_40[9],stage3_39[14],stage3_38[27],stage3_37[32]}
   );
   gpc615_5 gpc7523 (
      {stage2_37[54], stage2_37[55], stage2_37[56], stage2_37[57], stage2_37[58]},
      {stage2_38[44]},
      {stage2_39[18], stage2_39[19], stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23]},
      {stage3_41[3],stage3_40[10],stage3_39[15],stage3_38[28],stage3_37[33]}
   );
   gpc615_5 gpc7524 (
      {stage2_37[59], stage2_37[60], stage2_37[61], stage2_37[62], stage2_37[63]},
      {stage2_38[45]},
      {stage2_39[24], stage2_39[25], stage2_39[26], stage2_39[27], stage2_39[28], stage2_39[29]},
      {stage3_41[4],stage3_40[11],stage3_39[16],stage3_38[29],stage3_37[34]}
   );
   gpc615_5 gpc7525 (
      {stage2_37[64], stage2_37[65], stage2_37[66], stage2_37[67], stage2_37[68]},
      {stage2_38[46]},
      {stage2_39[30], stage2_39[31], stage2_39[32], stage2_39[33], stage2_39[34], stage2_39[35]},
      {stage3_41[5],stage3_40[12],stage3_39[17],stage3_38[30],stage3_37[35]}
   );
   gpc615_5 gpc7526 (
      {stage2_37[69], stage2_37[70], stage2_37[71], stage2_37[72], stage2_37[73]},
      {stage2_38[47]},
      {stage2_39[36], stage2_39[37], stage2_39[38], stage2_39[39], stage2_39[40], stage2_39[41]},
      {stage3_41[6],stage3_40[13],stage3_39[18],stage3_38[31],stage3_37[36]}
   );
   gpc606_5 gpc7527 (
      {stage2_38[48], stage2_38[49], stage2_38[50], stage2_38[51], stage2_38[52], stage2_38[53]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[7],stage3_40[14],stage3_39[19],stage3_38[32]}
   );
   gpc606_5 gpc7528 (
      {stage2_38[54], stage2_38[55], stage2_38[56], stage2_38[57], stage2_38[58], stage2_38[59]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[8],stage3_40[15],stage3_39[20],stage3_38[33]}
   );
   gpc606_5 gpc7529 (
      {stage2_38[60], stage2_38[61], stage2_38[62], stage2_38[63], stage2_38[64], stage2_38[65]},
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage3_42[2],stage3_41[9],stage3_40[16],stage3_39[21],stage3_38[34]}
   );
   gpc606_5 gpc7530 (
      {stage2_38[66], stage2_38[67], stage2_38[68], stage2_38[69], stage2_38[70], stage2_38[71]},
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage3_42[3],stage3_41[10],stage3_40[17],stage3_39[22],stage3_38[35]}
   );
   gpc606_5 gpc7531 (
      {stage2_38[72], stage2_38[73], stage2_38[74], stage2_38[75], stage2_38[76], stage2_38[77]},
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage3_42[4],stage3_41[11],stage3_40[18],stage3_39[23],stage3_38[36]}
   );
   gpc606_5 gpc7532 (
      {stage2_38[78], stage2_38[79], stage2_38[80], stage2_38[81], stage2_38[82], stage2_38[83]},
      {stage2_40[30], stage2_40[31], stage2_40[32], stage2_40[33], stage2_40[34], stage2_40[35]},
      {stage3_42[5],stage3_41[12],stage3_40[19],stage3_39[24],stage3_38[37]}
   );
   gpc606_5 gpc7533 (
      {stage2_38[84], stage2_38[85], stage2_38[86], stage2_38[87], stage2_38[88], stage2_38[89]},
      {stage2_40[36], stage2_40[37], stage2_40[38], stage2_40[39], stage2_40[40], stage2_40[41]},
      {stage3_42[6],stage3_41[13],stage3_40[20],stage3_39[25],stage3_38[38]}
   );
   gpc606_5 gpc7534 (
      {stage2_38[90], stage2_38[91], stage2_38[92], stage2_38[93], stage2_38[94], stage2_38[95]},
      {stage2_40[42], stage2_40[43], stage2_40[44], stage2_40[45], stage2_40[46], stage2_40[47]},
      {stage3_42[7],stage3_41[14],stage3_40[21],stage3_39[26],stage3_38[39]}
   );
   gpc606_5 gpc7535 (
      {stage2_38[96], stage2_38[97], stage2_38[98], stage2_38[99], stage2_38[100], stage2_38[101]},
      {stage2_40[48], stage2_40[49], stage2_40[50], stage2_40[51], stage2_40[52], stage2_40[53]},
      {stage3_42[8],stage3_41[15],stage3_40[22],stage3_39[27],stage3_38[40]}
   );
   gpc606_5 gpc7536 (
      {stage2_38[102], stage2_38[103], stage2_38[104], stage2_38[105], stage2_38[106], stage2_38[107]},
      {stage2_40[54], stage2_40[55], stage2_40[56], stage2_40[57], stage2_40[58], stage2_40[59]},
      {stage3_42[9],stage3_41[16],stage3_40[23],stage3_39[28],stage3_38[41]}
   );
   gpc606_5 gpc7537 (
      {stage2_38[108], stage2_38[109], stage2_38[110], stage2_38[111], stage2_38[112], stage2_38[113]},
      {stage2_40[60], stage2_40[61], stage2_40[62], stage2_40[63], stage2_40[64], stage2_40[65]},
      {stage3_42[10],stage3_41[17],stage3_40[24],stage3_39[29],stage3_38[42]}
   );
   gpc606_5 gpc7538 (
      {stage2_38[114], stage2_38[115], stage2_38[116], stage2_38[117], stage2_38[118], stage2_38[119]},
      {stage2_40[66], stage2_40[67], stage2_40[68], stage2_40[69], stage2_40[70], stage2_40[71]},
      {stage3_42[11],stage3_41[18],stage3_40[25],stage3_39[30],stage3_38[43]}
   );
   gpc615_5 gpc7539 (
      {stage2_38[120], stage2_38[121], stage2_38[122], stage2_38[123], stage2_38[124]},
      {stage2_39[42]},
      {stage2_40[72], stage2_40[73], stage2_40[74], stage2_40[75], stage2_40[76], stage2_40[77]},
      {stage3_42[12],stage3_41[19],stage3_40[26],stage3_39[31],stage3_38[44]}
   );
   gpc615_5 gpc7540 (
      {stage2_39[43], stage2_39[44], stage2_39[45], stage2_39[46], stage2_39[47]},
      {stage2_40[78]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[13],stage3_41[20],stage3_40[27],stage3_39[32]}
   );
   gpc615_5 gpc7541 (
      {stage2_39[48], stage2_39[49], stage2_39[50], stage2_39[51], stage2_39[52]},
      {stage2_40[79]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[14],stage3_41[21],stage3_40[28],stage3_39[33]}
   );
   gpc615_5 gpc7542 (
      {stage2_39[53], stage2_39[54], stage2_39[55], stage2_39[56], stage2_39[57]},
      {stage2_40[80]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[15],stage3_41[22],stage3_40[29],stage3_39[34]}
   );
   gpc615_5 gpc7543 (
      {stage2_39[58], stage2_39[59], stage2_39[60], stage2_39[61], stage2_39[62]},
      {stage2_40[81]},
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage3_43[3],stage3_42[16],stage3_41[23],stage3_40[30],stage3_39[35]}
   );
   gpc615_5 gpc7544 (
      {stage2_39[63], stage2_39[64], stage2_39[65], stage2_39[66], stage2_39[67]},
      {stage2_40[82]},
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage3_43[4],stage3_42[17],stage3_41[24],stage3_40[31],stage3_39[36]}
   );
   gpc615_5 gpc7545 (
      {stage2_39[68], stage2_39[69], stage2_39[70], stage2_39[71], stage2_39[72]},
      {stage2_40[83]},
      {stage2_41[30], stage2_41[31], stage2_41[32], stage2_41[33], stage2_41[34], stage2_41[35]},
      {stage3_43[5],stage3_42[18],stage3_41[25],stage3_40[32],stage3_39[37]}
   );
   gpc615_5 gpc7546 (
      {stage2_39[73], stage2_39[74], stage2_39[75], stage2_39[76], stage2_39[77]},
      {stage2_40[84]},
      {stage2_41[36], stage2_41[37], stage2_41[38], stage2_41[39], stage2_41[40], stage2_41[41]},
      {stage3_43[6],stage3_42[19],stage3_41[26],stage3_40[33],stage3_39[38]}
   );
   gpc615_5 gpc7547 (
      {stage2_39[78], stage2_39[79], stage2_39[80], stage2_39[81], stage2_39[82]},
      {stage2_40[85]},
      {stage2_41[42], stage2_41[43], stage2_41[44], stage2_41[45], stage2_41[46], stage2_41[47]},
      {stage3_43[7],stage3_42[20],stage3_41[27],stage3_40[34],stage3_39[39]}
   );
   gpc615_5 gpc7548 (
      {stage2_39[83], stage2_39[84], stage2_39[85], stage2_39[86], stage2_39[87]},
      {stage2_40[86]},
      {stage2_41[48], stage2_41[49], stage2_41[50], stage2_41[51], stage2_41[52], stage2_41[53]},
      {stage3_43[8],stage3_42[21],stage3_41[28],stage3_40[35],stage3_39[40]}
   );
   gpc615_5 gpc7549 (
      {stage2_39[88], stage2_39[89], stage2_39[90], stage2_39[91], stage2_39[92]},
      {stage2_40[87]},
      {stage2_41[54], stage2_41[55], stage2_41[56], stage2_41[57], stage2_41[58], stage2_41[59]},
      {stage3_43[9],stage3_42[22],stage3_41[29],stage3_40[36],stage3_39[41]}
   );
   gpc615_5 gpc7550 (
      {stage2_39[93], stage2_39[94], stage2_39[95], stage2_39[96], stage2_39[97]},
      {stage2_40[88]},
      {stage2_41[60], stage2_41[61], stage2_41[62], stage2_41[63], stage2_41[64], stage2_41[65]},
      {stage3_43[10],stage3_42[23],stage3_41[30],stage3_40[37],stage3_39[42]}
   );
   gpc615_5 gpc7551 (
      {stage2_39[98], stage2_39[99], stage2_39[100], stage2_39[101], stage2_39[102]},
      {stage2_40[89]},
      {stage2_41[66], stage2_41[67], stage2_41[68], stage2_41[69], stage2_41[70], stage2_41[71]},
      {stage3_43[11],stage3_42[24],stage3_41[31],stage3_40[38],stage3_39[43]}
   );
   gpc615_5 gpc7552 (
      {stage2_39[103], stage2_39[104], stage2_39[105], stage2_39[106], stage2_39[107]},
      {stage2_40[90]},
      {stage2_41[72], stage2_41[73], stage2_41[74], stage2_41[75], stage2_41[76], stage2_41[77]},
      {stage3_43[12],stage3_42[25],stage3_41[32],stage3_40[39],stage3_39[44]}
   );
   gpc615_5 gpc7553 (
      {stage2_39[108], stage2_39[109], stage2_39[110], stage2_39[111], stage2_39[112]},
      {stage2_40[91]},
      {stage2_41[78], stage2_41[79], stage2_41[80], stage2_41[81], stage2_41[82], stage2_41[83]},
      {stage3_43[13],stage3_42[26],stage3_41[33],stage3_40[40],stage3_39[45]}
   );
   gpc615_5 gpc7554 (
      {stage2_39[113], stage2_39[114], stage2_39[115], stage2_39[116], stage2_39[117]},
      {stage2_40[92]},
      {stage2_41[84], stage2_41[85], stage2_41[86], stage2_41[87], stage2_41[88], stage2_41[89]},
      {stage3_43[14],stage3_42[27],stage3_41[34],stage3_40[41],stage3_39[46]}
   );
   gpc615_5 gpc7555 (
      {stage2_39[118], stage2_39[119], stage2_39[120], stage2_39[121], stage2_39[122]},
      {stage2_40[93]},
      {stage2_41[90], stage2_41[91], stage2_41[92], stage2_41[93], stage2_41[94], stage2_41[95]},
      {stage3_43[15],stage3_42[28],stage3_41[35],stage3_40[42],stage3_39[47]}
   );
   gpc615_5 gpc7556 (
      {stage2_39[123], stage2_39[124], stage2_39[125], stage2_39[126], stage2_39[127]},
      {stage2_40[94]},
      {stage2_41[96], stage2_41[97], stage2_41[98], stage2_41[99], stage2_41[100], stage2_41[101]},
      {stage3_43[16],stage3_42[29],stage3_41[36],stage3_40[43],stage3_39[48]}
   );
   gpc606_5 gpc7557 (
      {stage2_40[95], stage2_40[96], stage2_40[97], stage2_40[98], stage2_40[99], stage2_40[100]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[17],stage3_42[30],stage3_41[37],stage3_40[44]}
   );
   gpc606_5 gpc7558 (
      {stage2_40[101], stage2_40[102], stage2_40[103], stage2_40[104], stage2_40[105], stage2_40[106]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[18],stage3_42[31],stage3_41[38],stage3_40[45]}
   );
   gpc615_5 gpc7559 (
      {stage2_42[12], stage2_42[13], stage2_42[14], stage2_42[15], stage2_42[16]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[0],stage3_44[2],stage3_43[19],stage3_42[32]}
   );
   gpc615_5 gpc7560 (
      {stage2_42[17], stage2_42[18], stage2_42[19], stage2_42[20], stage2_42[21]},
      {stage2_43[1]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[1],stage3_44[3],stage3_43[20],stage3_42[33]}
   );
   gpc615_5 gpc7561 (
      {stage2_42[22], stage2_42[23], stage2_42[24], stage2_42[25], stage2_42[26]},
      {stage2_43[2]},
      {stage2_44[12], stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17]},
      {stage3_46[2],stage3_45[2],stage3_44[4],stage3_43[21],stage3_42[34]}
   );
   gpc615_5 gpc7562 (
      {stage2_42[27], stage2_42[28], stage2_42[29], stage2_42[30], stage2_42[31]},
      {stage2_43[3]},
      {stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23]},
      {stage3_46[3],stage3_45[3],stage3_44[5],stage3_43[22],stage3_42[35]}
   );
   gpc615_5 gpc7563 (
      {stage2_42[32], stage2_42[33], stage2_42[34], stage2_42[35], stage2_42[36]},
      {stage2_43[4]},
      {stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage3_46[4],stage3_45[4],stage3_44[6],stage3_43[23],stage3_42[36]}
   );
   gpc615_5 gpc7564 (
      {stage2_42[37], stage2_42[38], stage2_42[39], stage2_42[40], stage2_42[41]},
      {stage2_43[5]},
      {stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33], stage2_44[34], stage2_44[35]},
      {stage3_46[5],stage3_45[5],stage3_44[7],stage3_43[24],stage3_42[37]}
   );
   gpc615_5 gpc7565 (
      {stage2_42[42], stage2_42[43], stage2_42[44], stage2_42[45], stage2_42[46]},
      {stage2_43[6]},
      {stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39], stage2_44[40], stage2_44[41]},
      {stage3_46[6],stage3_45[6],stage3_44[8],stage3_43[25],stage3_42[38]}
   );
   gpc615_5 gpc7566 (
      {stage2_42[47], stage2_42[48], stage2_42[49], stage2_42[50], stage2_42[51]},
      {stage2_43[7]},
      {stage2_44[42], stage2_44[43], stage2_44[44], stage2_44[45], stage2_44[46], stage2_44[47]},
      {stage3_46[7],stage3_45[7],stage3_44[9],stage3_43[26],stage3_42[39]}
   );
   gpc615_5 gpc7567 (
      {stage2_42[52], stage2_42[53], stage2_42[54], stage2_42[55], stage2_42[56]},
      {stage2_43[8]},
      {stage2_44[48], stage2_44[49], stage2_44[50], stage2_44[51], stage2_44[52], stage2_44[53]},
      {stage3_46[8],stage3_45[8],stage3_44[10],stage3_43[27],stage3_42[40]}
   );
   gpc615_5 gpc7568 (
      {stage2_42[57], stage2_42[58], stage2_42[59], stage2_42[60], stage2_42[61]},
      {stage2_43[9]},
      {stage2_44[54], stage2_44[55], stage2_44[56], stage2_44[57], stage2_44[58], stage2_44[59]},
      {stage3_46[9],stage3_45[9],stage3_44[11],stage3_43[28],stage3_42[41]}
   );
   gpc615_5 gpc7569 (
      {stage2_42[62], stage2_42[63], stage2_42[64], stage2_42[65], stage2_42[66]},
      {stage2_43[10]},
      {stage2_44[60], stage2_44[61], stage2_44[62], stage2_44[63], stage2_44[64], stage2_44[65]},
      {stage3_46[10],stage3_45[10],stage3_44[12],stage3_43[29],stage3_42[42]}
   );
   gpc615_5 gpc7570 (
      {stage2_42[67], stage2_42[68], stage2_42[69], stage2_42[70], stage2_42[71]},
      {stage2_43[11]},
      {stage2_44[66], stage2_44[67], stage2_44[68], stage2_44[69], stage2_44[70], stage2_44[71]},
      {stage3_46[11],stage3_45[11],stage3_44[13],stage3_43[30],stage3_42[43]}
   );
   gpc615_5 gpc7571 (
      {stage2_42[72], stage2_42[73], stage2_42[74], stage2_42[75], stage2_42[76]},
      {stage2_43[12]},
      {stage2_44[72], stage2_44[73], stage2_44[74], stage2_44[75], stage2_44[76], stage2_44[77]},
      {stage3_46[12],stage3_45[12],stage3_44[14],stage3_43[31],stage3_42[44]}
   );
   gpc615_5 gpc7572 (
      {stage2_42[77], stage2_42[78], stage2_42[79], stage2_42[80], stage2_42[81]},
      {stage2_43[13]},
      {stage2_44[78], stage2_44[79], stage2_44[80], stage2_44[81], stage2_44[82], stage2_44[83]},
      {stage3_46[13],stage3_45[13],stage3_44[15],stage3_43[32],stage3_42[45]}
   );
   gpc615_5 gpc7573 (
      {stage2_43[14], stage2_43[15], stage2_43[16], stage2_43[17], stage2_43[18]},
      {stage2_44[84]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[14],stage3_45[14],stage3_44[16],stage3_43[33]}
   );
   gpc615_5 gpc7574 (
      {stage2_43[19], stage2_43[20], stage2_43[21], stage2_43[22], stage2_43[23]},
      {stage2_44[85]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[15],stage3_45[15],stage3_44[17],stage3_43[34]}
   );
   gpc615_5 gpc7575 (
      {stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27], stage2_43[28]},
      {stage2_44[86]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[16],stage3_45[16],stage3_44[18],stage3_43[35]}
   );
   gpc615_5 gpc7576 (
      {stage2_43[29], stage2_43[30], stage2_43[31], stage2_43[32], stage2_43[33]},
      {stage2_44[87]},
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23]},
      {stage3_47[3],stage3_46[17],stage3_45[17],stage3_44[19],stage3_43[36]}
   );
   gpc615_5 gpc7577 (
      {stage2_43[34], stage2_43[35], stage2_43[36], stage2_43[37], stage2_43[38]},
      {stage2_44[88]},
      {stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27], stage2_45[28], stage2_45[29]},
      {stage3_47[4],stage3_46[18],stage3_45[18],stage3_44[20],stage3_43[37]}
   );
   gpc615_5 gpc7578 (
      {stage2_43[39], stage2_43[40], stage2_43[41], stage2_43[42], stage2_43[43]},
      {stage2_44[89]},
      {stage2_45[30], stage2_45[31], stage2_45[32], stage2_45[33], stage2_45[34], stage2_45[35]},
      {stage3_47[5],stage3_46[19],stage3_45[19],stage3_44[21],stage3_43[38]}
   );
   gpc615_5 gpc7579 (
      {stage2_43[44], stage2_43[45], stage2_43[46], stage2_43[47], stage2_43[48]},
      {stage2_44[90]},
      {stage2_45[36], stage2_45[37], stage2_45[38], stage2_45[39], stage2_45[40], stage2_45[41]},
      {stage3_47[6],stage3_46[20],stage3_45[20],stage3_44[22],stage3_43[39]}
   );
   gpc615_5 gpc7580 (
      {stage2_43[49], stage2_43[50], stage2_43[51], stage2_43[52], stage2_43[53]},
      {stage2_44[91]},
      {stage2_45[42], stage2_45[43], stage2_45[44], stage2_45[45], stage2_45[46], stage2_45[47]},
      {stage3_47[7],stage3_46[21],stage3_45[21],stage3_44[23],stage3_43[40]}
   );
   gpc615_5 gpc7581 (
      {stage2_43[54], stage2_43[55], stage2_43[56], stage2_43[57], stage2_43[58]},
      {stage2_44[92]},
      {stage2_45[48], stage2_45[49], stage2_45[50], stage2_45[51], stage2_45[52], stage2_45[53]},
      {stage3_47[8],stage3_46[22],stage3_45[22],stage3_44[24],stage3_43[41]}
   );
   gpc615_5 gpc7582 (
      {stage2_43[59], stage2_43[60], stage2_43[61], stage2_43[62], stage2_43[63]},
      {stage2_44[93]},
      {stage2_45[54], stage2_45[55], stage2_45[56], stage2_45[57], stage2_45[58], stage2_45[59]},
      {stage3_47[9],stage3_46[23],stage3_45[23],stage3_44[25],stage3_43[42]}
   );
   gpc615_5 gpc7583 (
      {stage2_43[64], stage2_43[65], stage2_43[66], stage2_43[67], stage2_43[68]},
      {stage2_44[94]},
      {stage2_45[60], stage2_45[61], stage2_45[62], stage2_45[63], stage2_45[64], stage2_45[65]},
      {stage3_47[10],stage3_46[24],stage3_45[24],stage3_44[26],stage3_43[43]}
   );
   gpc615_5 gpc7584 (
      {stage2_43[69], stage2_43[70], stage2_43[71], stage2_43[72], stage2_43[73]},
      {stage2_44[95]},
      {stage2_45[66], stage2_45[67], stage2_45[68], stage2_45[69], stage2_45[70], stage2_45[71]},
      {stage3_47[11],stage3_46[25],stage3_45[25],stage3_44[27],stage3_43[44]}
   );
   gpc615_5 gpc7585 (
      {stage2_43[74], stage2_43[75], stage2_43[76], stage2_43[77], stage2_43[78]},
      {stage2_44[96]},
      {stage2_45[72], stage2_45[73], stage2_45[74], stage2_45[75], stage2_45[76], stage2_45[77]},
      {stage3_47[12],stage3_46[26],stage3_45[26],stage3_44[28],stage3_43[45]}
   );
   gpc606_5 gpc7586 (
      {stage2_44[97], stage2_44[98], stage2_44[99], stage2_44[100], stage2_44[101], stage2_44[102]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[13],stage3_46[27],stage3_45[27],stage3_44[29]}
   );
   gpc606_5 gpc7587 (
      {stage2_44[103], stage2_44[104], stage2_44[105], stage2_44[106], stage2_44[107], stage2_44[108]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[14],stage3_46[28],stage3_45[28],stage3_44[30]}
   );
   gpc606_5 gpc7588 (
      {stage2_45[78], stage2_45[79], stage2_45[80], stage2_45[81], stage2_45[82], stage2_45[83]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[2],stage3_47[15],stage3_46[29],stage3_45[29]}
   );
   gpc606_5 gpc7589 (
      {stage2_45[84], stage2_45[85], stage2_45[86], stage2_45[87], stage2_45[88], stage2_45[89]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[3],stage3_47[16],stage3_46[30],stage3_45[30]}
   );
   gpc606_5 gpc7590 (
      {stage2_45[90], stage2_45[91], stage2_45[92], stage2_45[93], stage2_45[94], stage2_45[95]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[4],stage3_47[17],stage3_46[31],stage3_45[31]}
   );
   gpc606_5 gpc7591 (
      {stage2_45[96], stage2_45[97], stage2_45[98], stage2_45[99], stage2_45[100], stage2_45[101]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[5],stage3_47[18],stage3_46[32],stage3_45[32]}
   );
   gpc606_5 gpc7592 (
      {stage2_45[102], stage2_45[103], stage2_45[104], stage2_45[105], stage2_45[106], stage2_45[107]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[6],stage3_47[19],stage3_46[33],stage3_45[33]}
   );
   gpc1163_5 gpc7593 (
      {stage2_46[12], stage2_46[13], stage2_46[14]},
      {stage2_47[30], stage2_47[31], stage2_47[32], stage2_47[33], stage2_47[34], stage2_47[35]},
      {stage2_48[0]},
      {stage2_49[0]},
      {stage3_50[0],stage3_49[5],stage3_48[7],stage3_47[20],stage3_46[34]}
   );
   gpc1163_5 gpc7594 (
      {stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage2_47[36], stage2_47[37], stage2_47[38], stage2_47[39], stage2_47[40], stage2_47[41]},
      {stage2_48[1]},
      {stage2_49[1]},
      {stage3_50[1],stage3_49[6],stage3_48[8],stage3_47[21],stage3_46[35]}
   );
   gpc615_5 gpc7595 (
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22]},
      {stage2_47[42]},
      {stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5], stage2_48[6], stage2_48[7]},
      {stage3_50[2],stage3_49[7],stage3_48[9],stage3_47[22],stage3_46[36]}
   );
   gpc615_5 gpc7596 (
      {stage2_46[23], stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27]},
      {stage2_47[43]},
      {stage2_48[8], stage2_48[9], stage2_48[10], stage2_48[11], stage2_48[12], stage2_48[13]},
      {stage3_50[3],stage3_49[8],stage3_48[10],stage3_47[23],stage3_46[37]}
   );
   gpc615_5 gpc7597 (
      {stage2_46[28], stage2_46[29], stage2_46[30], stage2_46[31], stage2_46[32]},
      {stage2_47[44]},
      {stage2_48[14], stage2_48[15], stage2_48[16], stage2_48[17], stage2_48[18], stage2_48[19]},
      {stage3_50[4],stage3_49[9],stage3_48[11],stage3_47[24],stage3_46[38]}
   );
   gpc615_5 gpc7598 (
      {stage2_46[33], stage2_46[34], stage2_46[35], stage2_46[36], stage2_46[37]},
      {stage2_47[45]},
      {stage2_48[20], stage2_48[21], stage2_48[22], stage2_48[23], stage2_48[24], stage2_48[25]},
      {stage3_50[5],stage3_49[10],stage3_48[12],stage3_47[25],stage3_46[39]}
   );
   gpc615_5 gpc7599 (
      {stage2_46[38], stage2_46[39], stage2_46[40], stage2_46[41], stage2_46[42]},
      {stage2_47[46]},
      {stage2_48[26], stage2_48[27], stage2_48[28], stage2_48[29], stage2_48[30], stage2_48[31]},
      {stage3_50[6],stage3_49[11],stage3_48[13],stage3_47[26],stage3_46[40]}
   );
   gpc615_5 gpc7600 (
      {stage2_46[43], stage2_46[44], stage2_46[45], stage2_46[46], stage2_46[47]},
      {stage2_47[47]},
      {stage2_48[32], stage2_48[33], stage2_48[34], stage2_48[35], stage2_48[36], stage2_48[37]},
      {stage3_50[7],stage3_49[12],stage3_48[14],stage3_47[27],stage3_46[41]}
   );
   gpc615_5 gpc7601 (
      {stage2_46[48], stage2_46[49], stage2_46[50], stage2_46[51], stage2_46[52]},
      {stage2_47[48]},
      {stage2_48[38], stage2_48[39], stage2_48[40], stage2_48[41], stage2_48[42], stage2_48[43]},
      {stage3_50[8],stage3_49[13],stage3_48[15],stage3_47[28],stage3_46[42]}
   );
   gpc615_5 gpc7602 (
      {stage2_46[53], stage2_46[54], stage2_46[55], stage2_46[56], stage2_46[57]},
      {stage2_47[49]},
      {stage2_48[44], stage2_48[45], stage2_48[46], stage2_48[47], stage2_48[48], stage2_48[49]},
      {stage3_50[9],stage3_49[14],stage3_48[16],stage3_47[29],stage3_46[43]}
   );
   gpc615_5 gpc7603 (
      {stage2_46[58], stage2_46[59], stage2_46[60], stage2_46[61], stage2_46[62]},
      {stage2_47[50]},
      {stage2_48[50], stage2_48[51], stage2_48[52], stage2_48[53], stage2_48[54], stage2_48[55]},
      {stage3_50[10],stage3_49[15],stage3_48[17],stage3_47[30],stage3_46[44]}
   );
   gpc615_5 gpc7604 (
      {stage2_46[63], stage2_46[64], stage2_46[65], stage2_46[66], stage2_46[67]},
      {stage2_47[51]},
      {stage2_48[56], stage2_48[57], stage2_48[58], stage2_48[59], stage2_48[60], stage2_48[61]},
      {stage3_50[11],stage3_49[16],stage3_48[18],stage3_47[31],stage3_46[45]}
   );
   gpc615_5 gpc7605 (
      {stage2_46[68], stage2_46[69], stage2_46[70], stage2_46[71], stage2_46[72]},
      {stage2_47[52]},
      {stage2_48[62], stage2_48[63], stage2_48[64], stage2_48[65], stage2_48[66], stage2_48[67]},
      {stage3_50[12],stage3_49[17],stage3_48[19],stage3_47[32],stage3_46[46]}
   );
   gpc615_5 gpc7606 (
      {stage2_46[73], stage2_46[74], stage2_46[75], stage2_46[76], stage2_46[77]},
      {stage2_47[53]},
      {stage2_48[68], stage2_48[69], stage2_48[70], stage2_48[71], stage2_48[72], stage2_48[73]},
      {stage3_50[13],stage3_49[18],stage3_48[20],stage3_47[33],stage3_46[47]}
   );
   gpc615_5 gpc7607 (
      {stage2_47[54], stage2_47[55], stage2_47[56], stage2_47[57], stage2_47[58]},
      {stage2_48[74]},
      {stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5], stage2_49[6], stage2_49[7]},
      {stage3_51[0],stage3_50[14],stage3_49[19],stage3_48[21],stage3_47[34]}
   );
   gpc615_5 gpc7608 (
      {stage2_47[59], stage2_47[60], stage2_47[61], stage2_47[62], stage2_47[63]},
      {stage2_48[75]},
      {stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11], stage2_49[12], stage2_49[13]},
      {stage3_51[1],stage3_50[15],stage3_49[20],stage3_48[22],stage3_47[35]}
   );
   gpc615_5 gpc7609 (
      {stage2_47[64], stage2_47[65], stage2_47[66], stage2_47[67], stage2_47[68]},
      {stage2_48[76]},
      {stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17], stage2_49[18], stage2_49[19]},
      {stage3_51[2],stage3_50[16],stage3_49[21],stage3_48[23],stage3_47[36]}
   );
   gpc615_5 gpc7610 (
      {stage2_47[69], stage2_47[70], stage2_47[71], stage2_47[72], stage2_47[73]},
      {stage2_48[77]},
      {stage2_49[20], stage2_49[21], stage2_49[22], stage2_49[23], stage2_49[24], stage2_49[25]},
      {stage3_51[3],stage3_50[17],stage3_49[22],stage3_48[24],stage3_47[37]}
   );
   gpc615_5 gpc7611 (
      {stage2_47[74], stage2_47[75], stage2_47[76], stage2_47[77], stage2_47[78]},
      {stage2_48[78]},
      {stage2_49[26], stage2_49[27], stage2_49[28], stage2_49[29], stage2_49[30], stage2_49[31]},
      {stage3_51[4],stage3_50[18],stage3_49[23],stage3_48[25],stage3_47[38]}
   );
   gpc615_5 gpc7612 (
      {stage2_47[79], stage2_47[80], stage2_47[81], stage2_47[82], stage2_47[83]},
      {stage2_48[79]},
      {stage2_49[32], stage2_49[33], stage2_49[34], stage2_49[35], stage2_49[36], stage2_49[37]},
      {stage3_51[5],stage3_50[19],stage3_49[24],stage3_48[26],stage3_47[39]}
   );
   gpc615_5 gpc7613 (
      {stage2_47[84], stage2_47[85], stage2_47[86], stage2_47[87], stage2_47[88]},
      {stage2_48[80]},
      {stage2_49[38], stage2_49[39], stage2_49[40], stage2_49[41], stage2_49[42], stage2_49[43]},
      {stage3_51[6],stage3_50[20],stage3_49[25],stage3_48[27],stage3_47[40]}
   );
   gpc615_5 gpc7614 (
      {stage2_47[89], stage2_47[90], stage2_47[91], stage2_47[92], stage2_47[93]},
      {stage2_48[81]},
      {stage2_49[44], stage2_49[45], stage2_49[46], stage2_49[47], stage2_49[48], stage2_49[49]},
      {stage3_51[7],stage3_50[21],stage3_49[26],stage3_48[28],stage3_47[41]}
   );
   gpc615_5 gpc7615 (
      {stage2_47[94], stage2_47[95], stage2_47[96], stage2_47[97], stage2_47[98]},
      {stage2_48[82]},
      {stage2_49[50], stage2_49[51], stage2_49[52], stage2_49[53], stage2_49[54], stage2_49[55]},
      {stage3_51[8],stage3_50[22],stage3_49[27],stage3_48[29],stage3_47[42]}
   );
   gpc615_5 gpc7616 (
      {stage2_47[99], stage2_47[100], stage2_47[101], stage2_47[102], stage2_47[103]},
      {stage2_48[83]},
      {stage2_49[56], stage2_49[57], stage2_49[58], stage2_49[59], stage2_49[60], stage2_49[61]},
      {stage3_51[9],stage3_50[23],stage3_49[28],stage3_48[30],stage3_47[43]}
   );
   gpc606_5 gpc7617 (
      {stage2_48[84], stage2_48[85], stage2_48[86], stage2_48[87], stage2_48[88], stage2_48[89]},
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage3_52[0],stage3_51[10],stage3_50[24],stage3_49[29],stage3_48[31]}
   );
   gpc606_5 gpc7618 (
      {stage2_48[90], stage2_48[91], stage2_48[92], stage2_48[93], stage2_48[94], stage2_48[95]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[1],stage3_51[11],stage3_50[25],stage3_49[30],stage3_48[32]}
   );
   gpc606_5 gpc7619 (
      {stage2_48[96], stage2_48[97], stage2_48[98], stage2_48[99], stage2_48[100], stage2_48[101]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[2],stage3_51[12],stage3_50[26],stage3_49[31],stage3_48[33]}
   );
   gpc606_5 gpc7620 (
      {stage2_48[102], stage2_48[103], stage2_48[104], stage2_48[105], stage2_48[106], stage2_48[107]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[3],stage3_51[13],stage3_50[27],stage3_49[32],stage3_48[34]}
   );
   gpc606_5 gpc7621 (
      {stage2_48[108], stage2_48[109], stage2_48[110], stage2_48[111], stage2_48[112], stage2_48[113]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[4],stage3_51[14],stage3_50[28],stage3_49[33],stage3_48[35]}
   );
   gpc606_5 gpc7622 (
      {stage2_48[114], stage2_48[115], stage2_48[116], stage2_48[117], stage2_48[118], stage2_48[119]},
      {stage2_50[30], stage2_50[31], stage2_50[32], stage2_50[33], stage2_50[34], stage2_50[35]},
      {stage3_52[5],stage3_51[15],stage3_50[29],stage3_49[34],stage3_48[36]}
   );
   gpc606_5 gpc7623 (
      {stage2_48[120], stage2_48[121], stage2_48[122], stage2_48[123], stage2_48[124], stage2_48[125]},
      {stage2_50[36], stage2_50[37], stage2_50[38], stage2_50[39], stage2_50[40], stage2_50[41]},
      {stage3_52[6],stage3_51[16],stage3_50[30],stage3_49[35],stage3_48[37]}
   );
   gpc606_5 gpc7624 (
      {stage2_49[62], stage2_49[63], stage2_49[64], stage2_49[65], stage2_49[66], stage2_49[67]},
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage3_53[0],stage3_52[7],stage3_51[17],stage3_50[31],stage3_49[36]}
   );
   gpc606_5 gpc7625 (
      {stage2_49[68], stage2_49[69], stage2_49[70], stage2_49[71], stage2_49[72], stage2_49[73]},
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11]},
      {stage3_53[1],stage3_52[8],stage3_51[18],stage3_50[32],stage3_49[37]}
   );
   gpc606_5 gpc7626 (
      {stage2_49[74], stage2_49[75], stage2_49[76], stage2_49[77], stage2_49[78], stage2_49[79]},
      {stage2_51[12], stage2_51[13], stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17]},
      {stage3_53[2],stage3_52[9],stage3_51[19],stage3_50[33],stage3_49[38]}
   );
   gpc606_5 gpc7627 (
      {stage2_49[80], stage2_49[81], stage2_49[82], stage2_49[83], stage2_49[84], stage2_49[85]},
      {stage2_51[18], stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23]},
      {stage3_53[3],stage3_52[10],stage3_51[20],stage3_50[34],stage3_49[39]}
   );
   gpc615_5 gpc7628 (
      {stage2_49[86], stage2_49[87], stage2_49[88], stage2_49[89], stage2_49[90]},
      {stage2_50[42]},
      {stage2_51[24], stage2_51[25], stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29]},
      {stage3_53[4],stage3_52[11],stage3_51[21],stage3_50[35],stage3_49[40]}
   );
   gpc615_5 gpc7629 (
      {stage2_49[91], stage2_49[92], stage2_49[93], stage2_49[94], stage2_49[95]},
      {stage2_50[43]},
      {stage2_51[30], stage2_51[31], stage2_51[32], stage2_51[33], stage2_51[34], stage2_51[35]},
      {stage3_53[5],stage3_52[12],stage3_51[22],stage3_50[36],stage3_49[41]}
   );
   gpc615_5 gpc7630 (
      {stage2_50[44], stage2_50[45], stage2_50[46], stage2_50[47], stage2_50[48]},
      {stage2_51[36]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[6],stage3_52[13],stage3_51[23],stage3_50[37]}
   );
   gpc615_5 gpc7631 (
      {stage2_50[49], stage2_50[50], stage2_50[51], stage2_50[52], stage2_50[53]},
      {stage2_51[37]},
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11]},
      {stage3_54[1],stage3_53[7],stage3_52[14],stage3_51[24],stage3_50[38]}
   );
   gpc615_5 gpc7632 (
      {stage2_50[54], stage2_50[55], stage2_50[56], stage2_50[57], stage2_50[58]},
      {stage2_51[38]},
      {stage2_52[12], stage2_52[13], stage2_52[14], stage2_52[15], stage2_52[16], stage2_52[17]},
      {stage3_54[2],stage3_53[8],stage3_52[15],stage3_51[25],stage3_50[39]}
   );
   gpc615_5 gpc7633 (
      {stage2_50[59], stage2_50[60], stage2_50[61], stage2_50[62], stage2_50[63]},
      {stage2_51[39]},
      {stage2_52[18], stage2_52[19], stage2_52[20], stage2_52[21], stage2_52[22], stage2_52[23]},
      {stage3_54[3],stage3_53[9],stage3_52[16],stage3_51[26],stage3_50[40]}
   );
   gpc615_5 gpc7634 (
      {stage2_50[64], stage2_50[65], stage2_50[66], stage2_50[67], stage2_50[68]},
      {stage2_51[40]},
      {stage2_52[24], stage2_52[25], stage2_52[26], stage2_52[27], stage2_52[28], stage2_52[29]},
      {stage3_54[4],stage3_53[10],stage3_52[17],stage3_51[27],stage3_50[41]}
   );
   gpc615_5 gpc7635 (
      {stage2_50[69], stage2_50[70], stage2_50[71], stage2_50[72], stage2_50[73]},
      {stage2_51[41]},
      {stage2_52[30], stage2_52[31], stage2_52[32], stage2_52[33], stage2_52[34], stage2_52[35]},
      {stage3_54[5],stage3_53[11],stage3_52[18],stage3_51[28],stage3_50[42]}
   );
   gpc615_5 gpc7636 (
      {stage2_50[74], stage2_50[75], stage2_50[76], stage2_50[77], stage2_50[78]},
      {stage2_51[42]},
      {stage2_52[36], stage2_52[37], stage2_52[38], stage2_52[39], stage2_52[40], stage2_52[41]},
      {stage3_54[6],stage3_53[12],stage3_52[19],stage3_51[29],stage3_50[43]}
   );
   gpc615_5 gpc7637 (
      {stage2_50[79], stage2_50[80], stage2_50[81], stage2_50[82], stage2_50[83]},
      {stage2_51[43]},
      {stage2_52[42], stage2_52[43], stage2_52[44], stage2_52[45], stage2_52[46], stage2_52[47]},
      {stage3_54[7],stage3_53[13],stage3_52[20],stage3_51[30],stage3_50[44]}
   );
   gpc615_5 gpc7638 (
      {stage2_51[44], stage2_51[45], stage2_51[46], stage2_51[47], stage2_51[48]},
      {stage2_52[48]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[8],stage3_53[14],stage3_52[21],stage3_51[31]}
   );
   gpc615_5 gpc7639 (
      {stage2_51[49], stage2_51[50], stage2_51[51], stage2_51[52], stage2_51[53]},
      {stage2_52[49]},
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage3_55[1],stage3_54[9],stage3_53[15],stage3_52[22],stage3_51[32]}
   );
   gpc615_5 gpc7640 (
      {stage2_51[54], stage2_51[55], stage2_51[56], stage2_51[57], stage2_51[58]},
      {stage2_52[50]},
      {stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage3_55[2],stage3_54[10],stage3_53[16],stage3_52[23],stage3_51[33]}
   );
   gpc606_5 gpc7641 (
      {stage2_52[51], stage2_52[52], stage2_52[53], stage2_52[54], stage2_52[55], stage2_52[56]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[3],stage3_54[11],stage3_53[17],stage3_52[24]}
   );
   gpc606_5 gpc7642 (
      {stage2_52[57], stage2_52[58], stage2_52[59], stage2_52[60], stage2_52[61], stage2_52[62]},
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage3_56[1],stage3_55[4],stage3_54[12],stage3_53[18],stage3_52[25]}
   );
   gpc606_5 gpc7643 (
      {stage2_52[63], stage2_52[64], stage2_52[65], stage2_52[66], stage2_52[67], stage2_52[68]},
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage3_56[2],stage3_55[5],stage3_54[13],stage3_53[19],stage3_52[26]}
   );
   gpc606_5 gpc7644 (
      {stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22], stage2_53[23]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[3],stage3_55[6],stage3_54[14],stage3_53[20]}
   );
   gpc606_5 gpc7645 (
      {stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28], stage2_53[29]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[4],stage3_55[7],stage3_54[15],stage3_53[21]}
   );
   gpc606_5 gpc7646 (
      {stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34], stage2_53[35]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage3_57[2],stage3_56[5],stage3_55[8],stage3_54[16],stage3_53[22]}
   );
   gpc606_5 gpc7647 (
      {stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39], stage2_53[40], stage2_53[41]},
      {stage2_55[18], stage2_55[19], stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23]},
      {stage3_57[3],stage3_56[6],stage3_55[9],stage3_54[17],stage3_53[23]}
   );
   gpc606_5 gpc7648 (
      {stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45], stage2_53[46], stage2_53[47]},
      {stage2_55[24], stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage3_57[4],stage3_56[7],stage3_55[10],stage3_54[18],stage3_53[24]}
   );
   gpc606_5 gpc7649 (
      {stage2_53[48], stage2_53[49], stage2_53[50], stage2_53[51], stage2_53[52], stage2_53[53]},
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34], stage2_55[35]},
      {stage3_57[5],stage3_56[8],stage3_55[11],stage3_54[19],stage3_53[25]}
   );
   gpc615_5 gpc7650 (
      {stage2_53[54], stage2_53[55], stage2_53[56], stage2_53[57], stage2_53[58]},
      {stage2_54[18]},
      {stage2_55[36], stage2_55[37], stage2_55[38], stage2_55[39], stage2_55[40], stage2_55[41]},
      {stage3_57[6],stage3_56[9],stage3_55[12],stage3_54[20],stage3_53[26]}
   );
   gpc615_5 gpc7651 (
      {stage2_53[59], stage2_53[60], stage2_53[61], stage2_53[62], stage2_53[63]},
      {stage2_54[19]},
      {stage2_55[42], stage2_55[43], stage2_55[44], stage2_55[45], stage2_55[46], stage2_55[47]},
      {stage3_57[7],stage3_56[10],stage3_55[13],stage3_54[21],stage3_53[27]}
   );
   gpc615_5 gpc7652 (
      {stage2_53[64], stage2_53[65], stage2_53[66], stage2_53[67], stage2_53[68]},
      {stage2_54[20]},
      {stage2_55[48], stage2_55[49], stage2_55[50], stage2_55[51], stage2_55[52], stage2_55[53]},
      {stage3_57[8],stage3_56[11],stage3_55[14],stage3_54[22],stage3_53[28]}
   );
   gpc615_5 gpc7653 (
      {stage2_54[21], stage2_54[22], stage2_54[23], stage2_54[24], stage2_54[25]},
      {stage2_55[54]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[9],stage3_56[12],stage3_55[15],stage3_54[23]}
   );
   gpc615_5 gpc7654 (
      {stage2_54[26], stage2_54[27], stage2_54[28], stage2_54[29], stage2_54[30]},
      {stage2_55[55]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[10],stage3_56[13],stage3_55[16],stage3_54[24]}
   );
   gpc615_5 gpc7655 (
      {stage2_54[31], stage2_54[32], stage2_54[33], stage2_54[34], stage2_54[35]},
      {stage2_55[56]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[11],stage3_56[14],stage3_55[17],stage3_54[25]}
   );
   gpc615_5 gpc7656 (
      {stage2_54[36], stage2_54[37], stage2_54[38], stage2_54[39], stage2_54[40]},
      {stage2_55[57]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[12],stage3_56[15],stage3_55[18],stage3_54[26]}
   );
   gpc615_5 gpc7657 (
      {stage2_54[41], stage2_54[42], stage2_54[43], stage2_54[44], stage2_54[45]},
      {stage2_55[58]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[13],stage3_56[16],stage3_55[19],stage3_54[27]}
   );
   gpc615_5 gpc7658 (
      {stage2_54[46], stage2_54[47], stage2_54[48], stage2_54[49], stage2_54[50]},
      {stage2_55[59]},
      {stage2_56[30], stage2_56[31], stage2_56[32], stage2_56[33], stage2_56[34], stage2_56[35]},
      {stage3_58[5],stage3_57[14],stage3_56[17],stage3_55[20],stage3_54[28]}
   );
   gpc615_5 gpc7659 (
      {stage2_54[51], stage2_54[52], stage2_54[53], stage2_54[54], stage2_54[55]},
      {stage2_55[60]},
      {stage2_56[36], stage2_56[37], stage2_56[38], stage2_56[39], stage2_56[40], stage2_56[41]},
      {stage3_58[6],stage3_57[15],stage3_56[18],stage3_55[21],stage3_54[29]}
   );
   gpc615_5 gpc7660 (
      {stage2_54[56], stage2_54[57], stage2_54[58], stage2_54[59], stage2_54[60]},
      {stage2_55[61]},
      {stage2_56[42], stage2_56[43], stage2_56[44], stage2_56[45], stage2_56[46], stage2_56[47]},
      {stage3_58[7],stage3_57[16],stage3_56[19],stage3_55[22],stage3_54[30]}
   );
   gpc615_5 gpc7661 (
      {stage2_54[61], stage2_54[62], stage2_54[63], stage2_54[64], stage2_54[65]},
      {stage2_55[62]},
      {stage2_56[48], stage2_56[49], stage2_56[50], stage2_56[51], stage2_56[52], stage2_56[53]},
      {stage3_58[8],stage3_57[17],stage3_56[20],stage3_55[23],stage3_54[31]}
   );
   gpc615_5 gpc7662 (
      {stage2_54[66], stage2_54[67], stage2_54[68], stage2_54[69], stage2_54[70]},
      {stage2_55[63]},
      {stage2_56[54], stage2_56[55], stage2_56[56], stage2_56[57], stage2_56[58], stage2_56[59]},
      {stage3_58[9],stage3_57[18],stage3_56[21],stage3_55[24],stage3_54[32]}
   );
   gpc615_5 gpc7663 (
      {stage2_54[71], stage2_54[72], stage2_54[73], stage2_54[74], stage2_54[75]},
      {stage2_55[64]},
      {stage2_56[60], stage2_56[61], stage2_56[62], stage2_56[63], stage2_56[64], stage2_56[65]},
      {stage3_58[10],stage3_57[19],stage3_56[22],stage3_55[25],stage3_54[33]}
   );
   gpc615_5 gpc7664 (
      {stage2_54[76], stage2_54[77], stage2_54[78], stage2_54[79], stage2_54[80]},
      {stage2_55[65]},
      {stage2_56[66], stage2_56[67], stage2_56[68], stage2_56[69], stage2_56[70], stage2_56[71]},
      {stage3_58[11],stage3_57[20],stage3_56[23],stage3_55[26],stage3_54[34]}
   );
   gpc615_5 gpc7665 (
      {stage2_54[81], stage2_54[82], stage2_54[83], stage2_54[84], stage2_54[85]},
      {stage2_55[66]},
      {stage2_56[72], stage2_56[73], stage2_56[74], stage2_56[75], stage2_56[76], stage2_56[77]},
      {stage3_58[12],stage3_57[21],stage3_56[24],stage3_55[27],stage3_54[35]}
   );
   gpc615_5 gpc7666 (
      {stage2_54[86], stage2_54[87], stage2_54[88], stage2_54[89], stage2_54[90]},
      {stage2_55[67]},
      {stage2_56[78], stage2_56[79], stage2_56[80], stage2_56[81], stage2_56[82], stage2_56[83]},
      {stage3_58[13],stage3_57[22],stage3_56[25],stage3_55[28],stage3_54[36]}
   );
   gpc615_5 gpc7667 (
      {stage2_54[91], stage2_54[92], stage2_54[93], stage2_54[94], stage2_54[95]},
      {stage2_55[68]},
      {stage2_56[84], stage2_56[85], stage2_56[86], stage2_56[87], stage2_56[88], stage2_56[89]},
      {stage3_58[14],stage3_57[23],stage3_56[26],stage3_55[29],stage3_54[37]}
   );
   gpc615_5 gpc7668 (
      {stage2_54[96], stage2_54[97], stage2_54[98], stage2_54[99], 1'b0},
      {stage2_55[69]},
      {stage2_56[90], stage2_56[91], stage2_56[92], stage2_56[93], stage2_56[94], stage2_56[95]},
      {stage3_58[15],stage3_57[24],stage3_56[27],stage3_55[30],stage3_54[38]}
   );
   gpc615_5 gpc7669 (
      {stage2_56[96], stage2_56[97], stage2_56[98], stage2_56[99], stage2_56[100]},
      {stage2_57[0]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[16],stage3_57[25],stage3_56[28]}
   );
   gpc615_5 gpc7670 (
      {stage2_56[101], stage2_56[102], stage2_56[103], stage2_56[104], stage2_56[105]},
      {stage2_57[1]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[1],stage3_58[17],stage3_57[26],stage3_56[29]}
   );
   gpc615_5 gpc7671 (
      {stage2_56[106], stage2_56[107], stage2_56[108], stage2_56[109], stage2_56[110]},
      {stage2_57[2]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage3_60[2],stage3_59[2],stage3_58[18],stage3_57[27],stage3_56[30]}
   );
   gpc615_5 gpc7672 (
      {stage2_56[111], stage2_56[112], stage2_56[113], stage2_56[114], 1'b0},
      {stage2_57[3]},
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23]},
      {stage3_60[3],stage3_59[3],stage3_58[19],stage3_57[28],stage3_56[31]}
   );
   gpc207_4 gpc7673 (
      {stage2_57[4], stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10]},
      {stage2_59[0], stage2_59[1]},
      {stage3_60[4],stage3_59[4],stage3_58[20],stage3_57[29]}
   );
   gpc606_5 gpc7674 (
      {stage2_57[11], stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16]},
      {stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5], stage2_59[6], stage2_59[7]},
      {stage3_61[0],stage3_60[5],stage3_59[5],stage3_58[21],stage3_57[30]}
   );
   gpc606_5 gpc7675 (
      {stage2_57[17], stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22]},
      {stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11], stage2_59[12], stage2_59[13]},
      {stage3_61[1],stage3_60[6],stage3_59[6],stage3_58[22],stage3_57[31]}
   );
   gpc606_5 gpc7676 (
      {stage2_57[23], stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28]},
      {stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17], stage2_59[18], stage2_59[19]},
      {stage3_61[2],stage3_60[7],stage3_59[7],stage3_58[23],stage3_57[32]}
   );
   gpc615_5 gpc7677 (
      {stage2_57[29], stage2_57[30], stage2_57[31], stage2_57[32], stage2_57[33]},
      {stage2_58[24]},
      {stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23], stage2_59[24], stage2_59[25]},
      {stage3_61[3],stage3_60[8],stage3_59[8],stage3_58[24],stage3_57[33]}
   );
   gpc615_5 gpc7678 (
      {stage2_57[34], stage2_57[35], stage2_57[36], stage2_57[37], stage2_57[38]},
      {stage2_58[25]},
      {stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29], stage2_59[30], stage2_59[31]},
      {stage3_61[4],stage3_60[9],stage3_59[9],stage3_58[25],stage3_57[34]}
   );
   gpc615_5 gpc7679 (
      {stage2_57[39], stage2_57[40], stage2_57[41], stage2_57[42], stage2_57[43]},
      {stage2_58[26]},
      {stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35], stage2_59[36], stage2_59[37]},
      {stage3_61[5],stage3_60[10],stage3_59[10],stage3_58[26],stage3_57[35]}
   );
   gpc615_5 gpc7680 (
      {stage2_57[44], stage2_57[45], stage2_57[46], stage2_57[47], stage2_57[48]},
      {stage2_58[27]},
      {stage2_59[38], stage2_59[39], stage2_59[40], stage2_59[41], stage2_59[42], stage2_59[43]},
      {stage3_61[6],stage3_60[11],stage3_59[11],stage3_58[27],stage3_57[36]}
   );
   gpc615_5 gpc7681 (
      {stage2_58[28], stage2_58[29], stage2_58[30], stage2_58[31], stage2_58[32]},
      {stage2_59[44]},
      {stage2_60[0], stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage3_62[0],stage3_61[7],stage3_60[12],stage3_59[12],stage3_58[28]}
   );
   gpc615_5 gpc7682 (
      {stage2_58[33], stage2_58[34], stage2_58[35], stage2_58[36], stage2_58[37]},
      {stage2_59[45]},
      {stage2_60[6], stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11]},
      {stage3_62[1],stage3_61[8],stage3_60[13],stage3_59[13],stage3_58[29]}
   );
   gpc615_5 gpc7683 (
      {stage2_58[38], stage2_58[39], stage2_58[40], stage2_58[41], stage2_58[42]},
      {stage2_59[46]},
      {stage2_60[12], stage2_60[13], stage2_60[14], stage2_60[15], stage2_60[16], stage2_60[17]},
      {stage3_62[2],stage3_61[9],stage3_60[14],stage3_59[14],stage3_58[30]}
   );
   gpc615_5 gpc7684 (
      {stage2_58[43], stage2_58[44], stage2_58[45], stage2_58[46], stage2_58[47]},
      {stage2_59[47]},
      {stage2_60[18], stage2_60[19], stage2_60[20], stage2_60[21], stage2_60[22], stage2_60[23]},
      {stage3_62[3],stage3_61[10],stage3_60[15],stage3_59[15],stage3_58[31]}
   );
   gpc615_5 gpc7685 (
      {stage2_58[48], stage2_58[49], stage2_58[50], stage2_58[51], stage2_58[52]},
      {stage2_59[48]},
      {stage2_60[24], stage2_60[25], stage2_60[26], stage2_60[27], stage2_60[28], stage2_60[29]},
      {stage3_62[4],stage3_61[11],stage3_60[16],stage3_59[16],stage3_58[32]}
   );
   gpc615_5 gpc7686 (
      {stage2_58[53], stage2_58[54], stage2_58[55], stage2_58[56], stage2_58[57]},
      {stage2_59[49]},
      {stage2_60[30], stage2_60[31], stage2_60[32], stage2_60[33], stage2_60[34], stage2_60[35]},
      {stage3_62[5],stage3_61[12],stage3_60[17],stage3_59[17],stage3_58[33]}
   );
   gpc615_5 gpc7687 (
      {stage2_59[50], stage2_59[51], stage2_59[52], stage2_59[53], stage2_59[54]},
      {stage2_60[36]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[6],stage3_61[13],stage3_60[18],stage3_59[18]}
   );
   gpc615_5 gpc7688 (
      {stage2_59[55], stage2_59[56], stage2_59[57], stage2_59[58], stage2_59[59]},
      {stage2_60[37]},
      {stage2_61[6], stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11]},
      {stage3_63[1],stage3_62[7],stage3_61[14],stage3_60[19],stage3_59[19]}
   );
   gpc615_5 gpc7689 (
      {stage2_59[60], stage2_59[61], stage2_59[62], stage2_59[63], stage2_59[64]},
      {stage2_60[38]},
      {stage2_61[12], stage2_61[13], stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17]},
      {stage3_63[2],stage3_62[8],stage3_61[15],stage3_60[20],stage3_59[20]}
   );
   gpc615_5 gpc7690 (
      {stage2_59[65], stage2_59[66], stage2_59[67], stage2_59[68], stage2_59[69]},
      {stage2_60[39]},
      {stage2_61[18], stage2_61[19], stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23]},
      {stage3_63[3],stage3_62[9],stage3_61[16],stage3_60[21],stage3_59[21]}
   );
   gpc615_5 gpc7691 (
      {stage2_59[70], stage2_59[71], stage2_59[72], stage2_59[73], stage2_59[74]},
      {stage2_60[40]},
      {stage2_61[24], stage2_61[25], stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29]},
      {stage3_63[4],stage3_62[10],stage3_61[17],stage3_60[22],stage3_59[22]}
   );
   gpc615_5 gpc7692 (
      {stage2_59[75], stage2_59[76], stage2_59[77], stage2_59[78], stage2_59[79]},
      {stage2_60[41]},
      {stage2_61[30], stage2_61[31], stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35]},
      {stage3_63[5],stage3_62[11],stage3_61[18],stage3_60[23],stage3_59[23]}
   );
   gpc615_5 gpc7693 (
      {stage2_59[80], stage2_59[81], stage2_59[82], stage2_59[83], stage2_59[84]},
      {stage2_60[42]},
      {stage2_61[36], stage2_61[37], stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41]},
      {stage3_63[6],stage3_62[12],stage3_61[19],stage3_60[24],stage3_59[24]}
   );
   gpc606_5 gpc7694 (
      {stage2_60[43], stage2_60[44], stage2_60[45], stage2_60[46], stage2_60[47], stage2_60[48]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[7],stage3_62[13],stage3_61[20],stage3_60[25]}
   );
   gpc606_5 gpc7695 (
      {stage2_60[49], stage2_60[50], stage2_60[51], stage2_60[52], stage2_60[53], stage2_60[54]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[8],stage3_62[14],stage3_61[21],stage3_60[26]}
   );
   gpc606_5 gpc7696 (
      {stage2_60[55], stage2_60[56], stage2_60[57], stage2_60[58], stage2_60[59], stage2_60[60]},
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage3_64[2],stage3_63[9],stage3_62[15],stage3_61[22],stage3_60[27]}
   );
   gpc606_5 gpc7697 (
      {stage2_60[61], stage2_60[62], stage2_60[63], stage2_60[64], stage2_60[65], stage2_60[66]},
      {stage2_62[18], stage2_62[19], stage2_62[20], stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage3_64[3],stage3_63[10],stage3_62[16],stage3_61[23],stage3_60[28]}
   );
   gpc606_5 gpc7698 (
      {stage2_60[67], stage2_60[68], stage2_60[69], stage2_60[70], stage2_60[71], stage2_60[72]},
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage3_64[4],stage3_63[11],stage3_62[17],stage3_61[24],stage3_60[29]}
   );
   gpc606_5 gpc7699 (
      {stage2_61[42], stage2_61[43], stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[5],stage3_63[12],stage3_62[18],stage3_61[25]}
   );
   gpc615_5 gpc7700 (
      {stage2_62[30], stage2_62[31], stage2_62[32], stage2_62[33], stage2_62[34]},
      {stage2_63[6]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[1],stage3_64[6],stage3_63[13],stage3_62[19]}
   );
   gpc615_5 gpc7701 (
      {stage2_62[35], stage2_62[36], stage2_62[37], stage2_62[38], stage2_62[39]},
      {stage2_63[7]},
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10], stage2_64[11]},
      {stage3_66[1],stage3_65[2],stage3_64[7],stage3_63[14],stage3_62[20]}
   );
   gpc615_5 gpc7702 (
      {stage2_62[40], stage2_62[41], stage2_62[42], stage2_62[43], stage2_62[44]},
      {stage2_63[8]},
      {stage2_64[12], stage2_64[13], stage2_64[14], stage2_64[15], stage2_64[16], stage2_64[17]},
      {stage3_66[2],stage3_65[3],stage3_64[8],stage3_63[15],stage3_62[21]}
   );
   gpc615_5 gpc7703 (
      {stage2_62[45], stage2_62[46], stage2_62[47], stage2_62[48], stage2_62[49]},
      {stage2_63[9]},
      {stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21], stage2_64[22], stage2_64[23]},
      {stage3_66[3],stage3_65[4],stage3_64[9],stage3_63[16],stage3_62[22]}
   );
   gpc615_5 gpc7704 (
      {stage2_62[50], stage2_62[51], stage2_62[52], stage2_62[53], stage2_62[54]},
      {stage2_63[10]},
      {stage2_64[24], stage2_64[25], stage2_64[26], stage2_64[27], stage2_64[28], stage2_64[29]},
      {stage3_66[4],stage3_65[5],stage3_64[10],stage3_63[17],stage3_62[23]}
   );
   gpc615_5 gpc7705 (
      {stage2_62[55], stage2_62[56], stage2_62[57], stage2_62[58], stage2_62[59]},
      {stage2_63[11]},
      {stage2_64[30], stage2_64[31], stage2_64[32], stage2_64[33], stage2_64[34], stage2_64[35]},
      {stage3_66[5],stage3_65[6],stage3_64[11],stage3_63[18],stage3_62[24]}
   );
   gpc615_5 gpc7706 (
      {stage2_62[60], stage2_62[61], stage2_62[62], stage2_62[63], stage2_62[64]},
      {stage2_63[12]},
      {stage2_64[36], stage2_64[37], stage2_64[38], stage2_64[39], stage2_64[40], stage2_64[41]},
      {stage3_66[6],stage3_65[7],stage3_64[12],stage3_63[19],stage3_62[25]}
   );
   gpc615_5 gpc7707 (
      {stage2_62[65], stage2_62[66], stage2_62[67], stage2_62[68], stage2_62[69]},
      {stage2_63[13]},
      {stage2_64[42], stage2_64[43], stage2_64[44], stage2_64[45], stage2_64[46], stage2_64[47]},
      {stage3_66[7],stage3_65[8],stage3_64[13],stage3_63[20],stage3_62[26]}
   );
   gpc615_5 gpc7708 (
      {stage2_62[70], stage2_62[71], stage2_62[72], stage2_62[73], stage2_62[74]},
      {stage2_63[14]},
      {stage2_64[48], stage2_64[49], stage2_64[50], stage2_64[51], stage2_64[52], stage2_64[53]},
      {stage3_66[8],stage3_65[9],stage3_64[14],stage3_63[21],stage3_62[27]}
   );
   gpc615_5 gpc7709 (
      {stage2_62[75], stage2_62[76], stage2_62[77], stage2_62[78], stage2_62[79]},
      {stage2_63[15]},
      {stage2_64[54], stage2_64[55], stage2_64[56], stage2_64[57], stage2_64[58], stage2_64[59]},
      {stage3_66[9],stage3_65[10],stage3_64[15],stage3_63[22],stage3_62[28]}
   );
   gpc615_5 gpc7710 (
      {stage2_62[80], stage2_62[81], stage2_62[82], stage2_62[83], stage2_62[84]},
      {stage2_63[16]},
      {stage2_64[60], stage2_64[61], stage2_64[62], stage2_64[63], stage2_64[64], stage2_64[65]},
      {stage3_66[10],stage3_65[11],stage3_64[16],stage3_63[23],stage3_62[29]}
   );
   gpc615_5 gpc7711 (
      {stage2_62[85], stage2_62[86], stage2_62[87], stage2_62[88], stage2_62[89]},
      {stage2_63[17]},
      {stage2_64[66], stage2_64[67], stage2_64[68], stage2_64[69], stage2_64[70], stage2_64[71]},
      {stage3_66[11],stage3_65[12],stage3_64[17],stage3_63[24],stage3_62[30]}
   );
   gpc615_5 gpc7712 (
      {stage2_62[90], stage2_62[91], stage2_62[92], stage2_62[93], stage2_62[94]},
      {stage2_63[18]},
      {stage2_64[72], stage2_64[73], stage2_64[74], stage2_64[75], stage2_64[76], stage2_64[77]},
      {stage3_66[12],stage3_65[13],stage3_64[18],stage3_63[25],stage3_62[31]}
   );
   gpc615_5 gpc7713 (
      {stage2_62[95], stage2_62[96], stage2_62[97], stage2_62[98], stage2_62[99]},
      {stage2_63[19]},
      {stage2_64[78], stage2_64[79], stage2_64[80], stage2_64[81], stage2_64[82], stage2_64[83]},
      {stage3_66[13],stage3_65[14],stage3_64[19],stage3_63[26],stage3_62[32]}
   );
   gpc615_5 gpc7714 (
      {stage2_62[100], stage2_62[101], stage2_62[102], stage2_62[103], stage2_62[104]},
      {stage2_63[20]},
      {stage2_64[84], stage2_64[85], stage2_64[86], stage2_64[87], stage2_64[88], stage2_64[89]},
      {stage3_66[14],stage3_65[15],stage3_64[20],stage3_63[27],stage3_62[33]}
   );
   gpc117_4 gpc7715 (
      {stage2_63[21], stage2_63[22], stage2_63[23], stage2_63[24], stage2_63[25], stage2_63[26], stage2_63[27]},
      {stage2_64[90]},
      {stage2_65[0]},
      {stage3_66[15],stage3_65[16],stage3_64[21],stage3_63[28]}
   );
   gpc117_4 gpc7716 (
      {stage2_63[28], stage2_63[29], stage2_63[30], stage2_63[31], stage2_63[32], stage2_63[33], stage2_63[34]},
      {stage2_64[91]},
      {stage2_65[1]},
      {stage3_66[16],stage3_65[17],stage3_64[22],stage3_63[29]}
   );
   gpc117_4 gpc7717 (
      {stage2_63[35], stage2_63[36], stage2_63[37], stage2_63[38], stage2_63[39], stage2_63[40], stage2_63[41]},
      {stage2_64[92]},
      {stage2_65[2]},
      {stage3_66[17],stage3_65[18],stage3_64[23],stage3_63[30]}
   );
   gpc606_5 gpc7718 (
      {stage2_63[42], stage2_63[43], stage2_63[44], stage2_63[45], stage2_63[46], stage2_63[47]},
      {stage2_65[3], stage2_65[4], stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8]},
      {stage3_67[0],stage3_66[18],stage3_65[19],stage3_64[24],stage3_63[31]}
   );
   gpc606_5 gpc7719 (
      {stage2_63[48], stage2_63[49], stage2_63[50], stage2_63[51], stage2_63[52], stage2_63[53]},
      {stage2_65[9], stage2_65[10], stage2_65[11], stage2_65[12], stage2_65[13], stage2_65[14]},
      {stage3_67[1],stage3_66[19],stage3_65[20],stage3_64[25],stage3_63[32]}
   );
   gpc606_5 gpc7720 (
      {stage2_63[54], stage2_63[55], stage2_63[56], stage2_63[57], stage2_63[58], stage2_63[59]},
      {stage2_65[15], stage2_65[16], stage2_65[17], stage2_65[18], stage2_65[19], stage2_65[20]},
      {stage3_67[2],stage3_66[20],stage3_65[21],stage3_64[26],stage3_63[33]}
   );
   gpc606_5 gpc7721 (
      {stage2_63[60], stage2_63[61], stage2_63[62], stage2_63[63], stage2_63[64], stage2_63[65]},
      {stage2_65[21], stage2_65[22], stage2_65[23], stage2_65[24], stage2_65[25], stage2_65[26]},
      {stage3_67[3],stage3_66[21],stage3_65[22],stage3_64[27],stage3_63[34]}
   );
   gpc606_5 gpc7722 (
      {stage2_63[66], stage2_63[67], stage2_63[68], stage2_63[69], stage2_63[70], stage2_63[71]},
      {stage2_65[27], stage2_65[28], stage2_65[29], stage2_65[30], stage2_65[31], stage2_65[32]},
      {stage3_67[4],stage3_66[22],stage3_65[23],stage3_64[28],stage3_63[35]}
   );
   gpc606_5 gpc7723 (
      {stage2_63[72], stage2_63[73], stage2_63[74], stage2_63[75], stage2_63[76], stage2_63[77]},
      {stage2_65[33], stage2_65[34], stage2_65[35], stage2_65[36], stage2_65[37], stage2_65[38]},
      {stage3_67[5],stage3_66[23],stage3_65[24],stage3_64[29],stage3_63[36]}
   );
   gpc606_5 gpc7724 (
      {stage2_63[78], stage2_63[79], stage2_63[80], stage2_63[81], stage2_63[82], stage2_63[83]},
      {stage2_65[39], stage2_65[40], stage2_65[41], stage2_65[42], stage2_65[43], stage2_65[44]},
      {stage3_67[6],stage3_66[24],stage3_65[25],stage3_64[30],stage3_63[37]}
   );
   gpc606_5 gpc7725 (
      {stage2_63[84], stage2_63[85], stage2_63[86], stage2_63[87], stage2_63[88], stage2_63[89]},
      {stage2_65[45], stage2_65[46], stage2_65[47], stage2_65[48], stage2_65[49], stage2_65[50]},
      {stage3_67[7],stage3_66[25],stage3_65[26],stage3_64[31],stage3_63[38]}
   );
   gpc606_5 gpc7726 (
      {stage2_64[93], stage2_64[94], stage2_64[95], stage2_64[96], stage2_64[97], stage2_64[98]},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3], stage2_66[4], stage2_66[5]},
      {stage3_68[0],stage3_67[8],stage3_66[26],stage3_65[27],stage3_64[32]}
   );
   gpc606_5 gpc7727 (
      {stage2_64[99], stage2_64[100], stage2_64[101], stage2_64[102], stage2_64[103], stage2_64[104]},
      {stage2_66[6], stage2_66[7], stage2_66[8], stage2_66[9], stage2_66[10], stage2_66[11]},
      {stage3_68[1],stage3_67[9],stage3_66[27],stage3_65[28],stage3_64[33]}
   );
   gpc606_5 gpc7728 (
      {stage2_64[105], stage2_64[106], stage2_64[107], stage2_64[108], stage2_64[109], stage2_64[110]},
      {stage2_66[12], stage2_66[13], stage2_66[14], stage2_66[15], stage2_66[16], stage2_66[17]},
      {stage3_68[2],stage3_67[10],stage3_66[28],stage3_65[29],stage3_64[34]}
   );
   gpc606_5 gpc7729 (
      {stage2_64[111], stage2_64[112], stage2_64[113], stage2_64[114], stage2_64[115], stage2_64[116]},
      {stage2_66[18], stage2_66[19], stage2_66[20], stage2_66[21], stage2_66[22], stage2_66[23]},
      {stage3_68[3],stage3_67[11],stage3_66[29],stage3_65[30],stage3_64[35]}
   );
   gpc606_5 gpc7730 (
      {stage2_64[117], stage2_64[118], stage2_64[119], stage2_64[120], stage2_64[121], stage2_64[122]},
      {stage2_66[24], stage2_66[25], stage2_66[26], stage2_66[27], stage2_66[28], stage2_66[29]},
      {stage3_68[4],stage3_67[12],stage3_66[30],stage3_65[31],stage3_64[36]}
   );
   gpc606_5 gpc7731 (
      {stage2_64[123], stage2_64[124], stage2_64[125], stage2_64[126], stage2_64[127], stage2_64[128]},
      {stage2_66[30], stage2_66[31], stage2_66[32], stage2_66[33], stage2_66[34], stage2_66[35]},
      {stage3_68[5],stage3_67[13],stage3_66[31],stage3_65[32],stage3_64[37]}
   );
   gpc1_1 gpc7732 (
      {stage2_0[23]},
      {stage3_0[6]}
   );
   gpc1_1 gpc7733 (
      {stage2_0[24]},
      {stage3_0[7]}
   );
   gpc1_1 gpc7734 (
      {stage2_0[25]},
      {stage3_0[8]}
   );
   gpc1_1 gpc7735 (
      {stage2_0[26]},
      {stage3_0[9]}
   );
   gpc1_1 gpc7736 (
      {stage2_0[27]},
      {stage3_0[10]}
   );
   gpc1_1 gpc7737 (
      {stage2_0[28]},
      {stage3_0[11]}
   );
   gpc1_1 gpc7738 (
      {stage2_0[29]},
      {stage3_0[12]}
   );
   gpc1_1 gpc7739 (
      {stage2_0[30]},
      {stage3_0[13]}
   );
   gpc1_1 gpc7740 (
      {stage2_0[31]},
      {stage3_0[14]}
   );
   gpc1_1 gpc7741 (
      {stage2_0[32]},
      {stage3_0[15]}
   );
   gpc1_1 gpc7742 (
      {stage2_0[33]},
      {stage3_0[16]}
   );
   gpc1_1 gpc7743 (
      {stage2_0[34]},
      {stage3_0[17]}
   );
   gpc1_1 gpc7744 (
      {stage2_0[35]},
      {stage3_0[18]}
   );
   gpc1_1 gpc7745 (
      {stage2_0[36]},
      {stage3_0[19]}
   );
   gpc1_1 gpc7746 (
      {stage2_0[37]},
      {stage3_0[20]}
   );
   gpc1_1 gpc7747 (
      {stage2_1[42]},
      {stage3_1[10]}
   );
   gpc1_1 gpc7748 (
      {stage2_1[43]},
      {stage3_1[11]}
   );
   gpc1_1 gpc7749 (
      {stage2_1[44]},
      {stage3_1[12]}
   );
   gpc1_1 gpc7750 (
      {stage2_1[45]},
      {stage3_1[13]}
   );
   gpc1_1 gpc7751 (
      {stage2_1[46]},
      {stage3_1[14]}
   );
   gpc1_1 gpc7752 (
      {stage2_1[47]},
      {stage3_1[15]}
   );
   gpc1_1 gpc7753 (
      {stage2_1[48]},
      {stage3_1[16]}
   );
   gpc1_1 gpc7754 (
      {stage2_1[49]},
      {stage3_1[17]}
   );
   gpc1_1 gpc7755 (
      {stage2_1[50]},
      {stage3_1[18]}
   );
   gpc1_1 gpc7756 (
      {stage2_1[51]},
      {stage3_1[19]}
   );
   gpc1_1 gpc7757 (
      {stage2_1[52]},
      {stage3_1[20]}
   );
   gpc1_1 gpc7758 (
      {stage2_1[53]},
      {stage3_1[21]}
   );
   gpc1_1 gpc7759 (
      {stage2_2[32]},
      {stage3_2[12]}
   );
   gpc1_1 gpc7760 (
      {stage2_2[33]},
      {stage3_2[13]}
   );
   gpc1_1 gpc7761 (
      {stage2_2[34]},
      {stage3_2[14]}
   );
   gpc1_1 gpc7762 (
      {stage2_2[35]},
      {stage3_2[15]}
   );
   gpc1_1 gpc7763 (
      {stage2_2[36]},
      {stage3_2[16]}
   );
   gpc1_1 gpc7764 (
      {stage2_2[37]},
      {stage3_2[17]}
   );
   gpc1_1 gpc7765 (
      {stage2_2[38]},
      {stage3_2[18]}
   );
   gpc1_1 gpc7766 (
      {stage2_2[39]},
      {stage3_2[19]}
   );
   gpc1_1 gpc7767 (
      {stage2_2[40]},
      {stage3_2[20]}
   );
   gpc1_1 gpc7768 (
      {stage2_2[41]},
      {stage3_2[21]}
   );
   gpc1_1 gpc7769 (
      {stage2_2[42]},
      {stage3_2[22]}
   );
   gpc1_1 gpc7770 (
      {stage2_2[43]},
      {stage3_2[23]}
   );
   gpc1_1 gpc7771 (
      {stage2_2[44]},
      {stage3_2[24]}
   );
   gpc1_1 gpc7772 (
      {stage2_2[45]},
      {stage3_2[25]}
   );
   gpc1_1 gpc7773 (
      {stage2_2[46]},
      {stage3_2[26]}
   );
   gpc1_1 gpc7774 (
      {stage2_2[47]},
      {stage3_2[27]}
   );
   gpc1_1 gpc7775 (
      {stage2_2[48]},
      {stage3_2[28]}
   );
   gpc1_1 gpc7776 (
      {stage2_2[49]},
      {stage3_2[29]}
   );
   gpc1_1 gpc7777 (
      {stage2_2[50]},
      {stage3_2[30]}
   );
   gpc1_1 gpc7778 (
      {stage2_2[51]},
      {stage3_2[31]}
   );
   gpc1_1 gpc7779 (
      {stage2_2[52]},
      {stage3_2[32]}
   );
   gpc1_1 gpc7780 (
      {stage2_2[53]},
      {stage3_2[33]}
   );
   gpc1_1 gpc7781 (
      {stage2_2[54]},
      {stage3_2[34]}
   );
   gpc1_1 gpc7782 (
      {stage2_2[55]},
      {stage3_2[35]}
   );
   gpc1_1 gpc7783 (
      {stage2_2[56]},
      {stage3_2[36]}
   );
   gpc1_1 gpc7784 (
      {stage2_2[57]},
      {stage3_2[37]}
   );
   gpc1_1 gpc7785 (
      {stage2_2[58]},
      {stage3_2[38]}
   );
   gpc1_1 gpc7786 (
      {stage2_2[59]},
      {stage3_2[39]}
   );
   gpc1_1 gpc7787 (
      {stage2_2[60]},
      {stage3_2[40]}
   );
   gpc1_1 gpc7788 (
      {stage2_2[61]},
      {stage3_2[41]}
   );
   gpc1_1 gpc7789 (
      {stage2_2[62]},
      {stage3_2[42]}
   );
   gpc1_1 gpc7790 (
      {stage2_4[29]},
      {stage3_4[29]}
   );
   gpc1_1 gpc7791 (
      {stage2_4[30]},
      {stage3_4[30]}
   );
   gpc1_1 gpc7792 (
      {stage2_4[31]},
      {stage3_4[31]}
   );
   gpc1_1 gpc7793 (
      {stage2_4[32]},
      {stage3_4[32]}
   );
   gpc1_1 gpc7794 (
      {stage2_4[33]},
      {stage3_4[33]}
   );
   gpc1_1 gpc7795 (
      {stage2_4[34]},
      {stage3_4[34]}
   );
   gpc1_1 gpc7796 (
      {stage2_4[35]},
      {stage3_4[35]}
   );
   gpc1_1 gpc7797 (
      {stage2_4[36]},
      {stage3_4[36]}
   );
   gpc1_1 gpc7798 (
      {stage2_4[37]},
      {stage3_4[37]}
   );
   gpc1_1 gpc7799 (
      {stage2_4[38]},
      {stage3_4[38]}
   );
   gpc1_1 gpc7800 (
      {stage2_4[39]},
      {stage3_4[39]}
   );
   gpc1_1 gpc7801 (
      {stage2_4[40]},
      {stage3_4[40]}
   );
   gpc1_1 gpc7802 (
      {stage2_4[41]},
      {stage3_4[41]}
   );
   gpc1_1 gpc7803 (
      {stage2_4[42]},
      {stage3_4[42]}
   );
   gpc1_1 gpc7804 (
      {stage2_4[43]},
      {stage3_4[43]}
   );
   gpc1_1 gpc7805 (
      {stage2_4[44]},
      {stage3_4[44]}
   );
   gpc1_1 gpc7806 (
      {stage2_4[45]},
      {stage3_4[45]}
   );
   gpc1_1 gpc7807 (
      {stage2_4[46]},
      {stage3_4[46]}
   );
   gpc1_1 gpc7808 (
      {stage2_4[47]},
      {stage3_4[47]}
   );
   gpc1_1 gpc7809 (
      {stage2_4[48]},
      {stage3_4[48]}
   );
   gpc1_1 gpc7810 (
      {stage2_4[49]},
      {stage3_4[49]}
   );
   gpc1_1 gpc7811 (
      {stage2_4[50]},
      {stage3_4[50]}
   );
   gpc1_1 gpc7812 (
      {stage2_4[51]},
      {stage3_4[51]}
   );
   gpc1_1 gpc7813 (
      {stage2_4[52]},
      {stage3_4[52]}
   );
   gpc1_1 gpc7814 (
      {stage2_4[53]},
      {stage3_4[53]}
   );
   gpc1_1 gpc7815 (
      {stage2_4[54]},
      {stage3_4[54]}
   );
   gpc1_1 gpc7816 (
      {stage2_4[55]},
      {stage3_4[55]}
   );
   gpc1_1 gpc7817 (
      {stage2_4[56]},
      {stage3_4[56]}
   );
   gpc1_1 gpc7818 (
      {stage2_4[57]},
      {stage3_4[57]}
   );
   gpc1_1 gpc7819 (
      {stage2_4[58]},
      {stage3_4[58]}
   );
   gpc1_1 gpc7820 (
      {stage2_4[59]},
      {stage3_4[59]}
   );
   gpc1_1 gpc7821 (
      {stage2_4[60]},
      {stage3_4[60]}
   );
   gpc1_1 gpc7822 (
      {stage2_4[61]},
      {stage3_4[61]}
   );
   gpc1_1 gpc7823 (
      {stage2_4[62]},
      {stage3_4[62]}
   );
   gpc1_1 gpc7824 (
      {stage2_4[63]},
      {stage3_4[63]}
   );
   gpc1_1 gpc7825 (
      {stage2_4[64]},
      {stage3_4[64]}
   );
   gpc1_1 gpc7826 (
      {stage2_4[65]},
      {stage3_4[65]}
   );
   gpc1_1 gpc7827 (
      {stage2_4[66]},
      {stage3_4[66]}
   );
   gpc1_1 gpc7828 (
      {stage2_4[67]},
      {stage3_4[67]}
   );
   gpc1_1 gpc7829 (
      {stage2_4[68]},
      {stage3_4[68]}
   );
   gpc1_1 gpc7830 (
      {stage2_4[69]},
      {stage3_4[69]}
   );
   gpc1_1 gpc7831 (
      {stage2_4[70]},
      {stage3_4[70]}
   );
   gpc1_1 gpc7832 (
      {stage2_4[71]},
      {stage3_4[71]}
   );
   gpc1_1 gpc7833 (
      {stage2_4[72]},
      {stage3_4[72]}
   );
   gpc1_1 gpc7834 (
      {stage2_4[73]},
      {stage3_4[73]}
   );
   gpc1_1 gpc7835 (
      {stage2_4[74]},
      {stage3_4[74]}
   );
   gpc1_1 gpc7836 (
      {stage2_4[75]},
      {stage3_4[75]}
   );
   gpc1_1 gpc7837 (
      {stage2_4[76]},
      {stage3_4[76]}
   );
   gpc1_1 gpc7838 (
      {stage2_4[77]},
      {stage3_4[77]}
   );
   gpc1_1 gpc7839 (
      {stage2_4[78]},
      {stage3_4[78]}
   );
   gpc1_1 gpc7840 (
      {stage2_4[79]},
      {stage3_4[79]}
   );
   gpc1_1 gpc7841 (
      {stage2_4[80]},
      {stage3_4[80]}
   );
   gpc1_1 gpc7842 (
      {stage2_4[81]},
      {stage3_4[81]}
   );
   gpc1_1 gpc7843 (
      {stage2_4[82]},
      {stage3_4[82]}
   );
   gpc1_1 gpc7844 (
      {stage2_4[83]},
      {stage3_4[83]}
   );
   gpc1_1 gpc7845 (
      {stage2_4[84]},
      {stage3_4[84]}
   );
   gpc1_1 gpc7846 (
      {stage2_4[85]},
      {stage3_4[85]}
   );
   gpc1_1 gpc7847 (
      {stage2_4[86]},
      {stage3_4[86]}
   );
   gpc1_1 gpc7848 (
      {stage2_4[87]},
      {stage3_4[87]}
   );
   gpc1_1 gpc7849 (
      {stage2_4[88]},
      {stage3_4[88]}
   );
   gpc1_1 gpc7850 (
      {stage2_4[89]},
      {stage3_4[89]}
   );
   gpc1_1 gpc7851 (
      {stage2_4[90]},
      {stage3_4[90]}
   );
   gpc1_1 gpc7852 (
      {stage2_4[91]},
      {stage3_4[91]}
   );
   gpc1_1 gpc7853 (
      {stage2_4[92]},
      {stage3_4[92]}
   );
   gpc1_1 gpc7854 (
      {stage2_4[93]},
      {stage3_4[93]}
   );
   gpc1_1 gpc7855 (
      {stage2_4[94]},
      {stage3_4[94]}
   );
   gpc1_1 gpc7856 (
      {stage2_4[95]},
      {stage3_4[95]}
   );
   gpc1_1 gpc7857 (
      {stage2_4[96]},
      {stage3_4[96]}
   );
   gpc1_1 gpc7858 (
      {stage2_4[97]},
      {stage3_4[97]}
   );
   gpc1_1 gpc7859 (
      {stage2_4[98]},
      {stage3_4[98]}
   );
   gpc1_1 gpc7860 (
      {stage2_4[99]},
      {stage3_4[99]}
   );
   gpc1_1 gpc7861 (
      {stage2_4[100]},
      {stage3_4[100]}
   );
   gpc1_1 gpc7862 (
      {stage2_4[101]},
      {stage3_4[101]}
   );
   gpc1_1 gpc7863 (
      {stage2_4[102]},
      {stage3_4[102]}
   );
   gpc1_1 gpc7864 (
      {stage2_4[103]},
      {stage3_4[103]}
   );
   gpc1_1 gpc7865 (
      {stage2_4[104]},
      {stage3_4[104]}
   );
   gpc1_1 gpc7866 (
      {stage2_4[105]},
      {stage3_4[105]}
   );
   gpc1_1 gpc7867 (
      {stage2_4[106]},
      {stage3_4[106]}
   );
   gpc1_1 gpc7868 (
      {stage2_4[107]},
      {stage3_4[107]}
   );
   gpc1_1 gpc7869 (
      {stage2_4[108]},
      {stage3_4[108]}
   );
   gpc1_1 gpc7870 (
      {stage2_4[109]},
      {stage3_4[109]}
   );
   gpc1_1 gpc7871 (
      {stage2_4[110]},
      {stage3_4[110]}
   );
   gpc1_1 gpc7872 (
      {stage2_4[111]},
      {stage3_4[111]}
   );
   gpc1_1 gpc7873 (
      {stage2_5[126]},
      {stage3_5[27]}
   );
   gpc1_1 gpc7874 (
      {stage2_5[127]},
      {stage3_5[28]}
   );
   gpc1_1 gpc7875 (
      {stage2_5[128]},
      {stage3_5[29]}
   );
   gpc1_1 gpc7876 (
      {stage2_5[129]},
      {stage3_5[30]}
   );
   gpc1_1 gpc7877 (
      {stage2_5[130]},
      {stage3_5[31]}
   );
   gpc1_1 gpc7878 (
      {stage2_5[131]},
      {stage3_5[32]}
   );
   gpc1_1 gpc7879 (
      {stage2_5[132]},
      {stage3_5[33]}
   );
   gpc1_1 gpc7880 (
      {stage2_5[133]},
      {stage3_5[34]}
   );
   gpc1_1 gpc7881 (
      {stage2_5[134]},
      {stage3_5[35]}
   );
   gpc1_1 gpc7882 (
      {stage2_5[135]},
      {stage3_5[36]}
   );
   gpc1_1 gpc7883 (
      {stage2_5[136]},
      {stage3_5[37]}
   );
   gpc1_1 gpc7884 (
      {stage2_5[137]},
      {stage3_5[38]}
   );
   gpc1_1 gpc7885 (
      {stage2_5[138]},
      {stage3_5[39]}
   );
   gpc1_1 gpc7886 (
      {stage2_5[139]},
      {stage3_5[40]}
   );
   gpc1_1 gpc7887 (
      {stage2_5[140]},
      {stage3_5[41]}
   );
   gpc1_1 gpc7888 (
      {stage2_5[141]},
      {stage3_5[42]}
   );
   gpc1_1 gpc7889 (
      {stage2_5[142]},
      {stage3_5[43]}
   );
   gpc1_1 gpc7890 (
      {stage2_5[143]},
      {stage3_5[44]}
   );
   gpc1_1 gpc7891 (
      {stage2_5[144]},
      {stage3_5[45]}
   );
   gpc1_1 gpc7892 (
      {stage2_5[145]},
      {stage3_5[46]}
   );
   gpc1_1 gpc7893 (
      {stage2_5[146]},
      {stage3_5[47]}
   );
   gpc1_1 gpc7894 (
      {stage2_5[147]},
      {stage3_5[48]}
   );
   gpc1_1 gpc7895 (
      {stage2_5[148]},
      {stage3_5[49]}
   );
   gpc1_1 gpc7896 (
      {stage2_5[149]},
      {stage3_5[50]}
   );
   gpc1_1 gpc7897 (
      {stage2_5[150]},
      {stage3_5[51]}
   );
   gpc1_1 gpc7898 (
      {stage2_5[151]},
      {stage3_5[52]}
   );
   gpc1_1 gpc7899 (
      {stage2_6[46]},
      {stage3_6[32]}
   );
   gpc1_1 gpc7900 (
      {stage2_6[47]},
      {stage3_6[33]}
   );
   gpc1_1 gpc7901 (
      {stage2_6[48]},
      {stage3_6[34]}
   );
   gpc1_1 gpc7902 (
      {stage2_6[49]},
      {stage3_6[35]}
   );
   gpc1_1 gpc7903 (
      {stage2_6[50]},
      {stage3_6[36]}
   );
   gpc1_1 gpc7904 (
      {stage2_6[51]},
      {stage3_6[37]}
   );
   gpc1_1 gpc7905 (
      {stage2_6[52]},
      {stage3_6[38]}
   );
   gpc1_1 gpc7906 (
      {stage2_6[53]},
      {stage3_6[39]}
   );
   gpc1_1 gpc7907 (
      {stage2_6[54]},
      {stage3_6[40]}
   );
   gpc1_1 gpc7908 (
      {stage2_6[55]},
      {stage3_6[41]}
   );
   gpc1_1 gpc7909 (
      {stage2_6[56]},
      {stage3_6[42]}
   );
   gpc1_1 gpc7910 (
      {stage2_6[57]},
      {stage3_6[43]}
   );
   gpc1_1 gpc7911 (
      {stage2_6[58]},
      {stage3_6[44]}
   );
   gpc1_1 gpc7912 (
      {stage2_6[59]},
      {stage3_6[45]}
   );
   gpc1_1 gpc7913 (
      {stage2_6[60]},
      {stage3_6[46]}
   );
   gpc1_1 gpc7914 (
      {stage2_6[61]},
      {stage3_6[47]}
   );
   gpc1_1 gpc7915 (
      {stage2_6[62]},
      {stage3_6[48]}
   );
   gpc1_1 gpc7916 (
      {stage2_6[63]},
      {stage3_6[49]}
   );
   gpc1_1 gpc7917 (
      {stage2_6[64]},
      {stage3_6[50]}
   );
   gpc1_1 gpc7918 (
      {stage2_6[65]},
      {stage3_6[51]}
   );
   gpc1_1 gpc7919 (
      {stage2_6[66]},
      {stage3_6[52]}
   );
   gpc1_1 gpc7920 (
      {stage2_6[67]},
      {stage3_6[53]}
   );
   gpc1_1 gpc7921 (
      {stage2_6[68]},
      {stage3_6[54]}
   );
   gpc1_1 gpc7922 (
      {stage2_6[69]},
      {stage3_6[55]}
   );
   gpc1_1 gpc7923 (
      {stage2_6[70]},
      {stage3_6[56]}
   );
   gpc1_1 gpc7924 (
      {stage2_6[71]},
      {stage3_6[57]}
   );
   gpc1_1 gpc7925 (
      {stage2_6[72]},
      {stage3_6[58]}
   );
   gpc1_1 gpc7926 (
      {stage2_6[73]},
      {stage3_6[59]}
   );
   gpc1_1 gpc7927 (
      {stage2_6[74]},
      {stage3_6[60]}
   );
   gpc1_1 gpc7928 (
      {stage2_6[75]},
      {stage3_6[61]}
   );
   gpc1_1 gpc7929 (
      {stage2_6[76]},
      {stage3_6[62]}
   );
   gpc1_1 gpc7930 (
      {stage2_6[77]},
      {stage3_6[63]}
   );
   gpc1_1 gpc7931 (
      {stage2_6[78]},
      {stage3_6[64]}
   );
   gpc1_1 gpc7932 (
      {stage2_6[79]},
      {stage3_6[65]}
   );
   gpc1_1 gpc7933 (
      {stage2_6[80]},
      {stage3_6[66]}
   );
   gpc1_1 gpc7934 (
      {stage2_6[81]},
      {stage3_6[67]}
   );
   gpc1_1 gpc7935 (
      {stage2_6[82]},
      {stage3_6[68]}
   );
   gpc1_1 gpc7936 (
      {stage2_6[83]},
      {stage3_6[69]}
   );
   gpc1_1 gpc7937 (
      {stage2_6[84]},
      {stage3_6[70]}
   );
   gpc1_1 gpc7938 (
      {stage2_6[85]},
      {stage3_6[71]}
   );
   gpc1_1 gpc7939 (
      {stage2_6[86]},
      {stage3_6[72]}
   );
   gpc1_1 gpc7940 (
      {stage2_6[87]},
      {stage3_6[73]}
   );
   gpc1_1 gpc7941 (
      {stage2_6[88]},
      {stage3_6[74]}
   );
   gpc1_1 gpc7942 (
      {stage2_6[89]},
      {stage3_6[75]}
   );
   gpc1_1 gpc7943 (
      {stage2_6[90]},
      {stage3_6[76]}
   );
   gpc1_1 gpc7944 (
      {stage2_6[91]},
      {stage3_6[77]}
   );
   gpc1_1 gpc7945 (
      {stage2_7[57]},
      {stage3_7[35]}
   );
   gpc1_1 gpc7946 (
      {stage2_7[58]},
      {stage3_7[36]}
   );
   gpc1_1 gpc7947 (
      {stage2_7[59]},
      {stage3_7[37]}
   );
   gpc1_1 gpc7948 (
      {stage2_7[60]},
      {stage3_7[38]}
   );
   gpc1_1 gpc7949 (
      {stage2_7[61]},
      {stage3_7[39]}
   );
   gpc1_1 gpc7950 (
      {stage2_7[62]},
      {stage3_7[40]}
   );
   gpc1_1 gpc7951 (
      {stage2_7[63]},
      {stage3_7[41]}
   );
   gpc1_1 gpc7952 (
      {stage2_7[64]},
      {stage3_7[42]}
   );
   gpc1_1 gpc7953 (
      {stage2_7[65]},
      {stage3_7[43]}
   );
   gpc1_1 gpc7954 (
      {stage2_7[66]},
      {stage3_7[44]}
   );
   gpc1_1 gpc7955 (
      {stage2_7[67]},
      {stage3_7[45]}
   );
   gpc1_1 gpc7956 (
      {stage2_7[68]},
      {stage3_7[46]}
   );
   gpc1_1 gpc7957 (
      {stage2_7[69]},
      {stage3_7[47]}
   );
   gpc1_1 gpc7958 (
      {stage2_7[70]},
      {stage3_7[48]}
   );
   gpc1_1 gpc7959 (
      {stage2_7[71]},
      {stage3_7[49]}
   );
   gpc1_1 gpc7960 (
      {stage2_7[72]},
      {stage3_7[50]}
   );
   gpc1_1 gpc7961 (
      {stage2_10[117]},
      {stage3_10[53]}
   );
   gpc1_1 gpc7962 (
      {stage2_10[118]},
      {stage3_10[54]}
   );
   gpc1_1 gpc7963 (
      {stage2_10[119]},
      {stage3_10[55]}
   );
   gpc1_1 gpc7964 (
      {stage2_10[120]},
      {stage3_10[56]}
   );
   gpc1_1 gpc7965 (
      {stage2_10[121]},
      {stage3_10[57]}
   );
   gpc1_1 gpc7966 (
      {stage2_10[122]},
      {stage3_10[58]}
   );
   gpc1_1 gpc7967 (
      {stage2_10[123]},
      {stage3_10[59]}
   );
   gpc1_1 gpc7968 (
      {stage2_10[124]},
      {stage3_10[60]}
   );
   gpc1_1 gpc7969 (
      {stage2_10[125]},
      {stage3_10[61]}
   );
   gpc1_1 gpc7970 (
      {stage2_10[126]},
      {stage3_10[62]}
   );
   gpc1_1 gpc7971 (
      {stage2_10[127]},
      {stage3_10[63]}
   );
   gpc1_1 gpc7972 (
      {stage2_10[128]},
      {stage3_10[64]}
   );
   gpc1_1 gpc7973 (
      {stage2_10[129]},
      {stage3_10[65]}
   );
   gpc1_1 gpc7974 (
      {stage2_10[130]},
      {stage3_10[66]}
   );
   gpc1_1 gpc7975 (
      {stage2_10[131]},
      {stage3_10[67]}
   );
   gpc1_1 gpc7976 (
      {stage2_10[132]},
      {stage3_10[68]}
   );
   gpc1_1 gpc7977 (
      {stage2_10[133]},
      {stage3_10[69]}
   );
   gpc1_1 gpc7978 (
      {stage2_10[134]},
      {stage3_10[70]}
   );
   gpc1_1 gpc7979 (
      {stage2_10[135]},
      {stage3_10[71]}
   );
   gpc1_1 gpc7980 (
      {stage2_10[136]},
      {stage3_10[72]}
   );
   gpc1_1 gpc7981 (
      {stage2_10[137]},
      {stage3_10[73]}
   );
   gpc1_1 gpc7982 (
      {stage2_10[138]},
      {stage3_10[74]}
   );
   gpc1_1 gpc7983 (
      {stage2_10[139]},
      {stage3_10[75]}
   );
   gpc1_1 gpc7984 (
      {stage2_10[140]},
      {stage3_10[76]}
   );
   gpc1_1 gpc7985 (
      {stage2_10[141]},
      {stage3_10[77]}
   );
   gpc1_1 gpc7986 (
      {stage2_10[142]},
      {stage3_10[78]}
   );
   gpc1_1 gpc7987 (
      {stage2_10[143]},
      {stage3_10[79]}
   );
   gpc1_1 gpc7988 (
      {stage2_10[144]},
      {stage3_10[80]}
   );
   gpc1_1 gpc7989 (
      {stage2_10[145]},
      {stage3_10[81]}
   );
   gpc1_1 gpc7990 (
      {stage2_10[146]},
      {stage3_10[82]}
   );
   gpc1_1 gpc7991 (
      {stage2_10[147]},
      {stage3_10[83]}
   );
   gpc1_1 gpc7992 (
      {stage2_10[148]},
      {stage3_10[84]}
   );
   gpc1_1 gpc7993 (
      {stage2_10[149]},
      {stage3_10[85]}
   );
   gpc1_1 gpc7994 (
      {stage2_10[150]},
      {stage3_10[86]}
   );
   gpc1_1 gpc7995 (
      {stage2_10[151]},
      {stage3_10[87]}
   );
   gpc1_1 gpc7996 (
      {stage2_10[152]},
      {stage3_10[88]}
   );
   gpc1_1 gpc7997 (
      {stage2_10[153]},
      {stage3_10[89]}
   );
   gpc1_1 gpc7998 (
      {stage2_10[154]},
      {stage3_10[90]}
   );
   gpc1_1 gpc7999 (
      {stage2_10[155]},
      {stage3_10[91]}
   );
   gpc1_1 gpc8000 (
      {stage2_10[156]},
      {stage3_10[92]}
   );
   gpc1_1 gpc8001 (
      {stage2_10[157]},
      {stage3_10[93]}
   );
   gpc1_1 gpc8002 (
      {stage2_10[158]},
      {stage3_10[94]}
   );
   gpc1_1 gpc8003 (
      {stage2_10[159]},
      {stage3_10[95]}
   );
   gpc1_1 gpc8004 (
      {stage2_10[160]},
      {stage3_10[96]}
   );
   gpc1_1 gpc8005 (
      {stage2_10[161]},
      {stage3_10[97]}
   );
   gpc1_1 gpc8006 (
      {stage2_10[162]},
      {stage3_10[98]}
   );
   gpc1_1 gpc8007 (
      {stage2_10[163]},
      {stage3_10[99]}
   );
   gpc1_1 gpc8008 (
      {stage2_11[127]},
      {stage3_11[46]}
   );
   gpc1_1 gpc8009 (
      {stage2_11[128]},
      {stage3_11[47]}
   );
   gpc1_1 gpc8010 (
      {stage2_11[129]},
      {stage3_11[48]}
   );
   gpc1_1 gpc8011 (
      {stage2_11[130]},
      {stage3_11[49]}
   );
   gpc1_1 gpc8012 (
      {stage2_11[131]},
      {stage3_11[50]}
   );
   gpc1_1 gpc8013 (
      {stage2_11[132]},
      {stage3_11[51]}
   );
   gpc1_1 gpc8014 (
      {stage2_11[133]},
      {stage3_11[52]}
   );
   gpc1_1 gpc8015 (
      {stage2_11[134]},
      {stage3_11[53]}
   );
   gpc1_1 gpc8016 (
      {stage2_11[135]},
      {stage3_11[54]}
   );
   gpc1_1 gpc8017 (
      {stage2_11[136]},
      {stage3_11[55]}
   );
   gpc1_1 gpc8018 (
      {stage2_11[137]},
      {stage3_11[56]}
   );
   gpc1_1 gpc8019 (
      {stage2_11[138]},
      {stage3_11[57]}
   );
   gpc1_1 gpc8020 (
      {stage2_12[92]},
      {stage3_12[53]}
   );
   gpc1_1 gpc8021 (
      {stage2_12[93]},
      {stage3_12[54]}
   );
   gpc1_1 gpc8022 (
      {stage2_12[94]},
      {stage3_12[55]}
   );
   gpc1_1 gpc8023 (
      {stage2_12[95]},
      {stage3_12[56]}
   );
   gpc1_1 gpc8024 (
      {stage2_12[96]},
      {stage3_12[57]}
   );
   gpc1_1 gpc8025 (
      {stage2_12[97]},
      {stage3_12[58]}
   );
   gpc1_1 gpc8026 (
      {stage2_12[98]},
      {stage3_12[59]}
   );
   gpc1_1 gpc8027 (
      {stage2_12[99]},
      {stage3_12[60]}
   );
   gpc1_1 gpc8028 (
      {stage2_12[100]},
      {stage3_12[61]}
   );
   gpc1_1 gpc8029 (
      {stage2_12[101]},
      {stage3_12[62]}
   );
   gpc1_1 gpc8030 (
      {stage2_12[102]},
      {stage3_12[63]}
   );
   gpc1_1 gpc8031 (
      {stage2_12[103]},
      {stage3_12[64]}
   );
   gpc1_1 gpc8032 (
      {stage2_12[104]},
      {stage3_12[65]}
   );
   gpc1_1 gpc8033 (
      {stage2_12[105]},
      {stage3_12[66]}
   );
   gpc1_1 gpc8034 (
      {stage2_12[106]},
      {stage3_12[67]}
   );
   gpc1_1 gpc8035 (
      {stage2_13[66]},
      {stage3_13[45]}
   );
   gpc1_1 gpc8036 (
      {stage2_13[67]},
      {stage3_13[46]}
   );
   gpc1_1 gpc8037 (
      {stage2_13[68]},
      {stage3_13[47]}
   );
   gpc1_1 gpc8038 (
      {stage2_13[69]},
      {stage3_13[48]}
   );
   gpc1_1 gpc8039 (
      {stage2_13[70]},
      {stage3_13[49]}
   );
   gpc1_1 gpc8040 (
      {stage2_13[71]},
      {stage3_13[50]}
   );
   gpc1_1 gpc8041 (
      {stage2_13[72]},
      {stage3_13[51]}
   );
   gpc1_1 gpc8042 (
      {stage2_13[73]},
      {stage3_13[52]}
   );
   gpc1_1 gpc8043 (
      {stage2_13[74]},
      {stage3_13[53]}
   );
   gpc1_1 gpc8044 (
      {stage2_13[75]},
      {stage3_13[54]}
   );
   gpc1_1 gpc8045 (
      {stage2_13[76]},
      {stage3_13[55]}
   );
   gpc1_1 gpc8046 (
      {stage2_13[77]},
      {stage3_13[56]}
   );
   gpc1_1 gpc8047 (
      {stage2_15[138]},
      {stage3_15[45]}
   );
   gpc1_1 gpc8048 (
      {stage2_15[139]},
      {stage3_15[46]}
   );
   gpc1_1 gpc8049 (
      {stage2_15[140]},
      {stage3_15[47]}
   );
   gpc1_1 gpc8050 (
      {stage2_16[80]},
      {stage3_16[48]}
   );
   gpc1_1 gpc8051 (
      {stage2_16[81]},
      {stage3_16[49]}
   );
   gpc1_1 gpc8052 (
      {stage2_16[82]},
      {stage3_16[50]}
   );
   gpc1_1 gpc8053 (
      {stage2_18[100]},
      {stage3_18[41]}
   );
   gpc1_1 gpc8054 (
      {stage2_18[101]},
      {stage3_18[42]}
   );
   gpc1_1 gpc8055 (
      {stage2_18[102]},
      {stage3_18[43]}
   );
   gpc1_1 gpc8056 (
      {stage2_18[103]},
      {stage3_18[44]}
   );
   gpc1_1 gpc8057 (
      {stage2_18[104]},
      {stage3_18[45]}
   );
   gpc1_1 gpc8058 (
      {stage2_18[105]},
      {stage3_18[46]}
   );
   gpc1_1 gpc8059 (
      {stage2_18[106]},
      {stage3_18[47]}
   );
   gpc1_1 gpc8060 (
      {stage2_18[107]},
      {stage3_18[48]}
   );
   gpc1_1 gpc8061 (
      {stage2_18[108]},
      {stage3_18[49]}
   );
   gpc1_1 gpc8062 (
      {stage2_18[109]},
      {stage3_18[50]}
   );
   gpc1_1 gpc8063 (
      {stage2_18[110]},
      {stage3_18[51]}
   );
   gpc1_1 gpc8064 (
      {stage2_18[111]},
      {stage3_18[52]}
   );
   gpc1_1 gpc8065 (
      {stage2_18[112]},
      {stage3_18[53]}
   );
   gpc1_1 gpc8066 (
      {stage2_18[113]},
      {stage3_18[54]}
   );
   gpc1_1 gpc8067 (
      {stage2_18[114]},
      {stage3_18[55]}
   );
   gpc1_1 gpc8068 (
      {stage2_18[115]},
      {stage3_18[56]}
   );
   gpc1_1 gpc8069 (
      {stage2_18[116]},
      {stage3_18[57]}
   );
   gpc1_1 gpc8070 (
      {stage2_18[117]},
      {stage3_18[58]}
   );
   gpc1_1 gpc8071 (
      {stage2_18[118]},
      {stage3_18[59]}
   );
   gpc1_1 gpc8072 (
      {stage2_20[45]},
      {stage3_20[35]}
   );
   gpc1_1 gpc8073 (
      {stage2_20[46]},
      {stage3_20[36]}
   );
   gpc1_1 gpc8074 (
      {stage2_20[47]},
      {stage3_20[37]}
   );
   gpc1_1 gpc8075 (
      {stage2_20[48]},
      {stage3_20[38]}
   );
   gpc1_1 gpc8076 (
      {stage2_20[49]},
      {stage3_20[39]}
   );
   gpc1_1 gpc8077 (
      {stage2_20[50]},
      {stage3_20[40]}
   );
   gpc1_1 gpc8078 (
      {stage2_20[51]},
      {stage3_20[41]}
   );
   gpc1_1 gpc8079 (
      {stage2_20[52]},
      {stage3_20[42]}
   );
   gpc1_1 gpc8080 (
      {stage2_20[53]},
      {stage3_20[43]}
   );
   gpc1_1 gpc8081 (
      {stage2_20[54]},
      {stage3_20[44]}
   );
   gpc1_1 gpc8082 (
      {stage2_20[55]},
      {stage3_20[45]}
   );
   gpc1_1 gpc8083 (
      {stage2_20[56]},
      {stage3_20[46]}
   );
   gpc1_1 gpc8084 (
      {stage2_20[57]},
      {stage3_20[47]}
   );
   gpc1_1 gpc8085 (
      {stage2_20[58]},
      {stage3_20[48]}
   );
   gpc1_1 gpc8086 (
      {stage2_20[59]},
      {stage3_20[49]}
   );
   gpc1_1 gpc8087 (
      {stage2_20[60]},
      {stage3_20[50]}
   );
   gpc1_1 gpc8088 (
      {stage2_20[61]},
      {stage3_20[51]}
   );
   gpc1_1 gpc8089 (
      {stage2_20[62]},
      {stage3_20[52]}
   );
   gpc1_1 gpc8090 (
      {stage2_20[63]},
      {stage3_20[53]}
   );
   gpc1_1 gpc8091 (
      {stage2_20[64]},
      {stage3_20[54]}
   );
   gpc1_1 gpc8092 (
      {stage2_20[65]},
      {stage3_20[55]}
   );
   gpc1_1 gpc8093 (
      {stage2_20[66]},
      {stage3_20[56]}
   );
   gpc1_1 gpc8094 (
      {stage2_20[67]},
      {stage3_20[57]}
   );
   gpc1_1 gpc8095 (
      {stage2_20[68]},
      {stage3_20[58]}
   );
   gpc1_1 gpc8096 (
      {stage2_20[69]},
      {stage3_20[59]}
   );
   gpc1_1 gpc8097 (
      {stage2_20[70]},
      {stage3_20[60]}
   );
   gpc1_1 gpc8098 (
      {stage2_20[71]},
      {stage3_20[61]}
   );
   gpc1_1 gpc8099 (
      {stage2_20[72]},
      {stage3_20[62]}
   );
   gpc1_1 gpc8100 (
      {stage2_20[73]},
      {stage3_20[63]}
   );
   gpc1_1 gpc8101 (
      {stage2_20[74]},
      {stage3_20[64]}
   );
   gpc1_1 gpc8102 (
      {stage2_20[75]},
      {stage3_20[65]}
   );
   gpc1_1 gpc8103 (
      {stage2_20[76]},
      {stage3_20[66]}
   );
   gpc1_1 gpc8104 (
      {stage2_20[77]},
      {stage3_20[67]}
   );
   gpc1_1 gpc8105 (
      {stage2_20[78]},
      {stage3_20[68]}
   );
   gpc1_1 gpc8106 (
      {stage2_20[79]},
      {stage3_20[69]}
   );
   gpc1_1 gpc8107 (
      {stage2_20[80]},
      {stage3_20[70]}
   );
   gpc1_1 gpc8108 (
      {stage2_20[81]},
      {stage3_20[71]}
   );
   gpc1_1 gpc8109 (
      {stage2_20[82]},
      {stage3_20[72]}
   );
   gpc1_1 gpc8110 (
      {stage2_20[83]},
      {stage3_20[73]}
   );
   gpc1_1 gpc8111 (
      {stage2_20[84]},
      {stage3_20[74]}
   );
   gpc1_1 gpc8112 (
      {stage2_20[85]},
      {stage3_20[75]}
   );
   gpc1_1 gpc8113 (
      {stage2_20[86]},
      {stage3_20[76]}
   );
   gpc1_1 gpc8114 (
      {stage2_20[87]},
      {stage3_20[77]}
   );
   gpc1_1 gpc8115 (
      {stage2_20[88]},
      {stage3_20[78]}
   );
   gpc1_1 gpc8116 (
      {stage2_20[89]},
      {stage3_20[79]}
   );
   gpc1_1 gpc8117 (
      {stage2_20[90]},
      {stage3_20[80]}
   );
   gpc1_1 gpc8118 (
      {stage2_20[91]},
      {stage3_20[81]}
   );
   gpc1_1 gpc8119 (
      {stage2_20[92]},
      {stage3_20[82]}
   );
   gpc1_1 gpc8120 (
      {stage2_21[120]},
      {stage3_21[31]}
   );
   gpc1_1 gpc8121 (
      {stage2_21[121]},
      {stage3_21[32]}
   );
   gpc1_1 gpc8122 (
      {stage2_21[122]},
      {stage3_21[33]}
   );
   gpc1_1 gpc8123 (
      {stage2_21[123]},
      {stage3_21[34]}
   );
   gpc1_1 gpc8124 (
      {stage2_21[124]},
      {stage3_21[35]}
   );
   gpc1_1 gpc8125 (
      {stage2_21[125]},
      {stage3_21[36]}
   );
   gpc1_1 gpc8126 (
      {stage2_21[126]},
      {stage3_21[37]}
   );
   gpc1_1 gpc8127 (
      {stage2_21[127]},
      {stage3_21[38]}
   );
   gpc1_1 gpc8128 (
      {stage2_22[80]},
      {stage3_22[45]}
   );
   gpc1_1 gpc8129 (
      {stage2_22[81]},
      {stage3_22[46]}
   );
   gpc1_1 gpc8130 (
      {stage2_22[82]},
      {stage3_22[47]}
   );
   gpc1_1 gpc8131 (
      {stage2_22[83]},
      {stage3_22[48]}
   );
   gpc1_1 gpc8132 (
      {stage2_22[84]},
      {stage3_22[49]}
   );
   gpc1_1 gpc8133 (
      {stage2_22[85]},
      {stage3_22[50]}
   );
   gpc1_1 gpc8134 (
      {stage2_22[86]},
      {stage3_22[51]}
   );
   gpc1_1 gpc8135 (
      {stage2_22[87]},
      {stage3_22[52]}
   );
   gpc1_1 gpc8136 (
      {stage2_22[88]},
      {stage3_22[53]}
   );
   gpc1_1 gpc8137 (
      {stage2_22[89]},
      {stage3_22[54]}
   );
   gpc1_1 gpc8138 (
      {stage2_22[90]},
      {stage3_22[55]}
   );
   gpc1_1 gpc8139 (
      {stage2_22[91]},
      {stage3_22[56]}
   );
   gpc1_1 gpc8140 (
      {stage2_22[92]},
      {stage3_22[57]}
   );
   gpc1_1 gpc8141 (
      {stage2_22[93]},
      {stage3_22[58]}
   );
   gpc1_1 gpc8142 (
      {stage2_22[94]},
      {stage3_22[59]}
   );
   gpc1_1 gpc8143 (
      {stage2_22[95]},
      {stage3_22[60]}
   );
   gpc1_1 gpc8144 (
      {stage2_22[96]},
      {stage3_22[61]}
   );
   gpc1_1 gpc8145 (
      {stage2_22[97]},
      {stage3_22[62]}
   );
   gpc1_1 gpc8146 (
      {stage2_22[98]},
      {stage3_22[63]}
   );
   gpc1_1 gpc8147 (
      {stage2_22[99]},
      {stage3_22[64]}
   );
   gpc1_1 gpc8148 (
      {stage2_22[100]},
      {stage3_22[65]}
   );
   gpc1_1 gpc8149 (
      {stage2_22[101]},
      {stage3_22[66]}
   );
   gpc1_1 gpc8150 (
      {stage2_22[102]},
      {stage3_22[67]}
   );
   gpc1_1 gpc8151 (
      {stage2_22[103]},
      {stage3_22[68]}
   );
   gpc1_1 gpc8152 (
      {stage2_22[104]},
      {stage3_22[69]}
   );
   gpc1_1 gpc8153 (
      {stage2_22[105]},
      {stage3_22[70]}
   );
   gpc1_1 gpc8154 (
      {stage2_22[106]},
      {stage3_22[71]}
   );
   gpc1_1 gpc8155 (
      {stage2_22[107]},
      {stage3_22[72]}
   );
   gpc1_1 gpc8156 (
      {stage2_26[83]},
      {stage3_26[47]}
   );
   gpc1_1 gpc8157 (
      {stage2_26[84]},
      {stage3_26[48]}
   );
   gpc1_1 gpc8158 (
      {stage2_27[93]},
      {stage3_27[36]}
   );
   gpc1_1 gpc8159 (
      {stage2_27[94]},
      {stage3_27[37]}
   );
   gpc1_1 gpc8160 (
      {stage2_27[95]},
      {stage3_27[38]}
   );
   gpc1_1 gpc8161 (
      {stage2_27[96]},
      {stage3_27[39]}
   );
   gpc1_1 gpc8162 (
      {stage2_27[97]},
      {stage3_27[40]}
   );
   gpc1_1 gpc8163 (
      {stage2_27[98]},
      {stage3_27[41]}
   );
   gpc1_1 gpc8164 (
      {stage2_27[99]},
      {stage3_27[42]}
   );
   gpc1_1 gpc8165 (
      {stage2_27[100]},
      {stage3_27[43]}
   );
   gpc1_1 gpc8166 (
      {stage2_27[101]},
      {stage3_27[44]}
   );
   gpc1_1 gpc8167 (
      {stage2_27[102]},
      {stage3_27[45]}
   );
   gpc1_1 gpc8168 (
      {stage2_27[103]},
      {stage3_27[46]}
   );
   gpc1_1 gpc8169 (
      {stage2_27[104]},
      {stage3_27[47]}
   );
   gpc1_1 gpc8170 (
      {stage2_27[105]},
      {stage3_27[48]}
   );
   gpc1_1 gpc8171 (
      {stage2_28[69]},
      {stage3_28[34]}
   );
   gpc1_1 gpc8172 (
      {stage2_28[70]},
      {stage3_28[35]}
   );
   gpc1_1 gpc8173 (
      {stage2_28[71]},
      {stage3_28[36]}
   );
   gpc1_1 gpc8174 (
      {stage2_28[72]},
      {stage3_28[37]}
   );
   gpc1_1 gpc8175 (
      {stage2_28[73]},
      {stage3_28[38]}
   );
   gpc1_1 gpc8176 (
      {stage2_28[74]},
      {stage3_28[39]}
   );
   gpc1_1 gpc8177 (
      {stage2_28[75]},
      {stage3_28[40]}
   );
   gpc1_1 gpc8178 (
      {stage2_28[76]},
      {stage3_28[41]}
   );
   gpc1_1 gpc8179 (
      {stage2_28[77]},
      {stage3_28[42]}
   );
   gpc1_1 gpc8180 (
      {stage2_28[78]},
      {stage3_28[43]}
   );
   gpc1_1 gpc8181 (
      {stage2_28[79]},
      {stage3_28[44]}
   );
   gpc1_1 gpc8182 (
      {stage2_28[80]},
      {stage3_28[45]}
   );
   gpc1_1 gpc8183 (
      {stage2_28[81]},
      {stage3_28[46]}
   );
   gpc1_1 gpc8184 (
      {stage2_28[82]},
      {stage3_28[47]}
   );
   gpc1_1 gpc8185 (
      {stage2_28[83]},
      {stage3_28[48]}
   );
   gpc1_1 gpc8186 (
      {stage2_28[84]},
      {stage3_28[49]}
   );
   gpc1_1 gpc8187 (
      {stage2_28[85]},
      {stage3_28[50]}
   );
   gpc1_1 gpc8188 (
      {stage2_28[86]},
      {stage3_28[51]}
   );
   gpc1_1 gpc8189 (
      {stage2_28[87]},
      {stage3_28[52]}
   );
   gpc1_1 gpc8190 (
      {stage2_28[88]},
      {stage3_28[53]}
   );
   gpc1_1 gpc8191 (
      {stage2_28[89]},
      {stage3_28[54]}
   );
   gpc1_1 gpc8192 (
      {stage2_28[90]},
      {stage3_28[55]}
   );
   gpc1_1 gpc8193 (
      {stage2_28[91]},
      {stage3_28[56]}
   );
   gpc1_1 gpc8194 (
      {stage2_30[103]},
      {stage3_30[28]}
   );
   gpc1_1 gpc8195 (
      {stage2_30[104]},
      {stage3_30[29]}
   );
   gpc1_1 gpc8196 (
      {stage2_30[105]},
      {stage3_30[30]}
   );
   gpc1_1 gpc8197 (
      {stage2_30[106]},
      {stage3_30[31]}
   );
   gpc1_1 gpc8198 (
      {stage2_30[107]},
      {stage3_30[32]}
   );
   gpc1_1 gpc8199 (
      {stage2_30[108]},
      {stage3_30[33]}
   );
   gpc1_1 gpc8200 (
      {stage2_30[109]},
      {stage3_30[34]}
   );
   gpc1_1 gpc8201 (
      {stage2_30[110]},
      {stage3_30[35]}
   );
   gpc1_1 gpc8202 (
      {stage2_30[111]},
      {stage3_30[36]}
   );
   gpc1_1 gpc8203 (
      {stage2_30[112]},
      {stage3_30[37]}
   );
   gpc1_1 gpc8204 (
      {stage2_30[113]},
      {stage3_30[38]}
   );
   gpc1_1 gpc8205 (
      {stage2_30[114]},
      {stage3_30[39]}
   );
   gpc1_1 gpc8206 (
      {stage2_30[115]},
      {stage3_30[40]}
   );
   gpc1_1 gpc8207 (
      {stage2_30[116]},
      {stage3_30[41]}
   );
   gpc1_1 gpc8208 (
      {stage2_31[95]},
      {stage3_31[34]}
   );
   gpc1_1 gpc8209 (
      {stage2_31[96]},
      {stage3_31[35]}
   );
   gpc1_1 gpc8210 (
      {stage2_31[97]},
      {stage3_31[36]}
   );
   gpc1_1 gpc8211 (
      {stage2_31[98]},
      {stage3_31[37]}
   );
   gpc1_1 gpc8212 (
      {stage2_32[99]},
      {stage3_32[47]}
   );
   gpc1_1 gpc8213 (
      {stage2_32[100]},
      {stage3_32[48]}
   );
   gpc1_1 gpc8214 (
      {stage2_32[101]},
      {stage3_32[49]}
   );
   gpc1_1 gpc8215 (
      {stage2_32[102]},
      {stage3_32[50]}
   );
   gpc1_1 gpc8216 (
      {stage2_32[103]},
      {stage3_32[51]}
   );
   gpc1_1 gpc8217 (
      {stage2_32[104]},
      {stage3_32[52]}
   );
   gpc1_1 gpc8218 (
      {stage2_32[105]},
      {stage3_32[53]}
   );
   gpc1_1 gpc8219 (
      {stage2_33[72]},
      {stage3_33[42]}
   );
   gpc1_1 gpc8220 (
      {stage2_33[73]},
      {stage3_33[43]}
   );
   gpc1_1 gpc8221 (
      {stage2_33[74]},
      {stage3_33[44]}
   );
   gpc1_1 gpc8222 (
      {stage2_33[75]},
      {stage3_33[45]}
   );
   gpc1_1 gpc8223 (
      {stage2_34[129]},
      {stage3_34[39]}
   );
   gpc1_1 gpc8224 (
      {stage2_34[130]},
      {stage3_34[40]}
   );
   gpc1_1 gpc8225 (
      {stage2_34[131]},
      {stage3_34[41]}
   );
   gpc1_1 gpc8226 (
      {stage2_35[120]},
      {stage3_35[44]}
   );
   gpc1_1 gpc8227 (
      {stage2_35[121]},
      {stage3_35[45]}
   );
   gpc1_1 gpc8228 (
      {stage2_35[122]},
      {stage3_35[46]}
   );
   gpc1_1 gpc8229 (
      {stage2_35[123]},
      {stage3_35[47]}
   );
   gpc1_1 gpc8230 (
      {stage2_35[124]},
      {stage3_35[48]}
   );
   gpc1_1 gpc8231 (
      {stage2_35[125]},
      {stage3_35[49]}
   );
   gpc1_1 gpc8232 (
      {stage2_35[126]},
      {stage3_35[50]}
   );
   gpc1_1 gpc8233 (
      {stage2_35[127]},
      {stage3_35[51]}
   );
   gpc1_1 gpc8234 (
      {stage2_35[128]},
      {stage3_35[52]}
   );
   gpc1_1 gpc8235 (
      {stage2_35[129]},
      {stage3_35[53]}
   );
   gpc1_1 gpc8236 (
      {stage2_35[130]},
      {stage3_35[54]}
   );
   gpc1_1 gpc8237 (
      {stage2_35[131]},
      {stage3_35[55]}
   );
   gpc1_1 gpc8238 (
      {stage2_35[132]},
      {stage3_35[56]}
   );
   gpc1_1 gpc8239 (
      {stage2_36[73]},
      {stage3_36[44]}
   );
   gpc1_1 gpc8240 (
      {stage2_36[74]},
      {stage3_36[45]}
   );
   gpc1_1 gpc8241 (
      {stage2_37[74]},
      {stage3_37[37]}
   );
   gpc1_1 gpc8242 (
      {stage2_37[75]},
      {stage3_37[38]}
   );
   gpc1_1 gpc8243 (
      {stage2_37[76]},
      {stage3_37[39]}
   );
   gpc1_1 gpc8244 (
      {stage2_37[77]},
      {stage3_37[40]}
   );
   gpc1_1 gpc8245 (
      {stage2_37[78]},
      {stage3_37[41]}
   );
   gpc1_1 gpc8246 (
      {stage2_37[79]},
      {stage3_37[42]}
   );
   gpc1_1 gpc8247 (
      {stage2_37[80]},
      {stage3_37[43]}
   );
   gpc1_1 gpc8248 (
      {stage2_37[81]},
      {stage3_37[44]}
   );
   gpc1_1 gpc8249 (
      {stage2_37[82]},
      {stage3_37[45]}
   );
   gpc1_1 gpc8250 (
      {stage2_37[83]},
      {stage3_37[46]}
   );
   gpc1_1 gpc8251 (
      {stage2_37[84]},
      {stage3_37[47]}
   );
   gpc1_1 gpc8252 (
      {stage2_37[85]},
      {stage3_37[48]}
   );
   gpc1_1 gpc8253 (
      {stage2_37[86]},
      {stage3_37[49]}
   );
   gpc1_1 gpc8254 (
      {stage2_37[87]},
      {stage3_37[50]}
   );
   gpc1_1 gpc8255 (
      {stage2_37[88]},
      {stage3_37[51]}
   );
   gpc1_1 gpc8256 (
      {stage2_37[89]},
      {stage3_37[52]}
   );
   gpc1_1 gpc8257 (
      {stage2_38[125]},
      {stage3_38[45]}
   );
   gpc1_1 gpc8258 (
      {stage2_38[126]},
      {stage3_38[46]}
   );
   gpc1_1 gpc8259 (
      {stage2_38[127]},
      {stage3_38[47]}
   );
   gpc1_1 gpc8260 (
      {stage2_38[128]},
      {stage3_38[48]}
   );
   gpc1_1 gpc8261 (
      {stage2_38[129]},
      {stage3_38[49]}
   );
   gpc1_1 gpc8262 (
      {stage2_38[130]},
      {stage3_38[50]}
   );
   gpc1_1 gpc8263 (
      {stage2_38[131]},
      {stage3_38[51]}
   );
   gpc1_1 gpc8264 (
      {stage2_38[132]},
      {stage3_38[52]}
   );
   gpc1_1 gpc8265 (
      {stage2_38[133]},
      {stage3_38[53]}
   );
   gpc1_1 gpc8266 (
      {stage2_38[134]},
      {stage3_38[54]}
   );
   gpc1_1 gpc8267 (
      {stage2_38[135]},
      {stage3_38[55]}
   );
   gpc1_1 gpc8268 (
      {stage2_38[136]},
      {stage3_38[56]}
   );
   gpc1_1 gpc8269 (
      {stage2_38[137]},
      {stage3_38[57]}
   );
   gpc1_1 gpc8270 (
      {stage2_38[138]},
      {stage3_38[58]}
   );
   gpc1_1 gpc8271 (
      {stage2_38[139]},
      {stage3_38[59]}
   );
   gpc1_1 gpc8272 (
      {stage2_39[128]},
      {stage3_39[49]}
   );
   gpc1_1 gpc8273 (
      {stage2_39[129]},
      {stage3_39[50]}
   );
   gpc1_1 gpc8274 (
      {stage2_39[130]},
      {stage3_39[51]}
   );
   gpc1_1 gpc8275 (
      {stage2_39[131]},
      {stage3_39[52]}
   );
   gpc1_1 gpc8276 (
      {stage2_39[132]},
      {stage3_39[53]}
   );
   gpc1_1 gpc8277 (
      {stage2_39[133]},
      {stage3_39[54]}
   );
   gpc1_1 gpc8278 (
      {stage2_39[134]},
      {stage3_39[55]}
   );
   gpc1_1 gpc8279 (
      {stage2_39[135]},
      {stage3_39[56]}
   );
   gpc1_1 gpc8280 (
      {stage2_39[136]},
      {stage3_39[57]}
   );
   gpc1_1 gpc8281 (
      {stage2_40[107]},
      {stage3_40[46]}
   );
   gpc1_1 gpc8282 (
      {stage2_40[108]},
      {stage3_40[47]}
   );
   gpc1_1 gpc8283 (
      {stage2_40[109]},
      {stage3_40[48]}
   );
   gpc1_1 gpc8284 (
      {stage2_40[110]},
      {stage3_40[49]}
   );
   gpc1_1 gpc8285 (
      {stage2_40[111]},
      {stage3_40[50]}
   );
   gpc1_1 gpc8286 (
      {stage2_40[112]},
      {stage3_40[51]}
   );
   gpc1_1 gpc8287 (
      {stage2_41[102]},
      {stage3_41[39]}
   );
   gpc1_1 gpc8288 (
      {stage2_41[103]},
      {stage3_41[40]}
   );
   gpc1_1 gpc8289 (
      {stage2_41[104]},
      {stage3_41[41]}
   );
   gpc1_1 gpc8290 (
      {stage2_41[105]},
      {stage3_41[42]}
   );
   gpc1_1 gpc8291 (
      {stage2_42[82]},
      {stage3_42[46]}
   );
   gpc1_1 gpc8292 (
      {stage2_42[83]},
      {stage3_42[47]}
   );
   gpc1_1 gpc8293 (
      {stage2_42[84]},
      {stage3_42[48]}
   );
   gpc1_1 gpc8294 (
      {stage2_42[85]},
      {stage3_42[49]}
   );
   gpc1_1 gpc8295 (
      {stage2_44[109]},
      {stage3_44[31]}
   );
   gpc1_1 gpc8296 (
      {stage2_44[110]},
      {stage3_44[32]}
   );
   gpc1_1 gpc8297 (
      {stage2_44[111]},
      {stage3_44[33]}
   );
   gpc1_1 gpc8298 (
      {stage2_44[112]},
      {stage3_44[34]}
   );
   gpc1_1 gpc8299 (
      {stage2_44[113]},
      {stage3_44[35]}
   );
   gpc1_1 gpc8300 (
      {stage2_44[114]},
      {stage3_44[36]}
   );
   gpc1_1 gpc8301 (
      {stage2_44[115]},
      {stage3_44[37]}
   );
   gpc1_1 gpc8302 (
      {stage2_44[116]},
      {stage3_44[38]}
   );
   gpc1_1 gpc8303 (
      {stage2_44[117]},
      {stage3_44[39]}
   );
   gpc1_1 gpc8304 (
      {stage2_44[118]},
      {stage3_44[40]}
   );
   gpc1_1 gpc8305 (
      {stage2_45[108]},
      {stage3_45[34]}
   );
   gpc1_1 gpc8306 (
      {stage2_45[109]},
      {stage3_45[35]}
   );
   gpc1_1 gpc8307 (
      {stage2_45[110]},
      {stage3_45[36]}
   );
   gpc1_1 gpc8308 (
      {stage2_45[111]},
      {stage3_45[37]}
   );
   gpc1_1 gpc8309 (
      {stage2_45[112]},
      {stage3_45[38]}
   );
   gpc1_1 gpc8310 (
      {stage2_45[113]},
      {stage3_45[39]}
   );
   gpc1_1 gpc8311 (
      {stage2_45[114]},
      {stage3_45[40]}
   );
   gpc1_1 gpc8312 (
      {stage2_45[115]},
      {stage3_45[41]}
   );
   gpc1_1 gpc8313 (
      {stage2_45[116]},
      {stage3_45[42]}
   );
   gpc1_1 gpc8314 (
      {stage2_45[117]},
      {stage3_45[43]}
   );
   gpc1_1 gpc8315 (
      {stage2_46[78]},
      {stage3_46[48]}
   );
   gpc1_1 gpc8316 (
      {stage2_46[79]},
      {stage3_46[49]}
   );
   gpc1_1 gpc8317 (
      {stage2_46[80]},
      {stage3_46[50]}
   );
   gpc1_1 gpc8318 (
      {stage2_46[81]},
      {stage3_46[51]}
   );
   gpc1_1 gpc8319 (
      {stage2_46[82]},
      {stage3_46[52]}
   );
   gpc1_1 gpc8320 (
      {stage2_46[83]},
      {stage3_46[53]}
   );
   gpc1_1 gpc8321 (
      {stage2_46[84]},
      {stage3_46[54]}
   );
   gpc1_1 gpc8322 (
      {stage2_46[85]},
      {stage3_46[55]}
   );
   gpc1_1 gpc8323 (
      {stage2_46[86]},
      {stage3_46[56]}
   );
   gpc1_1 gpc8324 (
      {stage2_46[87]},
      {stage3_46[57]}
   );
   gpc1_1 gpc8325 (
      {stage2_48[126]},
      {stage3_48[38]}
   );
   gpc1_1 gpc8326 (
      {stage2_48[127]},
      {stage3_48[39]}
   );
   gpc1_1 gpc8327 (
      {stage2_48[128]},
      {stage3_48[40]}
   );
   gpc1_1 gpc8328 (
      {stage2_48[129]},
      {stage3_48[41]}
   );
   gpc1_1 gpc8329 (
      {stage2_50[84]},
      {stage3_50[45]}
   );
   gpc1_1 gpc8330 (
      {stage2_50[85]},
      {stage3_50[46]}
   );
   gpc1_1 gpc8331 (
      {stage2_51[59]},
      {stage3_51[34]}
   );
   gpc1_1 gpc8332 (
      {stage2_51[60]},
      {stage3_51[35]}
   );
   gpc1_1 gpc8333 (
      {stage2_51[61]},
      {stage3_51[36]}
   );
   gpc1_1 gpc8334 (
      {stage2_51[62]},
      {stage3_51[37]}
   );
   gpc1_1 gpc8335 (
      {stage2_51[63]},
      {stage3_51[38]}
   );
   gpc1_1 gpc8336 (
      {stage2_51[64]},
      {stage3_51[39]}
   );
   gpc1_1 gpc8337 (
      {stage2_51[65]},
      {stage3_51[40]}
   );
   gpc1_1 gpc8338 (
      {stage2_51[66]},
      {stage3_51[41]}
   );
   gpc1_1 gpc8339 (
      {stage2_51[67]},
      {stage3_51[42]}
   );
   gpc1_1 gpc8340 (
      {stage2_51[68]},
      {stage3_51[43]}
   );
   gpc1_1 gpc8341 (
      {stage2_51[69]},
      {stage3_51[44]}
   );
   gpc1_1 gpc8342 (
      {stage2_51[70]},
      {stage3_51[45]}
   );
   gpc1_1 gpc8343 (
      {stage2_51[71]},
      {stage3_51[46]}
   );
   gpc1_1 gpc8344 (
      {stage2_51[72]},
      {stage3_51[47]}
   );
   gpc1_1 gpc8345 (
      {stage2_51[73]},
      {stage3_51[48]}
   );
   gpc1_1 gpc8346 (
      {stage2_51[74]},
      {stage3_51[49]}
   );
   gpc1_1 gpc8347 (
      {stage2_51[75]},
      {stage3_51[50]}
   );
   gpc1_1 gpc8348 (
      {stage2_51[76]},
      {stage3_51[51]}
   );
   gpc1_1 gpc8349 (
      {stage2_51[77]},
      {stage3_51[52]}
   );
   gpc1_1 gpc8350 (
      {stage2_51[78]},
      {stage3_51[53]}
   );
   gpc1_1 gpc8351 (
      {stage2_51[79]},
      {stage3_51[54]}
   );
   gpc1_1 gpc8352 (
      {stage2_51[80]},
      {stage3_51[55]}
   );
   gpc1_1 gpc8353 (
      {stage2_51[81]},
      {stage3_51[56]}
   );
   gpc1_1 gpc8354 (
      {stage2_51[82]},
      {stage3_51[57]}
   );
   gpc1_1 gpc8355 (
      {stage2_51[83]},
      {stage3_51[58]}
   );
   gpc1_1 gpc8356 (
      {stage2_51[84]},
      {stage3_51[59]}
   );
   gpc1_1 gpc8357 (
      {stage2_51[85]},
      {stage3_51[60]}
   );
   gpc1_1 gpc8358 (
      {stage2_51[86]},
      {stage3_51[61]}
   );
   gpc1_1 gpc8359 (
      {stage2_51[87]},
      {stage3_51[62]}
   );
   gpc1_1 gpc8360 (
      {stage2_52[69]},
      {stage3_52[27]}
   );
   gpc1_1 gpc8361 (
      {stage2_52[70]},
      {stage3_52[28]}
   );
   gpc1_1 gpc8362 (
      {stage2_52[71]},
      {stage3_52[29]}
   );
   gpc1_1 gpc8363 (
      {stage2_52[72]},
      {stage3_52[30]}
   );
   gpc1_1 gpc8364 (
      {stage2_52[73]},
      {stage3_52[31]}
   );
   gpc1_1 gpc8365 (
      {stage2_52[74]},
      {stage3_52[32]}
   );
   gpc1_1 gpc8366 (
      {stage2_52[75]},
      {stage3_52[33]}
   );
   gpc1_1 gpc8367 (
      {stage2_52[76]},
      {stage3_52[34]}
   );
   gpc1_1 gpc8368 (
      {stage2_52[77]},
      {stage3_52[35]}
   );
   gpc1_1 gpc8369 (
      {stage2_52[78]},
      {stage3_52[36]}
   );
   gpc1_1 gpc8370 (
      {stage2_52[79]},
      {stage3_52[37]}
   );
   gpc1_1 gpc8371 (
      {stage2_52[80]},
      {stage3_52[38]}
   );
   gpc1_1 gpc8372 (
      {stage2_52[81]},
      {stage3_52[39]}
   );
   gpc1_1 gpc8373 (
      {stage2_52[82]},
      {stage3_52[40]}
   );
   gpc1_1 gpc8374 (
      {stage2_52[83]},
      {stage3_52[41]}
   );
   gpc1_1 gpc8375 (
      {stage2_52[84]},
      {stage3_52[42]}
   );
   gpc1_1 gpc8376 (
      {stage2_52[85]},
      {stage3_52[43]}
   );
   gpc1_1 gpc8377 (
      {stage2_52[86]},
      {stage3_52[44]}
   );
   gpc1_1 gpc8378 (
      {stage2_52[87]},
      {stage3_52[45]}
   );
   gpc1_1 gpc8379 (
      {stage2_52[88]},
      {stage3_52[46]}
   );
   gpc1_1 gpc8380 (
      {stage2_52[89]},
      {stage3_52[47]}
   );
   gpc1_1 gpc8381 (
      {stage2_52[90]},
      {stage3_52[48]}
   );
   gpc1_1 gpc8382 (
      {stage2_52[91]},
      {stage3_52[49]}
   );
   gpc1_1 gpc8383 (
      {stage2_52[92]},
      {stage3_52[50]}
   );
   gpc1_1 gpc8384 (
      {stage2_52[93]},
      {stage3_52[51]}
   );
   gpc1_1 gpc8385 (
      {stage2_52[94]},
      {stage3_52[52]}
   );
   gpc1_1 gpc8386 (
      {stage2_52[95]},
      {stage3_52[53]}
   );
   gpc1_1 gpc8387 (
      {stage2_52[96]},
      {stage3_52[54]}
   );
   gpc1_1 gpc8388 (
      {stage2_52[97]},
      {stage3_52[55]}
   );
   gpc1_1 gpc8389 (
      {stage2_52[98]},
      {stage3_52[56]}
   );
   gpc1_1 gpc8390 (
      {stage2_52[99]},
      {stage3_52[57]}
   );
   gpc1_1 gpc8391 (
      {stage2_52[100]},
      {stage3_52[58]}
   );
   gpc1_1 gpc8392 (
      {stage2_52[101]},
      {stage3_52[59]}
   );
   gpc1_1 gpc8393 (
      {stage2_52[102]},
      {stage3_52[60]}
   );
   gpc1_1 gpc8394 (
      {stage2_52[103]},
      {stage3_52[61]}
   );
   gpc1_1 gpc8395 (
      {stage2_52[104]},
      {stage3_52[62]}
   );
   gpc1_1 gpc8396 (
      {stage2_53[69]},
      {stage3_53[29]}
   );
   gpc1_1 gpc8397 (
      {stage2_53[70]},
      {stage3_53[30]}
   );
   gpc1_1 gpc8398 (
      {stage2_53[71]},
      {stage3_53[31]}
   );
   gpc1_1 gpc8399 (
      {stage2_53[72]},
      {stage3_53[32]}
   );
   gpc1_1 gpc8400 (
      {stage2_53[73]},
      {stage3_53[33]}
   );
   gpc1_1 gpc8401 (
      {stage2_53[74]},
      {stage3_53[34]}
   );
   gpc1_1 gpc8402 (
      {stage2_53[75]},
      {stage3_53[35]}
   );
   gpc1_1 gpc8403 (
      {stage2_53[76]},
      {stage3_53[36]}
   );
   gpc1_1 gpc8404 (
      {stage2_53[77]},
      {stage3_53[37]}
   );
   gpc1_1 gpc8405 (
      {stage2_53[78]},
      {stage3_53[38]}
   );
   gpc1_1 gpc8406 (
      {stage2_53[79]},
      {stage3_53[39]}
   );
   gpc1_1 gpc8407 (
      {stage2_53[80]},
      {stage3_53[40]}
   );
   gpc1_1 gpc8408 (
      {stage2_53[81]},
      {stage3_53[41]}
   );
   gpc1_1 gpc8409 (
      {stage2_53[82]},
      {stage3_53[42]}
   );
   gpc1_1 gpc8410 (
      {stage2_53[83]},
      {stage3_53[43]}
   );
   gpc1_1 gpc8411 (
      {stage2_53[84]},
      {stage3_53[44]}
   );
   gpc1_1 gpc8412 (
      {stage2_53[85]},
      {stage3_53[45]}
   );
   gpc1_1 gpc8413 (
      {stage2_53[86]},
      {stage3_53[46]}
   );
   gpc1_1 gpc8414 (
      {stage2_53[87]},
      {stage3_53[47]}
   );
   gpc1_1 gpc8415 (
      {stage2_53[88]},
      {stage3_53[48]}
   );
   gpc1_1 gpc8416 (
      {stage2_53[89]},
      {stage3_53[49]}
   );
   gpc1_1 gpc8417 (
      {stage2_53[90]},
      {stage3_53[50]}
   );
   gpc1_1 gpc8418 (
      {stage2_53[91]},
      {stage3_53[51]}
   );
   gpc1_1 gpc8419 (
      {stage2_53[92]},
      {stage3_53[52]}
   );
   gpc1_1 gpc8420 (
      {stage2_53[93]},
      {stage3_53[53]}
   );
   gpc1_1 gpc8421 (
      {stage2_53[94]},
      {stage3_53[54]}
   );
   gpc1_1 gpc8422 (
      {stage2_53[95]},
      {stage3_53[55]}
   );
   gpc1_1 gpc8423 (
      {stage2_53[96]},
      {stage3_53[56]}
   );
   gpc1_1 gpc8424 (
      {stage2_53[97]},
      {stage3_53[57]}
   );
   gpc1_1 gpc8425 (
      {stage2_53[98]},
      {stage3_53[58]}
   );
   gpc1_1 gpc8426 (
      {stage2_53[99]},
      {stage3_53[59]}
   );
   gpc1_1 gpc8427 (
      {stage2_53[100]},
      {stage3_53[60]}
   );
   gpc1_1 gpc8428 (
      {stage2_53[101]},
      {stage3_53[61]}
   );
   gpc1_1 gpc8429 (
      {stage2_53[102]},
      {stage3_53[62]}
   );
   gpc1_1 gpc8430 (
      {stage2_53[103]},
      {stage3_53[63]}
   );
   gpc1_1 gpc8431 (
      {stage2_53[104]},
      {stage3_53[64]}
   );
   gpc1_1 gpc8432 (
      {stage2_53[105]},
      {stage3_53[65]}
   );
   gpc1_1 gpc8433 (
      {stage2_53[106]},
      {stage3_53[66]}
   );
   gpc1_1 gpc8434 (
      {stage2_53[107]},
      {stage3_53[67]}
   );
   gpc1_1 gpc8435 (
      {stage2_53[108]},
      {stage3_53[68]}
   );
   gpc1_1 gpc8436 (
      {stage2_53[109]},
      {stage3_53[69]}
   );
   gpc1_1 gpc8437 (
      {stage2_53[110]},
      {stage3_53[70]}
   );
   gpc1_1 gpc8438 (
      {stage2_53[111]},
      {stage3_53[71]}
   );
   gpc1_1 gpc8439 (
      {stage2_53[112]},
      {stage3_53[72]}
   );
   gpc1_1 gpc8440 (
      {stage2_53[113]},
      {stage3_53[73]}
   );
   gpc1_1 gpc8441 (
      {stage2_53[114]},
      {stage3_53[74]}
   );
   gpc1_1 gpc8442 (
      {stage2_55[70]},
      {stage3_55[31]}
   );
   gpc1_1 gpc8443 (
      {stage2_55[71]},
      {stage3_55[32]}
   );
   gpc1_1 gpc8444 (
      {stage2_55[72]},
      {stage3_55[33]}
   );
   gpc1_1 gpc8445 (
      {stage2_55[73]},
      {stage3_55[34]}
   );
   gpc1_1 gpc8446 (
      {stage2_55[74]},
      {stage3_55[35]}
   );
   gpc1_1 gpc8447 (
      {stage2_55[75]},
      {stage3_55[36]}
   );
   gpc1_1 gpc8448 (
      {stage2_55[76]},
      {stage3_55[37]}
   );
   gpc1_1 gpc8449 (
      {stage2_55[77]},
      {stage3_55[38]}
   );
   gpc1_1 gpc8450 (
      {stage2_55[78]},
      {stage3_55[39]}
   );
   gpc1_1 gpc8451 (
      {stage2_55[79]},
      {stage3_55[40]}
   );
   gpc1_1 gpc8452 (
      {stage2_55[80]},
      {stage3_55[41]}
   );
   gpc1_1 gpc8453 (
      {stage2_55[81]},
      {stage3_55[42]}
   );
   gpc1_1 gpc8454 (
      {stage2_55[82]},
      {stage3_55[43]}
   );
   gpc1_1 gpc8455 (
      {stage2_55[83]},
      {stage3_55[44]}
   );
   gpc1_1 gpc8456 (
      {stage2_55[84]},
      {stage3_55[45]}
   );
   gpc1_1 gpc8457 (
      {stage2_55[85]},
      {stage3_55[46]}
   );
   gpc1_1 gpc8458 (
      {stage2_55[86]},
      {stage3_55[47]}
   );
   gpc1_1 gpc8459 (
      {stage2_55[87]},
      {stage3_55[48]}
   );
   gpc1_1 gpc8460 (
      {stage2_55[88]},
      {stage3_55[49]}
   );
   gpc1_1 gpc8461 (
      {stage2_55[89]},
      {stage3_55[50]}
   );
   gpc1_1 gpc8462 (
      {stage2_55[90]},
      {stage3_55[51]}
   );
   gpc1_1 gpc8463 (
      {stage2_55[91]},
      {stage3_55[52]}
   );
   gpc1_1 gpc8464 (
      {stage2_55[92]},
      {stage3_55[53]}
   );
   gpc1_1 gpc8465 (
      {stage2_55[93]},
      {stage3_55[54]}
   );
   gpc1_1 gpc8466 (
      {stage2_55[94]},
      {stage3_55[55]}
   );
   gpc1_1 gpc8467 (
      {stage2_55[95]},
      {stage3_55[56]}
   );
   gpc1_1 gpc8468 (
      {stage2_55[96]},
      {stage3_55[57]}
   );
   gpc1_1 gpc8469 (
      {stage2_55[97]},
      {stage3_55[58]}
   );
   gpc1_1 gpc8470 (
      {stage2_55[98]},
      {stage3_55[59]}
   );
   gpc1_1 gpc8471 (
      {stage2_55[99]},
      {stage3_55[60]}
   );
   gpc1_1 gpc8472 (
      {stage2_55[100]},
      {stage3_55[61]}
   );
   gpc1_1 gpc8473 (
      {stage2_55[101]},
      {stage3_55[62]}
   );
   gpc1_1 gpc8474 (
      {stage2_55[102]},
      {stage3_55[63]}
   );
   gpc1_1 gpc8475 (
      {stage2_55[103]},
      {stage3_55[64]}
   );
   gpc1_1 gpc8476 (
      {stage2_55[104]},
      {stage3_55[65]}
   );
   gpc1_1 gpc8477 (
      {stage2_55[105]},
      {stage3_55[66]}
   );
   gpc1_1 gpc8478 (
      {stage2_57[49]},
      {stage3_57[37]}
   );
   gpc1_1 gpc8479 (
      {stage2_57[50]},
      {stage3_57[38]}
   );
   gpc1_1 gpc8480 (
      {stage2_57[51]},
      {stage3_57[39]}
   );
   gpc1_1 gpc8481 (
      {stage2_57[52]},
      {stage3_57[40]}
   );
   gpc1_1 gpc8482 (
      {stage2_57[53]},
      {stage3_57[41]}
   );
   gpc1_1 gpc8483 (
      {stage2_57[54]},
      {stage3_57[42]}
   );
   gpc1_1 gpc8484 (
      {stage2_57[55]},
      {stage3_57[43]}
   );
   gpc1_1 gpc8485 (
      {stage2_57[56]},
      {stage3_57[44]}
   );
   gpc1_1 gpc8486 (
      {stage2_57[57]},
      {stage3_57[45]}
   );
   gpc1_1 gpc8487 (
      {stage2_57[58]},
      {stage3_57[46]}
   );
   gpc1_1 gpc8488 (
      {stage2_57[59]},
      {stage3_57[47]}
   );
   gpc1_1 gpc8489 (
      {stage2_57[60]},
      {stage3_57[48]}
   );
   gpc1_1 gpc8490 (
      {stage2_57[61]},
      {stage3_57[49]}
   );
   gpc1_1 gpc8491 (
      {stage2_57[62]},
      {stage3_57[50]}
   );
   gpc1_1 gpc8492 (
      {stage2_57[63]},
      {stage3_57[51]}
   );
   gpc1_1 gpc8493 (
      {stage2_57[64]},
      {stage3_57[52]}
   );
   gpc1_1 gpc8494 (
      {stage2_57[65]},
      {stage3_57[53]}
   );
   gpc1_1 gpc8495 (
      {stage2_58[58]},
      {stage3_58[34]}
   );
   gpc1_1 gpc8496 (
      {stage2_58[59]},
      {stage3_58[35]}
   );
   gpc1_1 gpc8497 (
      {stage2_58[60]},
      {stage3_58[36]}
   );
   gpc1_1 gpc8498 (
      {stage2_58[61]},
      {stage3_58[37]}
   );
   gpc1_1 gpc8499 (
      {stage2_58[62]},
      {stage3_58[38]}
   );
   gpc1_1 gpc8500 (
      {stage2_58[63]},
      {stage3_58[39]}
   );
   gpc1_1 gpc8501 (
      {stage2_58[64]},
      {stage3_58[40]}
   );
   gpc1_1 gpc8502 (
      {stage2_58[65]},
      {stage3_58[41]}
   );
   gpc1_1 gpc8503 (
      {stage2_58[66]},
      {stage3_58[42]}
   );
   gpc1_1 gpc8504 (
      {stage2_58[67]},
      {stage3_58[43]}
   );
   gpc1_1 gpc8505 (
      {stage2_58[68]},
      {stage3_58[44]}
   );
   gpc1_1 gpc8506 (
      {stage2_58[69]},
      {stage3_58[45]}
   );
   gpc1_1 gpc8507 (
      {stage2_58[70]},
      {stage3_58[46]}
   );
   gpc1_1 gpc8508 (
      {stage2_58[71]},
      {stage3_58[47]}
   );
   gpc1_1 gpc8509 (
      {stage2_58[72]},
      {stage3_58[48]}
   );
   gpc1_1 gpc8510 (
      {stage2_58[73]},
      {stage3_58[49]}
   );
   gpc1_1 gpc8511 (
      {stage2_58[74]},
      {stage3_58[50]}
   );
   gpc1_1 gpc8512 (
      {stage2_58[75]},
      {stage3_58[51]}
   );
   gpc1_1 gpc8513 (
      {stage2_58[76]},
      {stage3_58[52]}
   );
   gpc1_1 gpc8514 (
      {stage2_58[77]},
      {stage3_58[53]}
   );
   gpc1_1 gpc8515 (
      {stage2_58[78]},
      {stage3_58[54]}
   );
   gpc1_1 gpc8516 (
      {stage2_58[79]},
      {stage3_58[55]}
   );
   gpc1_1 gpc8517 (
      {stage2_58[80]},
      {stage3_58[56]}
   );
   gpc1_1 gpc8518 (
      {stage2_58[81]},
      {stage3_58[57]}
   );
   gpc1_1 gpc8519 (
      {stage2_58[82]},
      {stage3_58[58]}
   );
   gpc1_1 gpc8520 (
      {stage2_58[83]},
      {stage3_58[59]}
   );
   gpc1_1 gpc8521 (
      {stage2_58[84]},
      {stage3_58[60]}
   );
   gpc1_1 gpc8522 (
      {stage2_58[85]},
      {stage3_58[61]}
   );
   gpc1_1 gpc8523 (
      {stage2_59[85]},
      {stage3_59[25]}
   );
   gpc1_1 gpc8524 (
      {stage2_59[86]},
      {stage3_59[26]}
   );
   gpc1_1 gpc8525 (
      {stage2_59[87]},
      {stage3_59[27]}
   );
   gpc1_1 gpc8526 (
      {stage2_59[88]},
      {stage3_59[28]}
   );
   gpc1_1 gpc8527 (
      {stage2_59[89]},
      {stage3_59[29]}
   );
   gpc1_1 gpc8528 (
      {stage2_59[90]},
      {stage3_59[30]}
   );
   gpc1_1 gpc8529 (
      {stage2_59[91]},
      {stage3_59[31]}
   );
   gpc1_1 gpc8530 (
      {stage2_59[92]},
      {stage3_59[32]}
   );
   gpc1_1 gpc8531 (
      {stage2_59[93]},
      {stage3_59[33]}
   );
   gpc1_1 gpc8532 (
      {stage2_59[94]},
      {stage3_59[34]}
   );
   gpc1_1 gpc8533 (
      {stage2_59[95]},
      {stage3_59[35]}
   );
   gpc1_1 gpc8534 (
      {stage2_59[96]},
      {stage3_59[36]}
   );
   gpc1_1 gpc8535 (
      {stage2_59[97]},
      {stage3_59[37]}
   );
   gpc1_1 gpc8536 (
      {stage2_59[98]},
      {stage3_59[38]}
   );
   gpc1_1 gpc8537 (
      {stage2_59[99]},
      {stage3_59[39]}
   );
   gpc1_1 gpc8538 (
      {stage2_59[100]},
      {stage3_59[40]}
   );
   gpc1_1 gpc8539 (
      {stage2_59[101]},
      {stage3_59[41]}
   );
   gpc1_1 gpc8540 (
      {stage2_59[102]},
      {stage3_59[42]}
   );
   gpc1_1 gpc8541 (
      {stage2_59[103]},
      {stage3_59[43]}
   );
   gpc1_1 gpc8542 (
      {stage2_59[104]},
      {stage3_59[44]}
   );
   gpc1_1 gpc8543 (
      {stage2_59[105]},
      {stage3_59[45]}
   );
   gpc1_1 gpc8544 (
      {stage2_59[106]},
      {stage3_59[46]}
   );
   gpc1_1 gpc8545 (
      {stage2_59[107]},
      {stage3_59[47]}
   );
   gpc1_1 gpc8546 (
      {stage2_59[108]},
      {stage3_59[48]}
   );
   gpc1_1 gpc8547 (
      {stage2_59[109]},
      {stage3_59[49]}
   );
   gpc1_1 gpc8548 (
      {stage2_60[73]},
      {stage3_60[30]}
   );
   gpc1_1 gpc8549 (
      {stage2_60[74]},
      {stage3_60[31]}
   );
   gpc1_1 gpc8550 (
      {stage2_60[75]},
      {stage3_60[32]}
   );
   gpc1_1 gpc8551 (
      {stage2_60[76]},
      {stage3_60[33]}
   );
   gpc1_1 gpc8552 (
      {stage2_60[77]},
      {stage3_60[34]}
   );
   gpc1_1 gpc8553 (
      {stage2_60[78]},
      {stage3_60[35]}
   );
   gpc1_1 gpc8554 (
      {stage2_60[79]},
      {stage3_60[36]}
   );
   gpc1_1 gpc8555 (
      {stage2_60[80]},
      {stage3_60[37]}
   );
   gpc1_1 gpc8556 (
      {stage2_60[81]},
      {stage3_60[38]}
   );
   gpc1_1 gpc8557 (
      {stage2_60[82]},
      {stage3_60[39]}
   );
   gpc1_1 gpc8558 (
      {stage2_60[83]},
      {stage3_60[40]}
   );
   gpc1_1 gpc8559 (
      {stage2_60[84]},
      {stage3_60[41]}
   );
   gpc1_1 gpc8560 (
      {stage2_61[48]},
      {stage3_61[26]}
   );
   gpc1_1 gpc8561 (
      {stage2_61[49]},
      {stage3_61[27]}
   );
   gpc1_1 gpc8562 (
      {stage2_61[50]},
      {stage3_61[28]}
   );
   gpc1_1 gpc8563 (
      {stage2_61[51]},
      {stage3_61[29]}
   );
   gpc1_1 gpc8564 (
      {stage2_61[52]},
      {stage3_61[30]}
   );
   gpc1_1 gpc8565 (
      {stage2_61[53]},
      {stage3_61[31]}
   );
   gpc1_1 gpc8566 (
      {stage2_61[54]},
      {stage3_61[32]}
   );
   gpc1_1 gpc8567 (
      {stage2_61[55]},
      {stage3_61[33]}
   );
   gpc1_1 gpc8568 (
      {stage2_61[56]},
      {stage3_61[34]}
   );
   gpc1_1 gpc8569 (
      {stage2_61[57]},
      {stage3_61[35]}
   );
   gpc1_1 gpc8570 (
      {stage2_61[58]},
      {stage3_61[36]}
   );
   gpc1_1 gpc8571 (
      {stage2_61[59]},
      {stage3_61[37]}
   );
   gpc1_1 gpc8572 (
      {stage2_61[60]},
      {stage3_61[38]}
   );
   gpc1_1 gpc8573 (
      {stage2_61[61]},
      {stage3_61[39]}
   );
   gpc1_1 gpc8574 (
      {stage2_61[62]},
      {stage3_61[40]}
   );
   gpc1_1 gpc8575 (
      {stage2_61[63]},
      {stage3_61[41]}
   );
   gpc1_1 gpc8576 (
      {stage2_61[64]},
      {stage3_61[42]}
   );
   gpc1_1 gpc8577 (
      {stage2_61[65]},
      {stage3_61[43]}
   );
   gpc1_1 gpc8578 (
      {stage2_61[66]},
      {stage3_61[44]}
   );
   gpc1_1 gpc8579 (
      {stage2_61[67]},
      {stage3_61[45]}
   );
   gpc1_1 gpc8580 (
      {stage2_61[68]},
      {stage3_61[46]}
   );
   gpc1_1 gpc8581 (
      {stage2_61[69]},
      {stage3_61[47]}
   );
   gpc1_1 gpc8582 (
      {stage2_61[70]},
      {stage3_61[48]}
   );
   gpc1_1 gpc8583 (
      {stage2_61[71]},
      {stage3_61[49]}
   );
   gpc1_1 gpc8584 (
      {stage2_61[72]},
      {stage3_61[50]}
   );
   gpc1_1 gpc8585 (
      {stage2_61[73]},
      {stage3_61[51]}
   );
   gpc1_1 gpc8586 (
      {stage2_61[74]},
      {stage3_61[52]}
   );
   gpc1_1 gpc8587 (
      {stage2_63[90]},
      {stage3_63[39]}
   );
   gpc1_1 gpc8588 (
      {stage2_63[91]},
      {stage3_63[40]}
   );
   gpc1_1 gpc8589 (
      {stage2_63[92]},
      {stage3_63[41]}
   );
   gpc1_1 gpc8590 (
      {stage2_63[93]},
      {stage3_63[42]}
   );
   gpc1_1 gpc8591 (
      {stage2_63[94]},
      {stage3_63[43]}
   );
   gpc1_1 gpc8592 (
      {stage2_63[95]},
      {stage3_63[44]}
   );
   gpc1_1 gpc8593 (
      {stage2_63[96]},
      {stage3_63[45]}
   );
   gpc1_1 gpc8594 (
      {stage2_63[97]},
      {stage3_63[46]}
   );
   gpc1_1 gpc8595 (
      {stage2_63[98]},
      {stage3_63[47]}
   );
   gpc1_1 gpc8596 (
      {stage2_64[129]},
      {stage3_64[38]}
   );
   gpc1_1 gpc8597 (
      {stage2_64[130]},
      {stage3_64[39]}
   );
   gpc1_1 gpc8598 (
      {stage2_64[131]},
      {stage3_64[40]}
   );
   gpc1_1 gpc8599 (
      {stage2_64[132]},
      {stage3_64[41]}
   );
   gpc1_1 gpc8600 (
      {stage2_64[133]},
      {stage3_64[42]}
   );
   gpc1_1 gpc8601 (
      {stage2_64[134]},
      {stage3_64[43]}
   );
   gpc1_1 gpc8602 (
      {stage2_64[135]},
      {stage3_64[44]}
   );
   gpc1_1 gpc8603 (
      {stage2_64[136]},
      {stage3_64[45]}
   );
   gpc1_1 gpc8604 (
      {stage2_64[137]},
      {stage3_64[46]}
   );
   gpc1_1 gpc8605 (
      {stage2_64[138]},
      {stage3_64[47]}
   );
   gpc1_1 gpc8606 (
      {stage2_64[139]},
      {stage3_64[48]}
   );
   gpc1_1 gpc8607 (
      {stage2_64[140]},
      {stage3_64[49]}
   );
   gpc1_1 gpc8608 (
      {stage2_64[141]},
      {stage3_64[50]}
   );
   gpc1_1 gpc8609 (
      {stage2_65[51]},
      {stage3_65[33]}
   );
   gpc1_1 gpc8610 (
      {stage2_65[52]},
      {stage3_65[34]}
   );
   gpc1_1 gpc8611 (
      {stage2_65[53]},
      {stage3_65[35]}
   );
   gpc1_1 gpc8612 (
      {stage2_65[54]},
      {stage3_65[36]}
   );
   gpc1_1 gpc8613 (
      {stage2_65[55]},
      {stage3_65[37]}
   );
   gpc1_1 gpc8614 (
      {stage2_66[36]},
      {stage3_66[32]}
   );
   gpc1_1 gpc8615 (
      {stage2_66[37]},
      {stage3_66[33]}
   );
   gpc1_1 gpc8616 (
      {stage2_66[38]},
      {stage3_66[34]}
   );
   gpc1_1 gpc8617 (
      {stage2_66[39]},
      {stage3_66[35]}
   );
   gpc1_1 gpc8618 (
      {stage2_66[40]},
      {stage3_66[36]}
   );
   gpc1_1 gpc8619 (
      {stage2_66[41]},
      {stage3_66[37]}
   );
   gpc615_5 gpc8620 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4]},
      {stage3_1[0]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc8621 (
      {stage3_0[5], stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9]},
      {stage3_1[1]},
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc615_5 gpc8622 (
      {stage3_0[10], stage3_0[11], stage3_0[12], stage3_0[13], stage3_0[14]},
      {stage3_1[2]},
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2],stage4_0[2]}
   );
   gpc606_5 gpc8623 (
      {stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6], stage3_1[7], stage3_1[8]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc606_5 gpc8624 (
      {stage3_1[9], stage3_1[10], stage3_1[11], stage3_1[12], stage3_1[13], stage3_1[14]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[4],stage4_3[4],stage4_2[4],stage4_1[4]}
   );
   gpc606_5 gpc8625 (
      {stage3_1[15], stage3_1[16], stage3_1[17], stage3_1[18], stage3_1[19], stage3_1[20]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[5],stage4_3[5],stage4_2[5],stage4_1[5]}
   );
   gpc606_5 gpc8626 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[3],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc606_5 gpc8627 (
      {stage3_2[24], stage3_2[25], stage3_2[26], stage3_2[27], stage3_2[28], stage3_2[29]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[4],stage4_4[7],stage4_3[7],stage4_2[7]}
   );
   gpc606_5 gpc8628 (
      {stage3_2[30], stage3_2[31], stage3_2[32], stage3_2[33], stage3_2[34], stage3_2[35]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[5],stage4_4[8],stage4_3[8],stage4_2[8]}
   );
   gpc606_5 gpc8629 (
      {stage3_2[36], stage3_2[37], stage3_2[38], stage3_2[39], stage3_2[40], stage3_2[41]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[6],stage4_4[9],stage4_3[9],stage4_2[9]}
   );
   gpc615_5 gpc8630 (
      {stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22]},
      {stage3_4[24]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[4],stage4_5[7],stage4_4[10],stage4_3[10]}
   );
   gpc1163_5 gpc8631 (
      {stage3_4[25], stage3_4[26], stage3_4[27]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_6[0]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[1],stage4_6[5],stage4_5[8],stage4_4[11]}
   );
   gpc1163_5 gpc8632 (
      {stage3_4[28], stage3_4[29], stage3_4[30]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_6[1]},
      {stage3_7[1]},
      {stage4_8[1],stage4_7[2],stage4_6[6],stage4_5[9],stage4_4[12]}
   );
   gpc1163_5 gpc8633 (
      {stage3_4[31], stage3_4[32], stage3_4[33]},
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_6[2]},
      {stage3_7[2]},
      {stage4_8[2],stage4_7[3],stage4_6[7],stage4_5[10],stage4_4[13]}
   );
   gpc1163_5 gpc8634 (
      {stage3_4[34], stage3_4[35], stage3_4[36]},
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage3_6[3]},
      {stage3_7[3]},
      {stage4_8[3],stage4_7[4],stage4_6[8],stage4_5[11],stage4_4[14]}
   );
   gpc1163_5 gpc8635 (
      {stage3_4[37], stage3_4[38], stage3_4[39]},
      {stage3_5[30], stage3_5[31], stage3_5[32], stage3_5[33], stage3_5[34], stage3_5[35]},
      {stage3_6[4]},
      {stage3_7[4]},
      {stage4_8[4],stage4_7[5],stage4_6[9],stage4_5[12],stage4_4[15]}
   );
   gpc1163_5 gpc8636 (
      {stage3_4[40], stage3_4[41], stage3_4[42]},
      {stage3_5[36], stage3_5[37], stage3_5[38], stage3_5[39], stage3_5[40], stage3_5[41]},
      {stage3_6[5]},
      {stage3_7[5]},
      {stage4_8[5],stage4_7[6],stage4_6[10],stage4_5[13],stage4_4[16]}
   );
   gpc606_5 gpc8637 (
      {stage3_4[43], stage3_4[44], stage3_4[45], stage3_4[46], stage3_4[47], stage3_4[48]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[6],stage4_7[7],stage4_6[11],stage4_5[14],stage4_4[17]}
   );
   gpc606_5 gpc8638 (
      {stage3_4[49], stage3_4[50], stage3_4[51], stage3_4[52], stage3_4[53], stage3_4[54]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[7],stage4_7[8],stage4_6[12],stage4_5[15],stage4_4[18]}
   );
   gpc606_5 gpc8639 (
      {stage3_4[55], stage3_4[56], stage3_4[57], stage3_4[58], stage3_4[59], stage3_4[60]},
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage4_8[8],stage4_7[9],stage4_6[13],stage4_5[16],stage4_4[19]}
   );
   gpc606_5 gpc8640 (
      {stage3_4[61], stage3_4[62], stage3_4[63], stage3_4[64], stage3_4[65], stage3_4[66]},
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage4_8[9],stage4_7[10],stage4_6[14],stage4_5[17],stage4_4[20]}
   );
   gpc606_5 gpc8641 (
      {stage3_4[67], stage3_4[68], stage3_4[69], stage3_4[70], stage3_4[71], stage3_4[72]},
      {stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33], stage3_6[34], stage3_6[35]},
      {stage4_8[10],stage4_7[11],stage4_6[15],stage4_5[18],stage4_4[21]}
   );
   gpc606_5 gpc8642 (
      {stage3_4[73], stage3_4[74], stage3_4[75], stage3_4[76], stage3_4[77], stage3_4[78]},
      {stage3_6[36], stage3_6[37], stage3_6[38], stage3_6[39], stage3_6[40], stage3_6[41]},
      {stage4_8[11],stage4_7[12],stage4_6[16],stage4_5[19],stage4_4[22]}
   );
   gpc606_5 gpc8643 (
      {stage3_4[79], stage3_4[80], stage3_4[81], stage3_4[82], stage3_4[83], stage3_4[84]},
      {stage3_6[42], stage3_6[43], stage3_6[44], stage3_6[45], stage3_6[46], stage3_6[47]},
      {stage4_8[12],stage4_7[13],stage4_6[17],stage4_5[20],stage4_4[23]}
   );
   gpc606_5 gpc8644 (
      {stage3_4[85], stage3_4[86], stage3_4[87], stage3_4[88], stage3_4[89], stage3_4[90]},
      {stage3_6[48], stage3_6[49], stage3_6[50], stage3_6[51], stage3_6[52], stage3_6[53]},
      {stage4_8[13],stage4_7[14],stage4_6[18],stage4_5[21],stage4_4[24]}
   );
   gpc606_5 gpc8645 (
      {stage3_4[91], stage3_4[92], stage3_4[93], stage3_4[94], stage3_4[95], stage3_4[96]},
      {stage3_6[54], stage3_6[55], stage3_6[56], stage3_6[57], stage3_6[58], stage3_6[59]},
      {stage4_8[14],stage4_7[15],stage4_6[19],stage4_5[22],stage4_4[25]}
   );
   gpc606_5 gpc8646 (
      {stage3_4[97], stage3_4[98], stage3_4[99], stage3_4[100], stage3_4[101], stage3_4[102]},
      {stage3_6[60], stage3_6[61], stage3_6[62], stage3_6[63], stage3_6[64], stage3_6[65]},
      {stage4_8[15],stage4_7[16],stage4_6[20],stage4_5[23],stage4_4[26]}
   );
   gpc606_5 gpc8647 (
      {stage3_4[103], stage3_4[104], stage3_4[105], stage3_4[106], stage3_4[107], stage3_4[108]},
      {stage3_6[66], stage3_6[67], stage3_6[68], stage3_6[69], stage3_6[70], stage3_6[71]},
      {stage4_8[16],stage4_7[17],stage4_6[21],stage4_5[24],stage4_4[27]}
   );
   gpc615_5 gpc8648 (
      {stage3_6[72], stage3_6[73], stage3_6[74], stage3_6[75], stage3_6[76]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[17],stage4_7[18],stage4_6[22]}
   );
   gpc615_5 gpc8649 (
      {stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[18],stage4_7[19]}
   );
   gpc615_5 gpc8650 (
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16]},
      {stage3_8[7]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[19],stage4_7[20]}
   );
   gpc615_5 gpc8651 (
      {stage3_7[17], stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21]},
      {stage3_8[8]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[3],stage4_9[3],stage4_8[20],stage4_7[21]}
   );
   gpc615_5 gpc8652 (
      {stage3_7[22], stage3_7[23], stage3_7[24], stage3_7[25], stage3_7[26]},
      {stage3_8[9]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[4],stage4_9[4],stage4_8[21],stage4_7[22]}
   );
   gpc615_5 gpc8653 (
      {stage3_7[27], stage3_7[28], stage3_7[29], stage3_7[30], stage3_7[31]},
      {stage3_8[10]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[5],stage4_9[5],stage4_8[22],stage4_7[23]}
   );
   gpc615_5 gpc8654 (
      {stage3_7[32], stage3_7[33], stage3_7[34], stage3_7[35], stage3_7[36]},
      {stage3_8[11]},
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage4_11[5],stage4_10[6],stage4_9[6],stage4_8[23],stage4_7[24]}
   );
   gpc606_5 gpc8655 (
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[6],stage4_10[7],stage4_9[7],stage4_8[24]}
   );
   gpc606_5 gpc8656 (
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[7],stage4_10[8],stage4_9[8],stage4_8[25]}
   );
   gpc606_5 gpc8657 (
      {stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28], stage3_8[29]},
      {stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17]},
      {stage4_12[2],stage4_11[8],stage4_10[9],stage4_9[9],stage4_8[26]}
   );
   gpc606_5 gpc8658 (
      {stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33], stage3_8[34], 1'b0},
      {stage3_10[18], stage3_10[19], stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23]},
      {stage4_12[3],stage4_11[9],stage4_10[10],stage4_9[10],stage4_8[27]}
   );
   gpc606_5 gpc8659 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[4],stage4_11[10],stage4_10[11],stage4_9[11]}
   );
   gpc606_5 gpc8660 (
      {stage3_9[42], stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[5],stage4_11[11],stage4_10[12],stage4_9[12]}
   );
   gpc606_5 gpc8661 (
      {stage3_9[48], stage3_9[49], stage3_9[50], stage3_9[51], stage3_9[52], stage3_9[53]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[6],stage4_11[12],stage4_10[13],stage4_9[13]}
   );
   gpc615_5 gpc8662 (
      {stage3_10[24], stage3_10[25], stage3_10[26], stage3_10[27], stage3_10[28]},
      {stage3_11[18]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[3],stage4_12[7],stage4_11[13],stage4_10[14]}
   );
   gpc615_5 gpc8663 (
      {stage3_10[29], stage3_10[30], stage3_10[31], stage3_10[32], stage3_10[33]},
      {stage3_11[19]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[4],stage4_12[8],stage4_11[14],stage4_10[15]}
   );
   gpc615_5 gpc8664 (
      {stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37], stage3_10[38]},
      {stage3_11[20]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[5],stage4_12[9],stage4_11[15],stage4_10[16]}
   );
   gpc615_5 gpc8665 (
      {stage3_10[39], stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43]},
      {stage3_11[21]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[6],stage4_12[10],stage4_11[16],stage4_10[17]}
   );
   gpc615_5 gpc8666 (
      {stage3_10[44], stage3_10[45], stage3_10[46], stage3_10[47], stage3_10[48]},
      {stage3_11[22]},
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage4_14[4],stage4_13[7],stage4_12[11],stage4_11[17],stage4_10[18]}
   );
   gpc615_5 gpc8667 (
      {stage3_10[49], stage3_10[50], stage3_10[51], stage3_10[52], stage3_10[53]},
      {stage3_11[23]},
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage4_14[5],stage4_13[8],stage4_12[12],stage4_11[18],stage4_10[19]}
   );
   gpc615_5 gpc8668 (
      {stage3_10[54], stage3_10[55], stage3_10[56], stage3_10[57], stage3_10[58]},
      {stage3_11[24]},
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage4_14[6],stage4_13[9],stage4_12[13],stage4_11[19],stage4_10[20]}
   );
   gpc615_5 gpc8669 (
      {stage3_10[59], stage3_10[60], stage3_10[61], stage3_10[62], stage3_10[63]},
      {stage3_11[25]},
      {stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46], stage3_12[47]},
      {stage4_14[7],stage4_13[10],stage4_12[14],stage4_11[20],stage4_10[21]}
   );
   gpc615_5 gpc8670 (
      {stage3_10[64], stage3_10[65], stage3_10[66], stage3_10[67], stage3_10[68]},
      {stage3_11[26]},
      {stage3_12[48], stage3_12[49], stage3_12[50], stage3_12[51], stage3_12[52], stage3_12[53]},
      {stage4_14[8],stage4_13[11],stage4_12[15],stage4_11[21],stage4_10[22]}
   );
   gpc615_5 gpc8671 (
      {stage3_10[69], stage3_10[70], stage3_10[71], stage3_10[72], stage3_10[73]},
      {stage3_11[27]},
      {stage3_12[54], stage3_12[55], stage3_12[56], stage3_12[57], stage3_12[58], stage3_12[59]},
      {stage4_14[9],stage4_13[12],stage4_12[16],stage4_11[22],stage4_10[23]}
   );
   gpc1325_5 gpc8672 (
      {stage3_10[74], stage3_10[75], stage3_10[76], stage3_10[77], stage3_10[78]},
      {stage3_11[28], stage3_11[29]},
      {stage3_12[60], stage3_12[61], stage3_12[62]},
      {stage3_13[0]},
      {stage4_14[10],stage4_13[13],stage4_12[17],stage4_11[23],stage4_10[24]}
   );
   gpc1325_5 gpc8673 (
      {stage3_10[79], stage3_10[80], stage3_10[81], stage3_10[82], stage3_10[83]},
      {stage3_11[30], stage3_11[31]},
      {stage3_12[63], stage3_12[64], stage3_12[65]},
      {stage3_13[1]},
      {stage4_14[11],stage4_13[14],stage4_12[18],stage4_11[24],stage4_10[25]}
   );
   gpc207_4 gpc8674 (
      {stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35], stage3_11[36], stage3_11[37], stage3_11[38]},
      {stage3_13[2], stage3_13[3]},
      {stage4_14[12],stage4_13[15],stage4_12[19],stage4_11[25]}
   );
   gpc207_4 gpc8675 (
      {stage3_11[39], stage3_11[40], stage3_11[41], stage3_11[42], stage3_11[43], stage3_11[44], stage3_11[45]},
      {stage3_13[4], stage3_13[5]},
      {stage4_14[13],stage4_13[16],stage4_12[20],stage4_11[26]}
   );
   gpc207_4 gpc8676 (
      {stage3_11[46], stage3_11[47], stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51], stage3_11[52]},
      {stage3_13[6], stage3_13[7]},
      {stage4_14[14],stage4_13[17],stage4_12[21],stage4_11[27]}
   );
   gpc615_5 gpc8677 (
      {stage3_11[53], stage3_11[54], stage3_11[55], stage3_11[56], stage3_11[57]},
      {stage3_12[66]},
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13]},
      {stage4_15[0],stage4_14[15],stage4_13[18],stage4_12[22],stage4_11[28]}
   );
   gpc606_5 gpc8678 (
      {stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[16],stage4_13[19]}
   );
   gpc606_5 gpc8679 (
      {stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[1],stage4_15[2],stage4_14[17],stage4_13[20]}
   );
   gpc606_5 gpc8680 (
      {stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30], stage3_13[31]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[2],stage4_15[3],stage4_14[18],stage4_13[21]}
   );
   gpc606_5 gpc8681 (
      {stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35], stage3_13[36], stage3_13[37]},
      {stage3_15[18], stage3_15[19], stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23]},
      {stage4_17[3],stage4_16[3],stage4_15[4],stage4_14[19],stage4_13[22]}
   );
   gpc606_5 gpc8682 (
      {stage3_13[38], stage3_13[39], stage3_13[40], stage3_13[41], stage3_13[42], stage3_13[43]},
      {stage3_15[24], stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage4_17[4],stage4_16[4],stage4_15[5],stage4_14[20],stage4_13[23]}
   );
   gpc606_5 gpc8683 (
      {stage3_13[44], stage3_13[45], stage3_13[46], stage3_13[47], stage3_13[48], stage3_13[49]},
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34], stage3_15[35]},
      {stage4_17[5],stage4_16[5],stage4_15[6],stage4_14[21],stage4_13[24]}
   );
   gpc615_5 gpc8684 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4]},
      {stage3_15[36]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[6],stage4_16[6],stage4_15[7],stage4_14[22]}
   );
   gpc615_5 gpc8685 (
      {stage3_14[5], stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9]},
      {stage3_15[37]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[7],stage4_16[7],stage4_15[8],stage4_14[23]}
   );
   gpc615_5 gpc8686 (
      {stage3_14[10], stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14]},
      {stage3_15[38]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[8],stage4_16[8],stage4_15[9],stage4_14[24]}
   );
   gpc615_5 gpc8687 (
      {stage3_14[15], stage3_14[16], stage3_14[17], stage3_14[18], stage3_14[19]},
      {stage3_15[39]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[9],stage4_16[9],stage4_15[10],stage4_14[25]}
   );
   gpc615_5 gpc8688 (
      {stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24]},
      {stage3_15[40]},
      {stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29]},
      {stage4_18[4],stage4_17[10],stage4_16[10],stage4_15[11],stage4_14[26]}
   );
   gpc615_5 gpc8689 (
      {stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29]},
      {stage3_15[41]},
      {stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35]},
      {stage4_18[5],stage4_17[11],stage4_16[11],stage4_15[12],stage4_14[27]}
   );
   gpc615_5 gpc8690 (
      {stage3_15[42], stage3_15[43], stage3_15[44], stage3_15[45], stage3_15[46]},
      {stage3_16[36]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[6],stage4_17[12],stage4_16[12],stage4_15[13]}
   );
   gpc606_5 gpc8691 (
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[7],stage4_17[13]}
   );
   gpc606_5 gpc8692 (
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[1],stage4_19[2],stage4_18[8],stage4_17[14]}
   );
   gpc606_5 gpc8693 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage4_21[2],stage4_20[2],stage4_19[3],stage4_18[9],stage4_17[15]}
   );
   gpc606_5 gpc8694 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[18], stage3_19[19], stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23]},
      {stage4_21[3],stage4_20[3],stage4_19[4],stage4_18[10],stage4_17[16]}
   );
   gpc606_5 gpc8695 (
      {stage3_17[30], stage3_17[31], stage3_17[32], stage3_17[33], stage3_17[34], stage3_17[35]},
      {stage3_19[24], stage3_19[25], stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29]},
      {stage4_21[4],stage4_20[4],stage4_19[5],stage4_18[11],stage4_17[17]}
   );
   gpc207_4 gpc8696 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage3_20[0], stage3_20[1]},
      {stage4_21[5],stage4_20[5],stage4_19[6],stage4_18[12]}
   );
   gpc207_4 gpc8697 (
      {stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12], stage3_18[13]},
      {stage3_20[2], stage3_20[3]},
      {stage4_21[6],stage4_20[6],stage4_19[7],stage4_18[13]}
   );
   gpc207_4 gpc8698 (
      {stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17], stage3_18[18], stage3_18[19], stage3_18[20]},
      {stage3_20[4], stage3_20[5]},
      {stage4_21[7],stage4_20[7],stage4_19[8],stage4_18[14]}
   );
   gpc207_4 gpc8699 (
      {stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25], stage3_18[26], stage3_18[27]},
      {stage3_20[6], stage3_20[7]},
      {stage4_21[8],stage4_20[8],stage4_19[9],stage4_18[15]}
   );
   gpc207_4 gpc8700 (
      {stage3_18[28], stage3_18[29], stage3_18[30], stage3_18[31], stage3_18[32], stage3_18[33], stage3_18[34]},
      {stage3_20[8], stage3_20[9]},
      {stage4_21[9],stage4_20[9],stage4_19[10],stage4_18[16]}
   );
   gpc207_4 gpc8701 (
      {stage3_18[35], stage3_18[36], stage3_18[37], stage3_18[38], stage3_18[39], stage3_18[40], stage3_18[41]},
      {stage3_20[10], stage3_20[11]},
      {stage4_21[10],stage4_20[10],stage4_19[11],stage4_18[17]}
   );
   gpc207_4 gpc8702 (
      {stage3_18[42], stage3_18[43], stage3_18[44], stage3_18[45], stage3_18[46], stage3_18[47], stage3_18[48]},
      {stage3_20[12], stage3_20[13]},
      {stage4_21[11],stage4_20[11],stage4_19[12],stage4_18[18]}
   );
   gpc207_4 gpc8703 (
      {stage3_18[49], stage3_18[50], stage3_18[51], stage3_18[52], stage3_18[53], stage3_18[54], stage3_18[55]},
      {stage3_20[14], stage3_20[15]},
      {stage4_21[12],stage4_20[12],stage4_19[13],stage4_18[19]}
   );
   gpc207_4 gpc8704 (
      {stage3_18[56], stage3_18[57], stage3_18[58], stage3_18[59], 1'b0, 1'b0, 1'b0},
      {stage3_20[16], stage3_20[17]},
      {stage4_21[13],stage4_20[13],stage4_19[14],stage4_18[20]}
   );
   gpc615_5 gpc8705 (
      {stage3_19[30], stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34]},
      {stage3_20[18]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[14],stage4_20[14],stage4_19[15]}
   );
   gpc606_5 gpc8706 (
      {stage3_20[19], stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23], stage3_20[24]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[15],stage4_20[15]}
   );
   gpc606_5 gpc8707 (
      {stage3_20[25], stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29], stage3_20[30]},
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11]},
      {stage4_24[1],stage4_23[2],stage4_22[2],stage4_21[16],stage4_20[16]}
   );
   gpc606_5 gpc8708 (
      {stage3_20[31], stage3_20[32], stage3_20[33], stage3_20[34], stage3_20[35], stage3_20[36]},
      {stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17]},
      {stage4_24[2],stage4_23[3],stage4_22[3],stage4_21[17],stage4_20[17]}
   );
   gpc606_5 gpc8709 (
      {stage3_20[37], stage3_20[38], stage3_20[39], stage3_20[40], stage3_20[41], stage3_20[42]},
      {stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23]},
      {stage4_24[3],stage4_23[4],stage4_22[4],stage4_21[18],stage4_20[18]}
   );
   gpc606_5 gpc8710 (
      {stage3_20[43], stage3_20[44], stage3_20[45], stage3_20[46], stage3_20[47], stage3_20[48]},
      {stage3_22[24], stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28], stage3_22[29]},
      {stage4_24[4],stage4_23[5],stage4_22[5],stage4_21[19],stage4_20[19]}
   );
   gpc606_5 gpc8711 (
      {stage3_20[49], stage3_20[50], stage3_20[51], stage3_20[52], stage3_20[53], stage3_20[54]},
      {stage3_22[30], stage3_22[31], stage3_22[32], stage3_22[33], stage3_22[34], stage3_22[35]},
      {stage4_24[5],stage4_23[6],stage4_22[6],stage4_21[20],stage4_20[20]}
   );
   gpc606_5 gpc8712 (
      {stage3_20[55], stage3_20[56], stage3_20[57], stage3_20[58], stage3_20[59], stage3_20[60]},
      {stage3_22[36], stage3_22[37], stage3_22[38], stage3_22[39], stage3_22[40], stage3_22[41]},
      {stage4_24[6],stage4_23[7],stage4_22[7],stage4_21[21],stage4_20[21]}
   );
   gpc606_5 gpc8713 (
      {stage3_20[61], stage3_20[62], stage3_20[63], stage3_20[64], stage3_20[65], stage3_20[66]},
      {stage3_22[42], stage3_22[43], stage3_22[44], stage3_22[45], stage3_22[46], stage3_22[47]},
      {stage4_24[7],stage4_23[8],stage4_22[8],stage4_21[22],stage4_20[22]}
   );
   gpc606_5 gpc8714 (
      {stage3_20[67], stage3_20[68], stage3_20[69], stage3_20[70], stage3_20[71], stage3_20[72]},
      {stage3_22[48], stage3_22[49], stage3_22[50], stage3_22[51], stage3_22[52], stage3_22[53]},
      {stage4_24[8],stage4_23[9],stage4_22[9],stage4_21[23],stage4_20[23]}
   );
   gpc606_5 gpc8715 (
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[9],stage4_23[10],stage4_22[10],stage4_21[24]}
   );
   gpc606_5 gpc8716 (
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[10],stage4_23[11],stage4_22[11],stage4_21[25]}
   );
   gpc606_5 gpc8717 (
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage3_23[12], stage3_23[13], stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17]},
      {stage4_25[2],stage4_24[11],stage4_23[12],stage4_22[12],stage4_21[26]}
   );
   gpc606_5 gpc8718 (
      {stage3_21[24], stage3_21[25], stage3_21[26], stage3_21[27], stage3_21[28], stage3_21[29]},
      {stage3_23[18], stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23]},
      {stage4_25[3],stage4_24[12],stage4_23[13],stage4_22[13],stage4_21[27]}
   );
   gpc615_5 gpc8719 (
      {stage3_22[54], stage3_22[55], stage3_22[56], stage3_22[57], stage3_22[58]},
      {stage3_23[24]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[4],stage4_24[13],stage4_23[14],stage4_22[14]}
   );
   gpc615_5 gpc8720 (
      {stage3_22[59], stage3_22[60], stage3_22[61], stage3_22[62], stage3_22[63]},
      {stage3_23[25]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[5],stage4_24[14],stage4_23[15],stage4_22[15]}
   );
   gpc615_5 gpc8721 (
      {stage3_22[64], stage3_22[65], stage3_22[66], stage3_22[67], stage3_22[68]},
      {stage3_23[26]},
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17]},
      {stage4_26[2],stage4_25[6],stage4_24[15],stage4_23[16],stage4_22[16]}
   );
   gpc615_5 gpc8722 (
      {stage3_22[69], stage3_22[70], stage3_22[71], stage3_22[72], 1'b0},
      {stage3_23[27]},
      {stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23]},
      {stage4_26[3],stage4_25[7],stage4_24[16],stage4_23[17],stage4_22[17]}
   );
   gpc615_5 gpc8723 (
      {stage3_23[28], stage3_23[29], stage3_23[30], stage3_23[31], stage3_23[32]},
      {stage3_24[24]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[4],stage4_25[8],stage4_24[17],stage4_23[18]}
   );
   gpc615_5 gpc8724 (
      {stage3_23[33], stage3_23[34], stage3_23[35], stage3_23[36], stage3_23[37]},
      {stage3_24[25]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[5],stage4_25[9],stage4_24[18],stage4_23[19]}
   );
   gpc615_5 gpc8725 (
      {stage3_23[38], stage3_23[39], stage3_23[40], stage3_23[41], stage3_23[42]},
      {stage3_24[26]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[6],stage4_25[10],stage4_24[19],stage4_23[20]}
   );
   gpc606_5 gpc8726 (
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[3],stage4_26[7],stage4_25[11]}
   );
   gpc1163_5 gpc8727 (
      {stage3_26[0], stage3_26[1], stage3_26[2]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage3_28[0]},
      {stage3_29[0]},
      {stage4_30[0],stage4_29[1],stage4_28[1],stage4_27[4],stage4_26[8]}
   );
   gpc1163_5 gpc8728 (
      {stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage3_28[1]},
      {stage3_29[1]},
      {stage4_30[1],stage4_29[2],stage4_28[2],stage4_27[5],stage4_26[9]}
   );
   gpc1163_5 gpc8729 (
      {stage3_26[6], stage3_26[7], stage3_26[8]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage3_28[2]},
      {stage3_29[2]},
      {stage4_30[2],stage4_29[3],stage4_28[3],stage4_27[6],stage4_26[10]}
   );
   gpc615_5 gpc8730 (
      {stage3_26[9], stage3_26[10], stage3_26[11], stage3_26[12], stage3_26[13]},
      {stage3_27[24]},
      {stage3_28[3], stage3_28[4], stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8]},
      {stage4_30[3],stage4_29[4],stage4_28[4],stage4_27[7],stage4_26[11]}
   );
   gpc615_5 gpc8731 (
      {stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17], stage3_26[18]},
      {stage3_27[25]},
      {stage3_28[9], stage3_28[10], stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14]},
      {stage4_30[4],stage4_29[5],stage4_28[5],stage4_27[8],stage4_26[12]}
   );
   gpc615_5 gpc8732 (
      {stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage3_27[26]},
      {stage3_28[15], stage3_28[16], stage3_28[17], stage3_28[18], stage3_28[19], stage3_28[20]},
      {stage4_30[5],stage4_29[6],stage4_28[6],stage4_27[9],stage4_26[13]}
   );
   gpc615_5 gpc8733 (
      {stage3_26[24], stage3_26[25], stage3_26[26], stage3_26[27], stage3_26[28]},
      {stage3_27[27]},
      {stage3_28[21], stage3_28[22], stage3_28[23], stage3_28[24], stage3_28[25], stage3_28[26]},
      {stage4_30[6],stage4_29[7],stage4_28[7],stage4_27[10],stage4_26[14]}
   );
   gpc615_5 gpc8734 (
      {stage3_26[29], stage3_26[30], stage3_26[31], stage3_26[32], stage3_26[33]},
      {stage3_27[28]},
      {stage3_28[27], stage3_28[28], stage3_28[29], stage3_28[30], stage3_28[31], stage3_28[32]},
      {stage4_30[7],stage4_29[8],stage4_28[8],stage4_27[11],stage4_26[15]}
   );
   gpc615_5 gpc8735 (
      {stage3_26[34], stage3_26[35], stage3_26[36], stage3_26[37], stage3_26[38]},
      {stage3_27[29]},
      {stage3_28[33], stage3_28[34], stage3_28[35], stage3_28[36], stage3_28[37], stage3_28[38]},
      {stage4_30[8],stage4_29[9],stage4_28[9],stage4_27[12],stage4_26[16]}
   );
   gpc615_5 gpc8736 (
      {stage3_26[39], stage3_26[40], stage3_26[41], stage3_26[42], stage3_26[43]},
      {stage3_27[30]},
      {stage3_28[39], stage3_28[40], stage3_28[41], stage3_28[42], stage3_28[43], stage3_28[44]},
      {stage4_30[9],stage4_29[10],stage4_28[10],stage4_27[13],stage4_26[17]}
   );
   gpc615_5 gpc8737 (
      {stage3_26[44], stage3_26[45], stage3_26[46], stage3_26[47], stage3_26[48]},
      {stage3_27[31]},
      {stage3_28[45], stage3_28[46], stage3_28[47], stage3_28[48], stage3_28[49], stage3_28[50]},
      {stage4_30[10],stage4_29[11],stage4_28[11],stage4_27[14],stage4_26[18]}
   );
   gpc606_5 gpc8738 (
      {stage3_27[32], stage3_27[33], stage3_27[34], stage3_27[35], stage3_27[36], stage3_27[37]},
      {stage3_29[3], stage3_29[4], stage3_29[5], stage3_29[6], stage3_29[7], stage3_29[8]},
      {stage4_31[0],stage4_30[11],stage4_29[12],stage4_28[12],stage4_27[15]}
   );
   gpc1163_5 gpc8739 (
      {stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[0]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[1],stage4_30[12],stage4_29[13]}
   );
   gpc1163_5 gpc8740 (
      {stage3_29[12], stage3_29[13], stage3_29[14]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage3_31[1]},
      {stage3_32[1]},
      {stage4_33[1],stage4_32[1],stage4_31[2],stage4_30[13],stage4_29[14]}
   );
   gpc1163_5 gpc8741 (
      {stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage3_31[2]},
      {stage3_32[2]},
      {stage4_33[2],stage4_32[2],stage4_31[3],stage4_30[14],stage4_29[15]}
   );
   gpc1163_5 gpc8742 (
      {stage3_29[18], stage3_29[19], stage3_29[20]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage3_31[3]},
      {stage3_32[3]},
      {stage4_33[3],stage4_32[3],stage4_31[4],stage4_30[15],stage4_29[16]}
   );
   gpc1163_5 gpc8743 (
      {stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage3_31[4]},
      {stage3_32[4]},
      {stage4_33[4],stage4_32[4],stage4_31[5],stage4_30[16],stage4_29[17]}
   );
   gpc606_5 gpc8744 (
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10]},
      {stage4_33[5],stage4_32[5],stage4_31[6],stage4_30[17],stage4_29[18]}
   );
   gpc606_5 gpc8745 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34], stage3_29[35]},
      {stage3_31[11], stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16]},
      {stage4_33[6],stage4_32[6],stage4_31[7],stage4_30[18],stage4_29[19]}
   );
   gpc606_5 gpc8746 (
      {stage3_29[36], stage3_29[37], stage3_29[38], stage3_29[39], stage3_29[40], stage3_29[41]},
      {stage3_31[17], stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22]},
      {stage4_33[7],stage4_32[7],stage4_31[8],stage4_30[19],stage4_29[20]}
   );
   gpc606_5 gpc8747 (
      {stage3_29[42], stage3_29[43], stage3_29[44], stage3_29[45], stage3_29[46], stage3_29[47]},
      {stage3_31[23], stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28]},
      {stage4_33[8],stage4_32[8],stage4_31[9],stage4_30[20],stage4_29[21]}
   );
   gpc615_5 gpc8748 (
      {stage3_31[29], stage3_31[30], stage3_31[31], stage3_31[32], stage3_31[33]},
      {stage3_32[5]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[0],stage4_33[9],stage4_32[9],stage4_31[10]}
   );
   gpc2135_5 gpc8749 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10]},
      {stage3_33[6], stage3_33[7], stage3_33[8]},
      {stage3_34[0]},
      {stage3_35[0], stage3_35[1]},
      {stage4_36[0],stage4_35[1],stage4_34[1],stage4_33[10],stage4_32[10]}
   );
   gpc2135_5 gpc8750 (
      {stage3_32[11], stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15]},
      {stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_34[1]},
      {stage3_35[2], stage3_35[3]},
      {stage4_36[1],stage4_35[2],stage4_34[2],stage4_33[11],stage4_32[11]}
   );
   gpc615_5 gpc8751 (
      {stage3_32[16], stage3_32[17], stage3_32[18], stage3_32[19], stage3_32[20]},
      {stage3_33[12]},
      {stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5], stage3_34[6], stage3_34[7]},
      {stage4_36[2],stage4_35[3],stage4_34[3],stage4_33[12],stage4_32[12]}
   );
   gpc615_5 gpc8752 (
      {stage3_32[21], stage3_32[22], stage3_32[23], stage3_32[24], stage3_32[25]},
      {stage3_33[13]},
      {stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11], stage3_34[12], stage3_34[13]},
      {stage4_36[3],stage4_35[4],stage4_34[4],stage4_33[13],stage4_32[13]}
   );
   gpc615_5 gpc8753 (
      {stage3_32[26], stage3_32[27], stage3_32[28], stage3_32[29], stage3_32[30]},
      {stage3_33[14]},
      {stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17], stage3_34[18], stage3_34[19]},
      {stage4_36[4],stage4_35[5],stage4_34[5],stage4_33[14],stage4_32[14]}
   );
   gpc615_5 gpc8754 (
      {stage3_32[31], stage3_32[32], stage3_32[33], stage3_32[34], stage3_32[35]},
      {stage3_33[15]},
      {stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23], stage3_34[24], stage3_34[25]},
      {stage4_36[5],stage4_35[6],stage4_34[6],stage4_33[15],stage4_32[15]}
   );
   gpc615_5 gpc8755 (
      {stage3_32[36], stage3_32[37], stage3_32[38], stage3_32[39], stage3_32[40]},
      {stage3_33[16]},
      {stage3_34[26], stage3_34[27], stage3_34[28], stage3_34[29], stage3_34[30], stage3_34[31]},
      {stage4_36[6],stage4_35[7],stage4_34[7],stage4_33[16],stage4_32[16]}
   );
   gpc117_4 gpc8756 (
      {stage3_33[17], stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage3_34[32]},
      {stage3_35[4]},
      {stage4_36[7],stage4_35[8],stage4_34[8],stage4_33[17]}
   );
   gpc117_4 gpc8757 (
      {stage3_33[24], stage3_33[25], stage3_33[26], stage3_33[27], stage3_33[28], stage3_33[29], stage3_33[30]},
      {stage3_34[33]},
      {stage3_35[5]},
      {stage4_36[8],stage4_35[9],stage4_34[9],stage4_33[18]}
   );
   gpc606_5 gpc8758 (
      {stage3_33[31], stage3_33[32], stage3_33[33], stage3_33[34], stage3_33[35], stage3_33[36]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[0],stage4_36[9],stage4_35[10],stage4_34[10],stage4_33[19]}
   );
   gpc615_5 gpc8759 (
      {stage3_35[12], stage3_35[13], stage3_35[14], stage3_35[15], stage3_35[16]},
      {stage3_36[0]},
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage4_39[0],stage4_38[0],stage4_37[1],stage4_36[10],stage4_35[11]}
   );
   gpc615_5 gpc8760 (
      {stage3_35[17], stage3_35[18], stage3_35[19], stage3_35[20], stage3_35[21]},
      {stage3_36[1]},
      {stage3_37[6], stage3_37[7], stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage4_39[1],stage4_38[1],stage4_37[2],stage4_36[11],stage4_35[12]}
   );
   gpc615_5 gpc8761 (
      {stage3_35[22], stage3_35[23], stage3_35[24], stage3_35[25], stage3_35[26]},
      {stage3_36[2]},
      {stage3_37[12], stage3_37[13], stage3_37[14], stage3_37[15], stage3_37[16], stage3_37[17]},
      {stage4_39[2],stage4_38[2],stage4_37[3],stage4_36[12],stage4_35[13]}
   );
   gpc615_5 gpc8762 (
      {stage3_35[27], stage3_35[28], stage3_35[29], stage3_35[30], stage3_35[31]},
      {stage3_36[3]},
      {stage3_37[18], stage3_37[19], stage3_37[20], stage3_37[21], stage3_37[22], stage3_37[23]},
      {stage4_39[3],stage4_38[3],stage4_37[4],stage4_36[13],stage4_35[14]}
   );
   gpc615_5 gpc8763 (
      {stage3_35[32], stage3_35[33], stage3_35[34], stage3_35[35], stage3_35[36]},
      {stage3_36[4]},
      {stage3_37[24], stage3_37[25], stage3_37[26], stage3_37[27], stage3_37[28], stage3_37[29]},
      {stage4_39[4],stage4_38[4],stage4_37[5],stage4_36[14],stage4_35[15]}
   );
   gpc606_5 gpc8764 (
      {stage3_36[5], stage3_36[6], stage3_36[7], stage3_36[8], stage3_36[9], stage3_36[10]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[5],stage4_38[5],stage4_37[6],stage4_36[15]}
   );
   gpc606_5 gpc8765 (
      {stage3_36[11], stage3_36[12], stage3_36[13], stage3_36[14], stage3_36[15], stage3_36[16]},
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11]},
      {stage4_40[1],stage4_39[6],stage4_38[6],stage4_37[7],stage4_36[16]}
   );
   gpc606_5 gpc8766 (
      {stage3_36[17], stage3_36[18], stage3_36[19], stage3_36[20], stage3_36[21], stage3_36[22]},
      {stage3_38[12], stage3_38[13], stage3_38[14], stage3_38[15], stage3_38[16], stage3_38[17]},
      {stage4_40[2],stage4_39[7],stage4_38[7],stage4_37[8],stage4_36[17]}
   );
   gpc606_5 gpc8767 (
      {stage3_36[23], stage3_36[24], stage3_36[25], stage3_36[26], stage3_36[27], stage3_36[28]},
      {stage3_38[18], stage3_38[19], stage3_38[20], stage3_38[21], stage3_38[22], stage3_38[23]},
      {stage4_40[3],stage4_39[8],stage4_38[8],stage4_37[9],stage4_36[18]}
   );
   gpc606_5 gpc8768 (
      {stage3_37[30], stage3_37[31], stage3_37[32], stage3_37[33], stage3_37[34], stage3_37[35]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[4],stage4_39[9],stage4_38[9],stage4_37[10]}
   );
   gpc606_5 gpc8769 (
      {stage3_37[36], stage3_37[37], stage3_37[38], stage3_37[39], stage3_37[40], stage3_37[41]},
      {stage3_39[6], stage3_39[7], stage3_39[8], stage3_39[9], stage3_39[10], stage3_39[11]},
      {stage4_41[1],stage4_40[5],stage4_39[10],stage4_38[10],stage4_37[11]}
   );
   gpc606_5 gpc8770 (
      {stage3_37[42], stage3_37[43], stage3_37[44], stage3_37[45], stage3_37[46], stage3_37[47]},
      {stage3_39[12], stage3_39[13], stage3_39[14], stage3_39[15], stage3_39[16], stage3_39[17]},
      {stage4_41[2],stage4_40[6],stage4_39[11],stage4_38[11],stage4_37[12]}
   );
   gpc615_5 gpc8771 (
      {stage3_38[24], stage3_38[25], stage3_38[26], stage3_38[27], stage3_38[28]},
      {stage3_39[18]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[3],stage4_40[7],stage4_39[12],stage4_38[12]}
   );
   gpc615_5 gpc8772 (
      {stage3_38[29], stage3_38[30], stage3_38[31], stage3_38[32], stage3_38[33]},
      {stage3_39[19]},
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage4_42[1],stage4_41[4],stage4_40[8],stage4_39[13],stage4_38[13]}
   );
   gpc615_5 gpc8773 (
      {stage3_38[34], stage3_38[35], stage3_38[36], stage3_38[37], stage3_38[38]},
      {stage3_39[20]},
      {stage3_40[12], stage3_40[13], stage3_40[14], stage3_40[15], stage3_40[16], stage3_40[17]},
      {stage4_42[2],stage4_41[5],stage4_40[9],stage4_39[14],stage4_38[14]}
   );
   gpc615_5 gpc8774 (
      {stage3_38[39], stage3_38[40], stage3_38[41], stage3_38[42], stage3_38[43]},
      {stage3_39[21]},
      {stage3_40[18], stage3_40[19], stage3_40[20], stage3_40[21], stage3_40[22], stage3_40[23]},
      {stage4_42[3],stage4_41[6],stage4_40[10],stage4_39[15],stage4_38[15]}
   );
   gpc615_5 gpc8775 (
      {stage3_38[44], stage3_38[45], stage3_38[46], stage3_38[47], stage3_38[48]},
      {stage3_39[22]},
      {stage3_40[24], stage3_40[25], stage3_40[26], stage3_40[27], stage3_40[28], stage3_40[29]},
      {stage4_42[4],stage4_41[7],stage4_40[11],stage4_39[16],stage4_38[16]}
   );
   gpc615_5 gpc8776 (
      {stage3_38[49], stage3_38[50], stage3_38[51], stage3_38[52], stage3_38[53]},
      {stage3_39[23]},
      {stage3_40[30], stage3_40[31], stage3_40[32], stage3_40[33], stage3_40[34], stage3_40[35]},
      {stage4_42[5],stage4_41[8],stage4_40[12],stage4_39[17],stage4_38[17]}
   );
   gpc615_5 gpc8777 (
      {stage3_38[54], stage3_38[55], stage3_38[56], stage3_38[57], stage3_38[58]},
      {stage3_39[24]},
      {stage3_40[36], stage3_40[37], stage3_40[38], stage3_40[39], stage3_40[40], stage3_40[41]},
      {stage4_42[6],stage4_41[9],stage4_40[13],stage4_39[18],stage4_38[18]}
   );
   gpc207_4 gpc8778 (
      {stage3_39[25], stage3_39[26], stage3_39[27], stage3_39[28], stage3_39[29], stage3_39[30], stage3_39[31]},
      {stage3_41[0], stage3_41[1]},
      {stage4_42[7],stage4_41[10],stage4_40[14],stage4_39[19]}
   );
   gpc207_4 gpc8779 (
      {stage3_39[32], stage3_39[33], stage3_39[34], stage3_39[35], stage3_39[36], stage3_39[37], stage3_39[38]},
      {stage3_41[2], stage3_41[3]},
      {stage4_42[8],stage4_41[11],stage4_40[15],stage4_39[20]}
   );
   gpc207_4 gpc8780 (
      {stage3_39[39], stage3_39[40], stage3_39[41], stage3_39[42], stage3_39[43], stage3_39[44], stage3_39[45]},
      {stage3_41[4], stage3_41[5]},
      {stage4_42[9],stage4_41[12],stage4_40[16],stage4_39[21]}
   );
   gpc207_4 gpc8781 (
      {stage3_39[46], stage3_39[47], stage3_39[48], stage3_39[49], stage3_39[50], stage3_39[51], stage3_39[52]},
      {stage3_41[6], stage3_41[7]},
      {stage4_42[10],stage4_41[13],stage4_40[17],stage4_39[22]}
   );
   gpc615_5 gpc8782 (
      {stage3_39[53], stage3_39[54], stage3_39[55], stage3_39[56], stage3_39[57]},
      {stage3_40[42]},
      {stage3_41[8], stage3_41[9], stage3_41[10], stage3_41[11], stage3_41[12], stage3_41[13]},
      {stage4_43[0],stage4_42[11],stage4_41[14],stage4_40[18],stage4_39[23]}
   );
   gpc606_5 gpc8783 (
      {stage3_41[14], stage3_41[15], stage3_41[16], stage3_41[17], stage3_41[18], stage3_41[19]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[1],stage4_42[12],stage4_41[15]}
   );
   gpc606_5 gpc8784 (
      {stage3_41[20], stage3_41[21], stage3_41[22], stage3_41[23], stage3_41[24], stage3_41[25]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[1],stage4_43[2],stage4_42[13],stage4_41[16]}
   );
   gpc606_5 gpc8785 (
      {stage3_41[26], stage3_41[27], stage3_41[28], stage3_41[29], stage3_41[30], stage3_41[31]},
      {stage3_43[12], stage3_43[13], stage3_43[14], stage3_43[15], stage3_43[16], stage3_43[17]},
      {stage4_45[2],stage4_44[2],stage4_43[3],stage4_42[14],stage4_41[17]}
   );
   gpc606_5 gpc8786 (
      {stage3_41[32], stage3_41[33], stage3_41[34], stage3_41[35], stage3_41[36], stage3_41[37]},
      {stage3_43[18], stage3_43[19], stage3_43[20], stage3_43[21], stage3_43[22], stage3_43[23]},
      {stage4_45[3],stage4_44[3],stage4_43[4],stage4_42[15],stage4_41[18]}
   );
   gpc606_5 gpc8787 (
      {stage3_41[38], stage3_41[39], stage3_41[40], stage3_41[41], stage3_41[42], 1'b0},
      {stage3_43[24], stage3_43[25], stage3_43[26], stage3_43[27], stage3_43[28], stage3_43[29]},
      {stage4_45[4],stage4_44[4],stage4_43[5],stage4_42[16],stage4_41[19]}
   );
   gpc207_4 gpc8788 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5], stage3_42[6]},
      {stage3_44[0], stage3_44[1]},
      {stage4_45[5],stage4_44[5],stage4_43[6],stage4_42[17]}
   );
   gpc207_4 gpc8789 (
      {stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11], stage3_42[12], stage3_42[13]},
      {stage3_44[2], stage3_44[3]},
      {stage4_45[6],stage4_44[6],stage4_43[7],stage4_42[18]}
   );
   gpc207_4 gpc8790 (
      {stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17], stage3_42[18], stage3_42[19], stage3_42[20]},
      {stage3_44[4], stage3_44[5]},
      {stage4_45[7],stage4_44[7],stage4_43[8],stage4_42[19]}
   );
   gpc207_4 gpc8791 (
      {stage3_42[21], stage3_42[22], stage3_42[23], stage3_42[24], stage3_42[25], stage3_42[26], stage3_42[27]},
      {stage3_44[6], stage3_44[7]},
      {stage4_45[8],stage4_44[8],stage4_43[9],stage4_42[20]}
   );
   gpc606_5 gpc8792 (
      {stage3_42[28], stage3_42[29], stage3_42[30], stage3_42[31], stage3_42[32], stage3_42[33]},
      {stage3_44[8], stage3_44[9], stage3_44[10], stage3_44[11], stage3_44[12], stage3_44[13]},
      {stage4_46[0],stage4_45[9],stage4_44[9],stage4_43[10],stage4_42[21]}
   );
   gpc606_5 gpc8793 (
      {stage3_43[30], stage3_43[31], stage3_43[32], stage3_43[33], stage3_43[34], stage3_43[35]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[1],stage4_45[10],stage4_44[10],stage4_43[11]}
   );
   gpc606_5 gpc8794 (
      {stage3_43[36], stage3_43[37], stage3_43[38], stage3_43[39], stage3_43[40], stage3_43[41]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage4_47[1],stage4_46[2],stage4_45[11],stage4_44[11],stage4_43[12]}
   );
   gpc615_5 gpc8795 (
      {stage3_43[42], stage3_43[43], stage3_43[44], stage3_43[45], 1'b0},
      {stage3_44[14]},
      {stage3_45[12], stage3_45[13], stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage4_47[2],stage4_46[3],stage4_45[12],stage4_44[12],stage4_43[13]}
   );
   gpc606_5 gpc8796 (
      {stage3_44[15], stage3_44[16], stage3_44[17], stage3_44[18], stage3_44[19], stage3_44[20]},
      {stage3_46[0], stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage4_48[0],stage4_47[3],stage4_46[4],stage4_45[13],stage4_44[13]}
   );
   gpc606_5 gpc8797 (
      {stage3_44[21], stage3_44[22], stage3_44[23], stage3_44[24], stage3_44[25], stage3_44[26]},
      {stage3_46[6], stage3_46[7], stage3_46[8], stage3_46[9], stage3_46[10], stage3_46[11]},
      {stage4_48[1],stage4_47[4],stage4_46[5],stage4_45[14],stage4_44[14]}
   );
   gpc615_5 gpc8798 (
      {stage3_44[27], stage3_44[28], stage3_44[29], stage3_44[30], stage3_44[31]},
      {stage3_45[18]},
      {stage3_46[12], stage3_46[13], stage3_46[14], stage3_46[15], stage3_46[16], stage3_46[17]},
      {stage4_48[2],stage4_47[5],stage4_46[6],stage4_45[15],stage4_44[15]}
   );
   gpc135_4 gpc8799 (
      {stage3_45[19], stage3_45[20], stage3_45[21], stage3_45[22], stage3_45[23]},
      {stage3_46[18], stage3_46[19], stage3_46[20]},
      {stage3_47[0]},
      {stage4_48[3],stage4_47[6],stage4_46[7],stage4_45[16]}
   );
   gpc135_4 gpc8800 (
      {stage3_45[24], stage3_45[25], stage3_45[26], stage3_45[27], stage3_45[28]},
      {stage3_46[21], stage3_46[22], stage3_46[23]},
      {stage3_47[1]},
      {stage4_48[4],stage4_47[7],stage4_46[8],stage4_45[17]}
   );
   gpc135_4 gpc8801 (
      {stage3_45[29], stage3_45[30], stage3_45[31], stage3_45[32], stage3_45[33]},
      {stage3_46[24], stage3_46[25], stage3_46[26]},
      {stage3_47[2]},
      {stage4_48[5],stage4_47[8],stage4_46[9],stage4_45[18]}
   );
   gpc615_5 gpc8802 (
      {stage3_46[27], stage3_46[28], stage3_46[29], stage3_46[30], stage3_46[31]},
      {stage3_47[3]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[6],stage4_47[9],stage4_46[10]}
   );
   gpc615_5 gpc8803 (
      {stage3_46[32], stage3_46[33], stage3_46[34], stage3_46[35], stage3_46[36]},
      {stage3_47[4]},
      {stage3_48[6], stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11]},
      {stage4_50[1],stage4_49[1],stage4_48[7],stage4_47[10],stage4_46[11]}
   );
   gpc615_5 gpc8804 (
      {stage3_46[37], stage3_46[38], stage3_46[39], stage3_46[40], stage3_46[41]},
      {stage3_47[5]},
      {stage3_48[12], stage3_48[13], stage3_48[14], stage3_48[15], stage3_48[16], stage3_48[17]},
      {stage4_50[2],stage4_49[2],stage4_48[8],stage4_47[11],stage4_46[12]}
   );
   gpc615_5 gpc8805 (
      {stage3_46[42], stage3_46[43], stage3_46[44], stage3_46[45], stage3_46[46]},
      {stage3_47[6]},
      {stage3_48[18], stage3_48[19], stage3_48[20], stage3_48[21], stage3_48[22], stage3_48[23]},
      {stage4_50[3],stage4_49[3],stage4_48[9],stage4_47[12],stage4_46[13]}
   );
   gpc615_5 gpc8806 (
      {stage3_46[47], stage3_46[48], stage3_46[49], stage3_46[50], stage3_46[51]},
      {stage3_47[7]},
      {stage3_48[24], stage3_48[25], stage3_48[26], stage3_48[27], stage3_48[28], stage3_48[29]},
      {stage4_50[4],stage4_49[4],stage4_48[10],stage4_47[13],stage4_46[14]}
   );
   gpc615_5 gpc8807 (
      {stage3_46[52], stage3_46[53], stage3_46[54], stage3_46[55], stage3_46[56]},
      {stage3_47[8]},
      {stage3_48[30], stage3_48[31], stage3_48[32], stage3_48[33], stage3_48[34], stage3_48[35]},
      {stage4_50[5],stage4_49[5],stage4_48[11],stage4_47[14],stage4_46[15]}
   );
   gpc606_5 gpc8808 (
      {stage3_47[9], stage3_47[10], stage3_47[11], stage3_47[12], stage3_47[13], stage3_47[14]},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage4_51[0],stage4_50[6],stage4_49[6],stage4_48[12],stage4_47[15]}
   );
   gpc606_5 gpc8809 (
      {stage3_47[15], stage3_47[16], stage3_47[17], stage3_47[18], stage3_47[19], stage3_47[20]},
      {stage3_49[6], stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11]},
      {stage4_51[1],stage4_50[7],stage4_49[7],stage4_48[13],stage4_47[16]}
   );
   gpc606_5 gpc8810 (
      {stage3_47[21], stage3_47[22], stage3_47[23], stage3_47[24], stage3_47[25], stage3_47[26]},
      {stage3_49[12], stage3_49[13], stage3_49[14], stage3_49[15], stage3_49[16], stage3_49[17]},
      {stage4_51[2],stage4_50[8],stage4_49[8],stage4_48[14],stage4_47[17]}
   );
   gpc606_5 gpc8811 (
      {stage3_47[27], stage3_47[28], stage3_47[29], stage3_47[30], stage3_47[31], stage3_47[32]},
      {stage3_49[18], stage3_49[19], stage3_49[20], stage3_49[21], stage3_49[22], stage3_49[23]},
      {stage4_51[3],stage4_50[9],stage4_49[9],stage4_48[15],stage4_47[18]}
   );
   gpc606_5 gpc8812 (
      {stage3_47[33], stage3_47[34], stage3_47[35], stage3_47[36], stage3_47[37], stage3_47[38]},
      {stage3_49[24], stage3_49[25], stage3_49[26], stage3_49[27], stage3_49[28], stage3_49[29]},
      {stage4_51[4],stage4_50[10],stage4_49[10],stage4_48[16],stage4_47[19]}
   );
   gpc615_5 gpc8813 (
      {stage3_47[39], stage3_47[40], stage3_47[41], stage3_47[42], stage3_47[43]},
      {stage3_48[36]},
      {stage3_49[30], stage3_49[31], stage3_49[32], stage3_49[33], stage3_49[34], stage3_49[35]},
      {stage4_51[5],stage4_50[11],stage4_49[11],stage4_48[17],stage4_47[20]}
   );
   gpc606_5 gpc8814 (
      {stage3_49[36], stage3_49[37], stage3_49[38], stage3_49[39], stage3_49[40], stage3_49[41]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[0],stage4_51[6],stage4_50[12],stage4_49[12]}
   );
   gpc117_4 gpc8815 (
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6]},
      {stage3_51[6]},
      {stage3_52[0]},
      {stage4_53[1],stage4_52[1],stage4_51[7],stage4_50[13]}
   );
   gpc117_4 gpc8816 (
      {stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12], stage3_50[13]},
      {stage3_51[7]},
      {stage3_52[1]},
      {stage4_53[2],stage4_52[2],stage4_51[8],stage4_50[14]}
   );
   gpc615_5 gpc8817 (
      {stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17], stage3_50[18]},
      {stage3_51[8]},
      {stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5], stage3_52[6], stage3_52[7]},
      {stage4_54[0],stage4_53[3],stage4_52[3],stage4_51[9],stage4_50[15]}
   );
   gpc615_5 gpc8818 (
      {stage3_50[19], stage3_50[20], stage3_50[21], stage3_50[22], stage3_50[23]},
      {stage3_51[9]},
      {stage3_52[8], stage3_52[9], stage3_52[10], stage3_52[11], stage3_52[12], stage3_52[13]},
      {stage4_54[1],stage4_53[4],stage4_52[4],stage4_51[10],stage4_50[16]}
   );
   gpc615_5 gpc8819 (
      {stage3_50[24], stage3_50[25], stage3_50[26], stage3_50[27], stage3_50[28]},
      {stage3_51[10]},
      {stage3_52[14], stage3_52[15], stage3_52[16], stage3_52[17], stage3_52[18], stage3_52[19]},
      {stage4_54[2],stage4_53[5],stage4_52[5],stage4_51[11],stage4_50[17]}
   );
   gpc615_5 gpc8820 (
      {stage3_50[29], stage3_50[30], stage3_50[31], stage3_50[32], stage3_50[33]},
      {stage3_51[11]},
      {stage3_52[20], stage3_52[21], stage3_52[22], stage3_52[23], stage3_52[24], stage3_52[25]},
      {stage4_54[3],stage4_53[6],stage4_52[6],stage4_51[12],stage4_50[18]}
   );
   gpc615_5 gpc8821 (
      {stage3_50[34], stage3_50[35], stage3_50[36], stage3_50[37], stage3_50[38]},
      {stage3_51[12]},
      {stage3_52[26], stage3_52[27], stage3_52[28], stage3_52[29], stage3_52[30], stage3_52[31]},
      {stage4_54[4],stage4_53[7],stage4_52[7],stage4_51[13],stage4_50[19]}
   );
   gpc615_5 gpc8822 (
      {stage3_50[39], stage3_50[40], stage3_50[41], stage3_50[42], stage3_50[43]},
      {stage3_51[13]},
      {stage3_52[32], stage3_52[33], stage3_52[34], stage3_52[35], stage3_52[36], stage3_52[37]},
      {stage4_54[5],stage4_53[8],stage4_52[8],stage4_51[14],stage4_50[20]}
   );
   gpc615_5 gpc8823 (
      {stage3_50[44], stage3_50[45], stage3_50[46], 1'b0, 1'b0},
      {stage3_51[14]},
      {stage3_52[38], stage3_52[39], stage3_52[40], stage3_52[41], stage3_52[42], stage3_52[43]},
      {stage4_54[6],stage4_53[9],stage4_52[9],stage4_51[15],stage4_50[21]}
   );
   gpc2135_5 gpc8824 (
      {stage3_51[15], stage3_51[16], stage3_51[17], stage3_51[18], stage3_51[19]},
      {stage3_52[44], stage3_52[45], stage3_52[46]},
      {stage3_53[0]},
      {stage3_54[0], stage3_54[1]},
      {stage4_55[0],stage4_54[7],stage4_53[10],stage4_52[10],stage4_51[16]}
   );
   gpc2135_5 gpc8825 (
      {stage3_51[20], stage3_51[21], stage3_51[22], stage3_51[23], stage3_51[24]},
      {stage3_52[47], stage3_52[48], stage3_52[49]},
      {stage3_53[1]},
      {stage3_54[2], stage3_54[3]},
      {stage4_55[1],stage4_54[8],stage4_53[11],stage4_52[11],stage4_51[17]}
   );
   gpc2135_5 gpc8826 (
      {stage3_51[25], stage3_51[26], stage3_51[27], stage3_51[28], stage3_51[29]},
      {stage3_52[50], stage3_52[51], stage3_52[52]},
      {stage3_53[2]},
      {stage3_54[4], stage3_54[5]},
      {stage4_55[2],stage4_54[9],stage4_53[12],stage4_52[12],stage4_51[18]}
   );
   gpc2135_5 gpc8827 (
      {stage3_51[30], stage3_51[31], stage3_51[32], stage3_51[33], stage3_51[34]},
      {stage3_52[53], stage3_52[54], stage3_52[55]},
      {stage3_53[3]},
      {stage3_54[6], stage3_54[7]},
      {stage4_55[3],stage4_54[10],stage4_53[13],stage4_52[13],stage4_51[19]}
   );
   gpc2135_5 gpc8828 (
      {stage3_51[35], stage3_51[36], stage3_51[37], stage3_51[38], stage3_51[39]},
      {stage3_52[56], stage3_52[57], stage3_52[58]},
      {stage3_53[4]},
      {stage3_54[8], stage3_54[9]},
      {stage4_55[4],stage4_54[11],stage4_53[14],stage4_52[14],stage4_51[20]}
   );
   gpc615_5 gpc8829 (
      {stage3_51[40], stage3_51[41], stage3_51[42], stage3_51[43], stage3_51[44]},
      {stage3_52[59]},
      {stage3_53[5], stage3_53[6], stage3_53[7], stage3_53[8], stage3_53[9], stage3_53[10]},
      {stage4_55[5],stage4_54[12],stage4_53[15],stage4_52[15],stage4_51[21]}
   );
   gpc615_5 gpc8830 (
      {stage3_51[45], stage3_51[46], stage3_51[47], stage3_51[48], stage3_51[49]},
      {stage3_52[60]},
      {stage3_53[11], stage3_53[12], stage3_53[13], stage3_53[14], stage3_53[15], stage3_53[16]},
      {stage4_55[6],stage4_54[13],stage4_53[16],stage4_52[16],stage4_51[22]}
   );
   gpc606_5 gpc8831 (
      {stage3_53[17], stage3_53[18], stage3_53[19], stage3_53[20], stage3_53[21], stage3_53[22]},
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage4_57[0],stage4_56[0],stage4_55[7],stage4_54[14],stage4_53[17]}
   );
   gpc606_5 gpc8832 (
      {stage3_53[23], stage3_53[24], stage3_53[25], stage3_53[26], stage3_53[27], stage3_53[28]},
      {stage3_55[6], stage3_55[7], stage3_55[8], stage3_55[9], stage3_55[10], stage3_55[11]},
      {stage4_57[1],stage4_56[1],stage4_55[8],stage4_54[15],stage4_53[18]}
   );
   gpc606_5 gpc8833 (
      {stage3_53[29], stage3_53[30], stage3_53[31], stage3_53[32], stage3_53[33], stage3_53[34]},
      {stage3_55[12], stage3_55[13], stage3_55[14], stage3_55[15], stage3_55[16], stage3_55[17]},
      {stage4_57[2],stage4_56[2],stage4_55[9],stage4_54[16],stage4_53[19]}
   );
   gpc615_5 gpc8834 (
      {stage3_53[35], stage3_53[36], stage3_53[37], stage3_53[38], stage3_53[39]},
      {stage3_54[10]},
      {stage3_55[18], stage3_55[19], stage3_55[20], stage3_55[21], stage3_55[22], stage3_55[23]},
      {stage4_57[3],stage4_56[3],stage4_55[10],stage4_54[17],stage4_53[20]}
   );
   gpc615_5 gpc8835 (
      {stage3_53[40], stage3_53[41], stage3_53[42], stage3_53[43], stage3_53[44]},
      {stage3_54[11]},
      {stage3_55[24], stage3_55[25], stage3_55[26], stage3_55[27], stage3_55[28], stage3_55[29]},
      {stage4_57[4],stage4_56[4],stage4_55[11],stage4_54[18],stage4_53[21]}
   );
   gpc615_5 gpc8836 (
      {stage3_53[45], stage3_53[46], stage3_53[47], stage3_53[48], stage3_53[49]},
      {stage3_54[12]},
      {stage3_55[30], stage3_55[31], stage3_55[32], stage3_55[33], stage3_55[34], stage3_55[35]},
      {stage4_57[5],stage4_56[5],stage4_55[12],stage4_54[19],stage4_53[22]}
   );
   gpc615_5 gpc8837 (
      {stage3_53[50], stage3_53[51], stage3_53[52], stage3_53[53], stage3_53[54]},
      {stage3_54[13]},
      {stage3_55[36], stage3_55[37], stage3_55[38], stage3_55[39], stage3_55[40], stage3_55[41]},
      {stage4_57[6],stage4_56[6],stage4_55[13],stage4_54[20],stage4_53[23]}
   );
   gpc615_5 gpc8838 (
      {stage3_54[14], stage3_54[15], stage3_54[16], stage3_54[17], stage3_54[18]},
      {stage3_55[42]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage4_58[0],stage4_57[7],stage4_56[7],stage4_55[14],stage4_54[21]}
   );
   gpc615_5 gpc8839 (
      {stage3_54[19], stage3_54[20], stage3_54[21], stage3_54[22], stage3_54[23]},
      {stage3_55[43]},
      {stage3_56[6], stage3_56[7], stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11]},
      {stage4_58[1],stage4_57[8],stage4_56[8],stage4_55[15],stage4_54[22]}
   );
   gpc615_5 gpc8840 (
      {stage3_54[24], stage3_54[25], stage3_54[26], stage3_54[27], stage3_54[28]},
      {stage3_55[44]},
      {stage3_56[12], stage3_56[13], stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17]},
      {stage4_58[2],stage4_57[9],stage4_56[9],stage4_55[16],stage4_54[23]}
   );
   gpc615_5 gpc8841 (
      {stage3_54[29], stage3_54[30], stage3_54[31], stage3_54[32], stage3_54[33]},
      {stage3_55[45]},
      {stage3_56[18], stage3_56[19], stage3_56[20], stage3_56[21], stage3_56[22], stage3_56[23]},
      {stage4_58[3],stage4_57[10],stage4_56[10],stage4_55[17],stage4_54[24]}
   );
   gpc615_5 gpc8842 (
      {stage3_54[34], stage3_54[35], stage3_54[36], stage3_54[37], stage3_54[38]},
      {stage3_55[46]},
      {stage3_56[24], stage3_56[25], stage3_56[26], stage3_56[27], stage3_56[28], stage3_56[29]},
      {stage4_58[4],stage4_57[11],stage4_56[11],stage4_55[18],stage4_54[25]}
   );
   gpc1163_5 gpc8843 (
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage3_59[0]},
      {stage3_60[0]},
      {stage4_61[0],stage4_60[0],stage4_59[0],stage4_58[5],stage4_57[12]}
   );
   gpc1163_5 gpc8844 (
      {stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11]},
      {stage3_59[1]},
      {stage3_60[1]},
      {stage4_61[1],stage4_60[1],stage4_59[1],stage4_58[6],stage4_57[13]}
   );
   gpc1163_5 gpc8845 (
      {stage3_57[6], stage3_57[7], stage3_57[8]},
      {stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15], stage3_58[16], stage3_58[17]},
      {stage3_59[2]},
      {stage3_60[2]},
      {stage4_61[2],stage4_60[2],stage4_59[2],stage4_58[7],stage4_57[14]}
   );
   gpc1163_5 gpc8846 (
      {stage3_57[9], stage3_57[10], stage3_57[11]},
      {stage3_58[18], stage3_58[19], stage3_58[20], stage3_58[21], stage3_58[22], stage3_58[23]},
      {stage3_59[3]},
      {stage3_60[3]},
      {stage4_61[3],stage4_60[3],stage4_59[3],stage4_58[8],stage4_57[15]}
   );
   gpc1163_5 gpc8847 (
      {stage3_57[12], stage3_57[13], stage3_57[14]},
      {stage3_58[24], stage3_58[25], stage3_58[26], stage3_58[27], stage3_58[28], stage3_58[29]},
      {stage3_59[4]},
      {stage3_60[4]},
      {stage4_61[4],stage4_60[4],stage4_59[4],stage4_58[9],stage4_57[16]}
   );
   gpc1163_5 gpc8848 (
      {stage3_57[15], stage3_57[16], stage3_57[17]},
      {stage3_58[30], stage3_58[31], stage3_58[32], stage3_58[33], stage3_58[34], stage3_58[35]},
      {stage3_59[5]},
      {stage3_60[5]},
      {stage4_61[5],stage4_60[5],stage4_59[5],stage4_58[10],stage4_57[17]}
   );
   gpc1163_5 gpc8849 (
      {stage3_57[18], stage3_57[19], stage3_57[20]},
      {stage3_58[36], stage3_58[37], stage3_58[38], stage3_58[39], stage3_58[40], stage3_58[41]},
      {stage3_59[6]},
      {stage3_60[6]},
      {stage4_61[6],stage4_60[6],stage4_59[6],stage4_58[11],stage4_57[18]}
   );
   gpc1163_5 gpc8850 (
      {stage3_57[21], stage3_57[22], stage3_57[23]},
      {stage3_58[42], stage3_58[43], stage3_58[44], stage3_58[45], stage3_58[46], stage3_58[47]},
      {stage3_59[7]},
      {stage3_60[7]},
      {stage4_61[7],stage4_60[7],stage4_59[7],stage4_58[12],stage4_57[19]}
   );
   gpc1163_5 gpc8851 (
      {stage3_57[24], stage3_57[25], stage3_57[26]},
      {stage3_58[48], stage3_58[49], stage3_58[50], stage3_58[51], stage3_58[52], stage3_58[53]},
      {stage3_59[8]},
      {stage3_60[8]},
      {stage4_61[8],stage4_60[8],stage4_59[8],stage4_58[13],stage4_57[20]}
   );
   gpc606_5 gpc8852 (
      {stage3_57[27], stage3_57[28], stage3_57[29], stage3_57[30], stage3_57[31], stage3_57[32]},
      {stage3_59[9], stage3_59[10], stage3_59[11], stage3_59[12], stage3_59[13], stage3_59[14]},
      {stage4_61[9],stage4_60[9],stage4_59[9],stage4_58[14],stage4_57[21]}
   );
   gpc606_5 gpc8853 (
      {stage3_57[33], stage3_57[34], stage3_57[35], stage3_57[36], stage3_57[37], stage3_57[38]},
      {stage3_59[15], stage3_59[16], stage3_59[17], stage3_59[18], stage3_59[19], stage3_59[20]},
      {stage4_61[10],stage4_60[10],stage4_59[10],stage4_58[15],stage4_57[22]}
   );
   gpc615_5 gpc8854 (
      {stage3_57[39], stage3_57[40], stage3_57[41], stage3_57[42], stage3_57[43]},
      {stage3_58[54]},
      {stage3_59[21], stage3_59[22], stage3_59[23], stage3_59[24], stage3_59[25], stage3_59[26]},
      {stage4_61[11],stage4_60[11],stage4_59[11],stage4_58[16],stage4_57[23]}
   );
   gpc615_5 gpc8855 (
      {stage3_57[44], stage3_57[45], stage3_57[46], stage3_57[47], stage3_57[48]},
      {stage3_58[55]},
      {stage3_59[27], stage3_59[28], stage3_59[29], stage3_59[30], stage3_59[31], stage3_59[32]},
      {stage4_61[12],stage4_60[12],stage4_59[12],stage4_58[17],stage4_57[24]}
   );
   gpc615_5 gpc8856 (
      {stage3_57[49], stage3_57[50], stage3_57[51], stage3_57[52], stage3_57[53]},
      {stage3_58[56]},
      {stage3_59[33], stage3_59[34], stage3_59[35], stage3_59[36], stage3_59[37], stage3_59[38]},
      {stage4_61[13],stage4_60[13],stage4_59[13],stage4_58[18],stage4_57[25]}
   );
   gpc615_5 gpc8857 (
      {stage3_59[39], stage3_59[40], stage3_59[41], stage3_59[42], stage3_59[43]},
      {stage3_60[9]},
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {stage4_63[0],stage4_62[0],stage4_61[14],stage4_60[14],stage4_59[14]}
   );
   gpc606_5 gpc8858 (
      {stage3_60[10], stage3_60[11], stage3_60[12], stage3_60[13], stage3_60[14], stage3_60[15]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[1],stage4_62[1],stage4_61[15],stage4_60[15]}
   );
   gpc606_5 gpc8859 (
      {stage3_60[16], stage3_60[17], stage3_60[18], stage3_60[19], stage3_60[20], stage3_60[21]},
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage4_64[1],stage4_63[2],stage4_62[2],stage4_61[16],stage4_60[16]}
   );
   gpc606_5 gpc8860 (
      {stage3_60[22], stage3_60[23], stage3_60[24], stage3_60[25], stage3_60[26], stage3_60[27]},
      {stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15], stage3_62[16], stage3_62[17]},
      {stage4_64[2],stage4_63[3],stage4_62[3],stage4_61[17],stage4_60[17]}
   );
   gpc606_5 gpc8861 (
      {stage3_60[28], stage3_60[29], stage3_60[30], stage3_60[31], stage3_60[32], stage3_60[33]},
      {stage3_62[18], stage3_62[19], stage3_62[20], stage3_62[21], stage3_62[22], stage3_62[23]},
      {stage4_64[3],stage4_63[4],stage4_62[4],stage4_61[18],stage4_60[18]}
   );
   gpc606_5 gpc8862 (
      {stage3_60[34], stage3_60[35], stage3_60[36], stage3_60[37], stage3_60[38], stage3_60[39]},
      {stage3_62[24], stage3_62[25], stage3_62[26], stage3_62[27], stage3_62[28], stage3_62[29]},
      {stage4_64[4],stage4_63[5],stage4_62[5],stage4_61[19],stage4_60[19]}
   );
   gpc606_5 gpc8863 (
      {stage3_61[6], stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11]},
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage4_65[0],stage4_64[5],stage4_63[6],stage4_62[6],stage4_61[20]}
   );
   gpc606_5 gpc8864 (
      {stage3_61[12], stage3_61[13], stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17]},
      {stage3_63[6], stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11]},
      {stage4_65[1],stage4_64[6],stage4_63[7],stage4_62[7],stage4_61[21]}
   );
   gpc606_5 gpc8865 (
      {stage3_61[18], stage3_61[19], stage3_61[20], stage3_61[21], stage3_61[22], stage3_61[23]},
      {stage3_63[12], stage3_63[13], stage3_63[14], stage3_63[15], stage3_63[16], stage3_63[17]},
      {stage4_65[2],stage4_64[7],stage4_63[8],stage4_62[8],stage4_61[22]}
   );
   gpc606_5 gpc8866 (
      {stage3_61[24], stage3_61[25], stage3_61[26], stage3_61[27], stage3_61[28], stage3_61[29]},
      {stage3_63[18], stage3_63[19], stage3_63[20], stage3_63[21], stage3_63[22], stage3_63[23]},
      {stage4_65[3],stage4_64[8],stage4_63[9],stage4_62[9],stage4_61[23]}
   );
   gpc606_5 gpc8867 (
      {stage3_61[30], stage3_61[31], stage3_61[32], stage3_61[33], stage3_61[34], stage3_61[35]},
      {stage3_63[24], stage3_63[25], stage3_63[26], stage3_63[27], stage3_63[28], stage3_63[29]},
      {stage4_65[4],stage4_64[9],stage4_63[10],stage4_62[10],stage4_61[24]}
   );
   gpc606_5 gpc8868 (
      {stage3_61[36], stage3_61[37], stage3_61[38], stage3_61[39], stage3_61[40], stage3_61[41]},
      {stage3_63[30], stage3_63[31], stage3_63[32], stage3_63[33], stage3_63[34], stage3_63[35]},
      {stage4_65[5],stage4_64[10],stage4_63[11],stage4_62[11],stage4_61[25]}
   );
   gpc606_5 gpc8869 (
      {stage3_61[42], stage3_61[43], stage3_61[44], stage3_61[45], stage3_61[46], stage3_61[47]},
      {stage3_63[36], stage3_63[37], stage3_63[38], stage3_63[39], stage3_63[40], stage3_63[41]},
      {stage4_65[6],stage4_64[11],stage4_63[12],stage4_62[12],stage4_61[26]}
   );
   gpc606_5 gpc8870 (
      {stage3_63[42], stage3_63[43], stage3_63[44], stage3_63[45], stage3_63[46], stage3_63[47]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[0],stage4_65[7],stage4_64[12],stage4_63[13]}
   );
   gpc606_5 gpc8871 (
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[1],stage4_66[1],stage4_65[8],stage4_64[13]}
   );
   gpc606_5 gpc8872 (
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage3_66[6], stage3_66[7], stage3_66[8], stage3_66[9], stage3_66[10], stage3_66[11]},
      {stage4_68[1],stage4_67[2],stage4_66[2],stage4_65[9],stage4_64[14]}
   );
   gpc606_5 gpc8873 (
      {stage3_64[12], stage3_64[13], stage3_64[14], stage3_64[15], stage3_64[16], stage3_64[17]},
      {stage3_66[12], stage3_66[13], stage3_66[14], stage3_66[15], stage3_66[16], stage3_66[17]},
      {stage4_68[2],stage4_67[3],stage4_66[3],stage4_65[10],stage4_64[15]}
   );
   gpc606_5 gpc8874 (
      {stage3_64[18], stage3_64[19], stage3_64[20], stage3_64[21], stage3_64[22], stage3_64[23]},
      {stage3_66[18], stage3_66[19], stage3_66[20], stage3_66[21], stage3_66[22], stage3_66[23]},
      {stage4_68[3],stage4_67[4],stage4_66[4],stage4_65[11],stage4_64[16]}
   );
   gpc606_5 gpc8875 (
      {stage3_64[24], stage3_64[25], stage3_64[26], stage3_64[27], stage3_64[28], stage3_64[29]},
      {stage3_66[24], stage3_66[25], stage3_66[26], stage3_66[27], stage3_66[28], stage3_66[29]},
      {stage4_68[4],stage4_67[5],stage4_66[5],stage4_65[12],stage4_64[17]}
   );
   gpc606_5 gpc8876 (
      {stage3_64[30], stage3_64[31], stage3_64[32], stage3_64[33], stage3_64[34], stage3_64[35]},
      {stage3_66[30], stage3_66[31], stage3_66[32], stage3_66[33], stage3_66[34], stage3_66[35]},
      {stage4_68[5],stage4_67[6],stage4_66[6],stage4_65[13],stage4_64[18]}
   );
   gpc606_5 gpc8877 (
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage3_67[0], stage3_67[1], stage3_67[2], stage3_67[3], stage3_67[4], stage3_67[5]},
      {stage4_69[0],stage4_68[6],stage4_67[7],stage4_66[7],stage4_65[14]}
   );
   gpc606_5 gpc8878 (
      {stage3_65[12], stage3_65[13], stage3_65[14], stage3_65[15], stage3_65[16], stage3_65[17]},
      {stage3_67[6], stage3_67[7], stage3_67[8], stage3_67[9], stage3_67[10], stage3_67[11]},
      {stage4_69[1],stage4_68[7],stage4_67[8],stage4_66[8],stage4_65[15]}
   );
   gpc1_1 gpc8879 (
      {stage3_0[15]},
      {stage4_0[3]}
   );
   gpc1_1 gpc8880 (
      {stage3_0[16]},
      {stage4_0[4]}
   );
   gpc1_1 gpc8881 (
      {stage3_0[17]},
      {stage4_0[5]}
   );
   gpc1_1 gpc8882 (
      {stage3_0[18]},
      {stage4_0[6]}
   );
   gpc1_1 gpc8883 (
      {stage3_0[19]},
      {stage4_0[7]}
   );
   gpc1_1 gpc8884 (
      {stage3_0[20]},
      {stage4_0[8]}
   );
   gpc1_1 gpc8885 (
      {stage3_1[21]},
      {stage4_1[6]}
   );
   gpc1_1 gpc8886 (
      {stage3_2[42]},
      {stage4_2[10]}
   );
   gpc1_1 gpc8887 (
      {stage3_3[23]},
      {stage4_3[11]}
   );
   gpc1_1 gpc8888 (
      {stage3_3[24]},
      {stage4_3[12]}
   );
   gpc1_1 gpc8889 (
      {stage3_3[25]},
      {stage4_3[13]}
   );
   gpc1_1 gpc8890 (
      {stage3_3[26]},
      {stage4_3[14]}
   );
   gpc1_1 gpc8891 (
      {stage3_3[27]},
      {stage4_3[15]}
   );
   gpc1_1 gpc8892 (
      {stage3_3[28]},
      {stage4_3[16]}
   );
   gpc1_1 gpc8893 (
      {stage3_4[109]},
      {stage4_4[28]}
   );
   gpc1_1 gpc8894 (
      {stage3_4[110]},
      {stage4_4[29]}
   );
   gpc1_1 gpc8895 (
      {stage3_4[111]},
      {stage4_4[30]}
   );
   gpc1_1 gpc8896 (
      {stage3_5[42]},
      {stage4_5[25]}
   );
   gpc1_1 gpc8897 (
      {stage3_5[43]},
      {stage4_5[26]}
   );
   gpc1_1 gpc8898 (
      {stage3_5[44]},
      {stage4_5[27]}
   );
   gpc1_1 gpc8899 (
      {stage3_5[45]},
      {stage4_5[28]}
   );
   gpc1_1 gpc8900 (
      {stage3_5[46]},
      {stage4_5[29]}
   );
   gpc1_1 gpc8901 (
      {stage3_5[47]},
      {stage4_5[30]}
   );
   gpc1_1 gpc8902 (
      {stage3_5[48]},
      {stage4_5[31]}
   );
   gpc1_1 gpc8903 (
      {stage3_5[49]},
      {stage4_5[32]}
   );
   gpc1_1 gpc8904 (
      {stage3_5[50]},
      {stage4_5[33]}
   );
   gpc1_1 gpc8905 (
      {stage3_5[51]},
      {stage4_5[34]}
   );
   gpc1_1 gpc8906 (
      {stage3_5[52]},
      {stage4_5[35]}
   );
   gpc1_1 gpc8907 (
      {stage3_6[77]},
      {stage4_6[23]}
   );
   gpc1_1 gpc8908 (
      {stage3_7[37]},
      {stage4_7[25]}
   );
   gpc1_1 gpc8909 (
      {stage3_7[38]},
      {stage4_7[26]}
   );
   gpc1_1 gpc8910 (
      {stage3_7[39]},
      {stage4_7[27]}
   );
   gpc1_1 gpc8911 (
      {stage3_7[40]},
      {stage4_7[28]}
   );
   gpc1_1 gpc8912 (
      {stage3_7[41]},
      {stage4_7[29]}
   );
   gpc1_1 gpc8913 (
      {stage3_7[42]},
      {stage4_7[30]}
   );
   gpc1_1 gpc8914 (
      {stage3_7[43]},
      {stage4_7[31]}
   );
   gpc1_1 gpc8915 (
      {stage3_7[44]},
      {stage4_7[32]}
   );
   gpc1_1 gpc8916 (
      {stage3_7[45]},
      {stage4_7[33]}
   );
   gpc1_1 gpc8917 (
      {stage3_7[46]},
      {stage4_7[34]}
   );
   gpc1_1 gpc8918 (
      {stage3_7[47]},
      {stage4_7[35]}
   );
   gpc1_1 gpc8919 (
      {stage3_7[48]},
      {stage4_7[36]}
   );
   gpc1_1 gpc8920 (
      {stage3_7[49]},
      {stage4_7[37]}
   );
   gpc1_1 gpc8921 (
      {stage3_7[50]},
      {stage4_7[38]}
   );
   gpc1_1 gpc8922 (
      {stage3_10[84]},
      {stage4_10[26]}
   );
   gpc1_1 gpc8923 (
      {stage3_10[85]},
      {stage4_10[27]}
   );
   gpc1_1 gpc8924 (
      {stage3_10[86]},
      {stage4_10[28]}
   );
   gpc1_1 gpc8925 (
      {stage3_10[87]},
      {stage4_10[29]}
   );
   gpc1_1 gpc8926 (
      {stage3_10[88]},
      {stage4_10[30]}
   );
   gpc1_1 gpc8927 (
      {stage3_10[89]},
      {stage4_10[31]}
   );
   gpc1_1 gpc8928 (
      {stage3_10[90]},
      {stage4_10[32]}
   );
   gpc1_1 gpc8929 (
      {stage3_10[91]},
      {stage4_10[33]}
   );
   gpc1_1 gpc8930 (
      {stage3_10[92]},
      {stage4_10[34]}
   );
   gpc1_1 gpc8931 (
      {stage3_10[93]},
      {stage4_10[35]}
   );
   gpc1_1 gpc8932 (
      {stage3_10[94]},
      {stage4_10[36]}
   );
   gpc1_1 gpc8933 (
      {stage3_10[95]},
      {stage4_10[37]}
   );
   gpc1_1 gpc8934 (
      {stage3_10[96]},
      {stage4_10[38]}
   );
   gpc1_1 gpc8935 (
      {stage3_10[97]},
      {stage4_10[39]}
   );
   gpc1_1 gpc8936 (
      {stage3_10[98]},
      {stage4_10[40]}
   );
   gpc1_1 gpc8937 (
      {stage3_10[99]},
      {stage4_10[41]}
   );
   gpc1_1 gpc8938 (
      {stage3_12[67]},
      {stage4_12[23]}
   );
   gpc1_1 gpc8939 (
      {stage3_13[50]},
      {stage4_13[25]}
   );
   gpc1_1 gpc8940 (
      {stage3_13[51]},
      {stage4_13[26]}
   );
   gpc1_1 gpc8941 (
      {stage3_13[52]},
      {stage4_13[27]}
   );
   gpc1_1 gpc8942 (
      {stage3_13[53]},
      {stage4_13[28]}
   );
   gpc1_1 gpc8943 (
      {stage3_13[54]},
      {stage4_13[29]}
   );
   gpc1_1 gpc8944 (
      {stage3_13[55]},
      {stage4_13[30]}
   );
   gpc1_1 gpc8945 (
      {stage3_13[56]},
      {stage4_13[31]}
   );
   gpc1_1 gpc8946 (
      {stage3_14[30]},
      {stage4_14[28]}
   );
   gpc1_1 gpc8947 (
      {stage3_14[31]},
      {stage4_14[29]}
   );
   gpc1_1 gpc8948 (
      {stage3_15[47]},
      {stage4_15[14]}
   );
   gpc1_1 gpc8949 (
      {stage3_16[37]},
      {stage4_16[13]}
   );
   gpc1_1 gpc8950 (
      {stage3_16[38]},
      {stage4_16[14]}
   );
   gpc1_1 gpc8951 (
      {stage3_16[39]},
      {stage4_16[15]}
   );
   gpc1_1 gpc8952 (
      {stage3_16[40]},
      {stage4_16[16]}
   );
   gpc1_1 gpc8953 (
      {stage3_16[41]},
      {stage4_16[17]}
   );
   gpc1_1 gpc8954 (
      {stage3_16[42]},
      {stage4_16[18]}
   );
   gpc1_1 gpc8955 (
      {stage3_16[43]},
      {stage4_16[19]}
   );
   gpc1_1 gpc8956 (
      {stage3_16[44]},
      {stage4_16[20]}
   );
   gpc1_1 gpc8957 (
      {stage3_16[45]},
      {stage4_16[21]}
   );
   gpc1_1 gpc8958 (
      {stage3_16[46]},
      {stage4_16[22]}
   );
   gpc1_1 gpc8959 (
      {stage3_16[47]},
      {stage4_16[23]}
   );
   gpc1_1 gpc8960 (
      {stage3_16[48]},
      {stage4_16[24]}
   );
   gpc1_1 gpc8961 (
      {stage3_16[49]},
      {stage4_16[25]}
   );
   gpc1_1 gpc8962 (
      {stage3_16[50]},
      {stage4_16[26]}
   );
   gpc1_1 gpc8963 (
      {stage3_19[35]},
      {stage4_19[16]}
   );
   gpc1_1 gpc8964 (
      {stage3_19[36]},
      {stage4_19[17]}
   );
   gpc1_1 gpc8965 (
      {stage3_19[37]},
      {stage4_19[18]}
   );
   gpc1_1 gpc8966 (
      {stage3_19[38]},
      {stage4_19[19]}
   );
   gpc1_1 gpc8967 (
      {stage3_19[39]},
      {stage4_19[20]}
   );
   gpc1_1 gpc8968 (
      {stage3_19[40]},
      {stage4_19[21]}
   );
   gpc1_1 gpc8969 (
      {stage3_19[41]},
      {stage4_19[22]}
   );
   gpc1_1 gpc8970 (
      {stage3_19[42]},
      {stage4_19[23]}
   );
   gpc1_1 gpc8971 (
      {stage3_19[43]},
      {stage4_19[24]}
   );
   gpc1_1 gpc8972 (
      {stage3_19[44]},
      {stage4_19[25]}
   );
   gpc1_1 gpc8973 (
      {stage3_19[45]},
      {stage4_19[26]}
   );
   gpc1_1 gpc8974 (
      {stage3_19[46]},
      {stage4_19[27]}
   );
   gpc1_1 gpc8975 (
      {stage3_19[47]},
      {stage4_19[28]}
   );
   gpc1_1 gpc8976 (
      {stage3_20[73]},
      {stage4_20[24]}
   );
   gpc1_1 gpc8977 (
      {stage3_20[74]},
      {stage4_20[25]}
   );
   gpc1_1 gpc8978 (
      {stage3_20[75]},
      {stage4_20[26]}
   );
   gpc1_1 gpc8979 (
      {stage3_20[76]},
      {stage4_20[27]}
   );
   gpc1_1 gpc8980 (
      {stage3_20[77]},
      {stage4_20[28]}
   );
   gpc1_1 gpc8981 (
      {stage3_20[78]},
      {stage4_20[29]}
   );
   gpc1_1 gpc8982 (
      {stage3_20[79]},
      {stage4_20[30]}
   );
   gpc1_1 gpc8983 (
      {stage3_20[80]},
      {stage4_20[31]}
   );
   gpc1_1 gpc8984 (
      {stage3_20[81]},
      {stage4_20[32]}
   );
   gpc1_1 gpc8985 (
      {stage3_20[82]},
      {stage4_20[33]}
   );
   gpc1_1 gpc8986 (
      {stage3_21[30]},
      {stage4_21[28]}
   );
   gpc1_1 gpc8987 (
      {stage3_21[31]},
      {stage4_21[29]}
   );
   gpc1_1 gpc8988 (
      {stage3_21[32]},
      {stage4_21[30]}
   );
   gpc1_1 gpc8989 (
      {stage3_21[33]},
      {stage4_21[31]}
   );
   gpc1_1 gpc8990 (
      {stage3_21[34]},
      {stage4_21[32]}
   );
   gpc1_1 gpc8991 (
      {stage3_21[35]},
      {stage4_21[33]}
   );
   gpc1_1 gpc8992 (
      {stage3_21[36]},
      {stage4_21[34]}
   );
   gpc1_1 gpc8993 (
      {stage3_21[37]},
      {stage4_21[35]}
   );
   gpc1_1 gpc8994 (
      {stage3_21[38]},
      {stage4_21[36]}
   );
   gpc1_1 gpc8995 (
      {stage3_24[27]},
      {stage4_24[20]}
   );
   gpc1_1 gpc8996 (
      {stage3_24[28]},
      {stage4_24[21]}
   );
   gpc1_1 gpc8997 (
      {stage3_25[24]},
      {stage4_25[12]}
   );
   gpc1_1 gpc8998 (
      {stage3_25[25]},
      {stage4_25[13]}
   );
   gpc1_1 gpc8999 (
      {stage3_25[26]},
      {stage4_25[14]}
   );
   gpc1_1 gpc9000 (
      {stage3_25[27]},
      {stage4_25[15]}
   );
   gpc1_1 gpc9001 (
      {stage3_25[28]},
      {stage4_25[16]}
   );
   gpc1_1 gpc9002 (
      {stage3_25[29]},
      {stage4_25[17]}
   );
   gpc1_1 gpc9003 (
      {stage3_25[30]},
      {stage4_25[18]}
   );
   gpc1_1 gpc9004 (
      {stage3_25[31]},
      {stage4_25[19]}
   );
   gpc1_1 gpc9005 (
      {stage3_25[32]},
      {stage4_25[20]}
   );
   gpc1_1 gpc9006 (
      {stage3_27[38]},
      {stage4_27[16]}
   );
   gpc1_1 gpc9007 (
      {stage3_27[39]},
      {stage4_27[17]}
   );
   gpc1_1 gpc9008 (
      {stage3_27[40]},
      {stage4_27[18]}
   );
   gpc1_1 gpc9009 (
      {stage3_27[41]},
      {stage4_27[19]}
   );
   gpc1_1 gpc9010 (
      {stage3_27[42]},
      {stage4_27[20]}
   );
   gpc1_1 gpc9011 (
      {stage3_27[43]},
      {stage4_27[21]}
   );
   gpc1_1 gpc9012 (
      {stage3_27[44]},
      {stage4_27[22]}
   );
   gpc1_1 gpc9013 (
      {stage3_27[45]},
      {stage4_27[23]}
   );
   gpc1_1 gpc9014 (
      {stage3_27[46]},
      {stage4_27[24]}
   );
   gpc1_1 gpc9015 (
      {stage3_27[47]},
      {stage4_27[25]}
   );
   gpc1_1 gpc9016 (
      {stage3_27[48]},
      {stage4_27[26]}
   );
   gpc1_1 gpc9017 (
      {stage3_28[51]},
      {stage4_28[13]}
   );
   gpc1_1 gpc9018 (
      {stage3_28[52]},
      {stage4_28[14]}
   );
   gpc1_1 gpc9019 (
      {stage3_28[53]},
      {stage4_28[15]}
   );
   gpc1_1 gpc9020 (
      {stage3_28[54]},
      {stage4_28[16]}
   );
   gpc1_1 gpc9021 (
      {stage3_28[55]},
      {stage4_28[17]}
   );
   gpc1_1 gpc9022 (
      {stage3_28[56]},
      {stage4_28[18]}
   );
   gpc1_1 gpc9023 (
      {stage3_30[30]},
      {stage4_30[21]}
   );
   gpc1_1 gpc9024 (
      {stage3_30[31]},
      {stage4_30[22]}
   );
   gpc1_1 gpc9025 (
      {stage3_30[32]},
      {stage4_30[23]}
   );
   gpc1_1 gpc9026 (
      {stage3_30[33]},
      {stage4_30[24]}
   );
   gpc1_1 gpc9027 (
      {stage3_30[34]},
      {stage4_30[25]}
   );
   gpc1_1 gpc9028 (
      {stage3_30[35]},
      {stage4_30[26]}
   );
   gpc1_1 gpc9029 (
      {stage3_30[36]},
      {stage4_30[27]}
   );
   gpc1_1 gpc9030 (
      {stage3_30[37]},
      {stage4_30[28]}
   );
   gpc1_1 gpc9031 (
      {stage3_30[38]},
      {stage4_30[29]}
   );
   gpc1_1 gpc9032 (
      {stage3_30[39]},
      {stage4_30[30]}
   );
   gpc1_1 gpc9033 (
      {stage3_30[40]},
      {stage4_30[31]}
   );
   gpc1_1 gpc9034 (
      {stage3_30[41]},
      {stage4_30[32]}
   );
   gpc1_1 gpc9035 (
      {stage3_31[34]},
      {stage4_31[11]}
   );
   gpc1_1 gpc9036 (
      {stage3_31[35]},
      {stage4_31[12]}
   );
   gpc1_1 gpc9037 (
      {stage3_31[36]},
      {stage4_31[13]}
   );
   gpc1_1 gpc9038 (
      {stage3_31[37]},
      {stage4_31[14]}
   );
   gpc1_1 gpc9039 (
      {stage3_32[41]},
      {stage4_32[17]}
   );
   gpc1_1 gpc9040 (
      {stage3_32[42]},
      {stage4_32[18]}
   );
   gpc1_1 gpc9041 (
      {stage3_32[43]},
      {stage4_32[19]}
   );
   gpc1_1 gpc9042 (
      {stage3_32[44]},
      {stage4_32[20]}
   );
   gpc1_1 gpc9043 (
      {stage3_32[45]},
      {stage4_32[21]}
   );
   gpc1_1 gpc9044 (
      {stage3_32[46]},
      {stage4_32[22]}
   );
   gpc1_1 gpc9045 (
      {stage3_32[47]},
      {stage4_32[23]}
   );
   gpc1_1 gpc9046 (
      {stage3_32[48]},
      {stage4_32[24]}
   );
   gpc1_1 gpc9047 (
      {stage3_32[49]},
      {stage4_32[25]}
   );
   gpc1_1 gpc9048 (
      {stage3_32[50]},
      {stage4_32[26]}
   );
   gpc1_1 gpc9049 (
      {stage3_32[51]},
      {stage4_32[27]}
   );
   gpc1_1 gpc9050 (
      {stage3_32[52]},
      {stage4_32[28]}
   );
   gpc1_1 gpc9051 (
      {stage3_32[53]},
      {stage4_32[29]}
   );
   gpc1_1 gpc9052 (
      {stage3_33[37]},
      {stage4_33[20]}
   );
   gpc1_1 gpc9053 (
      {stage3_33[38]},
      {stage4_33[21]}
   );
   gpc1_1 gpc9054 (
      {stage3_33[39]},
      {stage4_33[22]}
   );
   gpc1_1 gpc9055 (
      {stage3_33[40]},
      {stage4_33[23]}
   );
   gpc1_1 gpc9056 (
      {stage3_33[41]},
      {stage4_33[24]}
   );
   gpc1_1 gpc9057 (
      {stage3_33[42]},
      {stage4_33[25]}
   );
   gpc1_1 gpc9058 (
      {stage3_33[43]},
      {stage4_33[26]}
   );
   gpc1_1 gpc9059 (
      {stage3_33[44]},
      {stage4_33[27]}
   );
   gpc1_1 gpc9060 (
      {stage3_33[45]},
      {stage4_33[28]}
   );
   gpc1_1 gpc9061 (
      {stage3_34[34]},
      {stage4_34[11]}
   );
   gpc1_1 gpc9062 (
      {stage3_34[35]},
      {stage4_34[12]}
   );
   gpc1_1 gpc9063 (
      {stage3_34[36]},
      {stage4_34[13]}
   );
   gpc1_1 gpc9064 (
      {stage3_34[37]},
      {stage4_34[14]}
   );
   gpc1_1 gpc9065 (
      {stage3_34[38]},
      {stage4_34[15]}
   );
   gpc1_1 gpc9066 (
      {stage3_34[39]},
      {stage4_34[16]}
   );
   gpc1_1 gpc9067 (
      {stage3_34[40]},
      {stage4_34[17]}
   );
   gpc1_1 gpc9068 (
      {stage3_34[41]},
      {stage4_34[18]}
   );
   gpc1_1 gpc9069 (
      {stage3_35[37]},
      {stage4_35[16]}
   );
   gpc1_1 gpc9070 (
      {stage3_35[38]},
      {stage4_35[17]}
   );
   gpc1_1 gpc9071 (
      {stage3_35[39]},
      {stage4_35[18]}
   );
   gpc1_1 gpc9072 (
      {stage3_35[40]},
      {stage4_35[19]}
   );
   gpc1_1 gpc9073 (
      {stage3_35[41]},
      {stage4_35[20]}
   );
   gpc1_1 gpc9074 (
      {stage3_35[42]},
      {stage4_35[21]}
   );
   gpc1_1 gpc9075 (
      {stage3_35[43]},
      {stage4_35[22]}
   );
   gpc1_1 gpc9076 (
      {stage3_35[44]},
      {stage4_35[23]}
   );
   gpc1_1 gpc9077 (
      {stage3_35[45]},
      {stage4_35[24]}
   );
   gpc1_1 gpc9078 (
      {stage3_35[46]},
      {stage4_35[25]}
   );
   gpc1_1 gpc9079 (
      {stage3_35[47]},
      {stage4_35[26]}
   );
   gpc1_1 gpc9080 (
      {stage3_35[48]},
      {stage4_35[27]}
   );
   gpc1_1 gpc9081 (
      {stage3_35[49]},
      {stage4_35[28]}
   );
   gpc1_1 gpc9082 (
      {stage3_35[50]},
      {stage4_35[29]}
   );
   gpc1_1 gpc9083 (
      {stage3_35[51]},
      {stage4_35[30]}
   );
   gpc1_1 gpc9084 (
      {stage3_35[52]},
      {stage4_35[31]}
   );
   gpc1_1 gpc9085 (
      {stage3_35[53]},
      {stage4_35[32]}
   );
   gpc1_1 gpc9086 (
      {stage3_35[54]},
      {stage4_35[33]}
   );
   gpc1_1 gpc9087 (
      {stage3_35[55]},
      {stage4_35[34]}
   );
   gpc1_1 gpc9088 (
      {stage3_35[56]},
      {stage4_35[35]}
   );
   gpc1_1 gpc9089 (
      {stage3_36[29]},
      {stage4_36[19]}
   );
   gpc1_1 gpc9090 (
      {stage3_36[30]},
      {stage4_36[20]}
   );
   gpc1_1 gpc9091 (
      {stage3_36[31]},
      {stage4_36[21]}
   );
   gpc1_1 gpc9092 (
      {stage3_36[32]},
      {stage4_36[22]}
   );
   gpc1_1 gpc9093 (
      {stage3_36[33]},
      {stage4_36[23]}
   );
   gpc1_1 gpc9094 (
      {stage3_36[34]},
      {stage4_36[24]}
   );
   gpc1_1 gpc9095 (
      {stage3_36[35]},
      {stage4_36[25]}
   );
   gpc1_1 gpc9096 (
      {stage3_36[36]},
      {stage4_36[26]}
   );
   gpc1_1 gpc9097 (
      {stage3_36[37]},
      {stage4_36[27]}
   );
   gpc1_1 gpc9098 (
      {stage3_36[38]},
      {stage4_36[28]}
   );
   gpc1_1 gpc9099 (
      {stage3_36[39]},
      {stage4_36[29]}
   );
   gpc1_1 gpc9100 (
      {stage3_36[40]},
      {stage4_36[30]}
   );
   gpc1_1 gpc9101 (
      {stage3_36[41]},
      {stage4_36[31]}
   );
   gpc1_1 gpc9102 (
      {stage3_36[42]},
      {stage4_36[32]}
   );
   gpc1_1 gpc9103 (
      {stage3_36[43]},
      {stage4_36[33]}
   );
   gpc1_1 gpc9104 (
      {stage3_36[44]},
      {stage4_36[34]}
   );
   gpc1_1 gpc9105 (
      {stage3_36[45]},
      {stage4_36[35]}
   );
   gpc1_1 gpc9106 (
      {stage3_37[48]},
      {stage4_37[13]}
   );
   gpc1_1 gpc9107 (
      {stage3_37[49]},
      {stage4_37[14]}
   );
   gpc1_1 gpc9108 (
      {stage3_37[50]},
      {stage4_37[15]}
   );
   gpc1_1 gpc9109 (
      {stage3_37[51]},
      {stage4_37[16]}
   );
   gpc1_1 gpc9110 (
      {stage3_37[52]},
      {stage4_37[17]}
   );
   gpc1_1 gpc9111 (
      {stage3_38[59]},
      {stage4_38[19]}
   );
   gpc1_1 gpc9112 (
      {stage3_40[43]},
      {stage4_40[19]}
   );
   gpc1_1 gpc9113 (
      {stage3_40[44]},
      {stage4_40[20]}
   );
   gpc1_1 gpc9114 (
      {stage3_40[45]},
      {stage4_40[21]}
   );
   gpc1_1 gpc9115 (
      {stage3_40[46]},
      {stage4_40[22]}
   );
   gpc1_1 gpc9116 (
      {stage3_40[47]},
      {stage4_40[23]}
   );
   gpc1_1 gpc9117 (
      {stage3_40[48]},
      {stage4_40[24]}
   );
   gpc1_1 gpc9118 (
      {stage3_40[49]},
      {stage4_40[25]}
   );
   gpc1_1 gpc9119 (
      {stage3_40[50]},
      {stage4_40[26]}
   );
   gpc1_1 gpc9120 (
      {stage3_40[51]},
      {stage4_40[27]}
   );
   gpc1_1 gpc9121 (
      {stage3_42[34]},
      {stage4_42[22]}
   );
   gpc1_1 gpc9122 (
      {stage3_42[35]},
      {stage4_42[23]}
   );
   gpc1_1 gpc9123 (
      {stage3_42[36]},
      {stage4_42[24]}
   );
   gpc1_1 gpc9124 (
      {stage3_42[37]},
      {stage4_42[25]}
   );
   gpc1_1 gpc9125 (
      {stage3_42[38]},
      {stage4_42[26]}
   );
   gpc1_1 gpc9126 (
      {stage3_42[39]},
      {stage4_42[27]}
   );
   gpc1_1 gpc9127 (
      {stage3_42[40]},
      {stage4_42[28]}
   );
   gpc1_1 gpc9128 (
      {stage3_42[41]},
      {stage4_42[29]}
   );
   gpc1_1 gpc9129 (
      {stage3_42[42]},
      {stage4_42[30]}
   );
   gpc1_1 gpc9130 (
      {stage3_42[43]},
      {stage4_42[31]}
   );
   gpc1_1 gpc9131 (
      {stage3_42[44]},
      {stage4_42[32]}
   );
   gpc1_1 gpc9132 (
      {stage3_42[45]},
      {stage4_42[33]}
   );
   gpc1_1 gpc9133 (
      {stage3_42[46]},
      {stage4_42[34]}
   );
   gpc1_1 gpc9134 (
      {stage3_42[47]},
      {stage4_42[35]}
   );
   gpc1_1 gpc9135 (
      {stage3_42[48]},
      {stage4_42[36]}
   );
   gpc1_1 gpc9136 (
      {stage3_42[49]},
      {stage4_42[37]}
   );
   gpc1_1 gpc9137 (
      {stage3_44[32]},
      {stage4_44[16]}
   );
   gpc1_1 gpc9138 (
      {stage3_44[33]},
      {stage4_44[17]}
   );
   gpc1_1 gpc9139 (
      {stage3_44[34]},
      {stage4_44[18]}
   );
   gpc1_1 gpc9140 (
      {stage3_44[35]},
      {stage4_44[19]}
   );
   gpc1_1 gpc9141 (
      {stage3_44[36]},
      {stage4_44[20]}
   );
   gpc1_1 gpc9142 (
      {stage3_44[37]},
      {stage4_44[21]}
   );
   gpc1_1 gpc9143 (
      {stage3_44[38]},
      {stage4_44[22]}
   );
   gpc1_1 gpc9144 (
      {stage3_44[39]},
      {stage4_44[23]}
   );
   gpc1_1 gpc9145 (
      {stage3_44[40]},
      {stage4_44[24]}
   );
   gpc1_1 gpc9146 (
      {stage3_45[34]},
      {stage4_45[19]}
   );
   gpc1_1 gpc9147 (
      {stage3_45[35]},
      {stage4_45[20]}
   );
   gpc1_1 gpc9148 (
      {stage3_45[36]},
      {stage4_45[21]}
   );
   gpc1_1 gpc9149 (
      {stage3_45[37]},
      {stage4_45[22]}
   );
   gpc1_1 gpc9150 (
      {stage3_45[38]},
      {stage4_45[23]}
   );
   gpc1_1 gpc9151 (
      {stage3_45[39]},
      {stage4_45[24]}
   );
   gpc1_1 gpc9152 (
      {stage3_45[40]},
      {stage4_45[25]}
   );
   gpc1_1 gpc9153 (
      {stage3_45[41]},
      {stage4_45[26]}
   );
   gpc1_1 gpc9154 (
      {stage3_45[42]},
      {stage4_45[27]}
   );
   gpc1_1 gpc9155 (
      {stage3_45[43]},
      {stage4_45[28]}
   );
   gpc1_1 gpc9156 (
      {stage3_46[57]},
      {stage4_46[16]}
   );
   gpc1_1 gpc9157 (
      {stage3_48[37]},
      {stage4_48[18]}
   );
   gpc1_1 gpc9158 (
      {stage3_48[38]},
      {stage4_48[19]}
   );
   gpc1_1 gpc9159 (
      {stage3_48[39]},
      {stage4_48[20]}
   );
   gpc1_1 gpc9160 (
      {stage3_48[40]},
      {stage4_48[21]}
   );
   gpc1_1 gpc9161 (
      {stage3_48[41]},
      {stage4_48[22]}
   );
   gpc1_1 gpc9162 (
      {stage3_51[50]},
      {stage4_51[23]}
   );
   gpc1_1 gpc9163 (
      {stage3_51[51]},
      {stage4_51[24]}
   );
   gpc1_1 gpc9164 (
      {stage3_51[52]},
      {stage4_51[25]}
   );
   gpc1_1 gpc9165 (
      {stage3_51[53]},
      {stage4_51[26]}
   );
   gpc1_1 gpc9166 (
      {stage3_51[54]},
      {stage4_51[27]}
   );
   gpc1_1 gpc9167 (
      {stage3_51[55]},
      {stage4_51[28]}
   );
   gpc1_1 gpc9168 (
      {stage3_51[56]},
      {stage4_51[29]}
   );
   gpc1_1 gpc9169 (
      {stage3_51[57]},
      {stage4_51[30]}
   );
   gpc1_1 gpc9170 (
      {stage3_51[58]},
      {stage4_51[31]}
   );
   gpc1_1 gpc9171 (
      {stage3_51[59]},
      {stage4_51[32]}
   );
   gpc1_1 gpc9172 (
      {stage3_51[60]},
      {stage4_51[33]}
   );
   gpc1_1 gpc9173 (
      {stage3_51[61]},
      {stage4_51[34]}
   );
   gpc1_1 gpc9174 (
      {stage3_51[62]},
      {stage4_51[35]}
   );
   gpc1_1 gpc9175 (
      {stage3_52[61]},
      {stage4_52[17]}
   );
   gpc1_1 gpc9176 (
      {stage3_52[62]},
      {stage4_52[18]}
   );
   gpc1_1 gpc9177 (
      {stage3_53[55]},
      {stage4_53[24]}
   );
   gpc1_1 gpc9178 (
      {stage3_53[56]},
      {stage4_53[25]}
   );
   gpc1_1 gpc9179 (
      {stage3_53[57]},
      {stage4_53[26]}
   );
   gpc1_1 gpc9180 (
      {stage3_53[58]},
      {stage4_53[27]}
   );
   gpc1_1 gpc9181 (
      {stage3_53[59]},
      {stage4_53[28]}
   );
   gpc1_1 gpc9182 (
      {stage3_53[60]},
      {stage4_53[29]}
   );
   gpc1_1 gpc9183 (
      {stage3_53[61]},
      {stage4_53[30]}
   );
   gpc1_1 gpc9184 (
      {stage3_53[62]},
      {stage4_53[31]}
   );
   gpc1_1 gpc9185 (
      {stage3_53[63]},
      {stage4_53[32]}
   );
   gpc1_1 gpc9186 (
      {stage3_53[64]},
      {stage4_53[33]}
   );
   gpc1_1 gpc9187 (
      {stage3_53[65]},
      {stage4_53[34]}
   );
   gpc1_1 gpc9188 (
      {stage3_53[66]},
      {stage4_53[35]}
   );
   gpc1_1 gpc9189 (
      {stage3_53[67]},
      {stage4_53[36]}
   );
   gpc1_1 gpc9190 (
      {stage3_53[68]},
      {stage4_53[37]}
   );
   gpc1_1 gpc9191 (
      {stage3_53[69]},
      {stage4_53[38]}
   );
   gpc1_1 gpc9192 (
      {stage3_53[70]},
      {stage4_53[39]}
   );
   gpc1_1 gpc9193 (
      {stage3_53[71]},
      {stage4_53[40]}
   );
   gpc1_1 gpc9194 (
      {stage3_53[72]},
      {stage4_53[41]}
   );
   gpc1_1 gpc9195 (
      {stage3_53[73]},
      {stage4_53[42]}
   );
   gpc1_1 gpc9196 (
      {stage3_53[74]},
      {stage4_53[43]}
   );
   gpc1_1 gpc9197 (
      {stage3_55[47]},
      {stage4_55[19]}
   );
   gpc1_1 gpc9198 (
      {stage3_55[48]},
      {stage4_55[20]}
   );
   gpc1_1 gpc9199 (
      {stage3_55[49]},
      {stage4_55[21]}
   );
   gpc1_1 gpc9200 (
      {stage3_55[50]},
      {stage4_55[22]}
   );
   gpc1_1 gpc9201 (
      {stage3_55[51]},
      {stage4_55[23]}
   );
   gpc1_1 gpc9202 (
      {stage3_55[52]},
      {stage4_55[24]}
   );
   gpc1_1 gpc9203 (
      {stage3_55[53]},
      {stage4_55[25]}
   );
   gpc1_1 gpc9204 (
      {stage3_55[54]},
      {stage4_55[26]}
   );
   gpc1_1 gpc9205 (
      {stage3_55[55]},
      {stage4_55[27]}
   );
   gpc1_1 gpc9206 (
      {stage3_55[56]},
      {stage4_55[28]}
   );
   gpc1_1 gpc9207 (
      {stage3_55[57]},
      {stage4_55[29]}
   );
   gpc1_1 gpc9208 (
      {stage3_55[58]},
      {stage4_55[30]}
   );
   gpc1_1 gpc9209 (
      {stage3_55[59]},
      {stage4_55[31]}
   );
   gpc1_1 gpc9210 (
      {stage3_55[60]},
      {stage4_55[32]}
   );
   gpc1_1 gpc9211 (
      {stage3_55[61]},
      {stage4_55[33]}
   );
   gpc1_1 gpc9212 (
      {stage3_55[62]},
      {stage4_55[34]}
   );
   gpc1_1 gpc9213 (
      {stage3_55[63]},
      {stage4_55[35]}
   );
   gpc1_1 gpc9214 (
      {stage3_55[64]},
      {stage4_55[36]}
   );
   gpc1_1 gpc9215 (
      {stage3_55[65]},
      {stage4_55[37]}
   );
   gpc1_1 gpc9216 (
      {stage3_55[66]},
      {stage4_55[38]}
   );
   gpc1_1 gpc9217 (
      {stage3_56[30]},
      {stage4_56[12]}
   );
   gpc1_1 gpc9218 (
      {stage3_56[31]},
      {stage4_56[13]}
   );
   gpc1_1 gpc9219 (
      {stage3_58[57]},
      {stage4_58[19]}
   );
   gpc1_1 gpc9220 (
      {stage3_58[58]},
      {stage4_58[20]}
   );
   gpc1_1 gpc9221 (
      {stage3_58[59]},
      {stage4_58[21]}
   );
   gpc1_1 gpc9222 (
      {stage3_58[60]},
      {stage4_58[22]}
   );
   gpc1_1 gpc9223 (
      {stage3_58[61]},
      {stage4_58[23]}
   );
   gpc1_1 gpc9224 (
      {stage3_59[44]},
      {stage4_59[15]}
   );
   gpc1_1 gpc9225 (
      {stage3_59[45]},
      {stage4_59[16]}
   );
   gpc1_1 gpc9226 (
      {stage3_59[46]},
      {stage4_59[17]}
   );
   gpc1_1 gpc9227 (
      {stage3_59[47]},
      {stage4_59[18]}
   );
   gpc1_1 gpc9228 (
      {stage3_59[48]},
      {stage4_59[19]}
   );
   gpc1_1 gpc9229 (
      {stage3_59[49]},
      {stage4_59[20]}
   );
   gpc1_1 gpc9230 (
      {stage3_60[40]},
      {stage4_60[20]}
   );
   gpc1_1 gpc9231 (
      {stage3_60[41]},
      {stage4_60[21]}
   );
   gpc1_1 gpc9232 (
      {stage3_61[48]},
      {stage4_61[27]}
   );
   gpc1_1 gpc9233 (
      {stage3_61[49]},
      {stage4_61[28]}
   );
   gpc1_1 gpc9234 (
      {stage3_61[50]},
      {stage4_61[29]}
   );
   gpc1_1 gpc9235 (
      {stage3_61[51]},
      {stage4_61[30]}
   );
   gpc1_1 gpc9236 (
      {stage3_61[52]},
      {stage4_61[31]}
   );
   gpc1_1 gpc9237 (
      {stage3_62[30]},
      {stage4_62[13]}
   );
   gpc1_1 gpc9238 (
      {stage3_62[31]},
      {stage4_62[14]}
   );
   gpc1_1 gpc9239 (
      {stage3_62[32]},
      {stage4_62[15]}
   );
   gpc1_1 gpc9240 (
      {stage3_62[33]},
      {stage4_62[16]}
   );
   gpc1_1 gpc9241 (
      {stage3_64[36]},
      {stage4_64[19]}
   );
   gpc1_1 gpc9242 (
      {stage3_64[37]},
      {stage4_64[20]}
   );
   gpc1_1 gpc9243 (
      {stage3_64[38]},
      {stage4_64[21]}
   );
   gpc1_1 gpc9244 (
      {stage3_64[39]},
      {stage4_64[22]}
   );
   gpc1_1 gpc9245 (
      {stage3_64[40]},
      {stage4_64[23]}
   );
   gpc1_1 gpc9246 (
      {stage3_64[41]},
      {stage4_64[24]}
   );
   gpc1_1 gpc9247 (
      {stage3_64[42]},
      {stage4_64[25]}
   );
   gpc1_1 gpc9248 (
      {stage3_64[43]},
      {stage4_64[26]}
   );
   gpc1_1 gpc9249 (
      {stage3_64[44]},
      {stage4_64[27]}
   );
   gpc1_1 gpc9250 (
      {stage3_64[45]},
      {stage4_64[28]}
   );
   gpc1_1 gpc9251 (
      {stage3_64[46]},
      {stage4_64[29]}
   );
   gpc1_1 gpc9252 (
      {stage3_64[47]},
      {stage4_64[30]}
   );
   gpc1_1 gpc9253 (
      {stage3_64[48]},
      {stage4_64[31]}
   );
   gpc1_1 gpc9254 (
      {stage3_64[49]},
      {stage4_64[32]}
   );
   gpc1_1 gpc9255 (
      {stage3_64[50]},
      {stage4_64[33]}
   );
   gpc1_1 gpc9256 (
      {stage3_65[18]},
      {stage4_65[16]}
   );
   gpc1_1 gpc9257 (
      {stage3_65[19]},
      {stage4_65[17]}
   );
   gpc1_1 gpc9258 (
      {stage3_65[20]},
      {stage4_65[18]}
   );
   gpc1_1 gpc9259 (
      {stage3_65[21]},
      {stage4_65[19]}
   );
   gpc1_1 gpc9260 (
      {stage3_65[22]},
      {stage4_65[20]}
   );
   gpc1_1 gpc9261 (
      {stage3_65[23]},
      {stage4_65[21]}
   );
   gpc1_1 gpc9262 (
      {stage3_65[24]},
      {stage4_65[22]}
   );
   gpc1_1 gpc9263 (
      {stage3_65[25]},
      {stage4_65[23]}
   );
   gpc1_1 gpc9264 (
      {stage3_65[26]},
      {stage4_65[24]}
   );
   gpc1_1 gpc9265 (
      {stage3_65[27]},
      {stage4_65[25]}
   );
   gpc1_1 gpc9266 (
      {stage3_65[28]},
      {stage4_65[26]}
   );
   gpc1_1 gpc9267 (
      {stage3_65[29]},
      {stage4_65[27]}
   );
   gpc1_1 gpc9268 (
      {stage3_65[30]},
      {stage4_65[28]}
   );
   gpc1_1 gpc9269 (
      {stage3_65[31]},
      {stage4_65[29]}
   );
   gpc1_1 gpc9270 (
      {stage3_65[32]},
      {stage4_65[30]}
   );
   gpc1_1 gpc9271 (
      {stage3_65[33]},
      {stage4_65[31]}
   );
   gpc1_1 gpc9272 (
      {stage3_65[34]},
      {stage4_65[32]}
   );
   gpc1_1 gpc9273 (
      {stage3_65[35]},
      {stage4_65[33]}
   );
   gpc1_1 gpc9274 (
      {stage3_65[36]},
      {stage4_65[34]}
   );
   gpc1_1 gpc9275 (
      {stage3_65[37]},
      {stage4_65[35]}
   );
   gpc1_1 gpc9276 (
      {stage3_66[36]},
      {stage4_66[9]}
   );
   gpc1_1 gpc9277 (
      {stage3_66[37]},
      {stage4_66[10]}
   );
   gpc1_1 gpc9278 (
      {stage3_67[12]},
      {stage4_67[9]}
   );
   gpc1_1 gpc9279 (
      {stage3_67[13]},
      {stage4_67[10]}
   );
   gpc1_1 gpc9280 (
      {stage3_68[0]},
      {stage4_68[8]}
   );
   gpc1_1 gpc9281 (
      {stage3_68[1]},
      {stage4_68[9]}
   );
   gpc1_1 gpc9282 (
      {stage3_68[2]},
      {stage4_68[10]}
   );
   gpc1_1 gpc9283 (
      {stage3_68[3]},
      {stage4_68[11]}
   );
   gpc1_1 gpc9284 (
      {stage3_68[4]},
      {stage4_68[12]}
   );
   gpc1_1 gpc9285 (
      {stage3_68[5]},
      {stage4_68[13]}
   );
   gpc615_5 gpc9286 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc9287 (
      {stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1163_5 gpc9288 (
      {stage4_2[6], stage4_2[7], stage4_2[8]},
      {stage4_3[6], stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[0]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[1],stage5_4[2],stage5_3[2],stage5_2[2]}
   );
   gpc1163_5 gpc9289 (
      {stage4_4[1], stage4_4[2], stage4_4[3]},
      {stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6]},
      {stage4_6[0]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[2],stage5_4[3]}
   );
   gpc606_5 gpc9290 (
      {stage4_4[4], stage4_4[5], stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9]},
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6]},
      {stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[3],stage5_4[4]}
   );
   gpc606_5 gpc9291 (
      {stage4_4[10], stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15]},
      {stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12]},
      {stage5_8[2],stage5_7[2],stage5_6[3],stage5_5[4],stage5_4[5]}
   );
   gpc606_5 gpc9292 (
      {stage4_4[16], stage4_4[17], stage4_4[18], stage4_4[19], stage4_4[20], stage4_4[21]},
      {stage4_6[13], stage4_6[14], stage4_6[15], stage4_6[16], stage4_6[17], stage4_6[18]},
      {stage5_8[3],stage5_7[3],stage5_6[4],stage5_5[5],stage5_4[6]}
   );
   gpc606_5 gpc9293 (
      {stage4_4[22], stage4_4[23], stage4_4[24], stage4_4[25], stage4_4[26], stage4_4[27]},
      {stage4_6[19], stage4_6[20], stage4_6[21], stage4_6[22], stage4_6[23], 1'b0},
      {stage5_8[4],stage5_7[4],stage5_6[5],stage5_5[6],stage5_4[7]}
   );
   gpc606_5 gpc9294 (
      {stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12]},
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6]},
      {stage5_9[0],stage5_8[5],stage5_7[5],stage5_6[6],stage5_5[7]}
   );
   gpc606_5 gpc9295 (
      {stage4_5[13], stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17], stage4_5[18]},
      {stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11], stage4_7[12]},
      {stage5_9[1],stage5_8[6],stage5_7[6],stage5_6[7],stage5_5[8]}
   );
   gpc606_5 gpc9296 (
      {stage4_5[19], stage4_5[20], stage4_5[21], stage4_5[22], stage4_5[23], stage4_5[24]},
      {stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17], stage4_7[18]},
      {stage5_9[2],stage5_8[7],stage5_7[7],stage5_6[8],stage5_5[9]}
   );
   gpc606_5 gpc9297 (
      {stage4_5[25], stage4_5[26], stage4_5[27], stage4_5[28], stage4_5[29], stage4_5[30]},
      {stage4_7[19], stage4_7[20], stage4_7[21], stage4_7[22], stage4_7[23], stage4_7[24]},
      {stage5_9[3],stage5_8[8],stage5_7[8],stage5_6[9],stage5_5[10]}
   );
   gpc207_4 gpc9298 (
      {stage4_7[25], stage4_7[26], stage4_7[27], stage4_7[28], stage4_7[29], stage4_7[30], stage4_7[31]},
      {stage4_9[0], stage4_9[1]},
      {stage5_10[0],stage5_9[4],stage5_8[9],stage5_7[9]}
   );
   gpc207_4 gpc9299 (
      {stage4_7[32], stage4_7[33], stage4_7[34], stage4_7[35], stage4_7[36], stage4_7[37], stage4_7[38]},
      {stage4_9[2], stage4_9[3]},
      {stage5_10[1],stage5_9[5],stage5_8[10],stage5_7[10]}
   );
   gpc135_4 gpc9300 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[2],stage5_9[6],stage5_8[11]}
   );
   gpc117_4 gpc9301 (
      {stage4_8[5], stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11]},
      {stage4_9[7]},
      {stage4_10[1]},
      {stage5_11[1],stage5_10[3],stage5_9[7],stage5_8[12]}
   );
   gpc606_5 gpc9302 (
      {stage4_8[12], stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17]},
      {stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[8],stage5_8[13]}
   );
   gpc606_5 gpc9303 (
      {stage4_8[18], stage4_8[19], stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23]},
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13]},
      {stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[9],stage5_8[14]}
   );
   gpc606_5 gpc9304 (
      {stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11], stage4_9[12], stage4_9[13]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[2],stage5_11[4],stage5_10[6],stage5_9[10]}
   );
   gpc2135_5 gpc9305 (
      {stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17], stage4_10[18]},
      {stage4_11[6], stage4_11[7], stage4_11[8]},
      {stage4_12[0]},
      {stage4_13[0], stage4_13[1]},
      {stage5_14[0],stage5_13[1],stage5_12[3],stage5_11[5],stage5_10[7]}
   );
   gpc606_5 gpc9306 (
      {stage4_10[19], stage4_10[20], stage4_10[21], stage4_10[22], stage4_10[23], stage4_10[24]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6]},
      {stage5_14[1],stage5_13[2],stage5_12[4],stage5_11[6],stage5_10[8]}
   );
   gpc606_5 gpc9307 (
      {stage4_10[25], stage4_10[26], stage4_10[27], stage4_10[28], stage4_10[29], stage4_10[30]},
      {stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11], stage4_12[12]},
      {stage5_14[2],stage5_13[3],stage5_12[5],stage5_11[7],stage5_10[9]}
   );
   gpc615_5 gpc9308 (
      {stage4_11[9], stage4_11[10], stage4_11[11], stage4_11[12], stage4_11[13]},
      {stage4_12[13]},
      {stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6], stage4_13[7]},
      {stage5_15[0],stage5_14[3],stage5_13[4],stage5_12[6],stage5_11[8]}
   );
   gpc615_5 gpc9309 (
      {stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17], stage4_11[18]},
      {stage4_12[14]},
      {stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13]},
      {stage5_15[1],stage5_14[4],stage5_13[5],stage5_12[7],stage5_11[9]}
   );
   gpc615_5 gpc9310 (
      {stage4_11[19], stage4_11[20], stage4_11[21], stage4_11[22], stage4_11[23]},
      {stage4_12[15]},
      {stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], stage4_13[19]},
      {stage5_15[2],stage5_14[5],stage5_13[6],stage5_12[8],stage5_11[10]}
   );
   gpc623_5 gpc9311 (
      {stage4_11[24], stage4_11[25], stage4_11[26]},
      {stage4_12[16], stage4_12[17]},
      {stage4_13[20], stage4_13[21], stage4_13[22], stage4_13[23], stage4_13[24], stage4_13[25]},
      {stage5_15[3],stage5_14[6],stage5_13[7],stage5_12[9],stage5_11[11]}
   );
   gpc606_5 gpc9312 (
      {stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21], stage4_12[22], stage4_12[23]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[4],stage5_14[7],stage5_13[8],stage5_12[10]}
   );
   gpc615_5 gpc9313 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[5],stage5_14[8]}
   );
   gpc615_5 gpc9314 (
      {stage4_14[11], stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15]},
      {stage4_15[1]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[1],stage5_16[2],stage5_15[6],stage5_14[9]}
   );
   gpc615_5 gpc9315 (
      {stage4_14[16], stage4_14[17], stage4_14[18], stage4_14[19], stage4_14[20]},
      {stage4_15[2]},
      {stage4_16[12], stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17]},
      {stage5_18[2],stage5_17[2],stage5_16[3],stage5_15[7],stage5_14[10]}
   );
   gpc615_5 gpc9316 (
      {stage4_14[21], stage4_14[22], stage4_14[23], stage4_14[24], stage4_14[25]},
      {stage4_15[3]},
      {stage4_16[18], stage4_16[19], stage4_16[20], stage4_16[21], stage4_16[22], stage4_16[23]},
      {stage5_18[3],stage5_17[3],stage5_16[4],stage5_15[8],stage5_14[11]}
   );
   gpc615_5 gpc9317 (
      {stage4_15[4], stage4_15[5], stage4_15[6], stage4_15[7], stage4_15[8]},
      {stage4_16[24]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[4],stage5_17[4],stage5_16[5],stage5_15[9]}
   );
   gpc615_5 gpc9318 (
      {stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12], stage4_15[13]},
      {stage4_16[25]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[5],stage5_17[5],stage5_16[6],stage5_15[10]}
   );
   gpc615_5 gpc9319 (
      {stage4_15[14], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage4_16[26]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[6],stage5_17[6],stage5_16[7],stage5_15[11]}
   );
   gpc615_5 gpc9320 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4]},
      {stage4_19[0]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[0],stage5_20[0],stage5_19[3],stage5_18[7]}
   );
   gpc615_5 gpc9321 (
      {stage4_18[5], stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9]},
      {stage4_19[1]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], stage4_20[11]},
      {stage5_22[1],stage5_21[1],stage5_20[1],stage5_19[4],stage5_18[8]}
   );
   gpc615_5 gpc9322 (
      {stage4_18[10], stage4_18[11], stage4_18[12], stage4_18[13], stage4_18[14]},
      {stage4_19[2]},
      {stage4_20[12], stage4_20[13], stage4_20[14], stage4_20[15], stage4_20[16], stage4_20[17]},
      {stage5_22[2],stage5_21[2],stage5_20[2],stage5_19[5],stage5_18[9]}
   );
   gpc615_5 gpc9323 (
      {stage4_18[15], stage4_18[16], stage4_18[17], stage4_18[18], stage4_18[19]},
      {stage4_19[3]},
      {stage4_20[18], stage4_20[19], stage4_20[20], stage4_20[21], stage4_20[22], stage4_20[23]},
      {stage5_22[3],stage5_21[3],stage5_20[3],stage5_19[6],stage5_18[10]}
   );
   gpc615_5 gpc9324 (
      {stage4_19[4], stage4_19[5], stage4_19[6], stage4_19[7], stage4_19[8]},
      {stage4_20[24]},
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5]},
      {stage5_23[0],stage5_22[4],stage5_21[4],stage5_20[4],stage5_19[7]}
   );
   gpc615_5 gpc9325 (
      {stage4_19[9], stage4_19[10], stage4_19[11], stage4_19[12], stage4_19[13]},
      {stage4_20[25]},
      {stage4_21[6], stage4_21[7], stage4_21[8], stage4_21[9], stage4_21[10], stage4_21[11]},
      {stage5_23[1],stage5_22[5],stage5_21[5],stage5_20[5],stage5_19[8]}
   );
   gpc615_5 gpc9326 (
      {stage4_19[14], stage4_19[15], stage4_19[16], stage4_19[17], stage4_19[18]},
      {stage4_20[26]},
      {stage4_21[12], stage4_21[13], stage4_21[14], stage4_21[15], stage4_21[16], stage4_21[17]},
      {stage5_23[2],stage5_22[6],stage5_21[6],stage5_20[6],stage5_19[9]}
   );
   gpc615_5 gpc9327 (
      {stage4_19[19], stage4_19[20], stage4_19[21], stage4_19[22], stage4_19[23]},
      {stage4_20[27]},
      {stage4_21[18], stage4_21[19], stage4_21[20], stage4_21[21], stage4_21[22], stage4_21[23]},
      {stage5_23[3],stage5_22[7],stage5_21[7],stage5_20[7],stage5_19[10]}
   );
   gpc606_5 gpc9328 (
      {stage4_21[24], stage4_21[25], stage4_21[26], stage4_21[27], stage4_21[28], stage4_21[29]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage5_25[0],stage5_24[0],stage5_23[4],stage5_22[8],stage5_21[8]}
   );
   gpc606_5 gpc9329 (
      {stage4_21[30], stage4_21[31], stage4_21[32], stage4_21[33], stage4_21[34], stage4_21[35]},
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10], stage4_23[11]},
      {stage5_25[1],stage5_24[1],stage5_23[5],stage5_22[9],stage5_21[9]}
   );
   gpc1163_5 gpc9330 (
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[12], stage4_23[13], stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17]},
      {stage4_24[0]},
      {stage4_25[0]},
      {stage5_26[0],stage5_25[2],stage5_24[2],stage5_23[6],stage5_22[10]}
   );
   gpc615_5 gpc9331 (
      {stage4_22[3], stage4_22[4], stage4_22[5], stage4_22[6], stage4_22[7]},
      {stage4_23[18]},
      {stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6]},
      {stage5_26[1],stage5_25[3],stage5_24[3],stage5_23[7],stage5_22[11]}
   );
   gpc615_5 gpc9332 (
      {stage4_22[8], stage4_22[9], stage4_22[10], stage4_22[11], stage4_22[12]},
      {stage4_23[19]},
      {stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11], stage4_24[12]},
      {stage5_26[2],stage5_25[4],stage5_24[4],stage5_23[8],stage5_22[12]}
   );
   gpc615_5 gpc9333 (
      {stage4_22[13], stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17]},
      {stage4_23[20]},
      {stage4_24[13], stage4_24[14], stage4_24[15], stage4_24[16], stage4_24[17], stage4_24[18]},
      {stage5_26[3],stage5_25[5],stage5_24[5],stage5_23[9],stage5_22[13]}
   );
   gpc606_5 gpc9334 (
      {stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5], stage4_25[6]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage5_29[0],stage5_28[0],stage5_27[0],stage5_26[4],stage5_25[6]}
   );
   gpc606_5 gpc9335 (
      {stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11], stage4_25[12]},
      {stage4_27[6], stage4_27[7], stage4_27[8], stage4_27[9], stage4_27[10], stage4_27[11]},
      {stage5_29[1],stage5_28[1],stage5_27[1],stage5_26[5],stage5_25[7]}
   );
   gpc606_5 gpc9336 (
      {stage4_25[13], stage4_25[14], stage4_25[15], stage4_25[16], stage4_25[17], stage4_25[18]},
      {stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16], stage4_27[17]},
      {stage5_29[2],stage5_28[2],stage5_27[2],stage5_26[6],stage5_25[8]}
   );
   gpc623_5 gpc9337 (
      {stage4_25[19], stage4_25[20], 1'b0},
      {stage4_26[0], stage4_26[1]},
      {stage4_27[18], stage4_27[19], stage4_27[20], stage4_27[21], stage4_27[22], stage4_27[23]},
      {stage5_29[3],stage5_28[3],stage5_27[3],stage5_26[7],stage5_25[9]}
   );
   gpc2135_5 gpc9338 (
      {stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5], stage4_26[6]},
      {stage4_27[24], stage4_27[25], stage4_27[26]},
      {stage4_28[0]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[0],stage5_29[4],stage5_28[4],stage5_27[4],stage5_26[8]}
   );
   gpc117_4 gpc9339 (
      {stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11], stage4_26[12], stage4_26[13]},
      {1'b0},
      {stage4_28[1]},
      {stage5_29[5],stage5_28[5],stage5_27[5],stage5_26[9]}
   );
   gpc606_5 gpc9340 (
      {stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5], stage4_28[6], stage4_28[7]},
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage5_32[0],stage5_31[0],stage5_30[1],stage5_29[6],stage5_28[6]}
   );
   gpc615_5 gpc9341 (
      {stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11], stage4_28[12]},
      {stage4_29[2]},
      {stage4_30[6], stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage5_32[1],stage5_31[1],stage5_30[2],stage5_29[7],stage5_28[7]}
   );
   gpc615_5 gpc9342 (
      {stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage4_29[3]},
      {stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15], stage4_30[16], stage4_30[17]},
      {stage5_32[2],stage5_31[2],stage5_30[3],stage5_29[8],stage5_28[8]}
   );
   gpc117_4 gpc9343 (
      {stage4_29[4], stage4_29[5], stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10]},
      {stage4_30[18]},
      {stage4_31[0]},
      {stage5_32[3],stage5_31[3],stage5_30[4],stage5_29[9]}
   );
   gpc117_4 gpc9344 (
      {stage4_29[11], stage4_29[12], stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17]},
      {stage4_30[19]},
      {stage4_31[1]},
      {stage5_32[4],stage5_31[4],stage5_30[5],stage5_29[10]}
   );
   gpc615_5 gpc9345 (
      {stage4_30[20], stage4_30[21], stage4_30[22], stage4_30[23], stage4_30[24]},
      {stage4_31[2]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[0],stage5_32[5],stage5_31[5],stage5_30[6]}
   );
   gpc615_5 gpc9346 (
      {stage4_30[25], stage4_30[26], stage4_30[27], stage4_30[28], stage4_30[29]},
      {stage4_31[3]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[1],stage5_32[6],stage5_31[6],stage5_30[7]}
   );
   gpc615_5 gpc9347 (
      {stage4_30[30], stage4_30[31], stage4_30[32], 1'b0, 1'b0},
      {stage4_31[4]},
      {stage4_32[12], stage4_32[13], stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17]},
      {stage5_34[2],stage5_33[2],stage5_32[7],stage5_31[7],stage5_30[8]}
   );
   gpc615_5 gpc9348 (
      {stage4_31[5], stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9]},
      {stage4_32[18]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[3],stage5_33[3],stage5_32[8],stage5_31[8]}
   );
   gpc615_5 gpc9349 (
      {stage4_31[10], stage4_31[11], stage4_31[12], stage4_31[13], stage4_31[14]},
      {stage4_32[19]},
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage5_35[1],stage5_34[4],stage5_33[4],stage5_32[9],stage5_31[9]}
   );
   gpc606_5 gpc9350 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], stage4_33[17]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[0],stage5_35[2],stage5_34[5],stage5_33[5]}
   );
   gpc606_5 gpc9351 (
      {stage4_33[18], stage4_33[19], stage4_33[20], stage4_33[21], stage4_33[22], stage4_33[23]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[1],stage5_35[3],stage5_34[6],stage5_33[6]}
   );
   gpc135_4 gpc9352 (
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4]},
      {stage4_35[12], stage4_35[13], stage4_35[14]},
      {stage4_36[0]},
      {stage5_37[2],stage5_36[2],stage5_35[4],stage5_34[7]}
   );
   gpc615_5 gpc9353 (
      {stage4_34[5], stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9]},
      {stage4_35[15]},
      {stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5], stage4_36[6]},
      {stage5_38[0],stage5_37[3],stage5_36[3],stage5_35[5],stage5_34[8]}
   );
   gpc615_5 gpc9354 (
      {stage4_34[10], stage4_34[11], stage4_34[12], stage4_34[13], stage4_34[14]},
      {stage4_35[16]},
      {stage4_36[7], stage4_36[8], stage4_36[9], stage4_36[10], stage4_36[11], stage4_36[12]},
      {stage5_38[1],stage5_37[4],stage5_36[4],stage5_35[6],stage5_34[9]}
   );
   gpc615_5 gpc9355 (
      {stage4_35[17], stage4_35[18], stage4_35[19], stage4_35[20], stage4_35[21]},
      {stage4_36[13]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage5_39[0],stage5_38[2],stage5_37[5],stage5_36[5],stage5_35[7]}
   );
   gpc615_5 gpc9356 (
      {stage4_35[22], stage4_35[23], stage4_35[24], stage4_35[25], stage4_35[26]},
      {stage4_36[14]},
      {stage4_37[6], stage4_37[7], stage4_37[8], stage4_37[9], stage4_37[10], stage4_37[11]},
      {stage5_39[1],stage5_38[3],stage5_37[6],stage5_36[6],stage5_35[8]}
   );
   gpc615_5 gpc9357 (
      {stage4_35[27], stage4_35[28], stage4_35[29], stage4_35[30], stage4_35[31]},
      {stage4_36[15]},
      {stage4_37[12], stage4_37[13], stage4_37[14], stage4_37[15], stage4_37[16], stage4_37[17]},
      {stage5_39[2],stage5_38[4],stage5_37[7],stage5_36[7],stage5_35[9]}
   );
   gpc606_5 gpc9358 (
      {stage4_36[16], stage4_36[17], stage4_36[18], stage4_36[19], stage4_36[20], stage4_36[21]},
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5]},
      {stage5_40[0],stage5_39[3],stage5_38[5],stage5_37[8],stage5_36[8]}
   );
   gpc606_5 gpc9359 (
      {stage4_36[22], stage4_36[23], stage4_36[24], stage4_36[25], stage4_36[26], stage4_36[27]},
      {stage4_38[6], stage4_38[7], stage4_38[8], stage4_38[9], stage4_38[10], stage4_38[11]},
      {stage5_40[1],stage5_39[4],stage5_38[6],stage5_37[9],stage5_36[9]}
   );
   gpc606_5 gpc9360 (
      {stage4_36[28], stage4_36[29], stage4_36[30], stage4_36[31], stage4_36[32], stage4_36[33]},
      {stage4_38[12], stage4_38[13], stage4_38[14], stage4_38[15], stage4_38[16], stage4_38[17]},
      {stage5_40[2],stage5_39[5],stage5_38[7],stage5_37[10],stage5_36[10]}
   );
   gpc117_4 gpc9361 (
      {stage4_39[0], stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5], stage4_39[6]},
      {stage4_40[0]},
      {stage4_41[0]},
      {stage5_42[0],stage5_41[0],stage5_40[3],stage5_39[6]}
   );
   gpc117_4 gpc9362 (
      {stage4_39[7], stage4_39[8], stage4_39[9], stage4_39[10], stage4_39[11], stage4_39[12], stage4_39[13]},
      {stage4_40[1]},
      {stage4_41[1]},
      {stage5_42[1],stage5_41[1],stage5_40[4],stage5_39[7]}
   );
   gpc615_5 gpc9363 (
      {stage4_39[14], stage4_39[15], stage4_39[16], stage4_39[17], stage4_39[18]},
      {stage4_40[2]},
      {stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5], stage4_41[6], stage4_41[7]},
      {stage5_43[0],stage5_42[2],stage5_41[2],stage5_40[5],stage5_39[8]}
   );
   gpc615_5 gpc9364 (
      {stage4_39[19], stage4_39[20], stage4_39[21], stage4_39[22], stage4_39[23]},
      {stage4_40[3]},
      {stage4_41[8], stage4_41[9], stage4_41[10], stage4_41[11], stage4_41[12], stage4_41[13]},
      {stage5_43[1],stage5_42[3],stage5_41[3],stage5_40[6],stage5_39[9]}
   );
   gpc606_5 gpc9365 (
      {stage4_40[4], stage4_40[5], stage4_40[6], stage4_40[7], stage4_40[8], stage4_40[9]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[2],stage5_42[4],stage5_41[4],stage5_40[7]}
   );
   gpc606_5 gpc9366 (
      {stage4_40[10], stage4_40[11], stage4_40[12], stage4_40[13], stage4_40[14], stage4_40[15]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[3],stage5_42[5],stage5_41[5],stage5_40[8]}
   );
   gpc606_5 gpc9367 (
      {stage4_40[16], stage4_40[17], stage4_40[18], stage4_40[19], stage4_40[20], stage4_40[21]},
      {stage4_42[12], stage4_42[13], stage4_42[14], stage4_42[15], stage4_42[16], stage4_42[17]},
      {stage5_44[2],stage5_43[4],stage5_42[6],stage5_41[6],stage5_40[9]}
   );
   gpc606_5 gpc9368 (
      {stage4_40[22], stage4_40[23], stage4_40[24], stage4_40[25], stage4_40[26], stage4_40[27]},
      {stage4_42[18], stage4_42[19], stage4_42[20], stage4_42[21], stage4_42[22], stage4_42[23]},
      {stage5_44[3],stage5_43[5],stage5_42[7],stage5_41[7],stage5_40[10]}
   );
   gpc606_5 gpc9369 (
      {stage4_41[14], stage4_41[15], stage4_41[16], stage4_41[17], stage4_41[18], stage4_41[19]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[4],stage5_43[6],stage5_42[8],stage5_41[8]}
   );
   gpc615_5 gpc9370 (
      {stage4_42[24], stage4_42[25], stage4_42[26], stage4_42[27], stage4_42[28]},
      {stage4_43[6]},
      {stage4_44[0], stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage5_46[0],stage5_45[1],stage5_44[5],stage5_43[7],stage5_42[9]}
   );
   gpc615_5 gpc9371 (
      {stage4_43[7], stage4_43[8], stage4_43[9], stage4_43[10], stage4_43[11]},
      {stage4_44[6]},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[1],stage5_45[2],stage5_44[6],stage5_43[8]}
   );
   gpc135_4 gpc9372 (
      {stage4_44[7], stage4_44[8], stage4_44[9], stage4_44[10], stage4_44[11]},
      {stage4_45[6], stage4_45[7], stage4_45[8]},
      {stage4_46[0]},
      {stage5_47[1],stage5_46[2],stage5_45[3],stage5_44[7]}
   );
   gpc135_4 gpc9373 (
      {stage4_44[12], stage4_44[13], stage4_44[14], stage4_44[15], stage4_44[16]},
      {stage4_45[9], stage4_45[10], stage4_45[11]},
      {stage4_46[1]},
      {stage5_47[2],stage5_46[3],stage5_45[4],stage5_44[8]}
   );
   gpc135_4 gpc9374 (
      {stage4_44[17], stage4_44[18], stage4_44[19], stage4_44[20], stage4_44[21]},
      {stage4_45[12], stage4_45[13], stage4_45[14]},
      {stage4_46[2]},
      {stage5_47[3],stage5_46[4],stage5_45[5],stage5_44[9]}
   );
   gpc606_5 gpc9375 (
      {stage4_45[15], stage4_45[16], stage4_45[17], stage4_45[18], stage4_45[19], stage4_45[20]},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4], stage4_47[5]},
      {stage5_49[0],stage5_48[0],stage5_47[4],stage5_46[5],stage5_45[6]}
   );
   gpc615_5 gpc9376 (
      {stage4_46[3], stage4_46[4], stage4_46[5], stage4_46[6], stage4_46[7]},
      {stage4_47[6]},
      {stage4_48[0], stage4_48[1], stage4_48[2], stage4_48[3], stage4_48[4], stage4_48[5]},
      {stage5_50[0],stage5_49[1],stage5_48[1],stage5_47[5],stage5_46[6]}
   );
   gpc615_5 gpc9377 (
      {stage4_46[8], stage4_46[9], stage4_46[10], stage4_46[11], stage4_46[12]},
      {stage4_47[7]},
      {stage4_48[6], stage4_48[7], stage4_48[8], stage4_48[9], stage4_48[10], stage4_48[11]},
      {stage5_50[1],stage5_49[2],stage5_48[2],stage5_47[6],stage5_46[7]}
   );
   gpc615_5 gpc9378 (
      {stage4_47[8], stage4_47[9], stage4_47[10], stage4_47[11], stage4_47[12]},
      {stage4_48[12]},
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4], stage4_49[5]},
      {stage5_51[0],stage5_50[2],stage5_49[3],stage5_48[3],stage5_47[7]}
   );
   gpc615_5 gpc9379 (
      {stage4_47[13], stage4_47[14], stage4_47[15], stage4_47[16], stage4_47[17]},
      {stage4_48[13]},
      {stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10], stage4_49[11]},
      {stage5_51[1],stage5_50[3],stage5_49[4],stage5_48[4],stage5_47[8]}
   );
   gpc7_3 gpc9380 (
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6]},
      {stage5_52[0],stage5_51[2],stage5_50[4]}
   );
   gpc615_5 gpc9381 (
      {stage4_50[7], stage4_50[8], stage4_50[9], stage4_50[10], stage4_50[11]},
      {stage4_51[0]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[0],stage5_52[1],stage5_51[3],stage5_50[5]}
   );
   gpc615_5 gpc9382 (
      {stage4_50[12], stage4_50[13], stage4_50[14], stage4_50[15], stage4_50[16]},
      {stage4_51[1]},
      {stage4_52[6], stage4_52[7], stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11]},
      {stage5_54[1],stage5_53[1],stage5_52[2],stage5_51[4],stage5_50[6]}
   );
   gpc615_5 gpc9383 (
      {stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5], stage4_51[6]},
      {stage4_52[12]},
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage5_55[0],stage5_54[2],stage5_53[2],stage5_52[3],stage5_51[5]}
   );
   gpc615_5 gpc9384 (
      {stage4_51[7], stage4_51[8], stage4_51[9], stage4_51[10], stage4_51[11]},
      {stage4_52[13]},
      {stage4_53[6], stage4_53[7], stage4_53[8], stage4_53[9], stage4_53[10], stage4_53[11]},
      {stage5_55[1],stage5_54[3],stage5_53[3],stage5_52[4],stage5_51[6]}
   );
   gpc615_5 gpc9385 (
      {stage4_51[12], stage4_51[13], stage4_51[14], stage4_51[15], stage4_51[16]},
      {stage4_52[14]},
      {stage4_53[12], stage4_53[13], stage4_53[14], stage4_53[15], stage4_53[16], stage4_53[17]},
      {stage5_55[2],stage5_54[4],stage5_53[4],stage5_52[5],stage5_51[7]}
   );
   gpc615_5 gpc9386 (
      {stage4_51[17], stage4_51[18], stage4_51[19], stage4_51[20], stage4_51[21]},
      {stage4_52[15]},
      {stage4_53[18], stage4_53[19], stage4_53[20], stage4_53[21], stage4_53[22], stage4_53[23]},
      {stage5_55[3],stage5_54[5],stage5_53[5],stage5_52[6],stage5_51[8]}
   );
   gpc615_5 gpc9387 (
      {stage4_51[22], stage4_51[23], stage4_51[24], stage4_51[25], stage4_51[26]},
      {stage4_52[16]},
      {stage4_53[24], stage4_53[25], stage4_53[26], stage4_53[27], stage4_53[28], stage4_53[29]},
      {stage5_55[4],stage5_54[6],stage5_53[6],stage5_52[7],stage5_51[9]}
   );
   gpc615_5 gpc9388 (
      {stage4_53[30], stage4_53[31], stage4_53[32], stage4_53[33], stage4_53[34]},
      {stage4_54[0]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[0],stage5_55[5],stage5_54[7],stage5_53[7]}
   );
   gpc615_5 gpc9389 (
      {stage4_53[35], stage4_53[36], stage4_53[37], stage4_53[38], stage4_53[39]},
      {stage4_54[1]},
      {stage4_55[6], stage4_55[7], stage4_55[8], stage4_55[9], stage4_55[10], stage4_55[11]},
      {stage5_57[1],stage5_56[1],stage5_55[6],stage5_54[8],stage5_53[8]}
   );
   gpc2135_5 gpc9390 (
      {stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5], stage4_54[6]},
      {stage4_55[12], stage4_55[13], stage4_55[14]},
      {stage4_56[0]},
      {stage4_57[0], stage4_57[1]},
      {stage5_58[0],stage5_57[2],stage5_56[2],stage5_55[7],stage5_54[9]}
   );
   gpc2135_5 gpc9391 (
      {stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10], stage4_54[11]},
      {stage4_55[15], stage4_55[16], stage4_55[17]},
      {stage4_56[1]},
      {stage4_57[2], stage4_57[3]},
      {stage5_58[1],stage5_57[3],stage5_56[3],stage5_55[8],stage5_54[10]}
   );
   gpc2135_5 gpc9392 (
      {stage4_54[12], stage4_54[13], stage4_54[14], stage4_54[15], stage4_54[16]},
      {stage4_55[18], stage4_55[19], stage4_55[20]},
      {stage4_56[2]},
      {stage4_57[4], stage4_57[5]},
      {stage5_58[2],stage5_57[4],stage5_56[4],stage5_55[9],stage5_54[11]}
   );
   gpc2135_5 gpc9393 (
      {stage4_54[17], stage4_54[18], stage4_54[19], stage4_54[20], stage4_54[21]},
      {stage4_55[21], stage4_55[22], stage4_55[23]},
      {stage4_56[3]},
      {stage4_57[6], stage4_57[7]},
      {stage5_58[3],stage5_57[5],stage5_56[5],stage5_55[10],stage5_54[12]}
   );
   gpc615_5 gpc9394 (
      {stage4_55[24], stage4_55[25], stage4_55[26], stage4_55[27], stage4_55[28]},
      {stage4_56[4]},
      {stage4_57[8], stage4_57[9], stage4_57[10], stage4_57[11], stage4_57[12], stage4_57[13]},
      {stage5_59[0],stage5_58[4],stage5_57[6],stage5_56[6],stage5_55[11]}
   );
   gpc606_5 gpc9395 (
      {stage4_56[5], stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10]},
      {stage4_58[0], stage4_58[1], stage4_58[2], stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage5_60[0],stage5_59[1],stage5_58[5],stage5_57[7],stage5_56[7]}
   );
   gpc623_5 gpc9396 (
      {stage4_56[11], stage4_56[12], stage4_56[13]},
      {stage4_57[14], stage4_57[15]},
      {stage4_58[6], stage4_58[7], stage4_58[8], stage4_58[9], stage4_58[10], stage4_58[11]},
      {stage5_60[1],stage5_59[2],stage5_58[6],stage5_57[8],stage5_56[8]}
   );
   gpc606_5 gpc9397 (
      {stage4_57[16], stage4_57[17], stage4_57[18], stage4_57[19], stage4_57[20], stage4_57[21]},
      {stage4_59[0], stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage5_61[0],stage5_60[2],stage5_59[3],stage5_58[7],stage5_57[9]}
   );
   gpc615_5 gpc9398 (
      {stage4_58[12], stage4_58[13], stage4_58[14], stage4_58[15], stage4_58[16]},
      {stage4_59[6]},
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage5_62[0],stage5_61[1],stage5_60[3],stage5_59[4],stage5_58[8]}
   );
   gpc615_5 gpc9399 (
      {stage4_59[7], stage4_59[8], stage4_59[9], stage4_59[10], stage4_59[11]},
      {stage4_60[6]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[1],stage5_61[2],stage5_60[4],stage5_59[5]}
   );
   gpc615_5 gpc9400 (
      {stage4_59[12], stage4_59[13], stage4_59[14], stage4_59[15], stage4_59[16]},
      {stage4_60[7]},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[2],stage5_61[3],stage5_60[5],stage5_59[6]}
   );
   gpc615_5 gpc9401 (
      {stage4_59[17], stage4_59[18], stage4_59[19], stage4_59[20], 1'b0},
      {stage4_60[8]},
      {stage4_61[12], stage4_61[13], stage4_61[14], stage4_61[15], stage4_61[16], stage4_61[17]},
      {stage5_63[2],stage5_62[3],stage5_61[4],stage5_60[6],stage5_59[7]}
   );
   gpc606_5 gpc9402 (
      {stage4_60[9], stage4_60[10], stage4_60[11], stage4_60[12], stage4_60[13], stage4_60[14]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[3],stage5_62[4],stage5_61[5],stage5_60[7]}
   );
   gpc615_5 gpc9403 (
      {stage4_61[18], stage4_61[19], stage4_61[20], stage4_61[21], stage4_61[22]},
      {stage4_62[6]},
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5]},
      {stage5_65[0],stage5_64[1],stage5_63[4],stage5_62[5],stage5_61[6]}
   );
   gpc615_5 gpc9404 (
      {stage4_62[7], stage4_62[8], stage4_62[9], stage4_62[10], stage4_62[11]},
      {stage4_63[6]},
      {stage4_64[0], stage4_64[1], stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5]},
      {stage5_66[0],stage5_65[1],stage5_64[2],stage5_63[5],stage5_62[6]}
   );
   gpc615_5 gpc9405 (
      {stage4_63[7], stage4_63[8], stage4_63[9], stage4_63[10], stage4_63[11]},
      {stage4_64[6]},
      {stage4_65[0], stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5]},
      {stage5_67[0],stage5_66[1],stage5_65[2],stage5_64[3],stage5_63[6]}
   );
   gpc2135_5 gpc9406 (
      {stage4_64[7], stage4_64[8], stage4_64[9], stage4_64[10], stage4_64[11]},
      {stage4_65[6], stage4_65[7], stage4_65[8]},
      {stage4_66[0]},
      {stage4_67[0], stage4_67[1]},
      {stage5_68[0],stage5_67[1],stage5_66[2],stage5_65[3],stage5_64[4]}
   );
   gpc2135_5 gpc9407 (
      {stage4_64[12], stage4_64[13], stage4_64[14], stage4_64[15], stage4_64[16]},
      {stage4_65[9], stage4_65[10], stage4_65[11]},
      {stage4_66[1]},
      {stage4_67[2], stage4_67[3]},
      {stage5_68[1],stage5_67[2],stage5_66[3],stage5_65[4],stage5_64[5]}
   );
   gpc1163_5 gpc9408 (
      {stage4_64[17], stage4_64[18], stage4_64[19]},
      {stage4_65[12], stage4_65[13], stage4_65[14], stage4_65[15], stage4_65[16], stage4_65[17]},
      {stage4_66[2]},
      {stage4_67[4]},
      {stage5_68[2],stage5_67[3],stage5_66[4],stage5_65[5],stage5_64[6]}
   );
   gpc1163_5 gpc9409 (
      {stage4_64[20], stage4_64[21], stage4_64[22]},
      {stage4_65[18], stage4_65[19], stage4_65[20], stage4_65[21], stage4_65[22], stage4_65[23]},
      {stage4_66[3]},
      {stage4_67[5]},
      {stage5_68[3],stage5_67[4],stage5_66[5],stage5_65[6],stage5_64[7]}
   );
   gpc1325_5 gpc9410 (
      {stage4_64[23], stage4_64[24], stage4_64[25], stage4_64[26], stage4_64[27]},
      {stage4_65[24], stage4_65[25]},
      {stage4_66[4], stage4_66[5], stage4_66[6]},
      {stage4_67[6]},
      {stage5_68[4],stage5_67[5],stage5_66[6],stage5_65[7],stage5_64[8]}
   );
   gpc606_5 gpc9411 (
      {stage4_66[7], stage4_66[8], stage4_66[9], stage4_66[10], 1'b0, 1'b0},
      {stage4_68[0], stage4_68[1], stage4_68[2], stage4_68[3], stage4_68[4], stage4_68[5]},
      {stage5_70[0],stage5_69[0],stage5_68[5],stage5_67[6],stage5_66[7]}
   );
   gpc1_1 gpc9412 (
      {stage4_0[5]},
      {stage5_0[1]}
   );
   gpc1_1 gpc9413 (
      {stage4_0[6]},
      {stage5_0[2]}
   );
   gpc1_1 gpc9414 (
      {stage4_0[7]},
      {stage5_0[3]}
   );
   gpc1_1 gpc9415 (
      {stage4_0[8]},
      {stage5_0[4]}
   );
   gpc1_1 gpc9416 (
      {stage4_2[9]},
      {stage5_2[3]}
   );
   gpc1_1 gpc9417 (
      {stage4_2[10]},
      {stage5_2[4]}
   );
   gpc1_1 gpc9418 (
      {stage4_3[12]},
      {stage5_3[3]}
   );
   gpc1_1 gpc9419 (
      {stage4_3[13]},
      {stage5_3[4]}
   );
   gpc1_1 gpc9420 (
      {stage4_3[14]},
      {stage5_3[5]}
   );
   gpc1_1 gpc9421 (
      {stage4_3[15]},
      {stage5_3[6]}
   );
   gpc1_1 gpc9422 (
      {stage4_3[16]},
      {stage5_3[7]}
   );
   gpc1_1 gpc9423 (
      {stage4_4[28]},
      {stage5_4[8]}
   );
   gpc1_1 gpc9424 (
      {stage4_4[29]},
      {stage5_4[9]}
   );
   gpc1_1 gpc9425 (
      {stage4_4[30]},
      {stage5_4[10]}
   );
   gpc1_1 gpc9426 (
      {stage4_5[31]},
      {stage5_5[11]}
   );
   gpc1_1 gpc9427 (
      {stage4_5[32]},
      {stage5_5[12]}
   );
   gpc1_1 gpc9428 (
      {stage4_5[33]},
      {stage5_5[13]}
   );
   gpc1_1 gpc9429 (
      {stage4_5[34]},
      {stage5_5[14]}
   );
   gpc1_1 gpc9430 (
      {stage4_5[35]},
      {stage5_5[15]}
   );
   gpc1_1 gpc9431 (
      {stage4_8[24]},
      {stage5_8[15]}
   );
   gpc1_1 gpc9432 (
      {stage4_8[25]},
      {stage5_8[16]}
   );
   gpc1_1 gpc9433 (
      {stage4_8[26]},
      {stage5_8[17]}
   );
   gpc1_1 gpc9434 (
      {stage4_8[27]},
      {stage5_8[18]}
   );
   gpc1_1 gpc9435 (
      {stage4_10[31]},
      {stage5_10[10]}
   );
   gpc1_1 gpc9436 (
      {stage4_10[32]},
      {stage5_10[11]}
   );
   gpc1_1 gpc9437 (
      {stage4_10[33]},
      {stage5_10[12]}
   );
   gpc1_1 gpc9438 (
      {stage4_10[34]},
      {stage5_10[13]}
   );
   gpc1_1 gpc9439 (
      {stage4_10[35]},
      {stage5_10[14]}
   );
   gpc1_1 gpc9440 (
      {stage4_10[36]},
      {stage5_10[15]}
   );
   gpc1_1 gpc9441 (
      {stage4_10[37]},
      {stage5_10[16]}
   );
   gpc1_1 gpc9442 (
      {stage4_10[38]},
      {stage5_10[17]}
   );
   gpc1_1 gpc9443 (
      {stage4_10[39]},
      {stage5_10[18]}
   );
   gpc1_1 gpc9444 (
      {stage4_10[40]},
      {stage5_10[19]}
   );
   gpc1_1 gpc9445 (
      {stage4_10[41]},
      {stage5_10[20]}
   );
   gpc1_1 gpc9446 (
      {stage4_11[27]},
      {stage5_11[12]}
   );
   gpc1_1 gpc9447 (
      {stage4_11[28]},
      {stage5_11[13]}
   );
   gpc1_1 gpc9448 (
      {stage4_13[26]},
      {stage5_13[9]}
   );
   gpc1_1 gpc9449 (
      {stage4_13[27]},
      {stage5_13[10]}
   );
   gpc1_1 gpc9450 (
      {stage4_13[28]},
      {stage5_13[11]}
   );
   gpc1_1 gpc9451 (
      {stage4_13[29]},
      {stage5_13[12]}
   );
   gpc1_1 gpc9452 (
      {stage4_13[30]},
      {stage5_13[13]}
   );
   gpc1_1 gpc9453 (
      {stage4_13[31]},
      {stage5_13[14]}
   );
   gpc1_1 gpc9454 (
      {stage4_14[26]},
      {stage5_14[12]}
   );
   gpc1_1 gpc9455 (
      {stage4_14[27]},
      {stage5_14[13]}
   );
   gpc1_1 gpc9456 (
      {stage4_14[28]},
      {stage5_14[14]}
   );
   gpc1_1 gpc9457 (
      {stage4_14[29]},
      {stage5_14[15]}
   );
   gpc1_1 gpc9458 (
      {stage4_18[20]},
      {stage5_18[11]}
   );
   gpc1_1 gpc9459 (
      {stage4_19[24]},
      {stage5_19[11]}
   );
   gpc1_1 gpc9460 (
      {stage4_19[25]},
      {stage5_19[12]}
   );
   gpc1_1 gpc9461 (
      {stage4_19[26]},
      {stage5_19[13]}
   );
   gpc1_1 gpc9462 (
      {stage4_19[27]},
      {stage5_19[14]}
   );
   gpc1_1 gpc9463 (
      {stage4_19[28]},
      {stage5_19[15]}
   );
   gpc1_1 gpc9464 (
      {stage4_20[28]},
      {stage5_20[8]}
   );
   gpc1_1 gpc9465 (
      {stage4_20[29]},
      {stage5_20[9]}
   );
   gpc1_1 gpc9466 (
      {stage4_20[30]},
      {stage5_20[10]}
   );
   gpc1_1 gpc9467 (
      {stage4_20[31]},
      {stage5_20[11]}
   );
   gpc1_1 gpc9468 (
      {stage4_20[32]},
      {stage5_20[12]}
   );
   gpc1_1 gpc9469 (
      {stage4_20[33]},
      {stage5_20[13]}
   );
   gpc1_1 gpc9470 (
      {stage4_21[36]},
      {stage5_21[10]}
   );
   gpc1_1 gpc9471 (
      {stage4_24[19]},
      {stage5_24[6]}
   );
   gpc1_1 gpc9472 (
      {stage4_24[20]},
      {stage5_24[7]}
   );
   gpc1_1 gpc9473 (
      {stage4_24[21]},
      {stage5_24[8]}
   );
   gpc1_1 gpc9474 (
      {stage4_26[14]},
      {stage5_26[10]}
   );
   gpc1_1 gpc9475 (
      {stage4_26[15]},
      {stage5_26[11]}
   );
   gpc1_1 gpc9476 (
      {stage4_26[16]},
      {stage5_26[12]}
   );
   gpc1_1 gpc9477 (
      {stage4_26[17]},
      {stage5_26[13]}
   );
   gpc1_1 gpc9478 (
      {stage4_26[18]},
      {stage5_26[14]}
   );
   gpc1_1 gpc9479 (
      {stage4_28[18]},
      {stage5_28[9]}
   );
   gpc1_1 gpc9480 (
      {stage4_29[18]},
      {stage5_29[11]}
   );
   gpc1_1 gpc9481 (
      {stage4_29[19]},
      {stage5_29[12]}
   );
   gpc1_1 gpc9482 (
      {stage4_29[20]},
      {stage5_29[13]}
   );
   gpc1_1 gpc9483 (
      {stage4_29[21]},
      {stage5_29[14]}
   );
   gpc1_1 gpc9484 (
      {stage4_32[20]},
      {stage5_32[10]}
   );
   gpc1_1 gpc9485 (
      {stage4_32[21]},
      {stage5_32[11]}
   );
   gpc1_1 gpc9486 (
      {stage4_32[22]},
      {stage5_32[12]}
   );
   gpc1_1 gpc9487 (
      {stage4_32[23]},
      {stage5_32[13]}
   );
   gpc1_1 gpc9488 (
      {stage4_32[24]},
      {stage5_32[14]}
   );
   gpc1_1 gpc9489 (
      {stage4_32[25]},
      {stage5_32[15]}
   );
   gpc1_1 gpc9490 (
      {stage4_32[26]},
      {stage5_32[16]}
   );
   gpc1_1 gpc9491 (
      {stage4_32[27]},
      {stage5_32[17]}
   );
   gpc1_1 gpc9492 (
      {stage4_32[28]},
      {stage5_32[18]}
   );
   gpc1_1 gpc9493 (
      {stage4_32[29]},
      {stage5_32[19]}
   );
   gpc1_1 gpc9494 (
      {stage4_33[24]},
      {stage5_33[7]}
   );
   gpc1_1 gpc9495 (
      {stage4_33[25]},
      {stage5_33[8]}
   );
   gpc1_1 gpc9496 (
      {stage4_33[26]},
      {stage5_33[9]}
   );
   gpc1_1 gpc9497 (
      {stage4_33[27]},
      {stage5_33[10]}
   );
   gpc1_1 gpc9498 (
      {stage4_33[28]},
      {stage5_33[11]}
   );
   gpc1_1 gpc9499 (
      {stage4_34[15]},
      {stage5_34[10]}
   );
   gpc1_1 gpc9500 (
      {stage4_34[16]},
      {stage5_34[11]}
   );
   gpc1_1 gpc9501 (
      {stage4_34[17]},
      {stage5_34[12]}
   );
   gpc1_1 gpc9502 (
      {stage4_34[18]},
      {stage5_34[13]}
   );
   gpc1_1 gpc9503 (
      {stage4_35[32]},
      {stage5_35[10]}
   );
   gpc1_1 gpc9504 (
      {stage4_35[33]},
      {stage5_35[11]}
   );
   gpc1_1 gpc9505 (
      {stage4_35[34]},
      {stage5_35[12]}
   );
   gpc1_1 gpc9506 (
      {stage4_35[35]},
      {stage5_35[13]}
   );
   gpc1_1 gpc9507 (
      {stage4_36[34]},
      {stage5_36[11]}
   );
   gpc1_1 gpc9508 (
      {stage4_36[35]},
      {stage5_36[12]}
   );
   gpc1_1 gpc9509 (
      {stage4_38[18]},
      {stage5_38[8]}
   );
   gpc1_1 gpc9510 (
      {stage4_38[19]},
      {stage5_38[9]}
   );
   gpc1_1 gpc9511 (
      {stage4_42[29]},
      {stage5_42[10]}
   );
   gpc1_1 gpc9512 (
      {stage4_42[30]},
      {stage5_42[11]}
   );
   gpc1_1 gpc9513 (
      {stage4_42[31]},
      {stage5_42[12]}
   );
   gpc1_1 gpc9514 (
      {stage4_42[32]},
      {stage5_42[13]}
   );
   gpc1_1 gpc9515 (
      {stage4_42[33]},
      {stage5_42[14]}
   );
   gpc1_1 gpc9516 (
      {stage4_42[34]},
      {stage5_42[15]}
   );
   gpc1_1 gpc9517 (
      {stage4_42[35]},
      {stage5_42[16]}
   );
   gpc1_1 gpc9518 (
      {stage4_42[36]},
      {stage5_42[17]}
   );
   gpc1_1 gpc9519 (
      {stage4_42[37]},
      {stage5_42[18]}
   );
   gpc1_1 gpc9520 (
      {stage4_43[12]},
      {stage5_43[9]}
   );
   gpc1_1 gpc9521 (
      {stage4_43[13]},
      {stage5_43[10]}
   );
   gpc1_1 gpc9522 (
      {stage4_44[22]},
      {stage5_44[10]}
   );
   gpc1_1 gpc9523 (
      {stage4_44[23]},
      {stage5_44[11]}
   );
   gpc1_1 gpc9524 (
      {stage4_44[24]},
      {stage5_44[12]}
   );
   gpc1_1 gpc9525 (
      {stage4_45[21]},
      {stage5_45[7]}
   );
   gpc1_1 gpc9526 (
      {stage4_45[22]},
      {stage5_45[8]}
   );
   gpc1_1 gpc9527 (
      {stage4_45[23]},
      {stage5_45[9]}
   );
   gpc1_1 gpc9528 (
      {stage4_45[24]},
      {stage5_45[10]}
   );
   gpc1_1 gpc9529 (
      {stage4_45[25]},
      {stage5_45[11]}
   );
   gpc1_1 gpc9530 (
      {stage4_45[26]},
      {stage5_45[12]}
   );
   gpc1_1 gpc9531 (
      {stage4_45[27]},
      {stage5_45[13]}
   );
   gpc1_1 gpc9532 (
      {stage4_45[28]},
      {stage5_45[14]}
   );
   gpc1_1 gpc9533 (
      {stage4_46[13]},
      {stage5_46[8]}
   );
   gpc1_1 gpc9534 (
      {stage4_46[14]},
      {stage5_46[9]}
   );
   gpc1_1 gpc9535 (
      {stage4_46[15]},
      {stage5_46[10]}
   );
   gpc1_1 gpc9536 (
      {stage4_46[16]},
      {stage5_46[11]}
   );
   gpc1_1 gpc9537 (
      {stage4_47[18]},
      {stage5_47[9]}
   );
   gpc1_1 gpc9538 (
      {stage4_47[19]},
      {stage5_47[10]}
   );
   gpc1_1 gpc9539 (
      {stage4_47[20]},
      {stage5_47[11]}
   );
   gpc1_1 gpc9540 (
      {stage4_48[14]},
      {stage5_48[5]}
   );
   gpc1_1 gpc9541 (
      {stage4_48[15]},
      {stage5_48[6]}
   );
   gpc1_1 gpc9542 (
      {stage4_48[16]},
      {stage5_48[7]}
   );
   gpc1_1 gpc9543 (
      {stage4_48[17]},
      {stage5_48[8]}
   );
   gpc1_1 gpc9544 (
      {stage4_48[18]},
      {stage5_48[9]}
   );
   gpc1_1 gpc9545 (
      {stage4_48[19]},
      {stage5_48[10]}
   );
   gpc1_1 gpc9546 (
      {stage4_48[20]},
      {stage5_48[11]}
   );
   gpc1_1 gpc9547 (
      {stage4_48[21]},
      {stage5_48[12]}
   );
   gpc1_1 gpc9548 (
      {stage4_48[22]},
      {stage5_48[13]}
   );
   gpc1_1 gpc9549 (
      {stage4_49[12]},
      {stage5_49[5]}
   );
   gpc1_1 gpc9550 (
      {stage4_50[17]},
      {stage5_50[7]}
   );
   gpc1_1 gpc9551 (
      {stage4_50[18]},
      {stage5_50[8]}
   );
   gpc1_1 gpc9552 (
      {stage4_50[19]},
      {stage5_50[9]}
   );
   gpc1_1 gpc9553 (
      {stage4_50[20]},
      {stage5_50[10]}
   );
   gpc1_1 gpc9554 (
      {stage4_50[21]},
      {stage5_50[11]}
   );
   gpc1_1 gpc9555 (
      {stage4_51[27]},
      {stage5_51[10]}
   );
   gpc1_1 gpc9556 (
      {stage4_51[28]},
      {stage5_51[11]}
   );
   gpc1_1 gpc9557 (
      {stage4_51[29]},
      {stage5_51[12]}
   );
   gpc1_1 gpc9558 (
      {stage4_51[30]},
      {stage5_51[13]}
   );
   gpc1_1 gpc9559 (
      {stage4_51[31]},
      {stage5_51[14]}
   );
   gpc1_1 gpc9560 (
      {stage4_51[32]},
      {stage5_51[15]}
   );
   gpc1_1 gpc9561 (
      {stage4_51[33]},
      {stage5_51[16]}
   );
   gpc1_1 gpc9562 (
      {stage4_51[34]},
      {stage5_51[17]}
   );
   gpc1_1 gpc9563 (
      {stage4_51[35]},
      {stage5_51[18]}
   );
   gpc1_1 gpc9564 (
      {stage4_52[17]},
      {stage5_52[8]}
   );
   gpc1_1 gpc9565 (
      {stage4_52[18]},
      {stage5_52[9]}
   );
   gpc1_1 gpc9566 (
      {stage4_53[40]},
      {stage5_53[9]}
   );
   gpc1_1 gpc9567 (
      {stage4_53[41]},
      {stage5_53[10]}
   );
   gpc1_1 gpc9568 (
      {stage4_53[42]},
      {stage5_53[11]}
   );
   gpc1_1 gpc9569 (
      {stage4_53[43]},
      {stage5_53[12]}
   );
   gpc1_1 gpc9570 (
      {stage4_54[22]},
      {stage5_54[13]}
   );
   gpc1_1 gpc9571 (
      {stage4_54[23]},
      {stage5_54[14]}
   );
   gpc1_1 gpc9572 (
      {stage4_54[24]},
      {stage5_54[15]}
   );
   gpc1_1 gpc9573 (
      {stage4_54[25]},
      {stage5_54[16]}
   );
   gpc1_1 gpc9574 (
      {stage4_55[29]},
      {stage5_55[12]}
   );
   gpc1_1 gpc9575 (
      {stage4_55[30]},
      {stage5_55[13]}
   );
   gpc1_1 gpc9576 (
      {stage4_55[31]},
      {stage5_55[14]}
   );
   gpc1_1 gpc9577 (
      {stage4_55[32]},
      {stage5_55[15]}
   );
   gpc1_1 gpc9578 (
      {stage4_55[33]},
      {stage5_55[16]}
   );
   gpc1_1 gpc9579 (
      {stage4_55[34]},
      {stage5_55[17]}
   );
   gpc1_1 gpc9580 (
      {stage4_55[35]},
      {stage5_55[18]}
   );
   gpc1_1 gpc9581 (
      {stage4_55[36]},
      {stage5_55[19]}
   );
   gpc1_1 gpc9582 (
      {stage4_55[37]},
      {stage5_55[20]}
   );
   gpc1_1 gpc9583 (
      {stage4_55[38]},
      {stage5_55[21]}
   );
   gpc1_1 gpc9584 (
      {stage4_57[22]},
      {stage5_57[10]}
   );
   gpc1_1 gpc9585 (
      {stage4_57[23]},
      {stage5_57[11]}
   );
   gpc1_1 gpc9586 (
      {stage4_57[24]},
      {stage5_57[12]}
   );
   gpc1_1 gpc9587 (
      {stage4_57[25]},
      {stage5_57[13]}
   );
   gpc1_1 gpc9588 (
      {stage4_58[17]},
      {stage5_58[9]}
   );
   gpc1_1 gpc9589 (
      {stage4_58[18]},
      {stage5_58[10]}
   );
   gpc1_1 gpc9590 (
      {stage4_58[19]},
      {stage5_58[11]}
   );
   gpc1_1 gpc9591 (
      {stage4_58[20]},
      {stage5_58[12]}
   );
   gpc1_1 gpc9592 (
      {stage4_58[21]},
      {stage5_58[13]}
   );
   gpc1_1 gpc9593 (
      {stage4_58[22]},
      {stage5_58[14]}
   );
   gpc1_1 gpc9594 (
      {stage4_58[23]},
      {stage5_58[15]}
   );
   gpc1_1 gpc9595 (
      {stage4_60[15]},
      {stage5_60[8]}
   );
   gpc1_1 gpc9596 (
      {stage4_60[16]},
      {stage5_60[9]}
   );
   gpc1_1 gpc9597 (
      {stage4_60[17]},
      {stage5_60[10]}
   );
   gpc1_1 gpc9598 (
      {stage4_60[18]},
      {stage5_60[11]}
   );
   gpc1_1 gpc9599 (
      {stage4_60[19]},
      {stage5_60[12]}
   );
   gpc1_1 gpc9600 (
      {stage4_60[20]},
      {stage5_60[13]}
   );
   gpc1_1 gpc9601 (
      {stage4_60[21]},
      {stage5_60[14]}
   );
   gpc1_1 gpc9602 (
      {stage4_61[23]},
      {stage5_61[7]}
   );
   gpc1_1 gpc9603 (
      {stage4_61[24]},
      {stage5_61[8]}
   );
   gpc1_1 gpc9604 (
      {stage4_61[25]},
      {stage5_61[9]}
   );
   gpc1_1 gpc9605 (
      {stage4_61[26]},
      {stage5_61[10]}
   );
   gpc1_1 gpc9606 (
      {stage4_61[27]},
      {stage5_61[11]}
   );
   gpc1_1 gpc9607 (
      {stage4_61[28]},
      {stage5_61[12]}
   );
   gpc1_1 gpc9608 (
      {stage4_61[29]},
      {stage5_61[13]}
   );
   gpc1_1 gpc9609 (
      {stage4_61[30]},
      {stage5_61[14]}
   );
   gpc1_1 gpc9610 (
      {stage4_61[31]},
      {stage5_61[15]}
   );
   gpc1_1 gpc9611 (
      {stage4_62[12]},
      {stage5_62[7]}
   );
   gpc1_1 gpc9612 (
      {stage4_62[13]},
      {stage5_62[8]}
   );
   gpc1_1 gpc9613 (
      {stage4_62[14]},
      {stage5_62[9]}
   );
   gpc1_1 gpc9614 (
      {stage4_62[15]},
      {stage5_62[10]}
   );
   gpc1_1 gpc9615 (
      {stage4_62[16]},
      {stage5_62[11]}
   );
   gpc1_1 gpc9616 (
      {stage4_63[12]},
      {stage5_63[7]}
   );
   gpc1_1 gpc9617 (
      {stage4_63[13]},
      {stage5_63[8]}
   );
   gpc1_1 gpc9618 (
      {stage4_64[28]},
      {stage5_64[9]}
   );
   gpc1_1 gpc9619 (
      {stage4_64[29]},
      {stage5_64[10]}
   );
   gpc1_1 gpc9620 (
      {stage4_64[30]},
      {stage5_64[11]}
   );
   gpc1_1 gpc9621 (
      {stage4_64[31]},
      {stage5_64[12]}
   );
   gpc1_1 gpc9622 (
      {stage4_64[32]},
      {stage5_64[13]}
   );
   gpc1_1 gpc9623 (
      {stage4_64[33]},
      {stage5_64[14]}
   );
   gpc1_1 gpc9624 (
      {stage4_65[26]},
      {stage5_65[8]}
   );
   gpc1_1 gpc9625 (
      {stage4_65[27]},
      {stage5_65[9]}
   );
   gpc1_1 gpc9626 (
      {stage4_65[28]},
      {stage5_65[10]}
   );
   gpc1_1 gpc9627 (
      {stage4_65[29]},
      {stage5_65[11]}
   );
   gpc1_1 gpc9628 (
      {stage4_65[30]},
      {stage5_65[12]}
   );
   gpc1_1 gpc9629 (
      {stage4_65[31]},
      {stage5_65[13]}
   );
   gpc1_1 gpc9630 (
      {stage4_65[32]},
      {stage5_65[14]}
   );
   gpc1_1 gpc9631 (
      {stage4_65[33]},
      {stage5_65[15]}
   );
   gpc1_1 gpc9632 (
      {stage4_65[34]},
      {stage5_65[16]}
   );
   gpc1_1 gpc9633 (
      {stage4_65[35]},
      {stage5_65[17]}
   );
   gpc1_1 gpc9634 (
      {stage4_67[7]},
      {stage5_67[7]}
   );
   gpc1_1 gpc9635 (
      {stage4_67[8]},
      {stage5_67[8]}
   );
   gpc1_1 gpc9636 (
      {stage4_67[9]},
      {stage5_67[9]}
   );
   gpc1_1 gpc9637 (
      {stage4_67[10]},
      {stage5_67[10]}
   );
   gpc1_1 gpc9638 (
      {stage4_68[6]},
      {stage5_68[6]}
   );
   gpc1_1 gpc9639 (
      {stage4_68[7]},
      {stage5_68[7]}
   );
   gpc1_1 gpc9640 (
      {stage4_68[8]},
      {stage5_68[8]}
   );
   gpc1_1 gpc9641 (
      {stage4_68[9]},
      {stage5_68[9]}
   );
   gpc1_1 gpc9642 (
      {stage4_68[10]},
      {stage5_68[10]}
   );
   gpc1_1 gpc9643 (
      {stage4_68[11]},
      {stage5_68[11]}
   );
   gpc1_1 gpc9644 (
      {stage4_68[12]},
      {stage5_68[12]}
   );
   gpc1_1 gpc9645 (
      {stage4_68[13]},
      {stage5_68[13]}
   );
   gpc1_1 gpc9646 (
      {stage4_69[0]},
      {stage5_69[1]}
   );
   gpc1_1 gpc9647 (
      {stage4_69[1]},
      {stage5_69[2]}
   );
   gpc615_5 gpc9648 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc615_5 gpc9649 (
      {stage5_3[5], stage5_3[6], stage5_3[7], 1'b0, 1'b0},
      {stage5_4[1]},
      {stage5_5[6], stage5_5[7], stage5_5[8], stage5_5[9], stage5_5[10], stage5_5[11]},
      {stage6_7[1],stage6_6[1],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc606_5 gpc9650 (
      {stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage6_8[0],stage6_7[2],stage6_6[2],stage6_5[2],stage6_4[2]}
   );
   gpc606_5 gpc9651 (
      {stage5_5[12], stage5_5[13], stage5_5[14], stage5_5[15], 1'b0, 1'b0},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[1],stage6_7[3],stage6_6[3],stage6_5[3]}
   );
   gpc615_5 gpc9652 (
      {stage5_7[6], stage5_7[7], stage5_7[8], stage5_7[9], stage5_7[10]},
      {stage5_8[0]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[2],stage6_7[4]}
   );
   gpc606_5 gpc9653 (
      {stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5], stage5_8[6]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[1],stage6_10[1],stage6_9[2],stage6_8[3]}
   );
   gpc606_5 gpc9654 (
      {stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11], stage5_8[12]},
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10], stage5_10[11]},
      {stage6_12[1],stage6_11[2],stage6_10[2],stage6_9[3],stage6_8[4]}
   );
   gpc606_5 gpc9655 (
      {stage5_8[13], stage5_8[14], stage5_8[15], stage5_8[16], stage5_8[17], stage5_8[18]},
      {stage5_10[12], stage5_10[13], stage5_10[14], stage5_10[15], stage5_10[16], stage5_10[17]},
      {stage6_12[2],stage6_11[3],stage6_10[3],stage6_9[4],stage6_8[5]}
   );
   gpc615_5 gpc9656 (
      {stage5_10[18], stage5_10[19], stage5_10[20], 1'b0, 1'b0},
      {stage5_11[0]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage6_14[0],stage6_13[0],stage6_12[3],stage6_11[4],stage6_10[4]}
   );
   gpc1406_5 gpc9657 (
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[1],stage6_13[1],stage6_12[4],stage6_11[5]}
   );
   gpc7_3 gpc9658 (
      {stage5_11[7], stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11], stage5_11[12], stage5_11[13]},
      {stage6_13[2],stage6_12[5],stage6_11[6]}
   );
   gpc606_5 gpc9659 (
      {stage5_12[6], stage5_12[7], stage5_12[8], stage5_12[9], stage5_12[10], 1'b0},
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5], stage5_14[6]},
      {stage6_16[0],stage6_15[1],stage6_14[2],stage6_13[3],stage6_12[6]}
   );
   gpc606_5 gpc9660 (
      {stage5_13[4], stage5_13[5], stage5_13[6], stage5_13[7], stage5_13[8], stage5_13[9]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[1],stage6_15[2],stage6_14[3],stage6_13[4]}
   );
   gpc1343_5 gpc9661 (
      {stage5_14[7], stage5_14[8], stage5_14[9]},
      {stage5_15[6], stage5_15[7], stage5_15[8], stage5_15[9]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[1],stage6_16[2],stage6_15[3],stage6_14[4]}
   );
   gpc615_5 gpc9662 (
      {stage5_14[10], stage5_14[11], stage5_14[12], stage5_14[13], stage5_14[14]},
      {stage5_15[10]},
      {stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7], 1'b0},
      {stage6_18[1],stage6_17[2],stage6_16[3],stage6_15[4],stage6_14[5]}
   );
   gpc615_5 gpc9663 (
      {stage5_14[15], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage5_15[11]},
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage6_18[2],stage6_17[3],stage6_16[4],stage6_15[5],stage6_14[6]}
   );
   gpc606_5 gpc9664 (
      {stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[3],stage6_17[4]}
   );
   gpc117_4 gpc9665 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage5_19[6]},
      {stage5_20[0]},
      {stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[4]}
   );
   gpc615_5 gpc9666 (
      {stage5_18[7], stage5_18[8], stage5_18[9], stage5_18[10], stage5_18[11]},
      {stage5_19[7]},
      {stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6]},
      {stage6_22[0],stage6_21[2],stage6_20[2],stage6_19[2],stage6_18[5]}
   );
   gpc615_5 gpc9667 (
      {stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12]},
      {stage5_20[7]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage6_23[0],stage6_22[1],stage6_21[3],stage6_20[3],stage6_19[3]}
   );
   gpc615_5 gpc9668 (
      {stage5_19[13], stage5_19[14], stage5_19[15], 1'b0, 1'b0},
      {stage5_20[8]},
      {stage5_21[6], stage5_21[7], stage5_21[8], stage5_21[9], stage5_21[10], 1'b0},
      {stage6_23[1],stage6_22[2],stage6_21[4],stage6_20[4],stage6_19[4]}
   );
   gpc606_5 gpc9669 (
      {stage5_20[9], stage5_20[10], stage5_20[11], stage5_20[12], stage5_20[13], 1'b0},
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage6_24[0],stage6_23[2],stage6_22[3],stage6_21[5],stage6_20[5]}
   );
   gpc15_3 gpc9670 (
      {stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9], stage5_22[10]},
      {stage5_23[0]},
      {stage6_24[1],stage6_23[3],stage6_22[4]}
   );
   gpc15_3 gpc9671 (
      {stage5_22[11], stage5_22[12], stage5_22[13], 1'b0, 1'b0},
      {stage5_23[1]},
      {stage6_24[2],stage6_23[4],stage6_22[5]}
   );
   gpc615_5 gpc9672 (
      {stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5], stage5_23[6]},
      {stage5_24[0]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3], stage5_25[4], stage5_25[5]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[3],stage6_23[5]}
   );
   gpc615_5 gpc9673 (
      {stage5_23[7], stage5_23[8], stage5_23[9], 1'b0, 1'b0},
      {stage5_24[1]},
      {stage5_25[6], stage5_25[7], stage5_25[8], stage5_25[9], 1'b0, 1'b0},
      {stage6_27[1],stage6_26[1],stage6_25[1],stage6_24[4],stage6_23[6]}
   );
   gpc606_5 gpc9674 (
      {stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6], stage5_24[7]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5]},
      {stage6_28[0],stage6_27[2],stage6_26[2],stage6_25[2],stage6_24[5]}
   );
   gpc615_5 gpc9675 (
      {stage5_26[6], stage5_26[7], stage5_26[8], stage5_26[9], stage5_26[10]},
      {stage5_27[0]},
      {stage5_28[0], stage5_28[1], stage5_28[2], stage5_28[3], stage5_28[4], stage5_28[5]},
      {stage6_30[0],stage6_29[0],stage6_28[1],stage6_27[3],stage6_26[3]}
   );
   gpc615_5 gpc9676 (
      {stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4], stage5_27[5]},
      {stage5_28[6]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[1],stage6_29[1],stage6_28[2],stage6_27[4]}
   );
   gpc606_5 gpc9677 (
      {stage5_29[6], stage5_29[7], stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[2],stage6_29[2]}
   );
   gpc615_5 gpc9678 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4]},
      {stage5_31[6]},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage6_34[0],stage6_33[1],stage6_32[1],stage6_31[2],stage6_30[3]}
   );
   gpc615_5 gpc9679 (
      {stage5_30[5], stage5_30[6], stage5_30[7], stage5_30[8], 1'b0},
      {stage5_31[7]},
      {stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9], stage5_32[10], stage5_32[11]},
      {stage6_34[1],stage6_33[2],stage6_32[2],stage6_31[3],stage6_30[4]}
   );
   gpc606_5 gpc9680 (
      {stage5_32[12], stage5_32[13], stage5_32[14], stage5_32[15], stage5_32[16], stage5_32[17]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[0],stage6_34[2],stage6_33[3],stage6_32[3]}
   );
   gpc606_5 gpc9681 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[1],stage6_35[1],stage6_34[3],stage6_33[4]}
   );
   gpc606_5 gpc9682 (
      {stage5_33[6], stage5_33[7], stage5_33[8], stage5_33[9], stage5_33[10], stage5_33[11]},
      {stage5_35[6], stage5_35[7], stage5_35[8], stage5_35[9], stage5_35[10], stage5_35[11]},
      {stage6_37[1],stage6_36[2],stage6_35[2],stage6_34[4],stage6_33[5]}
   );
   gpc615_5 gpc9683 (
      {stage5_34[6], stage5_34[7], stage5_34[8], stage5_34[9], stage5_34[10]},
      {stage5_35[12]},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5]},
      {stage6_38[0],stage6_37[2],stage6_36[3],stage6_35[3],stage6_34[5]}
   );
   gpc606_5 gpc9684 (
      {stage5_36[6], stage5_36[7], stage5_36[8], stage5_36[9], stage5_36[10], stage5_36[11]},
      {stage5_38[0], stage5_38[1], stage5_38[2], stage5_38[3], stage5_38[4], stage5_38[5]},
      {stage6_40[0],stage6_39[0],stage6_38[1],stage6_37[3],stage6_36[4]}
   );
   gpc2135_5 gpc9685 (
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4]},
      {stage5_38[6], stage5_38[7], stage5_38[8]},
      {stage5_39[0]},
      {stage5_40[0], stage5_40[1]},
      {stage6_41[0],stage6_40[1],stage6_39[1],stage6_38[2],stage6_37[4]}
   );
   gpc606_5 gpc9686 (
      {stage5_37[5], stage5_37[6], stage5_37[7], stage5_37[8], stage5_37[9], stage5_37[10]},
      {stage5_39[1], stage5_39[2], stage5_39[3], stage5_39[4], stage5_39[5], stage5_39[6]},
      {stage6_41[1],stage6_40[2],stage6_39[2],stage6_38[3],stage6_37[5]}
   );
   gpc23_3 gpc9687 (
      {stage5_39[7], stage5_39[8], stage5_39[9]},
      {stage5_40[2], stage5_40[3]},
      {stage6_41[2],stage6_40[3],stage6_39[3]}
   );
   gpc606_5 gpc9688 (
      {stage5_40[4], stage5_40[5], stage5_40[6], stage5_40[7], stage5_40[8], stage5_40[9]},
      {stage5_42[0], stage5_42[1], stage5_42[2], stage5_42[3], stage5_42[4], stage5_42[5]},
      {stage6_44[0],stage6_43[0],stage6_42[0],stage6_41[3],stage6_40[4]}
   );
   gpc606_5 gpc9689 (
      {stage5_41[0], stage5_41[1], stage5_41[2], stage5_41[3], stage5_41[4], stage5_41[5]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3], stage5_43[4], stage5_43[5]},
      {stage6_45[0],stage6_44[1],stage6_43[1],stage6_42[1],stage6_41[4]}
   );
   gpc615_5 gpc9690 (
      {stage5_42[6], stage5_42[7], stage5_42[8], stage5_42[9], stage5_42[10]},
      {stage5_43[6]},
      {stage5_44[0], stage5_44[1], stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5]},
      {stage6_46[0],stage6_45[1],stage6_44[2],stage6_43[2],stage6_42[2]}
   );
   gpc615_5 gpc9691 (
      {stage5_42[11], stage5_42[12], stage5_42[13], stage5_42[14], stage5_42[15]},
      {stage5_43[7]},
      {stage5_44[6], stage5_44[7], stage5_44[8], stage5_44[9], stage5_44[10], stage5_44[11]},
      {stage6_46[1],stage6_45[2],stage6_44[3],stage6_43[3],stage6_42[3]}
   );
   gpc1163_5 gpc9692 (
      {stage5_45[0], stage5_45[1], stage5_45[2]},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage5_47[0]},
      {stage5_48[0]},
      {stage6_49[0],stage6_48[0],stage6_47[0],stage6_46[2],stage6_45[3]}
   );
   gpc1163_5 gpc9693 (
      {stage5_45[3], stage5_45[4], stage5_45[5]},
      {stage5_46[6], stage5_46[7], stage5_46[8], stage5_46[9], stage5_46[10], stage5_46[11]},
      {stage5_47[1]},
      {stage5_48[1]},
      {stage6_49[1],stage6_48[1],stage6_47[1],stage6_46[3],stage6_45[4]}
   );
   gpc606_5 gpc9694 (
      {stage5_45[6], stage5_45[7], stage5_45[8], stage5_45[9], stage5_45[10], stage5_45[11]},
      {stage5_47[2], stage5_47[3], stage5_47[4], stage5_47[5], stage5_47[6], stage5_47[7]},
      {stage6_49[2],stage6_48[2],stage6_47[2],stage6_46[4],stage6_45[5]}
   );
   gpc606_5 gpc9695 (
      {stage5_48[2], stage5_48[3], stage5_48[4], stage5_48[5], stage5_48[6], stage5_48[7]},
      {stage5_50[0], stage5_50[1], stage5_50[2], stage5_50[3], stage5_50[4], stage5_50[5]},
      {stage6_52[0],stage6_51[0],stage6_50[0],stage6_49[3],stage6_48[3]}
   );
   gpc606_5 gpc9696 (
      {stage5_48[8], stage5_48[9], stage5_48[10], stage5_48[11], stage5_48[12], stage5_48[13]},
      {stage5_50[6], stage5_50[7], stage5_50[8], stage5_50[9], stage5_50[10], stage5_50[11]},
      {stage6_52[1],stage6_51[1],stage6_50[1],stage6_49[4],stage6_48[4]}
   );
   gpc606_5 gpc9697 (
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5]},
      {stage5_51[0], stage5_51[1], stage5_51[2], stage5_51[3], stage5_51[4], stage5_51[5]},
      {stage6_53[0],stage6_52[2],stage6_51[2],stage6_50[2],stage6_49[5]}
   );
   gpc7_3 gpc9698 (
      {stage5_51[6], stage5_51[7], stage5_51[8], stage5_51[9], stage5_51[10], stage5_51[11], stage5_51[12]},
      {stage6_53[1],stage6_52[3],stage6_51[3]}
   );
   gpc623_5 gpc9699 (
      {stage5_51[13], stage5_51[14], stage5_51[15]},
      {stage5_52[0], stage5_52[1]},
      {stage5_53[0], stage5_53[1], stage5_53[2], stage5_53[3], stage5_53[4], stage5_53[5]},
      {stage6_55[0],stage6_54[0],stage6_53[2],stage6_52[4],stage6_51[4]}
   );
   gpc117_4 gpc9700 (
      {stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5], stage5_52[6], stage5_52[7], stage5_52[8]},
      {stage5_53[6]},
      {stage5_54[0]},
      {stage6_55[1],stage6_54[1],stage6_53[3],stage6_52[5]}
   );
   gpc117_4 gpc9701 (
      {stage5_53[7], stage5_53[8], stage5_53[9], stage5_53[10], stage5_53[11], stage5_53[12], 1'b0},
      {stage5_54[1]},
      {stage5_55[0]},
      {stage6_56[0],stage6_55[2],stage6_54[2],stage6_53[4]}
   );
   gpc135_4 gpc9702 (
      {stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5], stage5_54[6]},
      {stage5_55[1], stage5_55[2], stage5_55[3]},
      {stage5_56[0]},
      {stage6_57[0],stage6_56[1],stage6_55[3],stage6_54[3]}
   );
   gpc135_4 gpc9703 (
      {stage5_54[7], stage5_54[8], stage5_54[9], stage5_54[10], stage5_54[11]},
      {stage5_55[4], stage5_55[5], stage5_55[6]},
      {stage5_56[1]},
      {stage6_57[1],stage6_56[2],stage6_55[4],stage6_54[4]}
   );
   gpc135_4 gpc9704 (
      {stage5_54[12], stage5_54[13], stage5_54[14], stage5_54[15], stage5_54[16]},
      {stage5_55[7], stage5_55[8], stage5_55[9]},
      {stage5_56[2]},
      {stage6_57[2],stage6_56[3],stage6_55[5],stage6_54[5]}
   );
   gpc615_5 gpc9705 (
      {stage5_55[10], stage5_55[11], stage5_55[12], stage5_55[13], stage5_55[14]},
      {stage5_56[3]},
      {stage5_57[0], stage5_57[1], stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5]},
      {stage6_59[0],stage6_58[0],stage6_57[3],stage6_56[4],stage6_55[6]}
   );
   gpc615_5 gpc9706 (
      {stage5_55[15], stage5_55[16], stage5_55[17], stage5_55[18], stage5_55[19]},
      {stage5_56[4]},
      {stage5_57[6], stage5_57[7], stage5_57[8], stage5_57[9], stage5_57[10], stage5_57[11]},
      {stage6_59[1],stage6_58[1],stage6_57[4],stage6_56[5],stage6_55[7]}
   );
   gpc2135_5 gpc9707 (
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4]},
      {stage5_59[0], stage5_59[1], stage5_59[2]},
      {stage5_60[0]},
      {stage5_61[0], stage5_61[1]},
      {stage6_62[0],stage6_61[0],stage6_60[0],stage6_59[2],stage6_58[2]}
   );
   gpc2135_5 gpc9708 (
      {stage5_58[5], stage5_58[6], stage5_58[7], stage5_58[8], stage5_58[9]},
      {stage5_59[3], stage5_59[4], stage5_59[5]},
      {stage5_60[1]},
      {stage5_61[2], stage5_61[3]},
      {stage6_62[1],stage6_61[1],stage6_60[1],stage6_59[3],stage6_58[3]}
   );
   gpc2135_5 gpc9709 (
      {stage5_58[10], stage5_58[11], stage5_58[12], stage5_58[13], stage5_58[14]},
      {stage5_59[6], stage5_59[7], 1'b0},
      {stage5_60[2]},
      {stage5_61[4], stage5_61[5]},
      {stage6_62[2],stage6_61[2],stage6_60[2],stage6_59[4],stage6_58[4]}
   );
   gpc606_5 gpc9710 (
      {stage5_60[3], stage5_60[4], stage5_60[5], stage5_60[6], stage5_60[7], stage5_60[8]},
      {stage5_62[0], stage5_62[1], stage5_62[2], stage5_62[3], stage5_62[4], stage5_62[5]},
      {stage6_64[0],stage6_63[0],stage6_62[3],stage6_61[3],stage6_60[3]}
   );
   gpc606_5 gpc9711 (
      {stage5_60[9], stage5_60[10], stage5_60[11], stage5_60[12], stage5_60[13], stage5_60[14]},
      {stage5_62[6], stage5_62[7], stage5_62[8], stage5_62[9], stage5_62[10], stage5_62[11]},
      {stage6_64[1],stage6_63[1],stage6_62[4],stage6_61[4],stage6_60[4]}
   );
   gpc207_4 gpc9712 (
      {stage5_61[6], stage5_61[7], stage5_61[8], stage5_61[9], stage5_61[10], stage5_61[11], stage5_61[12]},
      {stage5_63[0], stage5_63[1]},
      {stage6_64[2],stage6_63[2],stage6_62[5],stage6_61[5]}
   );
   gpc606_5 gpc9713 (
      {stage5_63[2], stage5_63[3], stage5_63[4], stage5_63[5], stage5_63[6], stage5_63[7]},
      {stage5_65[0], stage5_65[1], stage5_65[2], stage5_65[3], stage5_65[4], stage5_65[5]},
      {stage6_67[0],stage6_66[0],stage6_65[0],stage6_64[3],stage6_63[3]}
   );
   gpc1406_5 gpc9714 (
      {stage5_64[0], stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage5_66[0], stage5_66[1], stage5_66[2], stage5_66[3]},
      {stage5_67[0]},
      {stage6_68[0],stage6_67[1],stage6_66[1],stage6_65[1],stage6_64[4]}
   );
   gpc1406_5 gpc9715 (
      {stage5_64[6], stage5_64[7], stage5_64[8], stage5_64[9], stage5_64[10], stage5_64[11]},
      {stage5_66[4], stage5_66[5], stage5_66[6], stage5_66[7]},
      {stage5_67[1]},
      {stage6_68[1],stage6_67[2],stage6_66[2],stage6_65[2],stage6_64[5]}
   );
   gpc1406_5 gpc9716 (
      {stage5_65[6], stage5_65[7], stage5_65[8], stage5_65[9], stage5_65[10], stage5_65[11]},
      {stage5_67[2], stage5_67[3], stage5_67[4], stage5_67[5]},
      {stage5_68[0]},
      {stage6_69[0],stage6_68[2],stage6_67[3],stage6_66[3],stage6_65[3]}
   );
   gpc606_5 gpc9717 (
      {stage5_65[12], stage5_65[13], stage5_65[14], stage5_65[15], stage5_65[16], stage5_65[17]},
      {stage5_67[6], stage5_67[7], stage5_67[8], stage5_67[9], stage5_67[10], 1'b0},
      {stage6_69[1],stage6_68[3],stage6_67[4],stage6_66[4],stage6_65[4]}
   );
   gpc1_1 gpc9718 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc9719 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc9720 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc9721 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc9722 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc9723 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc9724 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc9725 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc9726 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc9727 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc9728 (
      {stage5_2[3]},
      {stage6_2[3]}
   );
   gpc1_1 gpc9729 (
      {stage5_2[4]},
      {stage6_2[4]}
   );
   gpc1_1 gpc9730 (
      {stage5_4[8]},
      {stage6_4[3]}
   );
   gpc1_1 gpc9731 (
      {stage5_4[9]},
      {stage6_4[4]}
   );
   gpc1_1 gpc9732 (
      {stage5_4[10]},
      {stage6_4[5]}
   );
   gpc1_1 gpc9733 (
      {stage5_6[6]},
      {stage6_6[4]}
   );
   gpc1_1 gpc9734 (
      {stage5_6[7]},
      {stage6_6[5]}
   );
   gpc1_1 gpc9735 (
      {stage5_6[8]},
      {stage6_6[6]}
   );
   gpc1_1 gpc9736 (
      {stage5_6[9]},
      {stage6_6[7]}
   );
   gpc1_1 gpc9737 (
      {stage5_9[6]},
      {stage6_9[5]}
   );
   gpc1_1 gpc9738 (
      {stage5_9[7]},
      {stage6_9[6]}
   );
   gpc1_1 gpc9739 (
      {stage5_9[8]},
      {stage6_9[7]}
   );
   gpc1_1 gpc9740 (
      {stage5_9[9]},
      {stage6_9[8]}
   );
   gpc1_1 gpc9741 (
      {stage5_9[10]},
      {stage6_9[9]}
   );
   gpc1_1 gpc9742 (
      {stage5_13[10]},
      {stage6_13[5]}
   );
   gpc1_1 gpc9743 (
      {stage5_13[11]},
      {stage6_13[6]}
   );
   gpc1_1 gpc9744 (
      {stage5_13[12]},
      {stage6_13[7]}
   );
   gpc1_1 gpc9745 (
      {stage5_13[13]},
      {stage6_13[8]}
   );
   gpc1_1 gpc9746 (
      {stage5_13[14]},
      {stage6_13[9]}
   );
   gpc1_1 gpc9747 (
      {stage5_24[8]},
      {stage6_24[6]}
   );
   gpc1_1 gpc9748 (
      {stage5_26[11]},
      {stage6_26[4]}
   );
   gpc1_1 gpc9749 (
      {stage5_26[12]},
      {stage6_26[5]}
   );
   gpc1_1 gpc9750 (
      {stage5_26[13]},
      {stage6_26[6]}
   );
   gpc1_1 gpc9751 (
      {stage5_26[14]},
      {stage6_26[7]}
   );
   gpc1_1 gpc9752 (
      {stage5_28[7]},
      {stage6_28[3]}
   );
   gpc1_1 gpc9753 (
      {stage5_28[8]},
      {stage6_28[4]}
   );
   gpc1_1 gpc9754 (
      {stage5_28[9]},
      {stage6_28[5]}
   );
   gpc1_1 gpc9755 (
      {stage5_29[12]},
      {stage6_29[3]}
   );
   gpc1_1 gpc9756 (
      {stage5_29[13]},
      {stage6_29[4]}
   );
   gpc1_1 gpc9757 (
      {stage5_29[14]},
      {stage6_29[5]}
   );
   gpc1_1 gpc9758 (
      {stage5_31[8]},
      {stage6_31[4]}
   );
   gpc1_1 gpc9759 (
      {stage5_31[9]},
      {stage6_31[5]}
   );
   gpc1_1 gpc9760 (
      {stage5_32[18]},
      {stage6_32[4]}
   );
   gpc1_1 gpc9761 (
      {stage5_32[19]},
      {stage6_32[5]}
   );
   gpc1_1 gpc9762 (
      {stage5_34[11]},
      {stage6_34[6]}
   );
   gpc1_1 gpc9763 (
      {stage5_34[12]},
      {stage6_34[7]}
   );
   gpc1_1 gpc9764 (
      {stage5_34[13]},
      {stage6_34[8]}
   );
   gpc1_1 gpc9765 (
      {stage5_35[13]},
      {stage6_35[4]}
   );
   gpc1_1 gpc9766 (
      {stage5_36[12]},
      {stage6_36[5]}
   );
   gpc1_1 gpc9767 (
      {stage5_38[9]},
      {stage6_38[4]}
   );
   gpc1_1 gpc9768 (
      {stage5_40[10]},
      {stage6_40[5]}
   );
   gpc1_1 gpc9769 (
      {stage5_41[6]},
      {stage6_41[5]}
   );
   gpc1_1 gpc9770 (
      {stage5_41[7]},
      {stage6_41[6]}
   );
   gpc1_1 gpc9771 (
      {stage5_41[8]},
      {stage6_41[7]}
   );
   gpc1_1 gpc9772 (
      {stage5_42[16]},
      {stage6_42[4]}
   );
   gpc1_1 gpc9773 (
      {stage5_42[17]},
      {stage6_42[5]}
   );
   gpc1_1 gpc9774 (
      {stage5_42[18]},
      {stage6_42[6]}
   );
   gpc1_1 gpc9775 (
      {stage5_43[8]},
      {stage6_43[4]}
   );
   gpc1_1 gpc9776 (
      {stage5_43[9]},
      {stage6_43[5]}
   );
   gpc1_1 gpc9777 (
      {stage5_43[10]},
      {stage6_43[6]}
   );
   gpc1_1 gpc9778 (
      {stage5_44[12]},
      {stage6_44[4]}
   );
   gpc1_1 gpc9779 (
      {stage5_45[12]},
      {stage6_45[6]}
   );
   gpc1_1 gpc9780 (
      {stage5_45[13]},
      {stage6_45[7]}
   );
   gpc1_1 gpc9781 (
      {stage5_45[14]},
      {stage6_45[8]}
   );
   gpc1_1 gpc9782 (
      {stage5_47[8]},
      {stage6_47[3]}
   );
   gpc1_1 gpc9783 (
      {stage5_47[9]},
      {stage6_47[4]}
   );
   gpc1_1 gpc9784 (
      {stage5_47[10]},
      {stage6_47[5]}
   );
   gpc1_1 gpc9785 (
      {stage5_47[11]},
      {stage6_47[6]}
   );
   gpc1_1 gpc9786 (
      {stage5_51[16]},
      {stage6_51[5]}
   );
   gpc1_1 gpc9787 (
      {stage5_51[17]},
      {stage6_51[6]}
   );
   gpc1_1 gpc9788 (
      {stage5_51[18]},
      {stage6_51[7]}
   );
   gpc1_1 gpc9789 (
      {stage5_52[9]},
      {stage6_52[6]}
   );
   gpc1_1 gpc9790 (
      {stage5_55[20]},
      {stage6_55[8]}
   );
   gpc1_1 gpc9791 (
      {stage5_55[21]},
      {stage6_55[9]}
   );
   gpc1_1 gpc9792 (
      {stage5_56[5]},
      {stage6_56[6]}
   );
   gpc1_1 gpc9793 (
      {stage5_56[6]},
      {stage6_56[7]}
   );
   gpc1_1 gpc9794 (
      {stage5_56[7]},
      {stage6_56[8]}
   );
   gpc1_1 gpc9795 (
      {stage5_56[8]},
      {stage6_56[9]}
   );
   gpc1_1 gpc9796 (
      {stage5_57[12]},
      {stage6_57[5]}
   );
   gpc1_1 gpc9797 (
      {stage5_57[13]},
      {stage6_57[6]}
   );
   gpc1_1 gpc9798 (
      {stage5_58[15]},
      {stage6_58[5]}
   );
   gpc1_1 gpc9799 (
      {stage5_61[13]},
      {stage6_61[6]}
   );
   gpc1_1 gpc9800 (
      {stage5_61[14]},
      {stage6_61[7]}
   );
   gpc1_1 gpc9801 (
      {stage5_61[15]},
      {stage6_61[8]}
   );
   gpc1_1 gpc9802 (
      {stage5_63[8]},
      {stage6_63[4]}
   );
   gpc1_1 gpc9803 (
      {stage5_64[12]},
      {stage6_64[6]}
   );
   gpc1_1 gpc9804 (
      {stage5_64[13]},
      {stage6_64[7]}
   );
   gpc1_1 gpc9805 (
      {stage5_64[14]},
      {stage6_64[8]}
   );
   gpc1_1 gpc9806 (
      {stage5_68[1]},
      {stage6_68[4]}
   );
   gpc1_1 gpc9807 (
      {stage5_68[2]},
      {stage6_68[5]}
   );
   gpc1_1 gpc9808 (
      {stage5_68[3]},
      {stage6_68[6]}
   );
   gpc1_1 gpc9809 (
      {stage5_68[4]},
      {stage6_68[7]}
   );
   gpc1_1 gpc9810 (
      {stage5_68[5]},
      {stage6_68[8]}
   );
   gpc1_1 gpc9811 (
      {stage5_68[6]},
      {stage6_68[9]}
   );
   gpc1_1 gpc9812 (
      {stage5_68[7]},
      {stage6_68[10]}
   );
   gpc1_1 gpc9813 (
      {stage5_68[8]},
      {stage6_68[11]}
   );
   gpc1_1 gpc9814 (
      {stage5_68[9]},
      {stage6_68[12]}
   );
   gpc1_1 gpc9815 (
      {stage5_68[10]},
      {stage6_68[13]}
   );
   gpc1_1 gpc9816 (
      {stage5_68[11]},
      {stage6_68[14]}
   );
   gpc1_1 gpc9817 (
      {stage5_68[12]},
      {stage6_68[15]}
   );
   gpc1_1 gpc9818 (
      {stage5_68[13]},
      {stage6_68[16]}
   );
   gpc1_1 gpc9819 (
      {stage5_69[0]},
      {stage6_69[2]}
   );
   gpc1_1 gpc9820 (
      {stage5_69[1]},
      {stage6_69[3]}
   );
   gpc1_1 gpc9821 (
      {stage5_69[2]},
      {stage6_69[4]}
   );
   gpc1_1 gpc9822 (
      {stage5_70[0]},
      {stage6_70[0]}
   );
   gpc1406_5 gpc9823 (
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3], stage6_4[4], stage6_4[5]},
      {stage6_6[0], stage6_6[1], stage6_6[2], stage6_6[3]},
      {stage6_7[0]},
      {stage7_8[0],stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0]}
   );
   gpc2135_5 gpc9824 (
      {stage6_5[0], stage6_5[1], stage6_5[2], stage6_5[3], 1'b0},
      {stage6_6[4], stage6_6[5], stage6_6[6]},
      {stage6_7[1]},
      {stage6_8[0], stage6_8[1]},
      {stage7_9[0],stage7_8[1],stage7_7[1],stage7_6[1],stage7_5[1]}
   );
   gpc623_5 gpc9825 (
      {stage6_7[2], stage6_7[3], stage6_7[4]},
      {stage6_8[2], stage6_8[3]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4], stage6_9[5]},
      {stage7_11[0],stage7_10[0],stage7_9[1],stage7_8[2],stage7_7[2]}
   );
   gpc615_5 gpc9826 (
      {stage6_10[0], stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4]},
      {stage6_11[0]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage7_14[0],stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[1]}
   );
   gpc615_5 gpc9827 (
      {stage6_11[1], stage6_11[2], stage6_11[3], stage6_11[4], stage6_11[5]},
      {stage6_12[6]},
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5]},
      {stage7_15[0],stage7_14[1],stage7_13[1],stage7_12[1],stage7_11[2]}
   );
   gpc7_3 gpc9828 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5], stage6_14[6]},
      {stage7_16[0],stage7_15[1],stage7_14[2]}
   );
   gpc623_5 gpc9829 (
      {stage6_15[0], stage6_15[1], stage6_15[2]},
      {stage6_16[0], stage6_16[1]},
      {stage6_17[0], stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4], 1'b0},
      {stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[2]}
   );
   gpc606_5 gpc9830 (
      {stage6_16[2], stage6_16[3], stage6_16[4], 1'b0, 1'b0, 1'b0},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage7_20[0],stage7_19[1],stage7_18[1],stage7_17[1],stage7_16[2]}
   );
   gpc15_3 gpc9831 (
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4]},
      {stage6_21[0]},
      {stage7_22[0],stage7_21[0],stage7_20[1]}
   );
   gpc207_4 gpc9832 (
      {stage6_23[0], stage6_23[1], stage6_23[2], stage6_23[3], stage6_23[4], stage6_23[5], stage6_23[6]},
      {stage6_25[0], stage6_25[1]},
      {stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[0]}
   );
   gpc15_3 gpc9833 (
      {stage6_24[0], stage6_24[1], stage6_24[2], stage6_24[3], stage6_24[4]},
      {stage6_25[2]},
      {stage7_26[1],stage7_25[1],stage7_24[1]}
   );
   gpc615_5 gpc9834 (
      {stage6_26[0], stage6_26[1], stage6_26[2], stage6_26[3], stage6_26[4]},
      {stage6_27[0]},
      {stage6_28[0], stage6_28[1], stage6_28[2], stage6_28[3], stage6_28[4], stage6_28[5]},
      {stage7_30[0],stage7_29[0],stage7_28[0],stage7_27[0],stage7_26[2]}
   );
   gpc3_2 gpc9835 (
      {stage6_29[0], stage6_29[1], stage6_29[2]},
      {stage7_30[1],stage7_29[1]}
   );
   gpc615_5 gpc9836 (
      {stage6_31[0], stage6_31[1], stage6_31[2], stage6_31[3], stage6_31[4]},
      {stage6_32[0]},
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3], stage6_33[4], stage6_33[5]},
      {stage7_35[0],stage7_34[0],stage7_33[0],stage7_32[0],stage7_31[0]}
   );
   gpc615_5 gpc9837 (
      {stage6_34[0], stage6_34[1], stage6_34[2], stage6_34[3], stage6_34[4]},
      {stage6_35[0]},
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5]},
      {stage7_38[0],stage7_37[0],stage7_36[0],stage7_35[1],stage7_34[1]}
   );
   gpc606_5 gpc9838 (
      {stage6_37[0], stage6_37[1], stage6_37[2], stage6_37[3], stage6_37[4], stage6_37[5]},
      {stage6_39[0], stage6_39[1], stage6_39[2], stage6_39[3], 1'b0, 1'b0},
      {stage7_41[0],stage7_40[0],stage7_39[0],stage7_38[1],stage7_37[1]}
   );
   gpc15_3 gpc9839 (
      {stage6_41[0], stage6_41[1], stage6_41[2], stage6_41[3], stage6_41[4]},
      {stage6_42[0]},
      {stage7_43[0],stage7_42[0],stage7_41[1]}
   );
   gpc615_5 gpc9840 (
      {stage6_42[1], stage6_42[2], stage6_42[3], stage6_42[4], stage6_42[5]},
      {stage6_43[0]},
      {stage6_44[0], stage6_44[1], stage6_44[2], stage6_44[3], stage6_44[4], 1'b0},
      {stage7_46[0],stage7_45[0],stage7_44[0],stage7_43[1],stage7_42[1]}
   );
   gpc615_5 gpc9841 (
      {stage6_43[1], stage6_43[2], stage6_43[3], stage6_43[4], stage6_43[5]},
      {1'b0},
      {stage6_45[0], stage6_45[1], stage6_45[2], stage6_45[3], stage6_45[4], stage6_45[5]},
      {stage7_47[0],stage7_46[1],stage7_45[1],stage7_44[1],stage7_43[2]}
   );
   gpc615_5 gpc9842 (
      {stage6_46[0], stage6_46[1], stage6_46[2], stage6_46[3], stage6_46[4]},
      {stage6_47[0]},
      {stage6_48[0], stage6_48[1], stage6_48[2], stage6_48[3], stage6_48[4], 1'b0},
      {stage7_50[0],stage7_49[0],stage7_48[0],stage7_47[1],stage7_46[2]}
   );
   gpc606_5 gpc9843 (
      {stage6_49[0], stage6_49[1], stage6_49[2], stage6_49[3], stage6_49[4], stage6_49[5]},
      {stage6_51[0], stage6_51[1], stage6_51[2], stage6_51[3], stage6_51[4], stage6_51[5]},
      {stage7_53[0],stage7_52[0],stage7_51[0],stage7_50[1],stage7_49[1]}
   );
   gpc3_2 gpc9844 (
      {stage6_50[0], stage6_50[1], stage6_50[2]},
      {stage7_51[1],stage7_50[2]}
   );
   gpc615_5 gpc9845 (
      {stage6_52[0], stage6_52[1], stage6_52[2], stage6_52[3], stage6_52[4]},
      {stage6_53[0]},
      {stage6_54[0], stage6_54[1], stage6_54[2], stage6_54[3], stage6_54[4], stage6_54[5]},
      {stage7_56[0],stage7_55[0],stage7_54[0],stage7_53[1],stage7_52[1]}
   );
   gpc615_5 gpc9846 (
      {stage6_55[0], stage6_55[1], stage6_55[2], stage6_55[3], stage6_55[4]},
      {stage6_56[0]},
      {stage6_57[0], stage6_57[1], stage6_57[2], stage6_57[3], stage6_57[4], stage6_57[5]},
      {stage7_59[0],stage7_58[0],stage7_57[0],stage7_56[1],stage7_55[1]}
   );
   gpc615_5 gpc9847 (
      {stage6_56[1], stage6_56[2], stage6_56[3], stage6_56[4], stage6_56[5]},
      {stage6_57[6]},
      {stage6_58[0], stage6_58[1], stage6_58[2], stage6_58[3], stage6_58[4], stage6_58[5]},
      {stage7_60[0],stage7_59[1],stage7_58[1],stage7_57[1],stage7_56[2]}
   );
   gpc135_4 gpc9848 (
      {stage6_61[0], stage6_61[1], stage6_61[2], stage6_61[3], stage6_61[4]},
      {stage6_62[0], stage6_62[1], stage6_62[2]},
      {stage6_63[0]},
      {stage7_64[0],stage7_63[0],stage7_62[0],stage7_61[0]}
   );
   gpc135_4 gpc9849 (
      {stage6_61[5], stage6_61[6], stage6_61[7], stage6_61[8], 1'b0},
      {stage6_62[3], stage6_62[4], stage6_62[5]},
      {stage6_63[1]},
      {stage7_64[1],stage7_63[1],stage7_62[1],stage7_61[1]}
   );
   gpc223_4 gpc9850 (
      {stage6_63[2], stage6_63[3], stage6_63[4]},
      {stage6_64[0], stage6_64[1]},
      {stage6_65[0], stage6_65[1]},
      {stage7_66[0],stage7_65[0],stage7_64[2],stage7_63[2]}
   );
   gpc7_3 gpc9851 (
      {stage6_64[2], stage6_64[3], stage6_64[4], stage6_64[5], stage6_64[6], stage6_64[7], stage6_64[8]},
      {stage7_66[1],stage7_65[1],stage7_64[3]}
   );
   gpc3_2 gpc9852 (
      {stage6_65[2], stage6_65[3], stage6_65[4]},
      {stage7_66[2],stage7_65[2]}
   );
   gpc1163_5 gpc9853 (
      {stage6_66[0], stage6_66[1], stage6_66[2]},
      {stage6_67[0], stage6_67[1], stage6_67[2], stage6_67[3], stage6_67[4], 1'b0},
      {stage6_68[0]},
      {stage6_69[0]},
      {stage7_70[0],stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[3]}
   );
   gpc117_4 gpc9854 (
      {stage6_68[1], stage6_68[2], stage6_68[3], stage6_68[4], stage6_68[5], stage6_68[6], stage6_68[7]},
      {stage6_69[1]},
      {stage6_70[0]},
      {stage7_71[0],stage7_70[1],stage7_69[1],stage7_68[1]}
   );
   gpc117_4 gpc9855 (
      {stage6_68[8], stage6_68[9], stage6_68[10], stage6_68[11], stage6_68[12], stage6_68[13], stage6_68[14]},
      {stage6_69[2]},
      {1'b0},
      {stage7_71[1],stage7_70[2],stage7_69[2],stage7_68[2]}
   );
   gpc1_1 gpc9856 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc9857 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc9858 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc9859 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc9860 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc9861 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc9862 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc9863 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc9864 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc9865 (
      {stage6_2[2]},
      {stage7_2[2]}
   );
   gpc1_1 gpc9866 (
      {stage6_2[3]},
      {stage7_2[3]}
   );
   gpc1_1 gpc9867 (
      {stage6_2[4]},
      {stage7_2[4]}
   );
   gpc1_1 gpc9868 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc9869 (
      {stage6_3[1]},
      {stage7_3[1]}
   );
   gpc1_1 gpc9870 (
      {stage6_6[7]},
      {stage7_6[2]}
   );
   gpc1_1 gpc9871 (
      {stage6_8[4]},
      {stage7_8[3]}
   );
   gpc1_1 gpc9872 (
      {stage6_8[5]},
      {stage7_8[4]}
   );
   gpc1_1 gpc9873 (
      {stage6_9[6]},
      {stage7_9[2]}
   );
   gpc1_1 gpc9874 (
      {stage6_9[7]},
      {stage7_9[3]}
   );
   gpc1_1 gpc9875 (
      {stage6_9[8]},
      {stage7_9[4]}
   );
   gpc1_1 gpc9876 (
      {stage6_9[9]},
      {stage7_9[5]}
   );
   gpc1_1 gpc9877 (
      {stage6_11[6]},
      {stage7_11[3]}
   );
   gpc1_1 gpc9878 (
      {stage6_13[6]},
      {stage7_13[2]}
   );
   gpc1_1 gpc9879 (
      {stage6_13[7]},
      {stage7_13[3]}
   );
   gpc1_1 gpc9880 (
      {stage6_13[8]},
      {stage7_13[4]}
   );
   gpc1_1 gpc9881 (
      {stage6_13[9]},
      {stage7_13[5]}
   );
   gpc1_1 gpc9882 (
      {stage6_15[3]},
      {stage7_15[3]}
   );
   gpc1_1 gpc9883 (
      {stage6_15[4]},
      {stage7_15[4]}
   );
   gpc1_1 gpc9884 (
      {stage6_15[5]},
      {stage7_15[5]}
   );
   gpc1_1 gpc9885 (
      {stage6_19[0]},
      {stage7_19[2]}
   );
   gpc1_1 gpc9886 (
      {stage6_19[1]},
      {stage7_19[3]}
   );
   gpc1_1 gpc9887 (
      {stage6_19[2]},
      {stage7_19[4]}
   );
   gpc1_1 gpc9888 (
      {stage6_19[3]},
      {stage7_19[5]}
   );
   gpc1_1 gpc9889 (
      {stage6_19[4]},
      {stage7_19[6]}
   );
   gpc1_1 gpc9890 (
      {stage6_20[5]},
      {stage7_20[2]}
   );
   gpc1_1 gpc9891 (
      {stage6_21[1]},
      {stage7_21[1]}
   );
   gpc1_1 gpc9892 (
      {stage6_21[2]},
      {stage7_21[2]}
   );
   gpc1_1 gpc9893 (
      {stage6_21[3]},
      {stage7_21[3]}
   );
   gpc1_1 gpc9894 (
      {stage6_21[4]},
      {stage7_21[4]}
   );
   gpc1_1 gpc9895 (
      {stage6_21[5]},
      {stage7_21[5]}
   );
   gpc1_1 gpc9896 (
      {stage6_22[0]},
      {stage7_22[1]}
   );
   gpc1_1 gpc9897 (
      {stage6_22[1]},
      {stage7_22[2]}
   );
   gpc1_1 gpc9898 (
      {stage6_22[2]},
      {stage7_22[3]}
   );
   gpc1_1 gpc9899 (
      {stage6_22[3]},
      {stage7_22[4]}
   );
   gpc1_1 gpc9900 (
      {stage6_22[4]},
      {stage7_22[5]}
   );
   gpc1_1 gpc9901 (
      {stage6_22[5]},
      {stage7_22[6]}
   );
   gpc1_1 gpc9902 (
      {stage6_24[5]},
      {stage7_24[2]}
   );
   gpc1_1 gpc9903 (
      {stage6_24[6]},
      {stage7_24[3]}
   );
   gpc1_1 gpc9904 (
      {stage6_26[5]},
      {stage7_26[3]}
   );
   gpc1_1 gpc9905 (
      {stage6_26[6]},
      {stage7_26[4]}
   );
   gpc1_1 gpc9906 (
      {stage6_26[7]},
      {stage7_26[5]}
   );
   gpc1_1 gpc9907 (
      {stage6_27[1]},
      {stage7_27[1]}
   );
   gpc1_1 gpc9908 (
      {stage6_27[2]},
      {stage7_27[2]}
   );
   gpc1_1 gpc9909 (
      {stage6_27[3]},
      {stage7_27[3]}
   );
   gpc1_1 gpc9910 (
      {stage6_27[4]},
      {stage7_27[4]}
   );
   gpc1_1 gpc9911 (
      {stage6_29[3]},
      {stage7_29[2]}
   );
   gpc1_1 gpc9912 (
      {stage6_29[4]},
      {stage7_29[3]}
   );
   gpc1_1 gpc9913 (
      {stage6_29[5]},
      {stage7_29[4]}
   );
   gpc1_1 gpc9914 (
      {stage6_30[0]},
      {stage7_30[2]}
   );
   gpc1_1 gpc9915 (
      {stage6_30[1]},
      {stage7_30[3]}
   );
   gpc1_1 gpc9916 (
      {stage6_30[2]},
      {stage7_30[4]}
   );
   gpc1_1 gpc9917 (
      {stage6_30[3]},
      {stage7_30[5]}
   );
   gpc1_1 gpc9918 (
      {stage6_30[4]},
      {stage7_30[6]}
   );
   gpc1_1 gpc9919 (
      {stage6_31[5]},
      {stage7_31[1]}
   );
   gpc1_1 gpc9920 (
      {stage6_32[1]},
      {stage7_32[1]}
   );
   gpc1_1 gpc9921 (
      {stage6_32[2]},
      {stage7_32[2]}
   );
   gpc1_1 gpc9922 (
      {stage6_32[3]},
      {stage7_32[3]}
   );
   gpc1_1 gpc9923 (
      {stage6_32[4]},
      {stage7_32[4]}
   );
   gpc1_1 gpc9924 (
      {stage6_32[5]},
      {stage7_32[5]}
   );
   gpc1_1 gpc9925 (
      {stage6_34[5]},
      {stage7_34[2]}
   );
   gpc1_1 gpc9926 (
      {stage6_34[6]},
      {stage7_34[3]}
   );
   gpc1_1 gpc9927 (
      {stage6_34[7]},
      {stage7_34[4]}
   );
   gpc1_1 gpc9928 (
      {stage6_34[8]},
      {stage7_34[5]}
   );
   gpc1_1 gpc9929 (
      {stage6_35[1]},
      {stage7_35[2]}
   );
   gpc1_1 gpc9930 (
      {stage6_35[2]},
      {stage7_35[3]}
   );
   gpc1_1 gpc9931 (
      {stage6_35[3]},
      {stage7_35[4]}
   );
   gpc1_1 gpc9932 (
      {stage6_35[4]},
      {stage7_35[5]}
   );
   gpc1_1 gpc9933 (
      {stage6_38[0]},
      {stage7_38[2]}
   );
   gpc1_1 gpc9934 (
      {stage6_38[1]},
      {stage7_38[3]}
   );
   gpc1_1 gpc9935 (
      {stage6_38[2]},
      {stage7_38[4]}
   );
   gpc1_1 gpc9936 (
      {stage6_38[3]},
      {stage7_38[5]}
   );
   gpc1_1 gpc9937 (
      {stage6_38[4]},
      {stage7_38[6]}
   );
   gpc1_1 gpc9938 (
      {stage6_40[0]},
      {stage7_40[1]}
   );
   gpc1_1 gpc9939 (
      {stage6_40[1]},
      {stage7_40[2]}
   );
   gpc1_1 gpc9940 (
      {stage6_40[2]},
      {stage7_40[3]}
   );
   gpc1_1 gpc9941 (
      {stage6_40[3]},
      {stage7_40[4]}
   );
   gpc1_1 gpc9942 (
      {stage6_40[4]},
      {stage7_40[5]}
   );
   gpc1_1 gpc9943 (
      {stage6_40[5]},
      {stage7_40[6]}
   );
   gpc1_1 gpc9944 (
      {stage6_41[5]},
      {stage7_41[2]}
   );
   gpc1_1 gpc9945 (
      {stage6_41[6]},
      {stage7_41[3]}
   );
   gpc1_1 gpc9946 (
      {stage6_41[7]},
      {stage7_41[4]}
   );
   gpc1_1 gpc9947 (
      {stage6_42[6]},
      {stage7_42[2]}
   );
   gpc1_1 gpc9948 (
      {stage6_43[6]},
      {stage7_43[3]}
   );
   gpc1_1 gpc9949 (
      {stage6_45[6]},
      {stage7_45[2]}
   );
   gpc1_1 gpc9950 (
      {stage6_45[7]},
      {stage7_45[3]}
   );
   gpc1_1 gpc9951 (
      {stage6_45[8]},
      {stage7_45[4]}
   );
   gpc1_1 gpc9952 (
      {stage6_47[1]},
      {stage7_47[2]}
   );
   gpc1_1 gpc9953 (
      {stage6_47[2]},
      {stage7_47[3]}
   );
   gpc1_1 gpc9954 (
      {stage6_47[3]},
      {stage7_47[4]}
   );
   gpc1_1 gpc9955 (
      {stage6_47[4]},
      {stage7_47[5]}
   );
   gpc1_1 gpc9956 (
      {stage6_47[5]},
      {stage7_47[6]}
   );
   gpc1_1 gpc9957 (
      {stage6_47[6]},
      {stage7_47[7]}
   );
   gpc1_1 gpc9958 (
      {stage6_51[6]},
      {stage7_51[2]}
   );
   gpc1_1 gpc9959 (
      {stage6_51[7]},
      {stage7_51[3]}
   );
   gpc1_1 gpc9960 (
      {stage6_52[5]},
      {stage7_52[2]}
   );
   gpc1_1 gpc9961 (
      {stage6_52[6]},
      {stage7_52[3]}
   );
   gpc1_1 gpc9962 (
      {stage6_53[1]},
      {stage7_53[2]}
   );
   gpc1_1 gpc9963 (
      {stage6_53[2]},
      {stage7_53[3]}
   );
   gpc1_1 gpc9964 (
      {stage6_53[3]},
      {stage7_53[4]}
   );
   gpc1_1 gpc9965 (
      {stage6_53[4]},
      {stage7_53[5]}
   );
   gpc1_1 gpc9966 (
      {stage6_55[5]},
      {stage7_55[2]}
   );
   gpc1_1 gpc9967 (
      {stage6_55[6]},
      {stage7_55[3]}
   );
   gpc1_1 gpc9968 (
      {stage6_55[7]},
      {stage7_55[4]}
   );
   gpc1_1 gpc9969 (
      {stage6_55[8]},
      {stage7_55[5]}
   );
   gpc1_1 gpc9970 (
      {stage6_55[9]},
      {stage7_55[6]}
   );
   gpc1_1 gpc9971 (
      {stage6_56[6]},
      {stage7_56[3]}
   );
   gpc1_1 gpc9972 (
      {stage6_56[7]},
      {stage7_56[4]}
   );
   gpc1_1 gpc9973 (
      {stage6_56[8]},
      {stage7_56[5]}
   );
   gpc1_1 gpc9974 (
      {stage6_56[9]},
      {stage7_56[6]}
   );
   gpc1_1 gpc9975 (
      {stage6_59[0]},
      {stage7_59[2]}
   );
   gpc1_1 gpc9976 (
      {stage6_59[1]},
      {stage7_59[3]}
   );
   gpc1_1 gpc9977 (
      {stage6_59[2]},
      {stage7_59[4]}
   );
   gpc1_1 gpc9978 (
      {stage6_59[3]},
      {stage7_59[5]}
   );
   gpc1_1 gpc9979 (
      {stage6_59[4]},
      {stage7_59[6]}
   );
   gpc1_1 gpc9980 (
      {stage6_60[0]},
      {stage7_60[1]}
   );
   gpc1_1 gpc9981 (
      {stage6_60[1]},
      {stage7_60[2]}
   );
   gpc1_1 gpc9982 (
      {stage6_60[2]},
      {stage7_60[3]}
   );
   gpc1_1 gpc9983 (
      {stage6_60[3]},
      {stage7_60[4]}
   );
   gpc1_1 gpc9984 (
      {stage6_60[4]},
      {stage7_60[5]}
   );
   gpc1_1 gpc9985 (
      {stage6_66[3]},
      {stage7_66[4]}
   );
   gpc1_1 gpc9986 (
      {stage6_66[4]},
      {stage7_66[5]}
   );
   gpc1_1 gpc9987 (
      {stage6_68[15]},
      {stage7_68[3]}
   );
   gpc1_1 gpc9988 (
      {stage6_68[16]},
      {stage7_68[4]}
   );
   gpc1_1 gpc9989 (
      {stage6_69[3]},
      {stage7_69[3]}
   );
   gpc1_1 gpc9990 (
      {stage6_69[4]},
      {stage7_69[4]}
   );
   gpc1415_5 gpc9991 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4]},
      {stage7_1[0]},
      {stage7_2[0], stage7_2[1], stage7_2[2], stage7_2[3]},
      {stage7_3[0]},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc3_2 gpc9992 (
      {stage7_6[0], stage7_6[1], stage7_6[2]},
      {stage8_7[0],stage8_6[0]}
   );
   gpc3_2 gpc9993 (
      {stage7_7[0], stage7_7[1], stage7_7[2]},
      {stage8_8[0],stage8_7[1]}
   );
   gpc215_4 gpc9994 (
      {stage7_8[0], stage7_8[1], stage7_8[2], stage7_8[3], stage7_8[4]},
      {stage7_9[0]},
      {stage7_10[0], stage7_10[1]},
      {stage8_11[0],stage8_10[0],stage8_9[0],stage8_8[1]}
   );
   gpc1415_5 gpc9995 (
      {stage7_9[1], stage7_9[2], stage7_9[3], stage7_9[4], stage7_9[5]},
      {1'b0},
      {stage7_11[0], stage7_11[1], stage7_11[2], stage7_11[3]},
      {stage7_12[0]},
      {stage8_13[0],stage8_12[0],stage8_11[1],stage8_10[1],stage8_9[1]}
   );
   gpc207_4 gpc9996 (
      {stage7_13[0], stage7_13[1], stage7_13[2], stage7_13[3], stage7_13[4], stage7_13[5], 1'b0},
      {stage7_15[0], stage7_15[1]},
      {stage8_16[0],stage8_15[0],stage8_14[0],stage8_13[1]}
   );
   gpc1343_5 gpc9997 (
      {stage7_14[0], stage7_14[1], stage7_14[2]},
      {stage7_15[2], stage7_15[3], stage7_15[4], stage7_15[5]},
      {stage7_16[0], stage7_16[1], stage7_16[2]},
      {stage7_17[0]},
      {stage8_18[0],stage8_17[0],stage8_16[1],stage8_15[1],stage8_14[1]}
   );
   gpc623_5 gpc9998 (
      {stage7_17[1], 1'b0, 1'b0},
      {stage7_18[0], stage7_18[1]},
      {stage7_19[0], stage7_19[1], stage7_19[2], stage7_19[3], stage7_19[4], stage7_19[5]},
      {stage8_21[0],stage8_20[0],stage8_19[0],stage8_18[1],stage8_17[1]}
   );
   gpc1163_5 gpc9999 (
      {stage7_20[0], stage7_20[1], stage7_20[2]},
      {stage7_21[0], stage7_21[1], stage7_21[2], stage7_21[3], stage7_21[4], stage7_21[5]},
      {stage7_22[0]},
      {stage7_23[0]},
      {stage8_24[0],stage8_23[0],stage8_22[0],stage8_21[1],stage8_20[1]}
   );
   gpc1406_5 gpc10000 (
      {stage7_22[1], stage7_22[2], stage7_22[3], stage7_22[4], stage7_22[5], stage7_22[6]},
      {stage7_24[0], stage7_24[1], stage7_24[2], stage7_24[3]},
      {stage7_25[0]},
      {stage8_26[0],stage8_25[0],stage8_24[1],stage8_23[1],stage8_22[1]}
   );
   gpc7_3 gpc10001 (
      {stage7_26[0], stage7_26[1], stage7_26[2], stage7_26[3], stage7_26[4], stage7_26[5], 1'b0},
      {stage8_28[0],stage8_27[0],stage8_26[1]}
   );
   gpc15_3 gpc10002 (
      {stage7_27[0], stage7_27[1], stage7_27[2], stage7_27[3], stage7_27[4]},
      {stage7_28[0]},
      {stage8_29[0],stage8_28[1],stage8_27[1]}
   );
   gpc135_4 gpc10003 (
      {stage7_29[0], stage7_29[1], stage7_29[2], stage7_29[3], stage7_29[4]},
      {stage7_30[0], stage7_30[1], stage7_30[2]},
      {stage7_31[0]},
      {stage8_32[0],stage8_31[0],stage8_30[0],stage8_29[1]}
   );
   gpc615_5 gpc10004 (
      {stage7_30[3], stage7_30[4], stage7_30[5], stage7_30[6], 1'b0},
      {stage7_31[1]},
      {stage7_32[0], stage7_32[1], stage7_32[2], stage7_32[3], stage7_32[4], stage7_32[5]},
      {stage8_34[0],stage8_33[0],stage8_32[1],stage8_31[1],stage8_30[1]}
   );
   gpc7_3 gpc10005 (
      {stage7_34[0], stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], 1'b0},
      {stage8_36[0],stage8_35[0],stage8_34[1]}
   );
   gpc117_4 gpc10006 (
      {stage7_35[0], stage7_35[1], stage7_35[2], stage7_35[3], stage7_35[4], stage7_35[5], 1'b0},
      {stage7_36[0]},
      {stage7_37[0]},
      {stage8_38[0],stage8_37[0],stage8_36[1],stage8_35[1]}
   );
   gpc7_3 gpc10007 (
      {stage7_38[0], stage7_38[1], stage7_38[2], stage7_38[3], stage7_38[4], stage7_38[5], stage7_38[6]},
      {stage8_40[0],stage8_39[0],stage8_38[1]}
   );
   gpc207_4 gpc10008 (
      {stage7_40[0], stage7_40[1], stage7_40[2], stage7_40[3], stage7_40[4], stage7_40[5], stage7_40[6]},
      {stage7_42[0], stage7_42[1]},
      {stage8_43[0],stage8_42[0],stage8_41[0],stage8_40[1]}
   );
   gpc1415_5 gpc10009 (
      {stage7_41[0], stage7_41[1], stage7_41[2], stage7_41[3], stage7_41[4]},
      {stage7_42[2]},
      {stage7_43[0], stage7_43[1], stage7_43[2], stage7_43[3]},
      {stage7_44[0]},
      {stage8_45[0],stage8_44[0],stage8_43[1],stage8_42[1],stage8_41[1]}
   );
   gpc2135_5 gpc10010 (
      {stage7_45[0], stage7_45[1], stage7_45[2], stage7_45[3], stage7_45[4]},
      {stage7_46[0], stage7_46[1], stage7_46[2]},
      {stage7_47[0]},
      {stage7_48[0], 1'b0},
      {stage8_49[0],stage8_48[0],stage8_47[0],stage8_46[0],stage8_45[1]}
   );
   gpc207_4 gpc10011 (
      {stage7_47[1], stage7_47[2], stage7_47[3], stage7_47[4], stage7_47[5], stage7_47[6], stage7_47[7]},
      {stage7_49[0], stage7_49[1]},
      {stage8_50[0],stage8_49[1],stage8_48[1],stage8_47[1]}
   );
   gpc3_2 gpc10012 (
      {stage7_50[0], stage7_50[1], stage7_50[2]},
      {stage8_51[0],stage8_50[1]}
   );
   gpc615_5 gpc10013 (
      {stage7_51[0], stage7_51[1], stage7_51[2], stage7_51[3], 1'b0},
      {stage7_52[0]},
      {stage7_53[0], stage7_53[1], stage7_53[2], stage7_53[3], stage7_53[4], stage7_53[5]},
      {stage8_55[0],stage8_54[0],stage8_53[0],stage8_52[0],stage8_51[1]}
   );
   gpc3_2 gpc10014 (
      {stage7_52[1], stage7_52[2], stage7_52[3]},
      {stage8_53[1],stage8_52[1]}
   );
   gpc207_4 gpc10015 (
      {stage7_55[0], stage7_55[1], stage7_55[2], stage7_55[3], stage7_55[4], stage7_55[5], stage7_55[6]},
      {stage7_57[0], stage7_57[1]},
      {stage8_58[0],stage8_57[0],stage8_56[0],stage8_55[1]}
   );
   gpc207_4 gpc10016 (
      {stage7_56[0], stage7_56[1], stage7_56[2], stage7_56[3], stage7_56[4], stage7_56[5], stage7_56[6]},
      {stage7_58[0], stage7_58[1]},
      {stage8_59[0],stage8_58[1],stage8_57[1],stage8_56[1]}
   );
   gpc117_4 gpc10017 (
      {stage7_59[0], stage7_59[1], stage7_59[2], stage7_59[3], stage7_59[4], stage7_59[5], stage7_59[6]},
      {stage7_60[0]},
      {stage7_61[0]},
      {stage8_62[0],stage8_61[0],stage8_60[0],stage8_59[1]}
   );
   gpc215_4 gpc10018 (
      {stage7_60[1], stage7_60[2], stage7_60[3], stage7_60[4], stage7_60[5]},
      {stage7_61[1]},
      {stage7_62[0], stage7_62[1]},
      {stage8_63[0],stage8_62[1],stage8_61[1],stage8_60[1]}
   );
   gpc3_2 gpc10019 (
      {stage7_63[0], stage7_63[1], stage7_63[2]},
      {stage8_64[0],stage8_63[1]}
   );
   gpc606_5 gpc10020 (
      {stage7_64[0], stage7_64[1], stage7_64[2], stage7_64[3], 1'b0, 1'b0},
      {stage7_66[0], stage7_66[1], stage7_66[2], stage7_66[3], stage7_66[4], stage7_66[5]},
      {stage8_68[0],stage8_67[0],stage8_66[0],stage8_65[0],stage8_64[1]}
   );
   gpc3_2 gpc10021 (
      {stage7_65[0], stage7_65[1], stage7_65[2]},
      {stage8_66[1],stage8_65[1]}
   );
   gpc615_5 gpc10022 (
      {stage7_68[0], stage7_68[1], stage7_68[2], stage7_68[3], stage7_68[4]},
      {stage7_69[0]},
      {stage7_70[0], stage7_70[1], stage7_70[2], 1'b0, 1'b0, 1'b0},
      {stage8_72[0],stage8_71[0],stage8_70[0],stage8_69[0],stage8_68[1]}
   );
   gpc606_5 gpc10023 (
      {stage7_69[1], stage7_69[2], stage7_69[3], stage7_69[4], 1'b0, 1'b0},
      {stage7_71[0], stage7_71[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage8_72[1],stage8_71[1],stage8_70[1],stage8_69[1]}
   );
   gpc1_1 gpc10024 (
      {stage7_1[1]},
      {stage8_1[1]}
   );
   gpc1_1 gpc10025 (
      {stage7_2[4]},
      {stage8_2[1]}
   );
   gpc1_1 gpc10026 (
      {stage7_3[1]},
      {stage8_3[1]}
   );
   gpc1_1 gpc10027 (
      {stage7_4[0]},
      {stage8_4[1]}
   );
   gpc1_1 gpc10028 (
      {stage7_5[0]},
      {stage8_5[0]}
   );
   gpc1_1 gpc10029 (
      {stage7_5[1]},
      {stage8_5[1]}
   );
   gpc1_1 gpc10030 (
      {stage7_12[1]},
      {stage8_12[1]}
   );
   gpc1_1 gpc10031 (
      {stage7_19[6]},
      {stage8_19[1]}
   );
   gpc1_1 gpc10032 (
      {stage7_25[1]},
      {stage8_25[1]}
   );
   gpc1_1 gpc10033 (
      {stage7_33[0]},
      {stage8_33[1]}
   );
   gpc1_1 gpc10034 (
      {stage7_37[1]},
      {stage8_37[1]}
   );
   gpc1_1 gpc10035 (
      {stage7_39[0]},
      {stage8_39[1]}
   );
   gpc1_1 gpc10036 (
      {stage7_44[1]},
      {stage8_44[1]}
   );
   gpc1_1 gpc10037 (
      {stage7_54[0]},
      {stage8_54[1]}
   );
   gpc1_1 gpc10038 (
      {stage7_67[0]},
      {stage8_67[1]}
   );
endmodule
module rowadder2_1_73(input [72:0] src0, input [72:0] src1, output [73:0] dst0);
    wire [72:0] gene;
    wire [72:0] prop;
    wire [75:0] out;
    wire [75:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_38_gene (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(gene[38])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_38_prop (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(prop[38])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_39_gene (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(gene[39])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_39_prop (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(prop[39])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_40_gene (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(gene[40])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_40_prop (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(prop[40])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_41_gene (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(gene[41])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_41_prop (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(prop[41])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_42_gene (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(gene[42])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_42_prop (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(prop[42])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_43_gene (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(gene[43])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_43_prop (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(prop[43])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_44_gene (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(gene[44])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_44_prop (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(prop[44])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_45_gene (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(gene[45])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_45_prop (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(prop[45])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_46_gene (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(gene[46])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_46_prop (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(prop[46])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_47_gene (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(gene[47])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_47_prop (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(prop[47])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_48_gene (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(gene[48])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_48_prop (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(prop[48])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_49_gene (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(gene[49])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_49_prop (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(prop[49])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_50_gene (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(gene[50])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_50_prop (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(prop[50])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_51_gene (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(gene[51])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_51_prop (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(prop[51])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_52_gene (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(gene[52])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_52_prop (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(prop[52])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_53_gene (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(gene[53])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_53_prop (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(prop[53])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_54_gene (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(gene[54])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_54_prop (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(prop[54])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_55_gene (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(gene[55])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_55_prop (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(prop[55])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_56_gene (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(gene[56])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_56_prop (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(prop[56])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_57_gene (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(gene[57])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_57_prop (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(prop[57])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_58_gene (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(gene[58])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_58_prop (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(prop[58])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_59_gene (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(gene[59])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_59_prop (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(prop[59])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_60_gene (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(gene[60])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_60_prop (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(prop[60])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_61_gene (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(gene[61])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_61_prop (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(prop[61])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_62_gene (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(gene[62])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_62_prop (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(prop[62])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_63_gene (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(gene[63])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_63_prop (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(prop[63])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_64_gene (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(gene[64])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_64_prop (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(prop[64])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_65_gene (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(gene[65])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_65_prop (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(prop[65])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_66_gene (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(gene[66])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_66_prop (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(prop[66])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_67_gene (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(gene[67])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_67_prop (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(prop[67])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_68_gene (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(gene[68])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_68_prop (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(prop[68])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_69_gene (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(gene[69])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_69_prop (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(prop[69])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_70_gene (
        .I0(src0[70]),
        .I1(src1[70]),
        .O(gene[70])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_70_prop (
        .I0(src0[70]),
        .I1(src1[70]),
        .O(prop[70])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_71_gene (
        .I0(src0[71]),
        .I1(src1[71]),
        .O(gene[71])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_71_prop (
        .I0(src0[71]),
        .I1(src1[71]),
        .O(prop[71])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_72_gene (
        .I0(src0[72]),
        .I1(src1[72]),
        .O(gene[72])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_72_prop (
        .I0(src0[72]),
        .I1(src1[72]),
        .O(prop[72])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI(gene[39:36]),
        .S(prop[39:36])
    );
    CARRY4 carry4_43_40 (
        .CO(carryout[43:40]),
        .O(out[43:40]),
        .CI(carryout[39]),
        .CYINIT(1'h0),
        .DI(gene[43:40]),
        .S(prop[43:40])
    );
    CARRY4 carry4_47_44 (
        .CO(carryout[47:44]),
        .O(out[47:44]),
        .CI(carryout[43]),
        .CYINIT(1'h0),
        .DI(gene[47:44]),
        .S(prop[47:44])
    );
    CARRY4 carry4_51_48 (
        .CO(carryout[51:48]),
        .O(out[51:48]),
        .CI(carryout[47]),
        .CYINIT(1'h0),
        .DI(gene[51:48]),
        .S(prop[51:48])
    );
    CARRY4 carry4_55_52 (
        .CO(carryout[55:52]),
        .O(out[55:52]),
        .CI(carryout[51]),
        .CYINIT(1'h0),
        .DI(gene[55:52]),
        .S(prop[55:52])
    );
    CARRY4 carry4_59_56 (
        .CO(carryout[59:56]),
        .O(out[59:56]),
        .CI(carryout[55]),
        .CYINIT(1'h0),
        .DI(gene[59:56]),
        .S(prop[59:56])
    );
    CARRY4 carry4_63_60 (
        .CO(carryout[63:60]),
        .O(out[63:60]),
        .CI(carryout[59]),
        .CYINIT(1'h0),
        .DI(gene[63:60]),
        .S(prop[63:60])
    );
    CARRY4 carry4_67_64 (
        .CO(carryout[67:64]),
        .O(out[67:64]),
        .CI(carryout[63]),
        .CYINIT(1'h0),
        .DI(gene[67:64]),
        .S(prop[67:64])
    );
    CARRY4 carry4_71_68 (
        .CO(carryout[71:68]),
        .O(out[71:68]),
        .CI(carryout[67]),
        .CYINIT(1'h0),
        .DI(gene[71:68]),
        .S(prop[71:68])
    );
    CARRY4 carry4_75_72 (
        .CO(carryout[75:72]),
        .O(out[75:72]),
        .CI(carryout[71]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[72:72]}),
        .S({3'h0, prop[72:72]})
    );
    assign dst0 = {carryout[72], out[72:0]};
endmodule


module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    reg [485:0] src32;
    reg [485:0] src33;
    reg [485:0] src34;
    reg [485:0] src35;
    reg [485:0] src36;
    reg [485:0] src37;
    reg [485:0] src38;
    reg [485:0] src39;
    reg [485:0] src40;
    reg [485:0] src41;
    reg [485:0] src42;
    reg [485:0] src43;
    reg [485:0] src44;
    reg [485:0] src45;
    reg [485:0] src46;
    reg [485:0] src47;
    reg [485:0] src48;
    reg [485:0] src49;
    reg [485:0] src50;
    reg [485:0] src51;
    reg [485:0] src52;
    reg [485:0] src53;
    reg [485:0] src54;
    reg [485:0] src55;
    reg [485:0] src56;
    reg [485:0] src57;
    reg [485:0] src58;
    reg [485:0] src59;
    reg [485:0] src60;
    reg [485:0] src61;
    reg [485:0] src62;
    reg [485:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [0:0] dst72;
    wire [72:0] srcsum;
    wire [72:0] dstsum;
    wire test;
    compressor2_1_486_64 compressor2_1_486_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71),
        .dst72(dst72));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161] + src32[162] + src32[163] + src32[164] + src32[165] + src32[166] + src32[167] + src32[168] + src32[169] + src32[170] + src32[171] + src32[172] + src32[173] + src32[174] + src32[175] + src32[176] + src32[177] + src32[178] + src32[179] + src32[180] + src32[181] + src32[182] + src32[183] + src32[184] + src32[185] + src32[186] + src32[187] + src32[188] + src32[189] + src32[190] + src32[191] + src32[192] + src32[193] + src32[194] + src32[195] + src32[196] + src32[197] + src32[198] + src32[199] + src32[200] + src32[201] + src32[202] + src32[203] + src32[204] + src32[205] + src32[206] + src32[207] + src32[208] + src32[209] + src32[210] + src32[211] + src32[212] + src32[213] + src32[214] + src32[215] + src32[216] + src32[217] + src32[218] + src32[219] + src32[220] + src32[221] + src32[222] + src32[223] + src32[224] + src32[225] + src32[226] + src32[227] + src32[228] + src32[229] + src32[230] + src32[231] + src32[232] + src32[233] + src32[234] + src32[235] + src32[236] + src32[237] + src32[238] + src32[239] + src32[240] + src32[241] + src32[242] + src32[243] + src32[244] + src32[245] + src32[246] + src32[247] + src32[248] + src32[249] + src32[250] + src32[251] + src32[252] + src32[253] + src32[254] + src32[255] + src32[256] + src32[257] + src32[258] + src32[259] + src32[260] + src32[261] + src32[262] + src32[263] + src32[264] + src32[265] + src32[266] + src32[267] + src32[268] + src32[269] + src32[270] + src32[271] + src32[272] + src32[273] + src32[274] + src32[275] + src32[276] + src32[277] + src32[278] + src32[279] + src32[280] + src32[281] + src32[282] + src32[283] + src32[284] + src32[285] + src32[286] + src32[287] + src32[288] + src32[289] + src32[290] + src32[291] + src32[292] + src32[293] + src32[294] + src32[295] + src32[296] + src32[297] + src32[298] + src32[299] + src32[300] + src32[301] + src32[302] + src32[303] + src32[304] + src32[305] + src32[306] + src32[307] + src32[308] + src32[309] + src32[310] + src32[311] + src32[312] + src32[313] + src32[314] + src32[315] + src32[316] + src32[317] + src32[318] + src32[319] + src32[320] + src32[321] + src32[322] + src32[323] + src32[324] + src32[325] + src32[326] + src32[327] + src32[328] + src32[329] + src32[330] + src32[331] + src32[332] + src32[333] + src32[334] + src32[335] + src32[336] + src32[337] + src32[338] + src32[339] + src32[340] + src32[341] + src32[342] + src32[343] + src32[344] + src32[345] + src32[346] + src32[347] + src32[348] + src32[349] + src32[350] + src32[351] + src32[352] + src32[353] + src32[354] + src32[355] + src32[356] + src32[357] + src32[358] + src32[359] + src32[360] + src32[361] + src32[362] + src32[363] + src32[364] + src32[365] + src32[366] + src32[367] + src32[368] + src32[369] + src32[370] + src32[371] + src32[372] + src32[373] + src32[374] + src32[375] + src32[376] + src32[377] + src32[378] + src32[379] + src32[380] + src32[381] + src32[382] + src32[383] + src32[384] + src32[385] + src32[386] + src32[387] + src32[388] + src32[389] + src32[390] + src32[391] + src32[392] + src32[393] + src32[394] + src32[395] + src32[396] + src32[397] + src32[398] + src32[399] + src32[400] + src32[401] + src32[402] + src32[403] + src32[404] + src32[405] + src32[406] + src32[407] + src32[408] + src32[409] + src32[410] + src32[411] + src32[412] + src32[413] + src32[414] + src32[415] + src32[416] + src32[417] + src32[418] + src32[419] + src32[420] + src32[421] + src32[422] + src32[423] + src32[424] + src32[425] + src32[426] + src32[427] + src32[428] + src32[429] + src32[430] + src32[431] + src32[432] + src32[433] + src32[434] + src32[435] + src32[436] + src32[437] + src32[438] + src32[439] + src32[440] + src32[441] + src32[442] + src32[443] + src32[444] + src32[445] + src32[446] + src32[447] + src32[448] + src32[449] + src32[450] + src32[451] + src32[452] + src32[453] + src32[454] + src32[455] + src32[456] + src32[457] + src32[458] + src32[459] + src32[460] + src32[461] + src32[462] + src32[463] + src32[464] + src32[465] + src32[466] + src32[467] + src32[468] + src32[469] + src32[470] + src32[471] + src32[472] + src32[473] + src32[474] + src32[475] + src32[476] + src32[477] + src32[478] + src32[479] + src32[480] + src32[481] + src32[482] + src32[483] + src32[484] + src32[485])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161] + src33[162] + src33[163] + src33[164] + src33[165] + src33[166] + src33[167] + src33[168] + src33[169] + src33[170] + src33[171] + src33[172] + src33[173] + src33[174] + src33[175] + src33[176] + src33[177] + src33[178] + src33[179] + src33[180] + src33[181] + src33[182] + src33[183] + src33[184] + src33[185] + src33[186] + src33[187] + src33[188] + src33[189] + src33[190] + src33[191] + src33[192] + src33[193] + src33[194] + src33[195] + src33[196] + src33[197] + src33[198] + src33[199] + src33[200] + src33[201] + src33[202] + src33[203] + src33[204] + src33[205] + src33[206] + src33[207] + src33[208] + src33[209] + src33[210] + src33[211] + src33[212] + src33[213] + src33[214] + src33[215] + src33[216] + src33[217] + src33[218] + src33[219] + src33[220] + src33[221] + src33[222] + src33[223] + src33[224] + src33[225] + src33[226] + src33[227] + src33[228] + src33[229] + src33[230] + src33[231] + src33[232] + src33[233] + src33[234] + src33[235] + src33[236] + src33[237] + src33[238] + src33[239] + src33[240] + src33[241] + src33[242] + src33[243] + src33[244] + src33[245] + src33[246] + src33[247] + src33[248] + src33[249] + src33[250] + src33[251] + src33[252] + src33[253] + src33[254] + src33[255] + src33[256] + src33[257] + src33[258] + src33[259] + src33[260] + src33[261] + src33[262] + src33[263] + src33[264] + src33[265] + src33[266] + src33[267] + src33[268] + src33[269] + src33[270] + src33[271] + src33[272] + src33[273] + src33[274] + src33[275] + src33[276] + src33[277] + src33[278] + src33[279] + src33[280] + src33[281] + src33[282] + src33[283] + src33[284] + src33[285] + src33[286] + src33[287] + src33[288] + src33[289] + src33[290] + src33[291] + src33[292] + src33[293] + src33[294] + src33[295] + src33[296] + src33[297] + src33[298] + src33[299] + src33[300] + src33[301] + src33[302] + src33[303] + src33[304] + src33[305] + src33[306] + src33[307] + src33[308] + src33[309] + src33[310] + src33[311] + src33[312] + src33[313] + src33[314] + src33[315] + src33[316] + src33[317] + src33[318] + src33[319] + src33[320] + src33[321] + src33[322] + src33[323] + src33[324] + src33[325] + src33[326] + src33[327] + src33[328] + src33[329] + src33[330] + src33[331] + src33[332] + src33[333] + src33[334] + src33[335] + src33[336] + src33[337] + src33[338] + src33[339] + src33[340] + src33[341] + src33[342] + src33[343] + src33[344] + src33[345] + src33[346] + src33[347] + src33[348] + src33[349] + src33[350] + src33[351] + src33[352] + src33[353] + src33[354] + src33[355] + src33[356] + src33[357] + src33[358] + src33[359] + src33[360] + src33[361] + src33[362] + src33[363] + src33[364] + src33[365] + src33[366] + src33[367] + src33[368] + src33[369] + src33[370] + src33[371] + src33[372] + src33[373] + src33[374] + src33[375] + src33[376] + src33[377] + src33[378] + src33[379] + src33[380] + src33[381] + src33[382] + src33[383] + src33[384] + src33[385] + src33[386] + src33[387] + src33[388] + src33[389] + src33[390] + src33[391] + src33[392] + src33[393] + src33[394] + src33[395] + src33[396] + src33[397] + src33[398] + src33[399] + src33[400] + src33[401] + src33[402] + src33[403] + src33[404] + src33[405] + src33[406] + src33[407] + src33[408] + src33[409] + src33[410] + src33[411] + src33[412] + src33[413] + src33[414] + src33[415] + src33[416] + src33[417] + src33[418] + src33[419] + src33[420] + src33[421] + src33[422] + src33[423] + src33[424] + src33[425] + src33[426] + src33[427] + src33[428] + src33[429] + src33[430] + src33[431] + src33[432] + src33[433] + src33[434] + src33[435] + src33[436] + src33[437] + src33[438] + src33[439] + src33[440] + src33[441] + src33[442] + src33[443] + src33[444] + src33[445] + src33[446] + src33[447] + src33[448] + src33[449] + src33[450] + src33[451] + src33[452] + src33[453] + src33[454] + src33[455] + src33[456] + src33[457] + src33[458] + src33[459] + src33[460] + src33[461] + src33[462] + src33[463] + src33[464] + src33[465] + src33[466] + src33[467] + src33[468] + src33[469] + src33[470] + src33[471] + src33[472] + src33[473] + src33[474] + src33[475] + src33[476] + src33[477] + src33[478] + src33[479] + src33[480] + src33[481] + src33[482] + src33[483] + src33[484] + src33[485])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161] + src34[162] + src34[163] + src34[164] + src34[165] + src34[166] + src34[167] + src34[168] + src34[169] + src34[170] + src34[171] + src34[172] + src34[173] + src34[174] + src34[175] + src34[176] + src34[177] + src34[178] + src34[179] + src34[180] + src34[181] + src34[182] + src34[183] + src34[184] + src34[185] + src34[186] + src34[187] + src34[188] + src34[189] + src34[190] + src34[191] + src34[192] + src34[193] + src34[194] + src34[195] + src34[196] + src34[197] + src34[198] + src34[199] + src34[200] + src34[201] + src34[202] + src34[203] + src34[204] + src34[205] + src34[206] + src34[207] + src34[208] + src34[209] + src34[210] + src34[211] + src34[212] + src34[213] + src34[214] + src34[215] + src34[216] + src34[217] + src34[218] + src34[219] + src34[220] + src34[221] + src34[222] + src34[223] + src34[224] + src34[225] + src34[226] + src34[227] + src34[228] + src34[229] + src34[230] + src34[231] + src34[232] + src34[233] + src34[234] + src34[235] + src34[236] + src34[237] + src34[238] + src34[239] + src34[240] + src34[241] + src34[242] + src34[243] + src34[244] + src34[245] + src34[246] + src34[247] + src34[248] + src34[249] + src34[250] + src34[251] + src34[252] + src34[253] + src34[254] + src34[255] + src34[256] + src34[257] + src34[258] + src34[259] + src34[260] + src34[261] + src34[262] + src34[263] + src34[264] + src34[265] + src34[266] + src34[267] + src34[268] + src34[269] + src34[270] + src34[271] + src34[272] + src34[273] + src34[274] + src34[275] + src34[276] + src34[277] + src34[278] + src34[279] + src34[280] + src34[281] + src34[282] + src34[283] + src34[284] + src34[285] + src34[286] + src34[287] + src34[288] + src34[289] + src34[290] + src34[291] + src34[292] + src34[293] + src34[294] + src34[295] + src34[296] + src34[297] + src34[298] + src34[299] + src34[300] + src34[301] + src34[302] + src34[303] + src34[304] + src34[305] + src34[306] + src34[307] + src34[308] + src34[309] + src34[310] + src34[311] + src34[312] + src34[313] + src34[314] + src34[315] + src34[316] + src34[317] + src34[318] + src34[319] + src34[320] + src34[321] + src34[322] + src34[323] + src34[324] + src34[325] + src34[326] + src34[327] + src34[328] + src34[329] + src34[330] + src34[331] + src34[332] + src34[333] + src34[334] + src34[335] + src34[336] + src34[337] + src34[338] + src34[339] + src34[340] + src34[341] + src34[342] + src34[343] + src34[344] + src34[345] + src34[346] + src34[347] + src34[348] + src34[349] + src34[350] + src34[351] + src34[352] + src34[353] + src34[354] + src34[355] + src34[356] + src34[357] + src34[358] + src34[359] + src34[360] + src34[361] + src34[362] + src34[363] + src34[364] + src34[365] + src34[366] + src34[367] + src34[368] + src34[369] + src34[370] + src34[371] + src34[372] + src34[373] + src34[374] + src34[375] + src34[376] + src34[377] + src34[378] + src34[379] + src34[380] + src34[381] + src34[382] + src34[383] + src34[384] + src34[385] + src34[386] + src34[387] + src34[388] + src34[389] + src34[390] + src34[391] + src34[392] + src34[393] + src34[394] + src34[395] + src34[396] + src34[397] + src34[398] + src34[399] + src34[400] + src34[401] + src34[402] + src34[403] + src34[404] + src34[405] + src34[406] + src34[407] + src34[408] + src34[409] + src34[410] + src34[411] + src34[412] + src34[413] + src34[414] + src34[415] + src34[416] + src34[417] + src34[418] + src34[419] + src34[420] + src34[421] + src34[422] + src34[423] + src34[424] + src34[425] + src34[426] + src34[427] + src34[428] + src34[429] + src34[430] + src34[431] + src34[432] + src34[433] + src34[434] + src34[435] + src34[436] + src34[437] + src34[438] + src34[439] + src34[440] + src34[441] + src34[442] + src34[443] + src34[444] + src34[445] + src34[446] + src34[447] + src34[448] + src34[449] + src34[450] + src34[451] + src34[452] + src34[453] + src34[454] + src34[455] + src34[456] + src34[457] + src34[458] + src34[459] + src34[460] + src34[461] + src34[462] + src34[463] + src34[464] + src34[465] + src34[466] + src34[467] + src34[468] + src34[469] + src34[470] + src34[471] + src34[472] + src34[473] + src34[474] + src34[475] + src34[476] + src34[477] + src34[478] + src34[479] + src34[480] + src34[481] + src34[482] + src34[483] + src34[484] + src34[485])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161] + src35[162] + src35[163] + src35[164] + src35[165] + src35[166] + src35[167] + src35[168] + src35[169] + src35[170] + src35[171] + src35[172] + src35[173] + src35[174] + src35[175] + src35[176] + src35[177] + src35[178] + src35[179] + src35[180] + src35[181] + src35[182] + src35[183] + src35[184] + src35[185] + src35[186] + src35[187] + src35[188] + src35[189] + src35[190] + src35[191] + src35[192] + src35[193] + src35[194] + src35[195] + src35[196] + src35[197] + src35[198] + src35[199] + src35[200] + src35[201] + src35[202] + src35[203] + src35[204] + src35[205] + src35[206] + src35[207] + src35[208] + src35[209] + src35[210] + src35[211] + src35[212] + src35[213] + src35[214] + src35[215] + src35[216] + src35[217] + src35[218] + src35[219] + src35[220] + src35[221] + src35[222] + src35[223] + src35[224] + src35[225] + src35[226] + src35[227] + src35[228] + src35[229] + src35[230] + src35[231] + src35[232] + src35[233] + src35[234] + src35[235] + src35[236] + src35[237] + src35[238] + src35[239] + src35[240] + src35[241] + src35[242] + src35[243] + src35[244] + src35[245] + src35[246] + src35[247] + src35[248] + src35[249] + src35[250] + src35[251] + src35[252] + src35[253] + src35[254] + src35[255] + src35[256] + src35[257] + src35[258] + src35[259] + src35[260] + src35[261] + src35[262] + src35[263] + src35[264] + src35[265] + src35[266] + src35[267] + src35[268] + src35[269] + src35[270] + src35[271] + src35[272] + src35[273] + src35[274] + src35[275] + src35[276] + src35[277] + src35[278] + src35[279] + src35[280] + src35[281] + src35[282] + src35[283] + src35[284] + src35[285] + src35[286] + src35[287] + src35[288] + src35[289] + src35[290] + src35[291] + src35[292] + src35[293] + src35[294] + src35[295] + src35[296] + src35[297] + src35[298] + src35[299] + src35[300] + src35[301] + src35[302] + src35[303] + src35[304] + src35[305] + src35[306] + src35[307] + src35[308] + src35[309] + src35[310] + src35[311] + src35[312] + src35[313] + src35[314] + src35[315] + src35[316] + src35[317] + src35[318] + src35[319] + src35[320] + src35[321] + src35[322] + src35[323] + src35[324] + src35[325] + src35[326] + src35[327] + src35[328] + src35[329] + src35[330] + src35[331] + src35[332] + src35[333] + src35[334] + src35[335] + src35[336] + src35[337] + src35[338] + src35[339] + src35[340] + src35[341] + src35[342] + src35[343] + src35[344] + src35[345] + src35[346] + src35[347] + src35[348] + src35[349] + src35[350] + src35[351] + src35[352] + src35[353] + src35[354] + src35[355] + src35[356] + src35[357] + src35[358] + src35[359] + src35[360] + src35[361] + src35[362] + src35[363] + src35[364] + src35[365] + src35[366] + src35[367] + src35[368] + src35[369] + src35[370] + src35[371] + src35[372] + src35[373] + src35[374] + src35[375] + src35[376] + src35[377] + src35[378] + src35[379] + src35[380] + src35[381] + src35[382] + src35[383] + src35[384] + src35[385] + src35[386] + src35[387] + src35[388] + src35[389] + src35[390] + src35[391] + src35[392] + src35[393] + src35[394] + src35[395] + src35[396] + src35[397] + src35[398] + src35[399] + src35[400] + src35[401] + src35[402] + src35[403] + src35[404] + src35[405] + src35[406] + src35[407] + src35[408] + src35[409] + src35[410] + src35[411] + src35[412] + src35[413] + src35[414] + src35[415] + src35[416] + src35[417] + src35[418] + src35[419] + src35[420] + src35[421] + src35[422] + src35[423] + src35[424] + src35[425] + src35[426] + src35[427] + src35[428] + src35[429] + src35[430] + src35[431] + src35[432] + src35[433] + src35[434] + src35[435] + src35[436] + src35[437] + src35[438] + src35[439] + src35[440] + src35[441] + src35[442] + src35[443] + src35[444] + src35[445] + src35[446] + src35[447] + src35[448] + src35[449] + src35[450] + src35[451] + src35[452] + src35[453] + src35[454] + src35[455] + src35[456] + src35[457] + src35[458] + src35[459] + src35[460] + src35[461] + src35[462] + src35[463] + src35[464] + src35[465] + src35[466] + src35[467] + src35[468] + src35[469] + src35[470] + src35[471] + src35[472] + src35[473] + src35[474] + src35[475] + src35[476] + src35[477] + src35[478] + src35[479] + src35[480] + src35[481] + src35[482] + src35[483] + src35[484] + src35[485])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161] + src36[162] + src36[163] + src36[164] + src36[165] + src36[166] + src36[167] + src36[168] + src36[169] + src36[170] + src36[171] + src36[172] + src36[173] + src36[174] + src36[175] + src36[176] + src36[177] + src36[178] + src36[179] + src36[180] + src36[181] + src36[182] + src36[183] + src36[184] + src36[185] + src36[186] + src36[187] + src36[188] + src36[189] + src36[190] + src36[191] + src36[192] + src36[193] + src36[194] + src36[195] + src36[196] + src36[197] + src36[198] + src36[199] + src36[200] + src36[201] + src36[202] + src36[203] + src36[204] + src36[205] + src36[206] + src36[207] + src36[208] + src36[209] + src36[210] + src36[211] + src36[212] + src36[213] + src36[214] + src36[215] + src36[216] + src36[217] + src36[218] + src36[219] + src36[220] + src36[221] + src36[222] + src36[223] + src36[224] + src36[225] + src36[226] + src36[227] + src36[228] + src36[229] + src36[230] + src36[231] + src36[232] + src36[233] + src36[234] + src36[235] + src36[236] + src36[237] + src36[238] + src36[239] + src36[240] + src36[241] + src36[242] + src36[243] + src36[244] + src36[245] + src36[246] + src36[247] + src36[248] + src36[249] + src36[250] + src36[251] + src36[252] + src36[253] + src36[254] + src36[255] + src36[256] + src36[257] + src36[258] + src36[259] + src36[260] + src36[261] + src36[262] + src36[263] + src36[264] + src36[265] + src36[266] + src36[267] + src36[268] + src36[269] + src36[270] + src36[271] + src36[272] + src36[273] + src36[274] + src36[275] + src36[276] + src36[277] + src36[278] + src36[279] + src36[280] + src36[281] + src36[282] + src36[283] + src36[284] + src36[285] + src36[286] + src36[287] + src36[288] + src36[289] + src36[290] + src36[291] + src36[292] + src36[293] + src36[294] + src36[295] + src36[296] + src36[297] + src36[298] + src36[299] + src36[300] + src36[301] + src36[302] + src36[303] + src36[304] + src36[305] + src36[306] + src36[307] + src36[308] + src36[309] + src36[310] + src36[311] + src36[312] + src36[313] + src36[314] + src36[315] + src36[316] + src36[317] + src36[318] + src36[319] + src36[320] + src36[321] + src36[322] + src36[323] + src36[324] + src36[325] + src36[326] + src36[327] + src36[328] + src36[329] + src36[330] + src36[331] + src36[332] + src36[333] + src36[334] + src36[335] + src36[336] + src36[337] + src36[338] + src36[339] + src36[340] + src36[341] + src36[342] + src36[343] + src36[344] + src36[345] + src36[346] + src36[347] + src36[348] + src36[349] + src36[350] + src36[351] + src36[352] + src36[353] + src36[354] + src36[355] + src36[356] + src36[357] + src36[358] + src36[359] + src36[360] + src36[361] + src36[362] + src36[363] + src36[364] + src36[365] + src36[366] + src36[367] + src36[368] + src36[369] + src36[370] + src36[371] + src36[372] + src36[373] + src36[374] + src36[375] + src36[376] + src36[377] + src36[378] + src36[379] + src36[380] + src36[381] + src36[382] + src36[383] + src36[384] + src36[385] + src36[386] + src36[387] + src36[388] + src36[389] + src36[390] + src36[391] + src36[392] + src36[393] + src36[394] + src36[395] + src36[396] + src36[397] + src36[398] + src36[399] + src36[400] + src36[401] + src36[402] + src36[403] + src36[404] + src36[405] + src36[406] + src36[407] + src36[408] + src36[409] + src36[410] + src36[411] + src36[412] + src36[413] + src36[414] + src36[415] + src36[416] + src36[417] + src36[418] + src36[419] + src36[420] + src36[421] + src36[422] + src36[423] + src36[424] + src36[425] + src36[426] + src36[427] + src36[428] + src36[429] + src36[430] + src36[431] + src36[432] + src36[433] + src36[434] + src36[435] + src36[436] + src36[437] + src36[438] + src36[439] + src36[440] + src36[441] + src36[442] + src36[443] + src36[444] + src36[445] + src36[446] + src36[447] + src36[448] + src36[449] + src36[450] + src36[451] + src36[452] + src36[453] + src36[454] + src36[455] + src36[456] + src36[457] + src36[458] + src36[459] + src36[460] + src36[461] + src36[462] + src36[463] + src36[464] + src36[465] + src36[466] + src36[467] + src36[468] + src36[469] + src36[470] + src36[471] + src36[472] + src36[473] + src36[474] + src36[475] + src36[476] + src36[477] + src36[478] + src36[479] + src36[480] + src36[481] + src36[482] + src36[483] + src36[484] + src36[485])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161] + src37[162] + src37[163] + src37[164] + src37[165] + src37[166] + src37[167] + src37[168] + src37[169] + src37[170] + src37[171] + src37[172] + src37[173] + src37[174] + src37[175] + src37[176] + src37[177] + src37[178] + src37[179] + src37[180] + src37[181] + src37[182] + src37[183] + src37[184] + src37[185] + src37[186] + src37[187] + src37[188] + src37[189] + src37[190] + src37[191] + src37[192] + src37[193] + src37[194] + src37[195] + src37[196] + src37[197] + src37[198] + src37[199] + src37[200] + src37[201] + src37[202] + src37[203] + src37[204] + src37[205] + src37[206] + src37[207] + src37[208] + src37[209] + src37[210] + src37[211] + src37[212] + src37[213] + src37[214] + src37[215] + src37[216] + src37[217] + src37[218] + src37[219] + src37[220] + src37[221] + src37[222] + src37[223] + src37[224] + src37[225] + src37[226] + src37[227] + src37[228] + src37[229] + src37[230] + src37[231] + src37[232] + src37[233] + src37[234] + src37[235] + src37[236] + src37[237] + src37[238] + src37[239] + src37[240] + src37[241] + src37[242] + src37[243] + src37[244] + src37[245] + src37[246] + src37[247] + src37[248] + src37[249] + src37[250] + src37[251] + src37[252] + src37[253] + src37[254] + src37[255] + src37[256] + src37[257] + src37[258] + src37[259] + src37[260] + src37[261] + src37[262] + src37[263] + src37[264] + src37[265] + src37[266] + src37[267] + src37[268] + src37[269] + src37[270] + src37[271] + src37[272] + src37[273] + src37[274] + src37[275] + src37[276] + src37[277] + src37[278] + src37[279] + src37[280] + src37[281] + src37[282] + src37[283] + src37[284] + src37[285] + src37[286] + src37[287] + src37[288] + src37[289] + src37[290] + src37[291] + src37[292] + src37[293] + src37[294] + src37[295] + src37[296] + src37[297] + src37[298] + src37[299] + src37[300] + src37[301] + src37[302] + src37[303] + src37[304] + src37[305] + src37[306] + src37[307] + src37[308] + src37[309] + src37[310] + src37[311] + src37[312] + src37[313] + src37[314] + src37[315] + src37[316] + src37[317] + src37[318] + src37[319] + src37[320] + src37[321] + src37[322] + src37[323] + src37[324] + src37[325] + src37[326] + src37[327] + src37[328] + src37[329] + src37[330] + src37[331] + src37[332] + src37[333] + src37[334] + src37[335] + src37[336] + src37[337] + src37[338] + src37[339] + src37[340] + src37[341] + src37[342] + src37[343] + src37[344] + src37[345] + src37[346] + src37[347] + src37[348] + src37[349] + src37[350] + src37[351] + src37[352] + src37[353] + src37[354] + src37[355] + src37[356] + src37[357] + src37[358] + src37[359] + src37[360] + src37[361] + src37[362] + src37[363] + src37[364] + src37[365] + src37[366] + src37[367] + src37[368] + src37[369] + src37[370] + src37[371] + src37[372] + src37[373] + src37[374] + src37[375] + src37[376] + src37[377] + src37[378] + src37[379] + src37[380] + src37[381] + src37[382] + src37[383] + src37[384] + src37[385] + src37[386] + src37[387] + src37[388] + src37[389] + src37[390] + src37[391] + src37[392] + src37[393] + src37[394] + src37[395] + src37[396] + src37[397] + src37[398] + src37[399] + src37[400] + src37[401] + src37[402] + src37[403] + src37[404] + src37[405] + src37[406] + src37[407] + src37[408] + src37[409] + src37[410] + src37[411] + src37[412] + src37[413] + src37[414] + src37[415] + src37[416] + src37[417] + src37[418] + src37[419] + src37[420] + src37[421] + src37[422] + src37[423] + src37[424] + src37[425] + src37[426] + src37[427] + src37[428] + src37[429] + src37[430] + src37[431] + src37[432] + src37[433] + src37[434] + src37[435] + src37[436] + src37[437] + src37[438] + src37[439] + src37[440] + src37[441] + src37[442] + src37[443] + src37[444] + src37[445] + src37[446] + src37[447] + src37[448] + src37[449] + src37[450] + src37[451] + src37[452] + src37[453] + src37[454] + src37[455] + src37[456] + src37[457] + src37[458] + src37[459] + src37[460] + src37[461] + src37[462] + src37[463] + src37[464] + src37[465] + src37[466] + src37[467] + src37[468] + src37[469] + src37[470] + src37[471] + src37[472] + src37[473] + src37[474] + src37[475] + src37[476] + src37[477] + src37[478] + src37[479] + src37[480] + src37[481] + src37[482] + src37[483] + src37[484] + src37[485])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161] + src38[162] + src38[163] + src38[164] + src38[165] + src38[166] + src38[167] + src38[168] + src38[169] + src38[170] + src38[171] + src38[172] + src38[173] + src38[174] + src38[175] + src38[176] + src38[177] + src38[178] + src38[179] + src38[180] + src38[181] + src38[182] + src38[183] + src38[184] + src38[185] + src38[186] + src38[187] + src38[188] + src38[189] + src38[190] + src38[191] + src38[192] + src38[193] + src38[194] + src38[195] + src38[196] + src38[197] + src38[198] + src38[199] + src38[200] + src38[201] + src38[202] + src38[203] + src38[204] + src38[205] + src38[206] + src38[207] + src38[208] + src38[209] + src38[210] + src38[211] + src38[212] + src38[213] + src38[214] + src38[215] + src38[216] + src38[217] + src38[218] + src38[219] + src38[220] + src38[221] + src38[222] + src38[223] + src38[224] + src38[225] + src38[226] + src38[227] + src38[228] + src38[229] + src38[230] + src38[231] + src38[232] + src38[233] + src38[234] + src38[235] + src38[236] + src38[237] + src38[238] + src38[239] + src38[240] + src38[241] + src38[242] + src38[243] + src38[244] + src38[245] + src38[246] + src38[247] + src38[248] + src38[249] + src38[250] + src38[251] + src38[252] + src38[253] + src38[254] + src38[255] + src38[256] + src38[257] + src38[258] + src38[259] + src38[260] + src38[261] + src38[262] + src38[263] + src38[264] + src38[265] + src38[266] + src38[267] + src38[268] + src38[269] + src38[270] + src38[271] + src38[272] + src38[273] + src38[274] + src38[275] + src38[276] + src38[277] + src38[278] + src38[279] + src38[280] + src38[281] + src38[282] + src38[283] + src38[284] + src38[285] + src38[286] + src38[287] + src38[288] + src38[289] + src38[290] + src38[291] + src38[292] + src38[293] + src38[294] + src38[295] + src38[296] + src38[297] + src38[298] + src38[299] + src38[300] + src38[301] + src38[302] + src38[303] + src38[304] + src38[305] + src38[306] + src38[307] + src38[308] + src38[309] + src38[310] + src38[311] + src38[312] + src38[313] + src38[314] + src38[315] + src38[316] + src38[317] + src38[318] + src38[319] + src38[320] + src38[321] + src38[322] + src38[323] + src38[324] + src38[325] + src38[326] + src38[327] + src38[328] + src38[329] + src38[330] + src38[331] + src38[332] + src38[333] + src38[334] + src38[335] + src38[336] + src38[337] + src38[338] + src38[339] + src38[340] + src38[341] + src38[342] + src38[343] + src38[344] + src38[345] + src38[346] + src38[347] + src38[348] + src38[349] + src38[350] + src38[351] + src38[352] + src38[353] + src38[354] + src38[355] + src38[356] + src38[357] + src38[358] + src38[359] + src38[360] + src38[361] + src38[362] + src38[363] + src38[364] + src38[365] + src38[366] + src38[367] + src38[368] + src38[369] + src38[370] + src38[371] + src38[372] + src38[373] + src38[374] + src38[375] + src38[376] + src38[377] + src38[378] + src38[379] + src38[380] + src38[381] + src38[382] + src38[383] + src38[384] + src38[385] + src38[386] + src38[387] + src38[388] + src38[389] + src38[390] + src38[391] + src38[392] + src38[393] + src38[394] + src38[395] + src38[396] + src38[397] + src38[398] + src38[399] + src38[400] + src38[401] + src38[402] + src38[403] + src38[404] + src38[405] + src38[406] + src38[407] + src38[408] + src38[409] + src38[410] + src38[411] + src38[412] + src38[413] + src38[414] + src38[415] + src38[416] + src38[417] + src38[418] + src38[419] + src38[420] + src38[421] + src38[422] + src38[423] + src38[424] + src38[425] + src38[426] + src38[427] + src38[428] + src38[429] + src38[430] + src38[431] + src38[432] + src38[433] + src38[434] + src38[435] + src38[436] + src38[437] + src38[438] + src38[439] + src38[440] + src38[441] + src38[442] + src38[443] + src38[444] + src38[445] + src38[446] + src38[447] + src38[448] + src38[449] + src38[450] + src38[451] + src38[452] + src38[453] + src38[454] + src38[455] + src38[456] + src38[457] + src38[458] + src38[459] + src38[460] + src38[461] + src38[462] + src38[463] + src38[464] + src38[465] + src38[466] + src38[467] + src38[468] + src38[469] + src38[470] + src38[471] + src38[472] + src38[473] + src38[474] + src38[475] + src38[476] + src38[477] + src38[478] + src38[479] + src38[480] + src38[481] + src38[482] + src38[483] + src38[484] + src38[485])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161] + src39[162] + src39[163] + src39[164] + src39[165] + src39[166] + src39[167] + src39[168] + src39[169] + src39[170] + src39[171] + src39[172] + src39[173] + src39[174] + src39[175] + src39[176] + src39[177] + src39[178] + src39[179] + src39[180] + src39[181] + src39[182] + src39[183] + src39[184] + src39[185] + src39[186] + src39[187] + src39[188] + src39[189] + src39[190] + src39[191] + src39[192] + src39[193] + src39[194] + src39[195] + src39[196] + src39[197] + src39[198] + src39[199] + src39[200] + src39[201] + src39[202] + src39[203] + src39[204] + src39[205] + src39[206] + src39[207] + src39[208] + src39[209] + src39[210] + src39[211] + src39[212] + src39[213] + src39[214] + src39[215] + src39[216] + src39[217] + src39[218] + src39[219] + src39[220] + src39[221] + src39[222] + src39[223] + src39[224] + src39[225] + src39[226] + src39[227] + src39[228] + src39[229] + src39[230] + src39[231] + src39[232] + src39[233] + src39[234] + src39[235] + src39[236] + src39[237] + src39[238] + src39[239] + src39[240] + src39[241] + src39[242] + src39[243] + src39[244] + src39[245] + src39[246] + src39[247] + src39[248] + src39[249] + src39[250] + src39[251] + src39[252] + src39[253] + src39[254] + src39[255] + src39[256] + src39[257] + src39[258] + src39[259] + src39[260] + src39[261] + src39[262] + src39[263] + src39[264] + src39[265] + src39[266] + src39[267] + src39[268] + src39[269] + src39[270] + src39[271] + src39[272] + src39[273] + src39[274] + src39[275] + src39[276] + src39[277] + src39[278] + src39[279] + src39[280] + src39[281] + src39[282] + src39[283] + src39[284] + src39[285] + src39[286] + src39[287] + src39[288] + src39[289] + src39[290] + src39[291] + src39[292] + src39[293] + src39[294] + src39[295] + src39[296] + src39[297] + src39[298] + src39[299] + src39[300] + src39[301] + src39[302] + src39[303] + src39[304] + src39[305] + src39[306] + src39[307] + src39[308] + src39[309] + src39[310] + src39[311] + src39[312] + src39[313] + src39[314] + src39[315] + src39[316] + src39[317] + src39[318] + src39[319] + src39[320] + src39[321] + src39[322] + src39[323] + src39[324] + src39[325] + src39[326] + src39[327] + src39[328] + src39[329] + src39[330] + src39[331] + src39[332] + src39[333] + src39[334] + src39[335] + src39[336] + src39[337] + src39[338] + src39[339] + src39[340] + src39[341] + src39[342] + src39[343] + src39[344] + src39[345] + src39[346] + src39[347] + src39[348] + src39[349] + src39[350] + src39[351] + src39[352] + src39[353] + src39[354] + src39[355] + src39[356] + src39[357] + src39[358] + src39[359] + src39[360] + src39[361] + src39[362] + src39[363] + src39[364] + src39[365] + src39[366] + src39[367] + src39[368] + src39[369] + src39[370] + src39[371] + src39[372] + src39[373] + src39[374] + src39[375] + src39[376] + src39[377] + src39[378] + src39[379] + src39[380] + src39[381] + src39[382] + src39[383] + src39[384] + src39[385] + src39[386] + src39[387] + src39[388] + src39[389] + src39[390] + src39[391] + src39[392] + src39[393] + src39[394] + src39[395] + src39[396] + src39[397] + src39[398] + src39[399] + src39[400] + src39[401] + src39[402] + src39[403] + src39[404] + src39[405] + src39[406] + src39[407] + src39[408] + src39[409] + src39[410] + src39[411] + src39[412] + src39[413] + src39[414] + src39[415] + src39[416] + src39[417] + src39[418] + src39[419] + src39[420] + src39[421] + src39[422] + src39[423] + src39[424] + src39[425] + src39[426] + src39[427] + src39[428] + src39[429] + src39[430] + src39[431] + src39[432] + src39[433] + src39[434] + src39[435] + src39[436] + src39[437] + src39[438] + src39[439] + src39[440] + src39[441] + src39[442] + src39[443] + src39[444] + src39[445] + src39[446] + src39[447] + src39[448] + src39[449] + src39[450] + src39[451] + src39[452] + src39[453] + src39[454] + src39[455] + src39[456] + src39[457] + src39[458] + src39[459] + src39[460] + src39[461] + src39[462] + src39[463] + src39[464] + src39[465] + src39[466] + src39[467] + src39[468] + src39[469] + src39[470] + src39[471] + src39[472] + src39[473] + src39[474] + src39[475] + src39[476] + src39[477] + src39[478] + src39[479] + src39[480] + src39[481] + src39[482] + src39[483] + src39[484] + src39[485])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161] + src40[162] + src40[163] + src40[164] + src40[165] + src40[166] + src40[167] + src40[168] + src40[169] + src40[170] + src40[171] + src40[172] + src40[173] + src40[174] + src40[175] + src40[176] + src40[177] + src40[178] + src40[179] + src40[180] + src40[181] + src40[182] + src40[183] + src40[184] + src40[185] + src40[186] + src40[187] + src40[188] + src40[189] + src40[190] + src40[191] + src40[192] + src40[193] + src40[194] + src40[195] + src40[196] + src40[197] + src40[198] + src40[199] + src40[200] + src40[201] + src40[202] + src40[203] + src40[204] + src40[205] + src40[206] + src40[207] + src40[208] + src40[209] + src40[210] + src40[211] + src40[212] + src40[213] + src40[214] + src40[215] + src40[216] + src40[217] + src40[218] + src40[219] + src40[220] + src40[221] + src40[222] + src40[223] + src40[224] + src40[225] + src40[226] + src40[227] + src40[228] + src40[229] + src40[230] + src40[231] + src40[232] + src40[233] + src40[234] + src40[235] + src40[236] + src40[237] + src40[238] + src40[239] + src40[240] + src40[241] + src40[242] + src40[243] + src40[244] + src40[245] + src40[246] + src40[247] + src40[248] + src40[249] + src40[250] + src40[251] + src40[252] + src40[253] + src40[254] + src40[255] + src40[256] + src40[257] + src40[258] + src40[259] + src40[260] + src40[261] + src40[262] + src40[263] + src40[264] + src40[265] + src40[266] + src40[267] + src40[268] + src40[269] + src40[270] + src40[271] + src40[272] + src40[273] + src40[274] + src40[275] + src40[276] + src40[277] + src40[278] + src40[279] + src40[280] + src40[281] + src40[282] + src40[283] + src40[284] + src40[285] + src40[286] + src40[287] + src40[288] + src40[289] + src40[290] + src40[291] + src40[292] + src40[293] + src40[294] + src40[295] + src40[296] + src40[297] + src40[298] + src40[299] + src40[300] + src40[301] + src40[302] + src40[303] + src40[304] + src40[305] + src40[306] + src40[307] + src40[308] + src40[309] + src40[310] + src40[311] + src40[312] + src40[313] + src40[314] + src40[315] + src40[316] + src40[317] + src40[318] + src40[319] + src40[320] + src40[321] + src40[322] + src40[323] + src40[324] + src40[325] + src40[326] + src40[327] + src40[328] + src40[329] + src40[330] + src40[331] + src40[332] + src40[333] + src40[334] + src40[335] + src40[336] + src40[337] + src40[338] + src40[339] + src40[340] + src40[341] + src40[342] + src40[343] + src40[344] + src40[345] + src40[346] + src40[347] + src40[348] + src40[349] + src40[350] + src40[351] + src40[352] + src40[353] + src40[354] + src40[355] + src40[356] + src40[357] + src40[358] + src40[359] + src40[360] + src40[361] + src40[362] + src40[363] + src40[364] + src40[365] + src40[366] + src40[367] + src40[368] + src40[369] + src40[370] + src40[371] + src40[372] + src40[373] + src40[374] + src40[375] + src40[376] + src40[377] + src40[378] + src40[379] + src40[380] + src40[381] + src40[382] + src40[383] + src40[384] + src40[385] + src40[386] + src40[387] + src40[388] + src40[389] + src40[390] + src40[391] + src40[392] + src40[393] + src40[394] + src40[395] + src40[396] + src40[397] + src40[398] + src40[399] + src40[400] + src40[401] + src40[402] + src40[403] + src40[404] + src40[405] + src40[406] + src40[407] + src40[408] + src40[409] + src40[410] + src40[411] + src40[412] + src40[413] + src40[414] + src40[415] + src40[416] + src40[417] + src40[418] + src40[419] + src40[420] + src40[421] + src40[422] + src40[423] + src40[424] + src40[425] + src40[426] + src40[427] + src40[428] + src40[429] + src40[430] + src40[431] + src40[432] + src40[433] + src40[434] + src40[435] + src40[436] + src40[437] + src40[438] + src40[439] + src40[440] + src40[441] + src40[442] + src40[443] + src40[444] + src40[445] + src40[446] + src40[447] + src40[448] + src40[449] + src40[450] + src40[451] + src40[452] + src40[453] + src40[454] + src40[455] + src40[456] + src40[457] + src40[458] + src40[459] + src40[460] + src40[461] + src40[462] + src40[463] + src40[464] + src40[465] + src40[466] + src40[467] + src40[468] + src40[469] + src40[470] + src40[471] + src40[472] + src40[473] + src40[474] + src40[475] + src40[476] + src40[477] + src40[478] + src40[479] + src40[480] + src40[481] + src40[482] + src40[483] + src40[484] + src40[485])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161] + src41[162] + src41[163] + src41[164] + src41[165] + src41[166] + src41[167] + src41[168] + src41[169] + src41[170] + src41[171] + src41[172] + src41[173] + src41[174] + src41[175] + src41[176] + src41[177] + src41[178] + src41[179] + src41[180] + src41[181] + src41[182] + src41[183] + src41[184] + src41[185] + src41[186] + src41[187] + src41[188] + src41[189] + src41[190] + src41[191] + src41[192] + src41[193] + src41[194] + src41[195] + src41[196] + src41[197] + src41[198] + src41[199] + src41[200] + src41[201] + src41[202] + src41[203] + src41[204] + src41[205] + src41[206] + src41[207] + src41[208] + src41[209] + src41[210] + src41[211] + src41[212] + src41[213] + src41[214] + src41[215] + src41[216] + src41[217] + src41[218] + src41[219] + src41[220] + src41[221] + src41[222] + src41[223] + src41[224] + src41[225] + src41[226] + src41[227] + src41[228] + src41[229] + src41[230] + src41[231] + src41[232] + src41[233] + src41[234] + src41[235] + src41[236] + src41[237] + src41[238] + src41[239] + src41[240] + src41[241] + src41[242] + src41[243] + src41[244] + src41[245] + src41[246] + src41[247] + src41[248] + src41[249] + src41[250] + src41[251] + src41[252] + src41[253] + src41[254] + src41[255] + src41[256] + src41[257] + src41[258] + src41[259] + src41[260] + src41[261] + src41[262] + src41[263] + src41[264] + src41[265] + src41[266] + src41[267] + src41[268] + src41[269] + src41[270] + src41[271] + src41[272] + src41[273] + src41[274] + src41[275] + src41[276] + src41[277] + src41[278] + src41[279] + src41[280] + src41[281] + src41[282] + src41[283] + src41[284] + src41[285] + src41[286] + src41[287] + src41[288] + src41[289] + src41[290] + src41[291] + src41[292] + src41[293] + src41[294] + src41[295] + src41[296] + src41[297] + src41[298] + src41[299] + src41[300] + src41[301] + src41[302] + src41[303] + src41[304] + src41[305] + src41[306] + src41[307] + src41[308] + src41[309] + src41[310] + src41[311] + src41[312] + src41[313] + src41[314] + src41[315] + src41[316] + src41[317] + src41[318] + src41[319] + src41[320] + src41[321] + src41[322] + src41[323] + src41[324] + src41[325] + src41[326] + src41[327] + src41[328] + src41[329] + src41[330] + src41[331] + src41[332] + src41[333] + src41[334] + src41[335] + src41[336] + src41[337] + src41[338] + src41[339] + src41[340] + src41[341] + src41[342] + src41[343] + src41[344] + src41[345] + src41[346] + src41[347] + src41[348] + src41[349] + src41[350] + src41[351] + src41[352] + src41[353] + src41[354] + src41[355] + src41[356] + src41[357] + src41[358] + src41[359] + src41[360] + src41[361] + src41[362] + src41[363] + src41[364] + src41[365] + src41[366] + src41[367] + src41[368] + src41[369] + src41[370] + src41[371] + src41[372] + src41[373] + src41[374] + src41[375] + src41[376] + src41[377] + src41[378] + src41[379] + src41[380] + src41[381] + src41[382] + src41[383] + src41[384] + src41[385] + src41[386] + src41[387] + src41[388] + src41[389] + src41[390] + src41[391] + src41[392] + src41[393] + src41[394] + src41[395] + src41[396] + src41[397] + src41[398] + src41[399] + src41[400] + src41[401] + src41[402] + src41[403] + src41[404] + src41[405] + src41[406] + src41[407] + src41[408] + src41[409] + src41[410] + src41[411] + src41[412] + src41[413] + src41[414] + src41[415] + src41[416] + src41[417] + src41[418] + src41[419] + src41[420] + src41[421] + src41[422] + src41[423] + src41[424] + src41[425] + src41[426] + src41[427] + src41[428] + src41[429] + src41[430] + src41[431] + src41[432] + src41[433] + src41[434] + src41[435] + src41[436] + src41[437] + src41[438] + src41[439] + src41[440] + src41[441] + src41[442] + src41[443] + src41[444] + src41[445] + src41[446] + src41[447] + src41[448] + src41[449] + src41[450] + src41[451] + src41[452] + src41[453] + src41[454] + src41[455] + src41[456] + src41[457] + src41[458] + src41[459] + src41[460] + src41[461] + src41[462] + src41[463] + src41[464] + src41[465] + src41[466] + src41[467] + src41[468] + src41[469] + src41[470] + src41[471] + src41[472] + src41[473] + src41[474] + src41[475] + src41[476] + src41[477] + src41[478] + src41[479] + src41[480] + src41[481] + src41[482] + src41[483] + src41[484] + src41[485])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161] + src42[162] + src42[163] + src42[164] + src42[165] + src42[166] + src42[167] + src42[168] + src42[169] + src42[170] + src42[171] + src42[172] + src42[173] + src42[174] + src42[175] + src42[176] + src42[177] + src42[178] + src42[179] + src42[180] + src42[181] + src42[182] + src42[183] + src42[184] + src42[185] + src42[186] + src42[187] + src42[188] + src42[189] + src42[190] + src42[191] + src42[192] + src42[193] + src42[194] + src42[195] + src42[196] + src42[197] + src42[198] + src42[199] + src42[200] + src42[201] + src42[202] + src42[203] + src42[204] + src42[205] + src42[206] + src42[207] + src42[208] + src42[209] + src42[210] + src42[211] + src42[212] + src42[213] + src42[214] + src42[215] + src42[216] + src42[217] + src42[218] + src42[219] + src42[220] + src42[221] + src42[222] + src42[223] + src42[224] + src42[225] + src42[226] + src42[227] + src42[228] + src42[229] + src42[230] + src42[231] + src42[232] + src42[233] + src42[234] + src42[235] + src42[236] + src42[237] + src42[238] + src42[239] + src42[240] + src42[241] + src42[242] + src42[243] + src42[244] + src42[245] + src42[246] + src42[247] + src42[248] + src42[249] + src42[250] + src42[251] + src42[252] + src42[253] + src42[254] + src42[255] + src42[256] + src42[257] + src42[258] + src42[259] + src42[260] + src42[261] + src42[262] + src42[263] + src42[264] + src42[265] + src42[266] + src42[267] + src42[268] + src42[269] + src42[270] + src42[271] + src42[272] + src42[273] + src42[274] + src42[275] + src42[276] + src42[277] + src42[278] + src42[279] + src42[280] + src42[281] + src42[282] + src42[283] + src42[284] + src42[285] + src42[286] + src42[287] + src42[288] + src42[289] + src42[290] + src42[291] + src42[292] + src42[293] + src42[294] + src42[295] + src42[296] + src42[297] + src42[298] + src42[299] + src42[300] + src42[301] + src42[302] + src42[303] + src42[304] + src42[305] + src42[306] + src42[307] + src42[308] + src42[309] + src42[310] + src42[311] + src42[312] + src42[313] + src42[314] + src42[315] + src42[316] + src42[317] + src42[318] + src42[319] + src42[320] + src42[321] + src42[322] + src42[323] + src42[324] + src42[325] + src42[326] + src42[327] + src42[328] + src42[329] + src42[330] + src42[331] + src42[332] + src42[333] + src42[334] + src42[335] + src42[336] + src42[337] + src42[338] + src42[339] + src42[340] + src42[341] + src42[342] + src42[343] + src42[344] + src42[345] + src42[346] + src42[347] + src42[348] + src42[349] + src42[350] + src42[351] + src42[352] + src42[353] + src42[354] + src42[355] + src42[356] + src42[357] + src42[358] + src42[359] + src42[360] + src42[361] + src42[362] + src42[363] + src42[364] + src42[365] + src42[366] + src42[367] + src42[368] + src42[369] + src42[370] + src42[371] + src42[372] + src42[373] + src42[374] + src42[375] + src42[376] + src42[377] + src42[378] + src42[379] + src42[380] + src42[381] + src42[382] + src42[383] + src42[384] + src42[385] + src42[386] + src42[387] + src42[388] + src42[389] + src42[390] + src42[391] + src42[392] + src42[393] + src42[394] + src42[395] + src42[396] + src42[397] + src42[398] + src42[399] + src42[400] + src42[401] + src42[402] + src42[403] + src42[404] + src42[405] + src42[406] + src42[407] + src42[408] + src42[409] + src42[410] + src42[411] + src42[412] + src42[413] + src42[414] + src42[415] + src42[416] + src42[417] + src42[418] + src42[419] + src42[420] + src42[421] + src42[422] + src42[423] + src42[424] + src42[425] + src42[426] + src42[427] + src42[428] + src42[429] + src42[430] + src42[431] + src42[432] + src42[433] + src42[434] + src42[435] + src42[436] + src42[437] + src42[438] + src42[439] + src42[440] + src42[441] + src42[442] + src42[443] + src42[444] + src42[445] + src42[446] + src42[447] + src42[448] + src42[449] + src42[450] + src42[451] + src42[452] + src42[453] + src42[454] + src42[455] + src42[456] + src42[457] + src42[458] + src42[459] + src42[460] + src42[461] + src42[462] + src42[463] + src42[464] + src42[465] + src42[466] + src42[467] + src42[468] + src42[469] + src42[470] + src42[471] + src42[472] + src42[473] + src42[474] + src42[475] + src42[476] + src42[477] + src42[478] + src42[479] + src42[480] + src42[481] + src42[482] + src42[483] + src42[484] + src42[485])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161] + src43[162] + src43[163] + src43[164] + src43[165] + src43[166] + src43[167] + src43[168] + src43[169] + src43[170] + src43[171] + src43[172] + src43[173] + src43[174] + src43[175] + src43[176] + src43[177] + src43[178] + src43[179] + src43[180] + src43[181] + src43[182] + src43[183] + src43[184] + src43[185] + src43[186] + src43[187] + src43[188] + src43[189] + src43[190] + src43[191] + src43[192] + src43[193] + src43[194] + src43[195] + src43[196] + src43[197] + src43[198] + src43[199] + src43[200] + src43[201] + src43[202] + src43[203] + src43[204] + src43[205] + src43[206] + src43[207] + src43[208] + src43[209] + src43[210] + src43[211] + src43[212] + src43[213] + src43[214] + src43[215] + src43[216] + src43[217] + src43[218] + src43[219] + src43[220] + src43[221] + src43[222] + src43[223] + src43[224] + src43[225] + src43[226] + src43[227] + src43[228] + src43[229] + src43[230] + src43[231] + src43[232] + src43[233] + src43[234] + src43[235] + src43[236] + src43[237] + src43[238] + src43[239] + src43[240] + src43[241] + src43[242] + src43[243] + src43[244] + src43[245] + src43[246] + src43[247] + src43[248] + src43[249] + src43[250] + src43[251] + src43[252] + src43[253] + src43[254] + src43[255] + src43[256] + src43[257] + src43[258] + src43[259] + src43[260] + src43[261] + src43[262] + src43[263] + src43[264] + src43[265] + src43[266] + src43[267] + src43[268] + src43[269] + src43[270] + src43[271] + src43[272] + src43[273] + src43[274] + src43[275] + src43[276] + src43[277] + src43[278] + src43[279] + src43[280] + src43[281] + src43[282] + src43[283] + src43[284] + src43[285] + src43[286] + src43[287] + src43[288] + src43[289] + src43[290] + src43[291] + src43[292] + src43[293] + src43[294] + src43[295] + src43[296] + src43[297] + src43[298] + src43[299] + src43[300] + src43[301] + src43[302] + src43[303] + src43[304] + src43[305] + src43[306] + src43[307] + src43[308] + src43[309] + src43[310] + src43[311] + src43[312] + src43[313] + src43[314] + src43[315] + src43[316] + src43[317] + src43[318] + src43[319] + src43[320] + src43[321] + src43[322] + src43[323] + src43[324] + src43[325] + src43[326] + src43[327] + src43[328] + src43[329] + src43[330] + src43[331] + src43[332] + src43[333] + src43[334] + src43[335] + src43[336] + src43[337] + src43[338] + src43[339] + src43[340] + src43[341] + src43[342] + src43[343] + src43[344] + src43[345] + src43[346] + src43[347] + src43[348] + src43[349] + src43[350] + src43[351] + src43[352] + src43[353] + src43[354] + src43[355] + src43[356] + src43[357] + src43[358] + src43[359] + src43[360] + src43[361] + src43[362] + src43[363] + src43[364] + src43[365] + src43[366] + src43[367] + src43[368] + src43[369] + src43[370] + src43[371] + src43[372] + src43[373] + src43[374] + src43[375] + src43[376] + src43[377] + src43[378] + src43[379] + src43[380] + src43[381] + src43[382] + src43[383] + src43[384] + src43[385] + src43[386] + src43[387] + src43[388] + src43[389] + src43[390] + src43[391] + src43[392] + src43[393] + src43[394] + src43[395] + src43[396] + src43[397] + src43[398] + src43[399] + src43[400] + src43[401] + src43[402] + src43[403] + src43[404] + src43[405] + src43[406] + src43[407] + src43[408] + src43[409] + src43[410] + src43[411] + src43[412] + src43[413] + src43[414] + src43[415] + src43[416] + src43[417] + src43[418] + src43[419] + src43[420] + src43[421] + src43[422] + src43[423] + src43[424] + src43[425] + src43[426] + src43[427] + src43[428] + src43[429] + src43[430] + src43[431] + src43[432] + src43[433] + src43[434] + src43[435] + src43[436] + src43[437] + src43[438] + src43[439] + src43[440] + src43[441] + src43[442] + src43[443] + src43[444] + src43[445] + src43[446] + src43[447] + src43[448] + src43[449] + src43[450] + src43[451] + src43[452] + src43[453] + src43[454] + src43[455] + src43[456] + src43[457] + src43[458] + src43[459] + src43[460] + src43[461] + src43[462] + src43[463] + src43[464] + src43[465] + src43[466] + src43[467] + src43[468] + src43[469] + src43[470] + src43[471] + src43[472] + src43[473] + src43[474] + src43[475] + src43[476] + src43[477] + src43[478] + src43[479] + src43[480] + src43[481] + src43[482] + src43[483] + src43[484] + src43[485])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161] + src44[162] + src44[163] + src44[164] + src44[165] + src44[166] + src44[167] + src44[168] + src44[169] + src44[170] + src44[171] + src44[172] + src44[173] + src44[174] + src44[175] + src44[176] + src44[177] + src44[178] + src44[179] + src44[180] + src44[181] + src44[182] + src44[183] + src44[184] + src44[185] + src44[186] + src44[187] + src44[188] + src44[189] + src44[190] + src44[191] + src44[192] + src44[193] + src44[194] + src44[195] + src44[196] + src44[197] + src44[198] + src44[199] + src44[200] + src44[201] + src44[202] + src44[203] + src44[204] + src44[205] + src44[206] + src44[207] + src44[208] + src44[209] + src44[210] + src44[211] + src44[212] + src44[213] + src44[214] + src44[215] + src44[216] + src44[217] + src44[218] + src44[219] + src44[220] + src44[221] + src44[222] + src44[223] + src44[224] + src44[225] + src44[226] + src44[227] + src44[228] + src44[229] + src44[230] + src44[231] + src44[232] + src44[233] + src44[234] + src44[235] + src44[236] + src44[237] + src44[238] + src44[239] + src44[240] + src44[241] + src44[242] + src44[243] + src44[244] + src44[245] + src44[246] + src44[247] + src44[248] + src44[249] + src44[250] + src44[251] + src44[252] + src44[253] + src44[254] + src44[255] + src44[256] + src44[257] + src44[258] + src44[259] + src44[260] + src44[261] + src44[262] + src44[263] + src44[264] + src44[265] + src44[266] + src44[267] + src44[268] + src44[269] + src44[270] + src44[271] + src44[272] + src44[273] + src44[274] + src44[275] + src44[276] + src44[277] + src44[278] + src44[279] + src44[280] + src44[281] + src44[282] + src44[283] + src44[284] + src44[285] + src44[286] + src44[287] + src44[288] + src44[289] + src44[290] + src44[291] + src44[292] + src44[293] + src44[294] + src44[295] + src44[296] + src44[297] + src44[298] + src44[299] + src44[300] + src44[301] + src44[302] + src44[303] + src44[304] + src44[305] + src44[306] + src44[307] + src44[308] + src44[309] + src44[310] + src44[311] + src44[312] + src44[313] + src44[314] + src44[315] + src44[316] + src44[317] + src44[318] + src44[319] + src44[320] + src44[321] + src44[322] + src44[323] + src44[324] + src44[325] + src44[326] + src44[327] + src44[328] + src44[329] + src44[330] + src44[331] + src44[332] + src44[333] + src44[334] + src44[335] + src44[336] + src44[337] + src44[338] + src44[339] + src44[340] + src44[341] + src44[342] + src44[343] + src44[344] + src44[345] + src44[346] + src44[347] + src44[348] + src44[349] + src44[350] + src44[351] + src44[352] + src44[353] + src44[354] + src44[355] + src44[356] + src44[357] + src44[358] + src44[359] + src44[360] + src44[361] + src44[362] + src44[363] + src44[364] + src44[365] + src44[366] + src44[367] + src44[368] + src44[369] + src44[370] + src44[371] + src44[372] + src44[373] + src44[374] + src44[375] + src44[376] + src44[377] + src44[378] + src44[379] + src44[380] + src44[381] + src44[382] + src44[383] + src44[384] + src44[385] + src44[386] + src44[387] + src44[388] + src44[389] + src44[390] + src44[391] + src44[392] + src44[393] + src44[394] + src44[395] + src44[396] + src44[397] + src44[398] + src44[399] + src44[400] + src44[401] + src44[402] + src44[403] + src44[404] + src44[405] + src44[406] + src44[407] + src44[408] + src44[409] + src44[410] + src44[411] + src44[412] + src44[413] + src44[414] + src44[415] + src44[416] + src44[417] + src44[418] + src44[419] + src44[420] + src44[421] + src44[422] + src44[423] + src44[424] + src44[425] + src44[426] + src44[427] + src44[428] + src44[429] + src44[430] + src44[431] + src44[432] + src44[433] + src44[434] + src44[435] + src44[436] + src44[437] + src44[438] + src44[439] + src44[440] + src44[441] + src44[442] + src44[443] + src44[444] + src44[445] + src44[446] + src44[447] + src44[448] + src44[449] + src44[450] + src44[451] + src44[452] + src44[453] + src44[454] + src44[455] + src44[456] + src44[457] + src44[458] + src44[459] + src44[460] + src44[461] + src44[462] + src44[463] + src44[464] + src44[465] + src44[466] + src44[467] + src44[468] + src44[469] + src44[470] + src44[471] + src44[472] + src44[473] + src44[474] + src44[475] + src44[476] + src44[477] + src44[478] + src44[479] + src44[480] + src44[481] + src44[482] + src44[483] + src44[484] + src44[485])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161] + src45[162] + src45[163] + src45[164] + src45[165] + src45[166] + src45[167] + src45[168] + src45[169] + src45[170] + src45[171] + src45[172] + src45[173] + src45[174] + src45[175] + src45[176] + src45[177] + src45[178] + src45[179] + src45[180] + src45[181] + src45[182] + src45[183] + src45[184] + src45[185] + src45[186] + src45[187] + src45[188] + src45[189] + src45[190] + src45[191] + src45[192] + src45[193] + src45[194] + src45[195] + src45[196] + src45[197] + src45[198] + src45[199] + src45[200] + src45[201] + src45[202] + src45[203] + src45[204] + src45[205] + src45[206] + src45[207] + src45[208] + src45[209] + src45[210] + src45[211] + src45[212] + src45[213] + src45[214] + src45[215] + src45[216] + src45[217] + src45[218] + src45[219] + src45[220] + src45[221] + src45[222] + src45[223] + src45[224] + src45[225] + src45[226] + src45[227] + src45[228] + src45[229] + src45[230] + src45[231] + src45[232] + src45[233] + src45[234] + src45[235] + src45[236] + src45[237] + src45[238] + src45[239] + src45[240] + src45[241] + src45[242] + src45[243] + src45[244] + src45[245] + src45[246] + src45[247] + src45[248] + src45[249] + src45[250] + src45[251] + src45[252] + src45[253] + src45[254] + src45[255] + src45[256] + src45[257] + src45[258] + src45[259] + src45[260] + src45[261] + src45[262] + src45[263] + src45[264] + src45[265] + src45[266] + src45[267] + src45[268] + src45[269] + src45[270] + src45[271] + src45[272] + src45[273] + src45[274] + src45[275] + src45[276] + src45[277] + src45[278] + src45[279] + src45[280] + src45[281] + src45[282] + src45[283] + src45[284] + src45[285] + src45[286] + src45[287] + src45[288] + src45[289] + src45[290] + src45[291] + src45[292] + src45[293] + src45[294] + src45[295] + src45[296] + src45[297] + src45[298] + src45[299] + src45[300] + src45[301] + src45[302] + src45[303] + src45[304] + src45[305] + src45[306] + src45[307] + src45[308] + src45[309] + src45[310] + src45[311] + src45[312] + src45[313] + src45[314] + src45[315] + src45[316] + src45[317] + src45[318] + src45[319] + src45[320] + src45[321] + src45[322] + src45[323] + src45[324] + src45[325] + src45[326] + src45[327] + src45[328] + src45[329] + src45[330] + src45[331] + src45[332] + src45[333] + src45[334] + src45[335] + src45[336] + src45[337] + src45[338] + src45[339] + src45[340] + src45[341] + src45[342] + src45[343] + src45[344] + src45[345] + src45[346] + src45[347] + src45[348] + src45[349] + src45[350] + src45[351] + src45[352] + src45[353] + src45[354] + src45[355] + src45[356] + src45[357] + src45[358] + src45[359] + src45[360] + src45[361] + src45[362] + src45[363] + src45[364] + src45[365] + src45[366] + src45[367] + src45[368] + src45[369] + src45[370] + src45[371] + src45[372] + src45[373] + src45[374] + src45[375] + src45[376] + src45[377] + src45[378] + src45[379] + src45[380] + src45[381] + src45[382] + src45[383] + src45[384] + src45[385] + src45[386] + src45[387] + src45[388] + src45[389] + src45[390] + src45[391] + src45[392] + src45[393] + src45[394] + src45[395] + src45[396] + src45[397] + src45[398] + src45[399] + src45[400] + src45[401] + src45[402] + src45[403] + src45[404] + src45[405] + src45[406] + src45[407] + src45[408] + src45[409] + src45[410] + src45[411] + src45[412] + src45[413] + src45[414] + src45[415] + src45[416] + src45[417] + src45[418] + src45[419] + src45[420] + src45[421] + src45[422] + src45[423] + src45[424] + src45[425] + src45[426] + src45[427] + src45[428] + src45[429] + src45[430] + src45[431] + src45[432] + src45[433] + src45[434] + src45[435] + src45[436] + src45[437] + src45[438] + src45[439] + src45[440] + src45[441] + src45[442] + src45[443] + src45[444] + src45[445] + src45[446] + src45[447] + src45[448] + src45[449] + src45[450] + src45[451] + src45[452] + src45[453] + src45[454] + src45[455] + src45[456] + src45[457] + src45[458] + src45[459] + src45[460] + src45[461] + src45[462] + src45[463] + src45[464] + src45[465] + src45[466] + src45[467] + src45[468] + src45[469] + src45[470] + src45[471] + src45[472] + src45[473] + src45[474] + src45[475] + src45[476] + src45[477] + src45[478] + src45[479] + src45[480] + src45[481] + src45[482] + src45[483] + src45[484] + src45[485])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161] + src46[162] + src46[163] + src46[164] + src46[165] + src46[166] + src46[167] + src46[168] + src46[169] + src46[170] + src46[171] + src46[172] + src46[173] + src46[174] + src46[175] + src46[176] + src46[177] + src46[178] + src46[179] + src46[180] + src46[181] + src46[182] + src46[183] + src46[184] + src46[185] + src46[186] + src46[187] + src46[188] + src46[189] + src46[190] + src46[191] + src46[192] + src46[193] + src46[194] + src46[195] + src46[196] + src46[197] + src46[198] + src46[199] + src46[200] + src46[201] + src46[202] + src46[203] + src46[204] + src46[205] + src46[206] + src46[207] + src46[208] + src46[209] + src46[210] + src46[211] + src46[212] + src46[213] + src46[214] + src46[215] + src46[216] + src46[217] + src46[218] + src46[219] + src46[220] + src46[221] + src46[222] + src46[223] + src46[224] + src46[225] + src46[226] + src46[227] + src46[228] + src46[229] + src46[230] + src46[231] + src46[232] + src46[233] + src46[234] + src46[235] + src46[236] + src46[237] + src46[238] + src46[239] + src46[240] + src46[241] + src46[242] + src46[243] + src46[244] + src46[245] + src46[246] + src46[247] + src46[248] + src46[249] + src46[250] + src46[251] + src46[252] + src46[253] + src46[254] + src46[255] + src46[256] + src46[257] + src46[258] + src46[259] + src46[260] + src46[261] + src46[262] + src46[263] + src46[264] + src46[265] + src46[266] + src46[267] + src46[268] + src46[269] + src46[270] + src46[271] + src46[272] + src46[273] + src46[274] + src46[275] + src46[276] + src46[277] + src46[278] + src46[279] + src46[280] + src46[281] + src46[282] + src46[283] + src46[284] + src46[285] + src46[286] + src46[287] + src46[288] + src46[289] + src46[290] + src46[291] + src46[292] + src46[293] + src46[294] + src46[295] + src46[296] + src46[297] + src46[298] + src46[299] + src46[300] + src46[301] + src46[302] + src46[303] + src46[304] + src46[305] + src46[306] + src46[307] + src46[308] + src46[309] + src46[310] + src46[311] + src46[312] + src46[313] + src46[314] + src46[315] + src46[316] + src46[317] + src46[318] + src46[319] + src46[320] + src46[321] + src46[322] + src46[323] + src46[324] + src46[325] + src46[326] + src46[327] + src46[328] + src46[329] + src46[330] + src46[331] + src46[332] + src46[333] + src46[334] + src46[335] + src46[336] + src46[337] + src46[338] + src46[339] + src46[340] + src46[341] + src46[342] + src46[343] + src46[344] + src46[345] + src46[346] + src46[347] + src46[348] + src46[349] + src46[350] + src46[351] + src46[352] + src46[353] + src46[354] + src46[355] + src46[356] + src46[357] + src46[358] + src46[359] + src46[360] + src46[361] + src46[362] + src46[363] + src46[364] + src46[365] + src46[366] + src46[367] + src46[368] + src46[369] + src46[370] + src46[371] + src46[372] + src46[373] + src46[374] + src46[375] + src46[376] + src46[377] + src46[378] + src46[379] + src46[380] + src46[381] + src46[382] + src46[383] + src46[384] + src46[385] + src46[386] + src46[387] + src46[388] + src46[389] + src46[390] + src46[391] + src46[392] + src46[393] + src46[394] + src46[395] + src46[396] + src46[397] + src46[398] + src46[399] + src46[400] + src46[401] + src46[402] + src46[403] + src46[404] + src46[405] + src46[406] + src46[407] + src46[408] + src46[409] + src46[410] + src46[411] + src46[412] + src46[413] + src46[414] + src46[415] + src46[416] + src46[417] + src46[418] + src46[419] + src46[420] + src46[421] + src46[422] + src46[423] + src46[424] + src46[425] + src46[426] + src46[427] + src46[428] + src46[429] + src46[430] + src46[431] + src46[432] + src46[433] + src46[434] + src46[435] + src46[436] + src46[437] + src46[438] + src46[439] + src46[440] + src46[441] + src46[442] + src46[443] + src46[444] + src46[445] + src46[446] + src46[447] + src46[448] + src46[449] + src46[450] + src46[451] + src46[452] + src46[453] + src46[454] + src46[455] + src46[456] + src46[457] + src46[458] + src46[459] + src46[460] + src46[461] + src46[462] + src46[463] + src46[464] + src46[465] + src46[466] + src46[467] + src46[468] + src46[469] + src46[470] + src46[471] + src46[472] + src46[473] + src46[474] + src46[475] + src46[476] + src46[477] + src46[478] + src46[479] + src46[480] + src46[481] + src46[482] + src46[483] + src46[484] + src46[485])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161] + src47[162] + src47[163] + src47[164] + src47[165] + src47[166] + src47[167] + src47[168] + src47[169] + src47[170] + src47[171] + src47[172] + src47[173] + src47[174] + src47[175] + src47[176] + src47[177] + src47[178] + src47[179] + src47[180] + src47[181] + src47[182] + src47[183] + src47[184] + src47[185] + src47[186] + src47[187] + src47[188] + src47[189] + src47[190] + src47[191] + src47[192] + src47[193] + src47[194] + src47[195] + src47[196] + src47[197] + src47[198] + src47[199] + src47[200] + src47[201] + src47[202] + src47[203] + src47[204] + src47[205] + src47[206] + src47[207] + src47[208] + src47[209] + src47[210] + src47[211] + src47[212] + src47[213] + src47[214] + src47[215] + src47[216] + src47[217] + src47[218] + src47[219] + src47[220] + src47[221] + src47[222] + src47[223] + src47[224] + src47[225] + src47[226] + src47[227] + src47[228] + src47[229] + src47[230] + src47[231] + src47[232] + src47[233] + src47[234] + src47[235] + src47[236] + src47[237] + src47[238] + src47[239] + src47[240] + src47[241] + src47[242] + src47[243] + src47[244] + src47[245] + src47[246] + src47[247] + src47[248] + src47[249] + src47[250] + src47[251] + src47[252] + src47[253] + src47[254] + src47[255] + src47[256] + src47[257] + src47[258] + src47[259] + src47[260] + src47[261] + src47[262] + src47[263] + src47[264] + src47[265] + src47[266] + src47[267] + src47[268] + src47[269] + src47[270] + src47[271] + src47[272] + src47[273] + src47[274] + src47[275] + src47[276] + src47[277] + src47[278] + src47[279] + src47[280] + src47[281] + src47[282] + src47[283] + src47[284] + src47[285] + src47[286] + src47[287] + src47[288] + src47[289] + src47[290] + src47[291] + src47[292] + src47[293] + src47[294] + src47[295] + src47[296] + src47[297] + src47[298] + src47[299] + src47[300] + src47[301] + src47[302] + src47[303] + src47[304] + src47[305] + src47[306] + src47[307] + src47[308] + src47[309] + src47[310] + src47[311] + src47[312] + src47[313] + src47[314] + src47[315] + src47[316] + src47[317] + src47[318] + src47[319] + src47[320] + src47[321] + src47[322] + src47[323] + src47[324] + src47[325] + src47[326] + src47[327] + src47[328] + src47[329] + src47[330] + src47[331] + src47[332] + src47[333] + src47[334] + src47[335] + src47[336] + src47[337] + src47[338] + src47[339] + src47[340] + src47[341] + src47[342] + src47[343] + src47[344] + src47[345] + src47[346] + src47[347] + src47[348] + src47[349] + src47[350] + src47[351] + src47[352] + src47[353] + src47[354] + src47[355] + src47[356] + src47[357] + src47[358] + src47[359] + src47[360] + src47[361] + src47[362] + src47[363] + src47[364] + src47[365] + src47[366] + src47[367] + src47[368] + src47[369] + src47[370] + src47[371] + src47[372] + src47[373] + src47[374] + src47[375] + src47[376] + src47[377] + src47[378] + src47[379] + src47[380] + src47[381] + src47[382] + src47[383] + src47[384] + src47[385] + src47[386] + src47[387] + src47[388] + src47[389] + src47[390] + src47[391] + src47[392] + src47[393] + src47[394] + src47[395] + src47[396] + src47[397] + src47[398] + src47[399] + src47[400] + src47[401] + src47[402] + src47[403] + src47[404] + src47[405] + src47[406] + src47[407] + src47[408] + src47[409] + src47[410] + src47[411] + src47[412] + src47[413] + src47[414] + src47[415] + src47[416] + src47[417] + src47[418] + src47[419] + src47[420] + src47[421] + src47[422] + src47[423] + src47[424] + src47[425] + src47[426] + src47[427] + src47[428] + src47[429] + src47[430] + src47[431] + src47[432] + src47[433] + src47[434] + src47[435] + src47[436] + src47[437] + src47[438] + src47[439] + src47[440] + src47[441] + src47[442] + src47[443] + src47[444] + src47[445] + src47[446] + src47[447] + src47[448] + src47[449] + src47[450] + src47[451] + src47[452] + src47[453] + src47[454] + src47[455] + src47[456] + src47[457] + src47[458] + src47[459] + src47[460] + src47[461] + src47[462] + src47[463] + src47[464] + src47[465] + src47[466] + src47[467] + src47[468] + src47[469] + src47[470] + src47[471] + src47[472] + src47[473] + src47[474] + src47[475] + src47[476] + src47[477] + src47[478] + src47[479] + src47[480] + src47[481] + src47[482] + src47[483] + src47[484] + src47[485])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161] + src48[162] + src48[163] + src48[164] + src48[165] + src48[166] + src48[167] + src48[168] + src48[169] + src48[170] + src48[171] + src48[172] + src48[173] + src48[174] + src48[175] + src48[176] + src48[177] + src48[178] + src48[179] + src48[180] + src48[181] + src48[182] + src48[183] + src48[184] + src48[185] + src48[186] + src48[187] + src48[188] + src48[189] + src48[190] + src48[191] + src48[192] + src48[193] + src48[194] + src48[195] + src48[196] + src48[197] + src48[198] + src48[199] + src48[200] + src48[201] + src48[202] + src48[203] + src48[204] + src48[205] + src48[206] + src48[207] + src48[208] + src48[209] + src48[210] + src48[211] + src48[212] + src48[213] + src48[214] + src48[215] + src48[216] + src48[217] + src48[218] + src48[219] + src48[220] + src48[221] + src48[222] + src48[223] + src48[224] + src48[225] + src48[226] + src48[227] + src48[228] + src48[229] + src48[230] + src48[231] + src48[232] + src48[233] + src48[234] + src48[235] + src48[236] + src48[237] + src48[238] + src48[239] + src48[240] + src48[241] + src48[242] + src48[243] + src48[244] + src48[245] + src48[246] + src48[247] + src48[248] + src48[249] + src48[250] + src48[251] + src48[252] + src48[253] + src48[254] + src48[255] + src48[256] + src48[257] + src48[258] + src48[259] + src48[260] + src48[261] + src48[262] + src48[263] + src48[264] + src48[265] + src48[266] + src48[267] + src48[268] + src48[269] + src48[270] + src48[271] + src48[272] + src48[273] + src48[274] + src48[275] + src48[276] + src48[277] + src48[278] + src48[279] + src48[280] + src48[281] + src48[282] + src48[283] + src48[284] + src48[285] + src48[286] + src48[287] + src48[288] + src48[289] + src48[290] + src48[291] + src48[292] + src48[293] + src48[294] + src48[295] + src48[296] + src48[297] + src48[298] + src48[299] + src48[300] + src48[301] + src48[302] + src48[303] + src48[304] + src48[305] + src48[306] + src48[307] + src48[308] + src48[309] + src48[310] + src48[311] + src48[312] + src48[313] + src48[314] + src48[315] + src48[316] + src48[317] + src48[318] + src48[319] + src48[320] + src48[321] + src48[322] + src48[323] + src48[324] + src48[325] + src48[326] + src48[327] + src48[328] + src48[329] + src48[330] + src48[331] + src48[332] + src48[333] + src48[334] + src48[335] + src48[336] + src48[337] + src48[338] + src48[339] + src48[340] + src48[341] + src48[342] + src48[343] + src48[344] + src48[345] + src48[346] + src48[347] + src48[348] + src48[349] + src48[350] + src48[351] + src48[352] + src48[353] + src48[354] + src48[355] + src48[356] + src48[357] + src48[358] + src48[359] + src48[360] + src48[361] + src48[362] + src48[363] + src48[364] + src48[365] + src48[366] + src48[367] + src48[368] + src48[369] + src48[370] + src48[371] + src48[372] + src48[373] + src48[374] + src48[375] + src48[376] + src48[377] + src48[378] + src48[379] + src48[380] + src48[381] + src48[382] + src48[383] + src48[384] + src48[385] + src48[386] + src48[387] + src48[388] + src48[389] + src48[390] + src48[391] + src48[392] + src48[393] + src48[394] + src48[395] + src48[396] + src48[397] + src48[398] + src48[399] + src48[400] + src48[401] + src48[402] + src48[403] + src48[404] + src48[405] + src48[406] + src48[407] + src48[408] + src48[409] + src48[410] + src48[411] + src48[412] + src48[413] + src48[414] + src48[415] + src48[416] + src48[417] + src48[418] + src48[419] + src48[420] + src48[421] + src48[422] + src48[423] + src48[424] + src48[425] + src48[426] + src48[427] + src48[428] + src48[429] + src48[430] + src48[431] + src48[432] + src48[433] + src48[434] + src48[435] + src48[436] + src48[437] + src48[438] + src48[439] + src48[440] + src48[441] + src48[442] + src48[443] + src48[444] + src48[445] + src48[446] + src48[447] + src48[448] + src48[449] + src48[450] + src48[451] + src48[452] + src48[453] + src48[454] + src48[455] + src48[456] + src48[457] + src48[458] + src48[459] + src48[460] + src48[461] + src48[462] + src48[463] + src48[464] + src48[465] + src48[466] + src48[467] + src48[468] + src48[469] + src48[470] + src48[471] + src48[472] + src48[473] + src48[474] + src48[475] + src48[476] + src48[477] + src48[478] + src48[479] + src48[480] + src48[481] + src48[482] + src48[483] + src48[484] + src48[485])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161] + src49[162] + src49[163] + src49[164] + src49[165] + src49[166] + src49[167] + src49[168] + src49[169] + src49[170] + src49[171] + src49[172] + src49[173] + src49[174] + src49[175] + src49[176] + src49[177] + src49[178] + src49[179] + src49[180] + src49[181] + src49[182] + src49[183] + src49[184] + src49[185] + src49[186] + src49[187] + src49[188] + src49[189] + src49[190] + src49[191] + src49[192] + src49[193] + src49[194] + src49[195] + src49[196] + src49[197] + src49[198] + src49[199] + src49[200] + src49[201] + src49[202] + src49[203] + src49[204] + src49[205] + src49[206] + src49[207] + src49[208] + src49[209] + src49[210] + src49[211] + src49[212] + src49[213] + src49[214] + src49[215] + src49[216] + src49[217] + src49[218] + src49[219] + src49[220] + src49[221] + src49[222] + src49[223] + src49[224] + src49[225] + src49[226] + src49[227] + src49[228] + src49[229] + src49[230] + src49[231] + src49[232] + src49[233] + src49[234] + src49[235] + src49[236] + src49[237] + src49[238] + src49[239] + src49[240] + src49[241] + src49[242] + src49[243] + src49[244] + src49[245] + src49[246] + src49[247] + src49[248] + src49[249] + src49[250] + src49[251] + src49[252] + src49[253] + src49[254] + src49[255] + src49[256] + src49[257] + src49[258] + src49[259] + src49[260] + src49[261] + src49[262] + src49[263] + src49[264] + src49[265] + src49[266] + src49[267] + src49[268] + src49[269] + src49[270] + src49[271] + src49[272] + src49[273] + src49[274] + src49[275] + src49[276] + src49[277] + src49[278] + src49[279] + src49[280] + src49[281] + src49[282] + src49[283] + src49[284] + src49[285] + src49[286] + src49[287] + src49[288] + src49[289] + src49[290] + src49[291] + src49[292] + src49[293] + src49[294] + src49[295] + src49[296] + src49[297] + src49[298] + src49[299] + src49[300] + src49[301] + src49[302] + src49[303] + src49[304] + src49[305] + src49[306] + src49[307] + src49[308] + src49[309] + src49[310] + src49[311] + src49[312] + src49[313] + src49[314] + src49[315] + src49[316] + src49[317] + src49[318] + src49[319] + src49[320] + src49[321] + src49[322] + src49[323] + src49[324] + src49[325] + src49[326] + src49[327] + src49[328] + src49[329] + src49[330] + src49[331] + src49[332] + src49[333] + src49[334] + src49[335] + src49[336] + src49[337] + src49[338] + src49[339] + src49[340] + src49[341] + src49[342] + src49[343] + src49[344] + src49[345] + src49[346] + src49[347] + src49[348] + src49[349] + src49[350] + src49[351] + src49[352] + src49[353] + src49[354] + src49[355] + src49[356] + src49[357] + src49[358] + src49[359] + src49[360] + src49[361] + src49[362] + src49[363] + src49[364] + src49[365] + src49[366] + src49[367] + src49[368] + src49[369] + src49[370] + src49[371] + src49[372] + src49[373] + src49[374] + src49[375] + src49[376] + src49[377] + src49[378] + src49[379] + src49[380] + src49[381] + src49[382] + src49[383] + src49[384] + src49[385] + src49[386] + src49[387] + src49[388] + src49[389] + src49[390] + src49[391] + src49[392] + src49[393] + src49[394] + src49[395] + src49[396] + src49[397] + src49[398] + src49[399] + src49[400] + src49[401] + src49[402] + src49[403] + src49[404] + src49[405] + src49[406] + src49[407] + src49[408] + src49[409] + src49[410] + src49[411] + src49[412] + src49[413] + src49[414] + src49[415] + src49[416] + src49[417] + src49[418] + src49[419] + src49[420] + src49[421] + src49[422] + src49[423] + src49[424] + src49[425] + src49[426] + src49[427] + src49[428] + src49[429] + src49[430] + src49[431] + src49[432] + src49[433] + src49[434] + src49[435] + src49[436] + src49[437] + src49[438] + src49[439] + src49[440] + src49[441] + src49[442] + src49[443] + src49[444] + src49[445] + src49[446] + src49[447] + src49[448] + src49[449] + src49[450] + src49[451] + src49[452] + src49[453] + src49[454] + src49[455] + src49[456] + src49[457] + src49[458] + src49[459] + src49[460] + src49[461] + src49[462] + src49[463] + src49[464] + src49[465] + src49[466] + src49[467] + src49[468] + src49[469] + src49[470] + src49[471] + src49[472] + src49[473] + src49[474] + src49[475] + src49[476] + src49[477] + src49[478] + src49[479] + src49[480] + src49[481] + src49[482] + src49[483] + src49[484] + src49[485])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161] + src50[162] + src50[163] + src50[164] + src50[165] + src50[166] + src50[167] + src50[168] + src50[169] + src50[170] + src50[171] + src50[172] + src50[173] + src50[174] + src50[175] + src50[176] + src50[177] + src50[178] + src50[179] + src50[180] + src50[181] + src50[182] + src50[183] + src50[184] + src50[185] + src50[186] + src50[187] + src50[188] + src50[189] + src50[190] + src50[191] + src50[192] + src50[193] + src50[194] + src50[195] + src50[196] + src50[197] + src50[198] + src50[199] + src50[200] + src50[201] + src50[202] + src50[203] + src50[204] + src50[205] + src50[206] + src50[207] + src50[208] + src50[209] + src50[210] + src50[211] + src50[212] + src50[213] + src50[214] + src50[215] + src50[216] + src50[217] + src50[218] + src50[219] + src50[220] + src50[221] + src50[222] + src50[223] + src50[224] + src50[225] + src50[226] + src50[227] + src50[228] + src50[229] + src50[230] + src50[231] + src50[232] + src50[233] + src50[234] + src50[235] + src50[236] + src50[237] + src50[238] + src50[239] + src50[240] + src50[241] + src50[242] + src50[243] + src50[244] + src50[245] + src50[246] + src50[247] + src50[248] + src50[249] + src50[250] + src50[251] + src50[252] + src50[253] + src50[254] + src50[255] + src50[256] + src50[257] + src50[258] + src50[259] + src50[260] + src50[261] + src50[262] + src50[263] + src50[264] + src50[265] + src50[266] + src50[267] + src50[268] + src50[269] + src50[270] + src50[271] + src50[272] + src50[273] + src50[274] + src50[275] + src50[276] + src50[277] + src50[278] + src50[279] + src50[280] + src50[281] + src50[282] + src50[283] + src50[284] + src50[285] + src50[286] + src50[287] + src50[288] + src50[289] + src50[290] + src50[291] + src50[292] + src50[293] + src50[294] + src50[295] + src50[296] + src50[297] + src50[298] + src50[299] + src50[300] + src50[301] + src50[302] + src50[303] + src50[304] + src50[305] + src50[306] + src50[307] + src50[308] + src50[309] + src50[310] + src50[311] + src50[312] + src50[313] + src50[314] + src50[315] + src50[316] + src50[317] + src50[318] + src50[319] + src50[320] + src50[321] + src50[322] + src50[323] + src50[324] + src50[325] + src50[326] + src50[327] + src50[328] + src50[329] + src50[330] + src50[331] + src50[332] + src50[333] + src50[334] + src50[335] + src50[336] + src50[337] + src50[338] + src50[339] + src50[340] + src50[341] + src50[342] + src50[343] + src50[344] + src50[345] + src50[346] + src50[347] + src50[348] + src50[349] + src50[350] + src50[351] + src50[352] + src50[353] + src50[354] + src50[355] + src50[356] + src50[357] + src50[358] + src50[359] + src50[360] + src50[361] + src50[362] + src50[363] + src50[364] + src50[365] + src50[366] + src50[367] + src50[368] + src50[369] + src50[370] + src50[371] + src50[372] + src50[373] + src50[374] + src50[375] + src50[376] + src50[377] + src50[378] + src50[379] + src50[380] + src50[381] + src50[382] + src50[383] + src50[384] + src50[385] + src50[386] + src50[387] + src50[388] + src50[389] + src50[390] + src50[391] + src50[392] + src50[393] + src50[394] + src50[395] + src50[396] + src50[397] + src50[398] + src50[399] + src50[400] + src50[401] + src50[402] + src50[403] + src50[404] + src50[405] + src50[406] + src50[407] + src50[408] + src50[409] + src50[410] + src50[411] + src50[412] + src50[413] + src50[414] + src50[415] + src50[416] + src50[417] + src50[418] + src50[419] + src50[420] + src50[421] + src50[422] + src50[423] + src50[424] + src50[425] + src50[426] + src50[427] + src50[428] + src50[429] + src50[430] + src50[431] + src50[432] + src50[433] + src50[434] + src50[435] + src50[436] + src50[437] + src50[438] + src50[439] + src50[440] + src50[441] + src50[442] + src50[443] + src50[444] + src50[445] + src50[446] + src50[447] + src50[448] + src50[449] + src50[450] + src50[451] + src50[452] + src50[453] + src50[454] + src50[455] + src50[456] + src50[457] + src50[458] + src50[459] + src50[460] + src50[461] + src50[462] + src50[463] + src50[464] + src50[465] + src50[466] + src50[467] + src50[468] + src50[469] + src50[470] + src50[471] + src50[472] + src50[473] + src50[474] + src50[475] + src50[476] + src50[477] + src50[478] + src50[479] + src50[480] + src50[481] + src50[482] + src50[483] + src50[484] + src50[485])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161] + src51[162] + src51[163] + src51[164] + src51[165] + src51[166] + src51[167] + src51[168] + src51[169] + src51[170] + src51[171] + src51[172] + src51[173] + src51[174] + src51[175] + src51[176] + src51[177] + src51[178] + src51[179] + src51[180] + src51[181] + src51[182] + src51[183] + src51[184] + src51[185] + src51[186] + src51[187] + src51[188] + src51[189] + src51[190] + src51[191] + src51[192] + src51[193] + src51[194] + src51[195] + src51[196] + src51[197] + src51[198] + src51[199] + src51[200] + src51[201] + src51[202] + src51[203] + src51[204] + src51[205] + src51[206] + src51[207] + src51[208] + src51[209] + src51[210] + src51[211] + src51[212] + src51[213] + src51[214] + src51[215] + src51[216] + src51[217] + src51[218] + src51[219] + src51[220] + src51[221] + src51[222] + src51[223] + src51[224] + src51[225] + src51[226] + src51[227] + src51[228] + src51[229] + src51[230] + src51[231] + src51[232] + src51[233] + src51[234] + src51[235] + src51[236] + src51[237] + src51[238] + src51[239] + src51[240] + src51[241] + src51[242] + src51[243] + src51[244] + src51[245] + src51[246] + src51[247] + src51[248] + src51[249] + src51[250] + src51[251] + src51[252] + src51[253] + src51[254] + src51[255] + src51[256] + src51[257] + src51[258] + src51[259] + src51[260] + src51[261] + src51[262] + src51[263] + src51[264] + src51[265] + src51[266] + src51[267] + src51[268] + src51[269] + src51[270] + src51[271] + src51[272] + src51[273] + src51[274] + src51[275] + src51[276] + src51[277] + src51[278] + src51[279] + src51[280] + src51[281] + src51[282] + src51[283] + src51[284] + src51[285] + src51[286] + src51[287] + src51[288] + src51[289] + src51[290] + src51[291] + src51[292] + src51[293] + src51[294] + src51[295] + src51[296] + src51[297] + src51[298] + src51[299] + src51[300] + src51[301] + src51[302] + src51[303] + src51[304] + src51[305] + src51[306] + src51[307] + src51[308] + src51[309] + src51[310] + src51[311] + src51[312] + src51[313] + src51[314] + src51[315] + src51[316] + src51[317] + src51[318] + src51[319] + src51[320] + src51[321] + src51[322] + src51[323] + src51[324] + src51[325] + src51[326] + src51[327] + src51[328] + src51[329] + src51[330] + src51[331] + src51[332] + src51[333] + src51[334] + src51[335] + src51[336] + src51[337] + src51[338] + src51[339] + src51[340] + src51[341] + src51[342] + src51[343] + src51[344] + src51[345] + src51[346] + src51[347] + src51[348] + src51[349] + src51[350] + src51[351] + src51[352] + src51[353] + src51[354] + src51[355] + src51[356] + src51[357] + src51[358] + src51[359] + src51[360] + src51[361] + src51[362] + src51[363] + src51[364] + src51[365] + src51[366] + src51[367] + src51[368] + src51[369] + src51[370] + src51[371] + src51[372] + src51[373] + src51[374] + src51[375] + src51[376] + src51[377] + src51[378] + src51[379] + src51[380] + src51[381] + src51[382] + src51[383] + src51[384] + src51[385] + src51[386] + src51[387] + src51[388] + src51[389] + src51[390] + src51[391] + src51[392] + src51[393] + src51[394] + src51[395] + src51[396] + src51[397] + src51[398] + src51[399] + src51[400] + src51[401] + src51[402] + src51[403] + src51[404] + src51[405] + src51[406] + src51[407] + src51[408] + src51[409] + src51[410] + src51[411] + src51[412] + src51[413] + src51[414] + src51[415] + src51[416] + src51[417] + src51[418] + src51[419] + src51[420] + src51[421] + src51[422] + src51[423] + src51[424] + src51[425] + src51[426] + src51[427] + src51[428] + src51[429] + src51[430] + src51[431] + src51[432] + src51[433] + src51[434] + src51[435] + src51[436] + src51[437] + src51[438] + src51[439] + src51[440] + src51[441] + src51[442] + src51[443] + src51[444] + src51[445] + src51[446] + src51[447] + src51[448] + src51[449] + src51[450] + src51[451] + src51[452] + src51[453] + src51[454] + src51[455] + src51[456] + src51[457] + src51[458] + src51[459] + src51[460] + src51[461] + src51[462] + src51[463] + src51[464] + src51[465] + src51[466] + src51[467] + src51[468] + src51[469] + src51[470] + src51[471] + src51[472] + src51[473] + src51[474] + src51[475] + src51[476] + src51[477] + src51[478] + src51[479] + src51[480] + src51[481] + src51[482] + src51[483] + src51[484] + src51[485])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161] + src52[162] + src52[163] + src52[164] + src52[165] + src52[166] + src52[167] + src52[168] + src52[169] + src52[170] + src52[171] + src52[172] + src52[173] + src52[174] + src52[175] + src52[176] + src52[177] + src52[178] + src52[179] + src52[180] + src52[181] + src52[182] + src52[183] + src52[184] + src52[185] + src52[186] + src52[187] + src52[188] + src52[189] + src52[190] + src52[191] + src52[192] + src52[193] + src52[194] + src52[195] + src52[196] + src52[197] + src52[198] + src52[199] + src52[200] + src52[201] + src52[202] + src52[203] + src52[204] + src52[205] + src52[206] + src52[207] + src52[208] + src52[209] + src52[210] + src52[211] + src52[212] + src52[213] + src52[214] + src52[215] + src52[216] + src52[217] + src52[218] + src52[219] + src52[220] + src52[221] + src52[222] + src52[223] + src52[224] + src52[225] + src52[226] + src52[227] + src52[228] + src52[229] + src52[230] + src52[231] + src52[232] + src52[233] + src52[234] + src52[235] + src52[236] + src52[237] + src52[238] + src52[239] + src52[240] + src52[241] + src52[242] + src52[243] + src52[244] + src52[245] + src52[246] + src52[247] + src52[248] + src52[249] + src52[250] + src52[251] + src52[252] + src52[253] + src52[254] + src52[255] + src52[256] + src52[257] + src52[258] + src52[259] + src52[260] + src52[261] + src52[262] + src52[263] + src52[264] + src52[265] + src52[266] + src52[267] + src52[268] + src52[269] + src52[270] + src52[271] + src52[272] + src52[273] + src52[274] + src52[275] + src52[276] + src52[277] + src52[278] + src52[279] + src52[280] + src52[281] + src52[282] + src52[283] + src52[284] + src52[285] + src52[286] + src52[287] + src52[288] + src52[289] + src52[290] + src52[291] + src52[292] + src52[293] + src52[294] + src52[295] + src52[296] + src52[297] + src52[298] + src52[299] + src52[300] + src52[301] + src52[302] + src52[303] + src52[304] + src52[305] + src52[306] + src52[307] + src52[308] + src52[309] + src52[310] + src52[311] + src52[312] + src52[313] + src52[314] + src52[315] + src52[316] + src52[317] + src52[318] + src52[319] + src52[320] + src52[321] + src52[322] + src52[323] + src52[324] + src52[325] + src52[326] + src52[327] + src52[328] + src52[329] + src52[330] + src52[331] + src52[332] + src52[333] + src52[334] + src52[335] + src52[336] + src52[337] + src52[338] + src52[339] + src52[340] + src52[341] + src52[342] + src52[343] + src52[344] + src52[345] + src52[346] + src52[347] + src52[348] + src52[349] + src52[350] + src52[351] + src52[352] + src52[353] + src52[354] + src52[355] + src52[356] + src52[357] + src52[358] + src52[359] + src52[360] + src52[361] + src52[362] + src52[363] + src52[364] + src52[365] + src52[366] + src52[367] + src52[368] + src52[369] + src52[370] + src52[371] + src52[372] + src52[373] + src52[374] + src52[375] + src52[376] + src52[377] + src52[378] + src52[379] + src52[380] + src52[381] + src52[382] + src52[383] + src52[384] + src52[385] + src52[386] + src52[387] + src52[388] + src52[389] + src52[390] + src52[391] + src52[392] + src52[393] + src52[394] + src52[395] + src52[396] + src52[397] + src52[398] + src52[399] + src52[400] + src52[401] + src52[402] + src52[403] + src52[404] + src52[405] + src52[406] + src52[407] + src52[408] + src52[409] + src52[410] + src52[411] + src52[412] + src52[413] + src52[414] + src52[415] + src52[416] + src52[417] + src52[418] + src52[419] + src52[420] + src52[421] + src52[422] + src52[423] + src52[424] + src52[425] + src52[426] + src52[427] + src52[428] + src52[429] + src52[430] + src52[431] + src52[432] + src52[433] + src52[434] + src52[435] + src52[436] + src52[437] + src52[438] + src52[439] + src52[440] + src52[441] + src52[442] + src52[443] + src52[444] + src52[445] + src52[446] + src52[447] + src52[448] + src52[449] + src52[450] + src52[451] + src52[452] + src52[453] + src52[454] + src52[455] + src52[456] + src52[457] + src52[458] + src52[459] + src52[460] + src52[461] + src52[462] + src52[463] + src52[464] + src52[465] + src52[466] + src52[467] + src52[468] + src52[469] + src52[470] + src52[471] + src52[472] + src52[473] + src52[474] + src52[475] + src52[476] + src52[477] + src52[478] + src52[479] + src52[480] + src52[481] + src52[482] + src52[483] + src52[484] + src52[485])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161] + src53[162] + src53[163] + src53[164] + src53[165] + src53[166] + src53[167] + src53[168] + src53[169] + src53[170] + src53[171] + src53[172] + src53[173] + src53[174] + src53[175] + src53[176] + src53[177] + src53[178] + src53[179] + src53[180] + src53[181] + src53[182] + src53[183] + src53[184] + src53[185] + src53[186] + src53[187] + src53[188] + src53[189] + src53[190] + src53[191] + src53[192] + src53[193] + src53[194] + src53[195] + src53[196] + src53[197] + src53[198] + src53[199] + src53[200] + src53[201] + src53[202] + src53[203] + src53[204] + src53[205] + src53[206] + src53[207] + src53[208] + src53[209] + src53[210] + src53[211] + src53[212] + src53[213] + src53[214] + src53[215] + src53[216] + src53[217] + src53[218] + src53[219] + src53[220] + src53[221] + src53[222] + src53[223] + src53[224] + src53[225] + src53[226] + src53[227] + src53[228] + src53[229] + src53[230] + src53[231] + src53[232] + src53[233] + src53[234] + src53[235] + src53[236] + src53[237] + src53[238] + src53[239] + src53[240] + src53[241] + src53[242] + src53[243] + src53[244] + src53[245] + src53[246] + src53[247] + src53[248] + src53[249] + src53[250] + src53[251] + src53[252] + src53[253] + src53[254] + src53[255] + src53[256] + src53[257] + src53[258] + src53[259] + src53[260] + src53[261] + src53[262] + src53[263] + src53[264] + src53[265] + src53[266] + src53[267] + src53[268] + src53[269] + src53[270] + src53[271] + src53[272] + src53[273] + src53[274] + src53[275] + src53[276] + src53[277] + src53[278] + src53[279] + src53[280] + src53[281] + src53[282] + src53[283] + src53[284] + src53[285] + src53[286] + src53[287] + src53[288] + src53[289] + src53[290] + src53[291] + src53[292] + src53[293] + src53[294] + src53[295] + src53[296] + src53[297] + src53[298] + src53[299] + src53[300] + src53[301] + src53[302] + src53[303] + src53[304] + src53[305] + src53[306] + src53[307] + src53[308] + src53[309] + src53[310] + src53[311] + src53[312] + src53[313] + src53[314] + src53[315] + src53[316] + src53[317] + src53[318] + src53[319] + src53[320] + src53[321] + src53[322] + src53[323] + src53[324] + src53[325] + src53[326] + src53[327] + src53[328] + src53[329] + src53[330] + src53[331] + src53[332] + src53[333] + src53[334] + src53[335] + src53[336] + src53[337] + src53[338] + src53[339] + src53[340] + src53[341] + src53[342] + src53[343] + src53[344] + src53[345] + src53[346] + src53[347] + src53[348] + src53[349] + src53[350] + src53[351] + src53[352] + src53[353] + src53[354] + src53[355] + src53[356] + src53[357] + src53[358] + src53[359] + src53[360] + src53[361] + src53[362] + src53[363] + src53[364] + src53[365] + src53[366] + src53[367] + src53[368] + src53[369] + src53[370] + src53[371] + src53[372] + src53[373] + src53[374] + src53[375] + src53[376] + src53[377] + src53[378] + src53[379] + src53[380] + src53[381] + src53[382] + src53[383] + src53[384] + src53[385] + src53[386] + src53[387] + src53[388] + src53[389] + src53[390] + src53[391] + src53[392] + src53[393] + src53[394] + src53[395] + src53[396] + src53[397] + src53[398] + src53[399] + src53[400] + src53[401] + src53[402] + src53[403] + src53[404] + src53[405] + src53[406] + src53[407] + src53[408] + src53[409] + src53[410] + src53[411] + src53[412] + src53[413] + src53[414] + src53[415] + src53[416] + src53[417] + src53[418] + src53[419] + src53[420] + src53[421] + src53[422] + src53[423] + src53[424] + src53[425] + src53[426] + src53[427] + src53[428] + src53[429] + src53[430] + src53[431] + src53[432] + src53[433] + src53[434] + src53[435] + src53[436] + src53[437] + src53[438] + src53[439] + src53[440] + src53[441] + src53[442] + src53[443] + src53[444] + src53[445] + src53[446] + src53[447] + src53[448] + src53[449] + src53[450] + src53[451] + src53[452] + src53[453] + src53[454] + src53[455] + src53[456] + src53[457] + src53[458] + src53[459] + src53[460] + src53[461] + src53[462] + src53[463] + src53[464] + src53[465] + src53[466] + src53[467] + src53[468] + src53[469] + src53[470] + src53[471] + src53[472] + src53[473] + src53[474] + src53[475] + src53[476] + src53[477] + src53[478] + src53[479] + src53[480] + src53[481] + src53[482] + src53[483] + src53[484] + src53[485])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161] + src54[162] + src54[163] + src54[164] + src54[165] + src54[166] + src54[167] + src54[168] + src54[169] + src54[170] + src54[171] + src54[172] + src54[173] + src54[174] + src54[175] + src54[176] + src54[177] + src54[178] + src54[179] + src54[180] + src54[181] + src54[182] + src54[183] + src54[184] + src54[185] + src54[186] + src54[187] + src54[188] + src54[189] + src54[190] + src54[191] + src54[192] + src54[193] + src54[194] + src54[195] + src54[196] + src54[197] + src54[198] + src54[199] + src54[200] + src54[201] + src54[202] + src54[203] + src54[204] + src54[205] + src54[206] + src54[207] + src54[208] + src54[209] + src54[210] + src54[211] + src54[212] + src54[213] + src54[214] + src54[215] + src54[216] + src54[217] + src54[218] + src54[219] + src54[220] + src54[221] + src54[222] + src54[223] + src54[224] + src54[225] + src54[226] + src54[227] + src54[228] + src54[229] + src54[230] + src54[231] + src54[232] + src54[233] + src54[234] + src54[235] + src54[236] + src54[237] + src54[238] + src54[239] + src54[240] + src54[241] + src54[242] + src54[243] + src54[244] + src54[245] + src54[246] + src54[247] + src54[248] + src54[249] + src54[250] + src54[251] + src54[252] + src54[253] + src54[254] + src54[255] + src54[256] + src54[257] + src54[258] + src54[259] + src54[260] + src54[261] + src54[262] + src54[263] + src54[264] + src54[265] + src54[266] + src54[267] + src54[268] + src54[269] + src54[270] + src54[271] + src54[272] + src54[273] + src54[274] + src54[275] + src54[276] + src54[277] + src54[278] + src54[279] + src54[280] + src54[281] + src54[282] + src54[283] + src54[284] + src54[285] + src54[286] + src54[287] + src54[288] + src54[289] + src54[290] + src54[291] + src54[292] + src54[293] + src54[294] + src54[295] + src54[296] + src54[297] + src54[298] + src54[299] + src54[300] + src54[301] + src54[302] + src54[303] + src54[304] + src54[305] + src54[306] + src54[307] + src54[308] + src54[309] + src54[310] + src54[311] + src54[312] + src54[313] + src54[314] + src54[315] + src54[316] + src54[317] + src54[318] + src54[319] + src54[320] + src54[321] + src54[322] + src54[323] + src54[324] + src54[325] + src54[326] + src54[327] + src54[328] + src54[329] + src54[330] + src54[331] + src54[332] + src54[333] + src54[334] + src54[335] + src54[336] + src54[337] + src54[338] + src54[339] + src54[340] + src54[341] + src54[342] + src54[343] + src54[344] + src54[345] + src54[346] + src54[347] + src54[348] + src54[349] + src54[350] + src54[351] + src54[352] + src54[353] + src54[354] + src54[355] + src54[356] + src54[357] + src54[358] + src54[359] + src54[360] + src54[361] + src54[362] + src54[363] + src54[364] + src54[365] + src54[366] + src54[367] + src54[368] + src54[369] + src54[370] + src54[371] + src54[372] + src54[373] + src54[374] + src54[375] + src54[376] + src54[377] + src54[378] + src54[379] + src54[380] + src54[381] + src54[382] + src54[383] + src54[384] + src54[385] + src54[386] + src54[387] + src54[388] + src54[389] + src54[390] + src54[391] + src54[392] + src54[393] + src54[394] + src54[395] + src54[396] + src54[397] + src54[398] + src54[399] + src54[400] + src54[401] + src54[402] + src54[403] + src54[404] + src54[405] + src54[406] + src54[407] + src54[408] + src54[409] + src54[410] + src54[411] + src54[412] + src54[413] + src54[414] + src54[415] + src54[416] + src54[417] + src54[418] + src54[419] + src54[420] + src54[421] + src54[422] + src54[423] + src54[424] + src54[425] + src54[426] + src54[427] + src54[428] + src54[429] + src54[430] + src54[431] + src54[432] + src54[433] + src54[434] + src54[435] + src54[436] + src54[437] + src54[438] + src54[439] + src54[440] + src54[441] + src54[442] + src54[443] + src54[444] + src54[445] + src54[446] + src54[447] + src54[448] + src54[449] + src54[450] + src54[451] + src54[452] + src54[453] + src54[454] + src54[455] + src54[456] + src54[457] + src54[458] + src54[459] + src54[460] + src54[461] + src54[462] + src54[463] + src54[464] + src54[465] + src54[466] + src54[467] + src54[468] + src54[469] + src54[470] + src54[471] + src54[472] + src54[473] + src54[474] + src54[475] + src54[476] + src54[477] + src54[478] + src54[479] + src54[480] + src54[481] + src54[482] + src54[483] + src54[484] + src54[485])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161] + src55[162] + src55[163] + src55[164] + src55[165] + src55[166] + src55[167] + src55[168] + src55[169] + src55[170] + src55[171] + src55[172] + src55[173] + src55[174] + src55[175] + src55[176] + src55[177] + src55[178] + src55[179] + src55[180] + src55[181] + src55[182] + src55[183] + src55[184] + src55[185] + src55[186] + src55[187] + src55[188] + src55[189] + src55[190] + src55[191] + src55[192] + src55[193] + src55[194] + src55[195] + src55[196] + src55[197] + src55[198] + src55[199] + src55[200] + src55[201] + src55[202] + src55[203] + src55[204] + src55[205] + src55[206] + src55[207] + src55[208] + src55[209] + src55[210] + src55[211] + src55[212] + src55[213] + src55[214] + src55[215] + src55[216] + src55[217] + src55[218] + src55[219] + src55[220] + src55[221] + src55[222] + src55[223] + src55[224] + src55[225] + src55[226] + src55[227] + src55[228] + src55[229] + src55[230] + src55[231] + src55[232] + src55[233] + src55[234] + src55[235] + src55[236] + src55[237] + src55[238] + src55[239] + src55[240] + src55[241] + src55[242] + src55[243] + src55[244] + src55[245] + src55[246] + src55[247] + src55[248] + src55[249] + src55[250] + src55[251] + src55[252] + src55[253] + src55[254] + src55[255] + src55[256] + src55[257] + src55[258] + src55[259] + src55[260] + src55[261] + src55[262] + src55[263] + src55[264] + src55[265] + src55[266] + src55[267] + src55[268] + src55[269] + src55[270] + src55[271] + src55[272] + src55[273] + src55[274] + src55[275] + src55[276] + src55[277] + src55[278] + src55[279] + src55[280] + src55[281] + src55[282] + src55[283] + src55[284] + src55[285] + src55[286] + src55[287] + src55[288] + src55[289] + src55[290] + src55[291] + src55[292] + src55[293] + src55[294] + src55[295] + src55[296] + src55[297] + src55[298] + src55[299] + src55[300] + src55[301] + src55[302] + src55[303] + src55[304] + src55[305] + src55[306] + src55[307] + src55[308] + src55[309] + src55[310] + src55[311] + src55[312] + src55[313] + src55[314] + src55[315] + src55[316] + src55[317] + src55[318] + src55[319] + src55[320] + src55[321] + src55[322] + src55[323] + src55[324] + src55[325] + src55[326] + src55[327] + src55[328] + src55[329] + src55[330] + src55[331] + src55[332] + src55[333] + src55[334] + src55[335] + src55[336] + src55[337] + src55[338] + src55[339] + src55[340] + src55[341] + src55[342] + src55[343] + src55[344] + src55[345] + src55[346] + src55[347] + src55[348] + src55[349] + src55[350] + src55[351] + src55[352] + src55[353] + src55[354] + src55[355] + src55[356] + src55[357] + src55[358] + src55[359] + src55[360] + src55[361] + src55[362] + src55[363] + src55[364] + src55[365] + src55[366] + src55[367] + src55[368] + src55[369] + src55[370] + src55[371] + src55[372] + src55[373] + src55[374] + src55[375] + src55[376] + src55[377] + src55[378] + src55[379] + src55[380] + src55[381] + src55[382] + src55[383] + src55[384] + src55[385] + src55[386] + src55[387] + src55[388] + src55[389] + src55[390] + src55[391] + src55[392] + src55[393] + src55[394] + src55[395] + src55[396] + src55[397] + src55[398] + src55[399] + src55[400] + src55[401] + src55[402] + src55[403] + src55[404] + src55[405] + src55[406] + src55[407] + src55[408] + src55[409] + src55[410] + src55[411] + src55[412] + src55[413] + src55[414] + src55[415] + src55[416] + src55[417] + src55[418] + src55[419] + src55[420] + src55[421] + src55[422] + src55[423] + src55[424] + src55[425] + src55[426] + src55[427] + src55[428] + src55[429] + src55[430] + src55[431] + src55[432] + src55[433] + src55[434] + src55[435] + src55[436] + src55[437] + src55[438] + src55[439] + src55[440] + src55[441] + src55[442] + src55[443] + src55[444] + src55[445] + src55[446] + src55[447] + src55[448] + src55[449] + src55[450] + src55[451] + src55[452] + src55[453] + src55[454] + src55[455] + src55[456] + src55[457] + src55[458] + src55[459] + src55[460] + src55[461] + src55[462] + src55[463] + src55[464] + src55[465] + src55[466] + src55[467] + src55[468] + src55[469] + src55[470] + src55[471] + src55[472] + src55[473] + src55[474] + src55[475] + src55[476] + src55[477] + src55[478] + src55[479] + src55[480] + src55[481] + src55[482] + src55[483] + src55[484] + src55[485])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161] + src56[162] + src56[163] + src56[164] + src56[165] + src56[166] + src56[167] + src56[168] + src56[169] + src56[170] + src56[171] + src56[172] + src56[173] + src56[174] + src56[175] + src56[176] + src56[177] + src56[178] + src56[179] + src56[180] + src56[181] + src56[182] + src56[183] + src56[184] + src56[185] + src56[186] + src56[187] + src56[188] + src56[189] + src56[190] + src56[191] + src56[192] + src56[193] + src56[194] + src56[195] + src56[196] + src56[197] + src56[198] + src56[199] + src56[200] + src56[201] + src56[202] + src56[203] + src56[204] + src56[205] + src56[206] + src56[207] + src56[208] + src56[209] + src56[210] + src56[211] + src56[212] + src56[213] + src56[214] + src56[215] + src56[216] + src56[217] + src56[218] + src56[219] + src56[220] + src56[221] + src56[222] + src56[223] + src56[224] + src56[225] + src56[226] + src56[227] + src56[228] + src56[229] + src56[230] + src56[231] + src56[232] + src56[233] + src56[234] + src56[235] + src56[236] + src56[237] + src56[238] + src56[239] + src56[240] + src56[241] + src56[242] + src56[243] + src56[244] + src56[245] + src56[246] + src56[247] + src56[248] + src56[249] + src56[250] + src56[251] + src56[252] + src56[253] + src56[254] + src56[255] + src56[256] + src56[257] + src56[258] + src56[259] + src56[260] + src56[261] + src56[262] + src56[263] + src56[264] + src56[265] + src56[266] + src56[267] + src56[268] + src56[269] + src56[270] + src56[271] + src56[272] + src56[273] + src56[274] + src56[275] + src56[276] + src56[277] + src56[278] + src56[279] + src56[280] + src56[281] + src56[282] + src56[283] + src56[284] + src56[285] + src56[286] + src56[287] + src56[288] + src56[289] + src56[290] + src56[291] + src56[292] + src56[293] + src56[294] + src56[295] + src56[296] + src56[297] + src56[298] + src56[299] + src56[300] + src56[301] + src56[302] + src56[303] + src56[304] + src56[305] + src56[306] + src56[307] + src56[308] + src56[309] + src56[310] + src56[311] + src56[312] + src56[313] + src56[314] + src56[315] + src56[316] + src56[317] + src56[318] + src56[319] + src56[320] + src56[321] + src56[322] + src56[323] + src56[324] + src56[325] + src56[326] + src56[327] + src56[328] + src56[329] + src56[330] + src56[331] + src56[332] + src56[333] + src56[334] + src56[335] + src56[336] + src56[337] + src56[338] + src56[339] + src56[340] + src56[341] + src56[342] + src56[343] + src56[344] + src56[345] + src56[346] + src56[347] + src56[348] + src56[349] + src56[350] + src56[351] + src56[352] + src56[353] + src56[354] + src56[355] + src56[356] + src56[357] + src56[358] + src56[359] + src56[360] + src56[361] + src56[362] + src56[363] + src56[364] + src56[365] + src56[366] + src56[367] + src56[368] + src56[369] + src56[370] + src56[371] + src56[372] + src56[373] + src56[374] + src56[375] + src56[376] + src56[377] + src56[378] + src56[379] + src56[380] + src56[381] + src56[382] + src56[383] + src56[384] + src56[385] + src56[386] + src56[387] + src56[388] + src56[389] + src56[390] + src56[391] + src56[392] + src56[393] + src56[394] + src56[395] + src56[396] + src56[397] + src56[398] + src56[399] + src56[400] + src56[401] + src56[402] + src56[403] + src56[404] + src56[405] + src56[406] + src56[407] + src56[408] + src56[409] + src56[410] + src56[411] + src56[412] + src56[413] + src56[414] + src56[415] + src56[416] + src56[417] + src56[418] + src56[419] + src56[420] + src56[421] + src56[422] + src56[423] + src56[424] + src56[425] + src56[426] + src56[427] + src56[428] + src56[429] + src56[430] + src56[431] + src56[432] + src56[433] + src56[434] + src56[435] + src56[436] + src56[437] + src56[438] + src56[439] + src56[440] + src56[441] + src56[442] + src56[443] + src56[444] + src56[445] + src56[446] + src56[447] + src56[448] + src56[449] + src56[450] + src56[451] + src56[452] + src56[453] + src56[454] + src56[455] + src56[456] + src56[457] + src56[458] + src56[459] + src56[460] + src56[461] + src56[462] + src56[463] + src56[464] + src56[465] + src56[466] + src56[467] + src56[468] + src56[469] + src56[470] + src56[471] + src56[472] + src56[473] + src56[474] + src56[475] + src56[476] + src56[477] + src56[478] + src56[479] + src56[480] + src56[481] + src56[482] + src56[483] + src56[484] + src56[485])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161] + src57[162] + src57[163] + src57[164] + src57[165] + src57[166] + src57[167] + src57[168] + src57[169] + src57[170] + src57[171] + src57[172] + src57[173] + src57[174] + src57[175] + src57[176] + src57[177] + src57[178] + src57[179] + src57[180] + src57[181] + src57[182] + src57[183] + src57[184] + src57[185] + src57[186] + src57[187] + src57[188] + src57[189] + src57[190] + src57[191] + src57[192] + src57[193] + src57[194] + src57[195] + src57[196] + src57[197] + src57[198] + src57[199] + src57[200] + src57[201] + src57[202] + src57[203] + src57[204] + src57[205] + src57[206] + src57[207] + src57[208] + src57[209] + src57[210] + src57[211] + src57[212] + src57[213] + src57[214] + src57[215] + src57[216] + src57[217] + src57[218] + src57[219] + src57[220] + src57[221] + src57[222] + src57[223] + src57[224] + src57[225] + src57[226] + src57[227] + src57[228] + src57[229] + src57[230] + src57[231] + src57[232] + src57[233] + src57[234] + src57[235] + src57[236] + src57[237] + src57[238] + src57[239] + src57[240] + src57[241] + src57[242] + src57[243] + src57[244] + src57[245] + src57[246] + src57[247] + src57[248] + src57[249] + src57[250] + src57[251] + src57[252] + src57[253] + src57[254] + src57[255] + src57[256] + src57[257] + src57[258] + src57[259] + src57[260] + src57[261] + src57[262] + src57[263] + src57[264] + src57[265] + src57[266] + src57[267] + src57[268] + src57[269] + src57[270] + src57[271] + src57[272] + src57[273] + src57[274] + src57[275] + src57[276] + src57[277] + src57[278] + src57[279] + src57[280] + src57[281] + src57[282] + src57[283] + src57[284] + src57[285] + src57[286] + src57[287] + src57[288] + src57[289] + src57[290] + src57[291] + src57[292] + src57[293] + src57[294] + src57[295] + src57[296] + src57[297] + src57[298] + src57[299] + src57[300] + src57[301] + src57[302] + src57[303] + src57[304] + src57[305] + src57[306] + src57[307] + src57[308] + src57[309] + src57[310] + src57[311] + src57[312] + src57[313] + src57[314] + src57[315] + src57[316] + src57[317] + src57[318] + src57[319] + src57[320] + src57[321] + src57[322] + src57[323] + src57[324] + src57[325] + src57[326] + src57[327] + src57[328] + src57[329] + src57[330] + src57[331] + src57[332] + src57[333] + src57[334] + src57[335] + src57[336] + src57[337] + src57[338] + src57[339] + src57[340] + src57[341] + src57[342] + src57[343] + src57[344] + src57[345] + src57[346] + src57[347] + src57[348] + src57[349] + src57[350] + src57[351] + src57[352] + src57[353] + src57[354] + src57[355] + src57[356] + src57[357] + src57[358] + src57[359] + src57[360] + src57[361] + src57[362] + src57[363] + src57[364] + src57[365] + src57[366] + src57[367] + src57[368] + src57[369] + src57[370] + src57[371] + src57[372] + src57[373] + src57[374] + src57[375] + src57[376] + src57[377] + src57[378] + src57[379] + src57[380] + src57[381] + src57[382] + src57[383] + src57[384] + src57[385] + src57[386] + src57[387] + src57[388] + src57[389] + src57[390] + src57[391] + src57[392] + src57[393] + src57[394] + src57[395] + src57[396] + src57[397] + src57[398] + src57[399] + src57[400] + src57[401] + src57[402] + src57[403] + src57[404] + src57[405] + src57[406] + src57[407] + src57[408] + src57[409] + src57[410] + src57[411] + src57[412] + src57[413] + src57[414] + src57[415] + src57[416] + src57[417] + src57[418] + src57[419] + src57[420] + src57[421] + src57[422] + src57[423] + src57[424] + src57[425] + src57[426] + src57[427] + src57[428] + src57[429] + src57[430] + src57[431] + src57[432] + src57[433] + src57[434] + src57[435] + src57[436] + src57[437] + src57[438] + src57[439] + src57[440] + src57[441] + src57[442] + src57[443] + src57[444] + src57[445] + src57[446] + src57[447] + src57[448] + src57[449] + src57[450] + src57[451] + src57[452] + src57[453] + src57[454] + src57[455] + src57[456] + src57[457] + src57[458] + src57[459] + src57[460] + src57[461] + src57[462] + src57[463] + src57[464] + src57[465] + src57[466] + src57[467] + src57[468] + src57[469] + src57[470] + src57[471] + src57[472] + src57[473] + src57[474] + src57[475] + src57[476] + src57[477] + src57[478] + src57[479] + src57[480] + src57[481] + src57[482] + src57[483] + src57[484] + src57[485])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161] + src58[162] + src58[163] + src58[164] + src58[165] + src58[166] + src58[167] + src58[168] + src58[169] + src58[170] + src58[171] + src58[172] + src58[173] + src58[174] + src58[175] + src58[176] + src58[177] + src58[178] + src58[179] + src58[180] + src58[181] + src58[182] + src58[183] + src58[184] + src58[185] + src58[186] + src58[187] + src58[188] + src58[189] + src58[190] + src58[191] + src58[192] + src58[193] + src58[194] + src58[195] + src58[196] + src58[197] + src58[198] + src58[199] + src58[200] + src58[201] + src58[202] + src58[203] + src58[204] + src58[205] + src58[206] + src58[207] + src58[208] + src58[209] + src58[210] + src58[211] + src58[212] + src58[213] + src58[214] + src58[215] + src58[216] + src58[217] + src58[218] + src58[219] + src58[220] + src58[221] + src58[222] + src58[223] + src58[224] + src58[225] + src58[226] + src58[227] + src58[228] + src58[229] + src58[230] + src58[231] + src58[232] + src58[233] + src58[234] + src58[235] + src58[236] + src58[237] + src58[238] + src58[239] + src58[240] + src58[241] + src58[242] + src58[243] + src58[244] + src58[245] + src58[246] + src58[247] + src58[248] + src58[249] + src58[250] + src58[251] + src58[252] + src58[253] + src58[254] + src58[255] + src58[256] + src58[257] + src58[258] + src58[259] + src58[260] + src58[261] + src58[262] + src58[263] + src58[264] + src58[265] + src58[266] + src58[267] + src58[268] + src58[269] + src58[270] + src58[271] + src58[272] + src58[273] + src58[274] + src58[275] + src58[276] + src58[277] + src58[278] + src58[279] + src58[280] + src58[281] + src58[282] + src58[283] + src58[284] + src58[285] + src58[286] + src58[287] + src58[288] + src58[289] + src58[290] + src58[291] + src58[292] + src58[293] + src58[294] + src58[295] + src58[296] + src58[297] + src58[298] + src58[299] + src58[300] + src58[301] + src58[302] + src58[303] + src58[304] + src58[305] + src58[306] + src58[307] + src58[308] + src58[309] + src58[310] + src58[311] + src58[312] + src58[313] + src58[314] + src58[315] + src58[316] + src58[317] + src58[318] + src58[319] + src58[320] + src58[321] + src58[322] + src58[323] + src58[324] + src58[325] + src58[326] + src58[327] + src58[328] + src58[329] + src58[330] + src58[331] + src58[332] + src58[333] + src58[334] + src58[335] + src58[336] + src58[337] + src58[338] + src58[339] + src58[340] + src58[341] + src58[342] + src58[343] + src58[344] + src58[345] + src58[346] + src58[347] + src58[348] + src58[349] + src58[350] + src58[351] + src58[352] + src58[353] + src58[354] + src58[355] + src58[356] + src58[357] + src58[358] + src58[359] + src58[360] + src58[361] + src58[362] + src58[363] + src58[364] + src58[365] + src58[366] + src58[367] + src58[368] + src58[369] + src58[370] + src58[371] + src58[372] + src58[373] + src58[374] + src58[375] + src58[376] + src58[377] + src58[378] + src58[379] + src58[380] + src58[381] + src58[382] + src58[383] + src58[384] + src58[385] + src58[386] + src58[387] + src58[388] + src58[389] + src58[390] + src58[391] + src58[392] + src58[393] + src58[394] + src58[395] + src58[396] + src58[397] + src58[398] + src58[399] + src58[400] + src58[401] + src58[402] + src58[403] + src58[404] + src58[405] + src58[406] + src58[407] + src58[408] + src58[409] + src58[410] + src58[411] + src58[412] + src58[413] + src58[414] + src58[415] + src58[416] + src58[417] + src58[418] + src58[419] + src58[420] + src58[421] + src58[422] + src58[423] + src58[424] + src58[425] + src58[426] + src58[427] + src58[428] + src58[429] + src58[430] + src58[431] + src58[432] + src58[433] + src58[434] + src58[435] + src58[436] + src58[437] + src58[438] + src58[439] + src58[440] + src58[441] + src58[442] + src58[443] + src58[444] + src58[445] + src58[446] + src58[447] + src58[448] + src58[449] + src58[450] + src58[451] + src58[452] + src58[453] + src58[454] + src58[455] + src58[456] + src58[457] + src58[458] + src58[459] + src58[460] + src58[461] + src58[462] + src58[463] + src58[464] + src58[465] + src58[466] + src58[467] + src58[468] + src58[469] + src58[470] + src58[471] + src58[472] + src58[473] + src58[474] + src58[475] + src58[476] + src58[477] + src58[478] + src58[479] + src58[480] + src58[481] + src58[482] + src58[483] + src58[484] + src58[485])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161] + src59[162] + src59[163] + src59[164] + src59[165] + src59[166] + src59[167] + src59[168] + src59[169] + src59[170] + src59[171] + src59[172] + src59[173] + src59[174] + src59[175] + src59[176] + src59[177] + src59[178] + src59[179] + src59[180] + src59[181] + src59[182] + src59[183] + src59[184] + src59[185] + src59[186] + src59[187] + src59[188] + src59[189] + src59[190] + src59[191] + src59[192] + src59[193] + src59[194] + src59[195] + src59[196] + src59[197] + src59[198] + src59[199] + src59[200] + src59[201] + src59[202] + src59[203] + src59[204] + src59[205] + src59[206] + src59[207] + src59[208] + src59[209] + src59[210] + src59[211] + src59[212] + src59[213] + src59[214] + src59[215] + src59[216] + src59[217] + src59[218] + src59[219] + src59[220] + src59[221] + src59[222] + src59[223] + src59[224] + src59[225] + src59[226] + src59[227] + src59[228] + src59[229] + src59[230] + src59[231] + src59[232] + src59[233] + src59[234] + src59[235] + src59[236] + src59[237] + src59[238] + src59[239] + src59[240] + src59[241] + src59[242] + src59[243] + src59[244] + src59[245] + src59[246] + src59[247] + src59[248] + src59[249] + src59[250] + src59[251] + src59[252] + src59[253] + src59[254] + src59[255] + src59[256] + src59[257] + src59[258] + src59[259] + src59[260] + src59[261] + src59[262] + src59[263] + src59[264] + src59[265] + src59[266] + src59[267] + src59[268] + src59[269] + src59[270] + src59[271] + src59[272] + src59[273] + src59[274] + src59[275] + src59[276] + src59[277] + src59[278] + src59[279] + src59[280] + src59[281] + src59[282] + src59[283] + src59[284] + src59[285] + src59[286] + src59[287] + src59[288] + src59[289] + src59[290] + src59[291] + src59[292] + src59[293] + src59[294] + src59[295] + src59[296] + src59[297] + src59[298] + src59[299] + src59[300] + src59[301] + src59[302] + src59[303] + src59[304] + src59[305] + src59[306] + src59[307] + src59[308] + src59[309] + src59[310] + src59[311] + src59[312] + src59[313] + src59[314] + src59[315] + src59[316] + src59[317] + src59[318] + src59[319] + src59[320] + src59[321] + src59[322] + src59[323] + src59[324] + src59[325] + src59[326] + src59[327] + src59[328] + src59[329] + src59[330] + src59[331] + src59[332] + src59[333] + src59[334] + src59[335] + src59[336] + src59[337] + src59[338] + src59[339] + src59[340] + src59[341] + src59[342] + src59[343] + src59[344] + src59[345] + src59[346] + src59[347] + src59[348] + src59[349] + src59[350] + src59[351] + src59[352] + src59[353] + src59[354] + src59[355] + src59[356] + src59[357] + src59[358] + src59[359] + src59[360] + src59[361] + src59[362] + src59[363] + src59[364] + src59[365] + src59[366] + src59[367] + src59[368] + src59[369] + src59[370] + src59[371] + src59[372] + src59[373] + src59[374] + src59[375] + src59[376] + src59[377] + src59[378] + src59[379] + src59[380] + src59[381] + src59[382] + src59[383] + src59[384] + src59[385] + src59[386] + src59[387] + src59[388] + src59[389] + src59[390] + src59[391] + src59[392] + src59[393] + src59[394] + src59[395] + src59[396] + src59[397] + src59[398] + src59[399] + src59[400] + src59[401] + src59[402] + src59[403] + src59[404] + src59[405] + src59[406] + src59[407] + src59[408] + src59[409] + src59[410] + src59[411] + src59[412] + src59[413] + src59[414] + src59[415] + src59[416] + src59[417] + src59[418] + src59[419] + src59[420] + src59[421] + src59[422] + src59[423] + src59[424] + src59[425] + src59[426] + src59[427] + src59[428] + src59[429] + src59[430] + src59[431] + src59[432] + src59[433] + src59[434] + src59[435] + src59[436] + src59[437] + src59[438] + src59[439] + src59[440] + src59[441] + src59[442] + src59[443] + src59[444] + src59[445] + src59[446] + src59[447] + src59[448] + src59[449] + src59[450] + src59[451] + src59[452] + src59[453] + src59[454] + src59[455] + src59[456] + src59[457] + src59[458] + src59[459] + src59[460] + src59[461] + src59[462] + src59[463] + src59[464] + src59[465] + src59[466] + src59[467] + src59[468] + src59[469] + src59[470] + src59[471] + src59[472] + src59[473] + src59[474] + src59[475] + src59[476] + src59[477] + src59[478] + src59[479] + src59[480] + src59[481] + src59[482] + src59[483] + src59[484] + src59[485])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161] + src60[162] + src60[163] + src60[164] + src60[165] + src60[166] + src60[167] + src60[168] + src60[169] + src60[170] + src60[171] + src60[172] + src60[173] + src60[174] + src60[175] + src60[176] + src60[177] + src60[178] + src60[179] + src60[180] + src60[181] + src60[182] + src60[183] + src60[184] + src60[185] + src60[186] + src60[187] + src60[188] + src60[189] + src60[190] + src60[191] + src60[192] + src60[193] + src60[194] + src60[195] + src60[196] + src60[197] + src60[198] + src60[199] + src60[200] + src60[201] + src60[202] + src60[203] + src60[204] + src60[205] + src60[206] + src60[207] + src60[208] + src60[209] + src60[210] + src60[211] + src60[212] + src60[213] + src60[214] + src60[215] + src60[216] + src60[217] + src60[218] + src60[219] + src60[220] + src60[221] + src60[222] + src60[223] + src60[224] + src60[225] + src60[226] + src60[227] + src60[228] + src60[229] + src60[230] + src60[231] + src60[232] + src60[233] + src60[234] + src60[235] + src60[236] + src60[237] + src60[238] + src60[239] + src60[240] + src60[241] + src60[242] + src60[243] + src60[244] + src60[245] + src60[246] + src60[247] + src60[248] + src60[249] + src60[250] + src60[251] + src60[252] + src60[253] + src60[254] + src60[255] + src60[256] + src60[257] + src60[258] + src60[259] + src60[260] + src60[261] + src60[262] + src60[263] + src60[264] + src60[265] + src60[266] + src60[267] + src60[268] + src60[269] + src60[270] + src60[271] + src60[272] + src60[273] + src60[274] + src60[275] + src60[276] + src60[277] + src60[278] + src60[279] + src60[280] + src60[281] + src60[282] + src60[283] + src60[284] + src60[285] + src60[286] + src60[287] + src60[288] + src60[289] + src60[290] + src60[291] + src60[292] + src60[293] + src60[294] + src60[295] + src60[296] + src60[297] + src60[298] + src60[299] + src60[300] + src60[301] + src60[302] + src60[303] + src60[304] + src60[305] + src60[306] + src60[307] + src60[308] + src60[309] + src60[310] + src60[311] + src60[312] + src60[313] + src60[314] + src60[315] + src60[316] + src60[317] + src60[318] + src60[319] + src60[320] + src60[321] + src60[322] + src60[323] + src60[324] + src60[325] + src60[326] + src60[327] + src60[328] + src60[329] + src60[330] + src60[331] + src60[332] + src60[333] + src60[334] + src60[335] + src60[336] + src60[337] + src60[338] + src60[339] + src60[340] + src60[341] + src60[342] + src60[343] + src60[344] + src60[345] + src60[346] + src60[347] + src60[348] + src60[349] + src60[350] + src60[351] + src60[352] + src60[353] + src60[354] + src60[355] + src60[356] + src60[357] + src60[358] + src60[359] + src60[360] + src60[361] + src60[362] + src60[363] + src60[364] + src60[365] + src60[366] + src60[367] + src60[368] + src60[369] + src60[370] + src60[371] + src60[372] + src60[373] + src60[374] + src60[375] + src60[376] + src60[377] + src60[378] + src60[379] + src60[380] + src60[381] + src60[382] + src60[383] + src60[384] + src60[385] + src60[386] + src60[387] + src60[388] + src60[389] + src60[390] + src60[391] + src60[392] + src60[393] + src60[394] + src60[395] + src60[396] + src60[397] + src60[398] + src60[399] + src60[400] + src60[401] + src60[402] + src60[403] + src60[404] + src60[405] + src60[406] + src60[407] + src60[408] + src60[409] + src60[410] + src60[411] + src60[412] + src60[413] + src60[414] + src60[415] + src60[416] + src60[417] + src60[418] + src60[419] + src60[420] + src60[421] + src60[422] + src60[423] + src60[424] + src60[425] + src60[426] + src60[427] + src60[428] + src60[429] + src60[430] + src60[431] + src60[432] + src60[433] + src60[434] + src60[435] + src60[436] + src60[437] + src60[438] + src60[439] + src60[440] + src60[441] + src60[442] + src60[443] + src60[444] + src60[445] + src60[446] + src60[447] + src60[448] + src60[449] + src60[450] + src60[451] + src60[452] + src60[453] + src60[454] + src60[455] + src60[456] + src60[457] + src60[458] + src60[459] + src60[460] + src60[461] + src60[462] + src60[463] + src60[464] + src60[465] + src60[466] + src60[467] + src60[468] + src60[469] + src60[470] + src60[471] + src60[472] + src60[473] + src60[474] + src60[475] + src60[476] + src60[477] + src60[478] + src60[479] + src60[480] + src60[481] + src60[482] + src60[483] + src60[484] + src60[485])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161] + src61[162] + src61[163] + src61[164] + src61[165] + src61[166] + src61[167] + src61[168] + src61[169] + src61[170] + src61[171] + src61[172] + src61[173] + src61[174] + src61[175] + src61[176] + src61[177] + src61[178] + src61[179] + src61[180] + src61[181] + src61[182] + src61[183] + src61[184] + src61[185] + src61[186] + src61[187] + src61[188] + src61[189] + src61[190] + src61[191] + src61[192] + src61[193] + src61[194] + src61[195] + src61[196] + src61[197] + src61[198] + src61[199] + src61[200] + src61[201] + src61[202] + src61[203] + src61[204] + src61[205] + src61[206] + src61[207] + src61[208] + src61[209] + src61[210] + src61[211] + src61[212] + src61[213] + src61[214] + src61[215] + src61[216] + src61[217] + src61[218] + src61[219] + src61[220] + src61[221] + src61[222] + src61[223] + src61[224] + src61[225] + src61[226] + src61[227] + src61[228] + src61[229] + src61[230] + src61[231] + src61[232] + src61[233] + src61[234] + src61[235] + src61[236] + src61[237] + src61[238] + src61[239] + src61[240] + src61[241] + src61[242] + src61[243] + src61[244] + src61[245] + src61[246] + src61[247] + src61[248] + src61[249] + src61[250] + src61[251] + src61[252] + src61[253] + src61[254] + src61[255] + src61[256] + src61[257] + src61[258] + src61[259] + src61[260] + src61[261] + src61[262] + src61[263] + src61[264] + src61[265] + src61[266] + src61[267] + src61[268] + src61[269] + src61[270] + src61[271] + src61[272] + src61[273] + src61[274] + src61[275] + src61[276] + src61[277] + src61[278] + src61[279] + src61[280] + src61[281] + src61[282] + src61[283] + src61[284] + src61[285] + src61[286] + src61[287] + src61[288] + src61[289] + src61[290] + src61[291] + src61[292] + src61[293] + src61[294] + src61[295] + src61[296] + src61[297] + src61[298] + src61[299] + src61[300] + src61[301] + src61[302] + src61[303] + src61[304] + src61[305] + src61[306] + src61[307] + src61[308] + src61[309] + src61[310] + src61[311] + src61[312] + src61[313] + src61[314] + src61[315] + src61[316] + src61[317] + src61[318] + src61[319] + src61[320] + src61[321] + src61[322] + src61[323] + src61[324] + src61[325] + src61[326] + src61[327] + src61[328] + src61[329] + src61[330] + src61[331] + src61[332] + src61[333] + src61[334] + src61[335] + src61[336] + src61[337] + src61[338] + src61[339] + src61[340] + src61[341] + src61[342] + src61[343] + src61[344] + src61[345] + src61[346] + src61[347] + src61[348] + src61[349] + src61[350] + src61[351] + src61[352] + src61[353] + src61[354] + src61[355] + src61[356] + src61[357] + src61[358] + src61[359] + src61[360] + src61[361] + src61[362] + src61[363] + src61[364] + src61[365] + src61[366] + src61[367] + src61[368] + src61[369] + src61[370] + src61[371] + src61[372] + src61[373] + src61[374] + src61[375] + src61[376] + src61[377] + src61[378] + src61[379] + src61[380] + src61[381] + src61[382] + src61[383] + src61[384] + src61[385] + src61[386] + src61[387] + src61[388] + src61[389] + src61[390] + src61[391] + src61[392] + src61[393] + src61[394] + src61[395] + src61[396] + src61[397] + src61[398] + src61[399] + src61[400] + src61[401] + src61[402] + src61[403] + src61[404] + src61[405] + src61[406] + src61[407] + src61[408] + src61[409] + src61[410] + src61[411] + src61[412] + src61[413] + src61[414] + src61[415] + src61[416] + src61[417] + src61[418] + src61[419] + src61[420] + src61[421] + src61[422] + src61[423] + src61[424] + src61[425] + src61[426] + src61[427] + src61[428] + src61[429] + src61[430] + src61[431] + src61[432] + src61[433] + src61[434] + src61[435] + src61[436] + src61[437] + src61[438] + src61[439] + src61[440] + src61[441] + src61[442] + src61[443] + src61[444] + src61[445] + src61[446] + src61[447] + src61[448] + src61[449] + src61[450] + src61[451] + src61[452] + src61[453] + src61[454] + src61[455] + src61[456] + src61[457] + src61[458] + src61[459] + src61[460] + src61[461] + src61[462] + src61[463] + src61[464] + src61[465] + src61[466] + src61[467] + src61[468] + src61[469] + src61[470] + src61[471] + src61[472] + src61[473] + src61[474] + src61[475] + src61[476] + src61[477] + src61[478] + src61[479] + src61[480] + src61[481] + src61[482] + src61[483] + src61[484] + src61[485])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161] + src62[162] + src62[163] + src62[164] + src62[165] + src62[166] + src62[167] + src62[168] + src62[169] + src62[170] + src62[171] + src62[172] + src62[173] + src62[174] + src62[175] + src62[176] + src62[177] + src62[178] + src62[179] + src62[180] + src62[181] + src62[182] + src62[183] + src62[184] + src62[185] + src62[186] + src62[187] + src62[188] + src62[189] + src62[190] + src62[191] + src62[192] + src62[193] + src62[194] + src62[195] + src62[196] + src62[197] + src62[198] + src62[199] + src62[200] + src62[201] + src62[202] + src62[203] + src62[204] + src62[205] + src62[206] + src62[207] + src62[208] + src62[209] + src62[210] + src62[211] + src62[212] + src62[213] + src62[214] + src62[215] + src62[216] + src62[217] + src62[218] + src62[219] + src62[220] + src62[221] + src62[222] + src62[223] + src62[224] + src62[225] + src62[226] + src62[227] + src62[228] + src62[229] + src62[230] + src62[231] + src62[232] + src62[233] + src62[234] + src62[235] + src62[236] + src62[237] + src62[238] + src62[239] + src62[240] + src62[241] + src62[242] + src62[243] + src62[244] + src62[245] + src62[246] + src62[247] + src62[248] + src62[249] + src62[250] + src62[251] + src62[252] + src62[253] + src62[254] + src62[255] + src62[256] + src62[257] + src62[258] + src62[259] + src62[260] + src62[261] + src62[262] + src62[263] + src62[264] + src62[265] + src62[266] + src62[267] + src62[268] + src62[269] + src62[270] + src62[271] + src62[272] + src62[273] + src62[274] + src62[275] + src62[276] + src62[277] + src62[278] + src62[279] + src62[280] + src62[281] + src62[282] + src62[283] + src62[284] + src62[285] + src62[286] + src62[287] + src62[288] + src62[289] + src62[290] + src62[291] + src62[292] + src62[293] + src62[294] + src62[295] + src62[296] + src62[297] + src62[298] + src62[299] + src62[300] + src62[301] + src62[302] + src62[303] + src62[304] + src62[305] + src62[306] + src62[307] + src62[308] + src62[309] + src62[310] + src62[311] + src62[312] + src62[313] + src62[314] + src62[315] + src62[316] + src62[317] + src62[318] + src62[319] + src62[320] + src62[321] + src62[322] + src62[323] + src62[324] + src62[325] + src62[326] + src62[327] + src62[328] + src62[329] + src62[330] + src62[331] + src62[332] + src62[333] + src62[334] + src62[335] + src62[336] + src62[337] + src62[338] + src62[339] + src62[340] + src62[341] + src62[342] + src62[343] + src62[344] + src62[345] + src62[346] + src62[347] + src62[348] + src62[349] + src62[350] + src62[351] + src62[352] + src62[353] + src62[354] + src62[355] + src62[356] + src62[357] + src62[358] + src62[359] + src62[360] + src62[361] + src62[362] + src62[363] + src62[364] + src62[365] + src62[366] + src62[367] + src62[368] + src62[369] + src62[370] + src62[371] + src62[372] + src62[373] + src62[374] + src62[375] + src62[376] + src62[377] + src62[378] + src62[379] + src62[380] + src62[381] + src62[382] + src62[383] + src62[384] + src62[385] + src62[386] + src62[387] + src62[388] + src62[389] + src62[390] + src62[391] + src62[392] + src62[393] + src62[394] + src62[395] + src62[396] + src62[397] + src62[398] + src62[399] + src62[400] + src62[401] + src62[402] + src62[403] + src62[404] + src62[405] + src62[406] + src62[407] + src62[408] + src62[409] + src62[410] + src62[411] + src62[412] + src62[413] + src62[414] + src62[415] + src62[416] + src62[417] + src62[418] + src62[419] + src62[420] + src62[421] + src62[422] + src62[423] + src62[424] + src62[425] + src62[426] + src62[427] + src62[428] + src62[429] + src62[430] + src62[431] + src62[432] + src62[433] + src62[434] + src62[435] + src62[436] + src62[437] + src62[438] + src62[439] + src62[440] + src62[441] + src62[442] + src62[443] + src62[444] + src62[445] + src62[446] + src62[447] + src62[448] + src62[449] + src62[450] + src62[451] + src62[452] + src62[453] + src62[454] + src62[455] + src62[456] + src62[457] + src62[458] + src62[459] + src62[460] + src62[461] + src62[462] + src62[463] + src62[464] + src62[465] + src62[466] + src62[467] + src62[468] + src62[469] + src62[470] + src62[471] + src62[472] + src62[473] + src62[474] + src62[475] + src62[476] + src62[477] + src62[478] + src62[479] + src62[480] + src62[481] + src62[482] + src62[483] + src62[484] + src62[485])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161] + src63[162] + src63[163] + src63[164] + src63[165] + src63[166] + src63[167] + src63[168] + src63[169] + src63[170] + src63[171] + src63[172] + src63[173] + src63[174] + src63[175] + src63[176] + src63[177] + src63[178] + src63[179] + src63[180] + src63[181] + src63[182] + src63[183] + src63[184] + src63[185] + src63[186] + src63[187] + src63[188] + src63[189] + src63[190] + src63[191] + src63[192] + src63[193] + src63[194] + src63[195] + src63[196] + src63[197] + src63[198] + src63[199] + src63[200] + src63[201] + src63[202] + src63[203] + src63[204] + src63[205] + src63[206] + src63[207] + src63[208] + src63[209] + src63[210] + src63[211] + src63[212] + src63[213] + src63[214] + src63[215] + src63[216] + src63[217] + src63[218] + src63[219] + src63[220] + src63[221] + src63[222] + src63[223] + src63[224] + src63[225] + src63[226] + src63[227] + src63[228] + src63[229] + src63[230] + src63[231] + src63[232] + src63[233] + src63[234] + src63[235] + src63[236] + src63[237] + src63[238] + src63[239] + src63[240] + src63[241] + src63[242] + src63[243] + src63[244] + src63[245] + src63[246] + src63[247] + src63[248] + src63[249] + src63[250] + src63[251] + src63[252] + src63[253] + src63[254] + src63[255] + src63[256] + src63[257] + src63[258] + src63[259] + src63[260] + src63[261] + src63[262] + src63[263] + src63[264] + src63[265] + src63[266] + src63[267] + src63[268] + src63[269] + src63[270] + src63[271] + src63[272] + src63[273] + src63[274] + src63[275] + src63[276] + src63[277] + src63[278] + src63[279] + src63[280] + src63[281] + src63[282] + src63[283] + src63[284] + src63[285] + src63[286] + src63[287] + src63[288] + src63[289] + src63[290] + src63[291] + src63[292] + src63[293] + src63[294] + src63[295] + src63[296] + src63[297] + src63[298] + src63[299] + src63[300] + src63[301] + src63[302] + src63[303] + src63[304] + src63[305] + src63[306] + src63[307] + src63[308] + src63[309] + src63[310] + src63[311] + src63[312] + src63[313] + src63[314] + src63[315] + src63[316] + src63[317] + src63[318] + src63[319] + src63[320] + src63[321] + src63[322] + src63[323] + src63[324] + src63[325] + src63[326] + src63[327] + src63[328] + src63[329] + src63[330] + src63[331] + src63[332] + src63[333] + src63[334] + src63[335] + src63[336] + src63[337] + src63[338] + src63[339] + src63[340] + src63[341] + src63[342] + src63[343] + src63[344] + src63[345] + src63[346] + src63[347] + src63[348] + src63[349] + src63[350] + src63[351] + src63[352] + src63[353] + src63[354] + src63[355] + src63[356] + src63[357] + src63[358] + src63[359] + src63[360] + src63[361] + src63[362] + src63[363] + src63[364] + src63[365] + src63[366] + src63[367] + src63[368] + src63[369] + src63[370] + src63[371] + src63[372] + src63[373] + src63[374] + src63[375] + src63[376] + src63[377] + src63[378] + src63[379] + src63[380] + src63[381] + src63[382] + src63[383] + src63[384] + src63[385] + src63[386] + src63[387] + src63[388] + src63[389] + src63[390] + src63[391] + src63[392] + src63[393] + src63[394] + src63[395] + src63[396] + src63[397] + src63[398] + src63[399] + src63[400] + src63[401] + src63[402] + src63[403] + src63[404] + src63[405] + src63[406] + src63[407] + src63[408] + src63[409] + src63[410] + src63[411] + src63[412] + src63[413] + src63[414] + src63[415] + src63[416] + src63[417] + src63[418] + src63[419] + src63[420] + src63[421] + src63[422] + src63[423] + src63[424] + src63[425] + src63[426] + src63[427] + src63[428] + src63[429] + src63[430] + src63[431] + src63[432] + src63[433] + src63[434] + src63[435] + src63[436] + src63[437] + src63[438] + src63[439] + src63[440] + src63[441] + src63[442] + src63[443] + src63[444] + src63[445] + src63[446] + src63[447] + src63[448] + src63[449] + src63[450] + src63[451] + src63[452] + src63[453] + src63[454] + src63[455] + src63[456] + src63[457] + src63[458] + src63[459] + src63[460] + src63[461] + src63[462] + src63[463] + src63[464] + src63[465] + src63[466] + src63[467] + src63[468] + src63[469] + src63[470] + src63[471] + src63[472] + src63[473] + src63[474] + src63[475] + src63[476] + src63[477] + src63[478] + src63[479] + src63[480] + src63[481] + src63[482] + src63[483] + src63[484] + src63[485])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71) + ((dst72[0])<<72);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha6049419e2dfeeb138ec22eb54fa2a42b1088130f85240b760e03c1600cf7e59a27665f4bfa594f5aaf8efd4ec381db0c02a1bff027ede02ddfcce1c78a49a03d2ad8a204028d26fe02689755f9de6617209e7798df5f2330c498aa3cba834209d8e5e3e941ecf4c7d9ad73c0afb95ea69c71093d453a64f764f1663a54f2ecdbf63ccbf0c9a3c92f117fece9c9560f3e67e7789793db38d756a3ab93af991bbaf267eeb0e109793384092801e763b063331b6996843d124367b10889d51b7785ea17320e9f90627ceb7949175adc7c882efb288d8ed0da3225131db8965a469796f41edf52a0670355c5a81455a419b2015a868d7c49284e58d386f232f310f7f94765ffe9913c6426fd6d01bcf5dc15a775f56688cf79f87fe26d94c08331289f93d1251f34c46e467409fffa4a00f79c29b320f6f4b06bfc9d374e89795d21d7dc9015226c29f643605be7b649011a50ccb71e4cd401c27ea37173bb7f3e3bd246dbb852760558ec009eb8a5adac8d0825c886125e007a8c35d275e4cb838dc603b4736cd0cce4ac9783038617a3167e1176a191781811f57f71f0ba28a6de6735b694573febe3aceda8f0b9740b1c6151e43e6b1df39d700a30f6cfed4b37244ff4f219e6560e2246d44e28fa3a9a1f08e84ac3dd296449d01d1622d73bad63a448cca192f8fcbed2c9caeca92044a7feeddda37137af05216362698ba02073f12997dd49839c285ca7b7e45a006454ec362d0c2f92be48bec33824ac542b49f4b591d0c38d1fbf2db894205fc4807a2d7de707c784f93c063a22fe44c77bc304fb3beea5e588e4fad3a608256de9ec1157aad7dc1d877d5cee025ebac767caa510c7ea0d5428b7744108d60901b2955daa2a222caf23c1120369362ae4af8e47231c687355f8b8f35e7d87a6416a9f97a9758e167fb09849b39cc07a9b77a1940ab96289b3e2244107c67e5b39943d7f70dc720690fe733611ead500f4c0d05ea3ea33615169f89c896131b63968432e0eea830790fe1981ea95f127e925a7cdb6df13799ed564ffc16e0c21dfddd7113277dbd26e429953fbc9824e10b1e68e0a2d40d504095b7b00bced09f0f045f691dfce94ac5cb8b5e20d0f65becc750cec420aaafc80112990798bafd21afc3296f13b39235ea21a93d1daca136944f4b35da480a067103faa01cdd5b24c71084fa6898ea219bf7f997ae2428193fc5dc607db6b900e74edc44df57a6e4c359e141ae005a34389193439b45968647af9be55c1ee4c79020c1ea952a5b4415c41c7a476e7e88720c02c1f443159bb922e5e7176bbd04af18b2bd0693149acd7f947631693cce759b3447ffedb9bb0366a1b2dab192ac258d165296ade86ad704dc24437b7f56da2acd3b541ef3cc8051c25924dceb60502834a0b2975e737b9ff57bf0037cbcb2ff35f465a7bc4d89a34e360dd8823e5eced2defd3dadeb711593bd952b5f73efc49031256ac81fab80834383d07c7f05352afe2a9462d6cd70c553a8f5c02000e1050c57f938b0576a9e5b5494d1d43dc108ed77e7769e2c96fc2e33642a6672f38f77035b4af2679ea44db8bf778fd85f4c5708518140aad335e6a93fdb4023f71d2ca908d1b62693b82276e7b07bf05a360814d404c40470f83ef85226a7d94b993b88abd964c1bd848f78645814baf57ec697b45ebcf326c0da6f6d9886356a8f889106fba05c80080ac243ab4d571547d8716050e11b1ab354a9333af5b40cefe535b5c86aca348d1b74a7669c833233d670e3488cefa1795e8745465c0b02bf4cf141112753002c6caa2730b12934afef4d118709e902da84fa8c5744922c67722a592e1e0a6e043147fb78c4eb37689352e522756ed253d037eb3ecfb34b8ac7fbbeb85cf3e7102f8d765ac9552966c94a2684efe1bb9a183163795566a98f40c6d12c5c65ef054338ddb79678822d1b88fbe12ff032370a31b5b841bdb7f5af0f5573f82e531f5450bf8276215363c5bc77b2f15980ffed4940f211e9c0310812d6778ac98c0e25a304c1f05e3533dc0a59837b104cc819e8a867b5e0d64ad6520eec1f76b09165f9227f91cfca3ceebc52838cc78759e9b0b6a94cce67d91c23eb52d59a4c79a964f664a7429d0ad13cc028182e4c2290591a219de1dd6d746dbc64abfc333be7e69ff9882ea3ee0333095e7bf12a7155f909e133af14ddb901b8821577776153060c5b0734f070d3e5cf3a5bea987439e619fa0f4a5fd1a84d34ad85657726c1d6f1ff56623cb59967d792d7900de2cf2d8b8b6e9f9f96e9421c035a11392adf7054e0443ad50c019bd465f88567e47a042645cf3a533ef0c39692554c715201828765f180d49f5d08a28a2ad3b6e3b378186739db31294877261c79f168e2f527919a79043d61dc7370aa9579dd6a2e4e9233ab63af9e98d56c52108e6d8059c5d61c74214d078a0830080b5962aa44fcecbc685faaf45a3b92f0a813cd190d108818b4da9051d731a2504b4d7729482f8d0ee787555572e0d642820cbb2b774865d826fb5b65bdf4eafd6854e0965fed446115ace7c44812633f505f1ddc56b432cfa8e0181b6dafd93788ed3eb46577e88df0d83809071a2f4387ac300f129097b6c56a3519889d2c6fc617a5f8c996f52a9b8c3605549e3253875567ab6dba575c3307cfd732e1637ac026deda410e9adbab04b36192967f337bfc59046e1be991c0c44c2911223c0dc4959c6936c0f7ab1a2707a86c2bad85a15ba94a8038d8eb603305ad99199fa0b7173311f612dc8ca89c5e01023475f09f004f2a22830e5c0f5f01cbd96848944c537f0babed591f73ba798a7fecfd868fb8aa2105f8ac5ef54bcb926afab1a3ccbc3c9890607393173f58cf709d0110bc544a925c3079a5756d64807a52e43df7f13786f02472d4aa12071f141753a71e29bc3371197a75b82cb3e16bb5c4af7a89ff275345c4f496a054ff1fcaf2452271c3e9666ea44c47355792cabbd8f7155c2ac470e569cca0d98e08d81d994a14ffeb2e84259ab1913473e3ed492140468d60765ac65e07bde22773744590f65376945236ee9bdc7d0c872fcec849b069f4e8e87819cbc400e586c4dea36b44ac3dc9025b3c9f5355269a41c58483e752b0c304439414d35c890b7b8ad4cd2786da2f574dee9049e1ebbb52eb108f412ac57cbd9cd6481a8704263d9010ac2c031893ac7d912830d81d4e9d449d863342a04c3a1f92719db9964680e5fc371805b14d838f1316efea59cb1e57b95c6a42874585ceaf7849e64f29489abb462dd371bb46b9524161b5850d7f91a36d4c5b5e36403ab15fff2da7ba6d9f8d3dc70c36c4945944f5985e470ef97d0e5ce689a2c22f513a879a2a9b6d553a9074c441b45c39077dbc50474f39165d4569a9428aad8ae1f8e979f8d49bca9e6af5dc4a45b999286fc521a092291517f8d210496d7d6c06f8dc0e7f3b410b4786e4dcc598c883cfe42812685c1371bdeb7f97d82e4b6538c1df312897bf23ef030f156ea3af3ff1de21d01cc8c24a4cabf83b1f109966bfbaa4845a32ec300b91ff24439160ad326d490aae979c2158de6b5d71dfb15992fe1c66c0ec7af5ba3b99c161cc9f87343f1821bc4bacb585d76a3f3b6ebafea899ef70a43d834032504b6b967dd04fdadd61c4159134c0e1dfa7aae4eff227e51c73aa6c7fd1e99331e9cf6ee6331195b11bef226272b1a3c5189ff3c8bedb6c71afe129a0fff3535737ddfdac4b94b01e82e3ba87771a113abcd80bff35ecb47feaac27d1f52a9e7b466a0faa6a8d2df9253e4f8ca0d9f8fa1c7e3bde466ae6b285e5edbc11a765b13b778a96da05e7136f10e8c212a2bc23f6a6cfde8f0ad763ff8b637a94a39019997e624d95fb602fd42d975a54463099be2176ed3ed176be4d655719140d93db3247b60803e3d329aba4dc076f6821600a8ec511afbb173a497837a2d85a71fc4e3ace56bf313510b7752a133dd580c2d6cf5e5c3ba37c2bd2d8c5fa6ff2b32f9865ebb25281c07bab34d4ebb663c84b4cc2ec22fe08e9449503e9226c9508940664b73873f46ea75ace9d2319d4759e4e69a72e1a00494149d3b2d302b965b7a43c9bbd75e2d0551431c53faa65fa36e7ae53c3d80463d75730e22b05f95ea80b1ae0c3283c3b49fe937e6208e3c3d98433d31be68fa89dd4c549a74093456531eeeb248cae3d911fbbd1a9ca9c9a657889939f3af6a09971a5aad21735ef913ce0a96aabe53b8f540d6231f10ea2044f498eec866309b6cd16613d98ee7770cca306e2fd470e519b8fb2d3ad22bf4a22e5dc8575e96f760e1b14ab1e29626553221a0294d9f090aefb3a1961b5aef6f48d77f72c0c23a81a1f8a77607abeadeaf3e7a782e4a0382fdd34d40fb902e565d4beb5c7f153ddb57057163a62fca64e25f1c6dac3740ddd629d481e49fc0a3656ba1d43b75877ba21c4165712a66f78205528cf41651bfbd0b7bc2d45a6028682c18a443727fb6e41393f7074d31faf79c330320ab0c8dbf75484f4b41379c3010e04d30b8270d7338889fc17bb84db47496112dac36292e2b02cba097c31f2297810ba6702ce6fb89aa48eb37622aeec5ef46ca3b3b8e72f0ad97deba02acc63c79cd442868ddf06c927c01575a62b012b2c6197ef893d1856e572fb25128d7c1866a18b0ca46c87e11ea3d4a07ded152a46fefb3dbd78d7b914495954f4f1ba4ad74397a353b36b146c9eb1605c6ed9ed567c367c1982b7d459634ff5ec3f4d4ff8aae471df57a2764ae69fd2e7319667a41eeb4983589e082fb2b10121fc0e78fa91b5a1ffbc473065518d06148498110b8e9d0b57c79500db13b2b94401744ac01ff081d05e61866b92b27d73504e0b2a28984b3f85dfdc58fc3a9d61c0aabff0d244de8229a1a49fcc4d66e86249203c132e550887d06f780452d1c7e9b30a4673450790a9c9c8dd460c0e3c392f37faa65e880acf9734446f9d9b7c22ac6cfc15c3b0e57e36f263d522dcaea8c64c2ca1c859c4ffdee66092e6e8736161505bdedd3df4a236d868e44805f5690e7618a0d331e94cc523d8dc48a90658af615f1bb774eba82ed3d76d18227c3094196dad7c150f10494184e737ce206d9054070e2c41fc37fcf8877ab37013a3fdf9546ac065581911d7b8e67af1f10a63922f706186941ef40a325bc497504812452a114ed58d0bd07aa0ccc896fbd2437c42f637aa0122f1a2c80babed44ceb633b0b7fd70c1a87fb7e409bc155277055d04c522ac518c71416afebfd2eda41b4a5b7878318c5b3a65fd40c8435dd75d774dcc59cebf572b681f77fffea2d66d08b562aa3e842d5db891eb668d5272dc6a40f013a0e3ac0c7cbf7c9d8858874f912ebc403d16f1ce33955f98cde7fedddc44eda44f2204933248da1ec8c389dbcec1b3094378d4351993bf0a90ca217cb56f1296fece0f4ff29be55207344c86a416df7b6c7b4e73fc50395ad73a205c94;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8664c5cba7164c66092663eeb546730a2cf51504667cf512ead31934d714c39884b40dd9a4d91a23ff3a07d1387c48139e5ae32546e92d083a5869bd132c495f5177e0d32ab69a6141cb7a987560b4c872ff6c07a646680e9383096dd71e31d89be2e887ddd27567880f77bf2c1ce23382863d57263c3262f8f4013e62bad2033fe0cc20ff97766955674f06820d29b3dfee1e4e2e4109066ad0ffb35cc8fccf9cbaf323f604aa6e51e58556656c2b178c5330c23ec4f4db37a81d3508259e079e2cb08a3364ed45567ac6775630a41b7e6b53615342c370af79331f8f86912fe39f9069fbdd553039cfa8d48aab8e4973bf6bb8e44f342971f64b43429252b55ca0bec2e4b5dbe4fb389de5b5fa330f5f51b78462080bda4b1c3f6ce99e8ee4ba2c75c0ce12a64f917df8c6809e1289e44ca02b5e3d227488caf88e0cfa681c56b8681fa7ba1a0d1be4b11a7834706f2a97e6b8c12d064ceb8dfb574971ec6ff00357eb6e650fc8ae3cace3d97cb3956a77aa895c120b490f91eb2137c1fbbec66c2eb990eb3a2ec5c7ff42e3aab49af2e047ef5d08c5737364f0d88b9bc9fefd7e692a2b3fc9a197a80ef32f705cd5ef34c29ee02e2cf826fa29121d3fed20c107e1cde469bef874d7a7afb1f93f8d17ccc3bf7a33e6d2f93b11a30e012b90cf4b50b381c1d249dd040902d12b1f6b1244b298a8ca8424c4ba47133dd6799e79b3449a3fc029e7df3f4d5b4b7de9cd0798f3dcb513b6f271f1d36f566eb9ae5a765e10f09cbd9e2a44d8058e5a7930ffac29dd3ed9a1feb482bf5b330ab06409ac15a079eb442b8f55b1af06f8f2cf1764758b3ccc3e5a31164677ac827d1179f660239b54bd63d907685eb8aa193b501e56107a233e67835acda267fb7d57ef44d35ae3a034086a298a6607c3c9f9d5328c6f2f2777da2f8937db9e251a400b8390b586246ac7614ea9c660271b4aaa3343075b6cfbe407789c0211dc307068dc177058c7ad5ea5883783582f132227d73795e073fc369cb0f3bd6ce2a39cdc17f86f63d45e9991cf3527366bb4b0e81c4c272687a55cac577f8897a343c4d0b2d62634f7ebfb39d4df0b585e47ab17559b28e71fbf129b2e2c81b1f3e69cb26e1d87f1267e6e3a3e69a8688ffe712cac552d97d131f1243656a4a7d51cc58b44a7780579f31b83e247de0c3b4b99f2111b8645ce18f8f90c9101aabe0a565695ac5c7f2416b2b1ab71a7bfcf13af0e62008e012d6d007841f9a228476ec0604270c2463bfcaf0d79dbcc4b4fe82ab6ea032ae84eb5299cab49f0ac68130c73c348af76195120a10f8ea75bc79654c330f5778a546476a6156d71cc5395d11c9ce17581b9c357fa6242372ebdac901fbc4f59281d4880da5755df0bcabc216bb89b4578bfd0116e2e6a5a8af20b02acab8d79fff2b6a77d34c9adcc9b0b25a65d6519f27d94b71781e8353ccccc7e47827391cbb13e8069126bb000f9be1a3f5d6d182020d80a9ee67000674d7e78a95f5e1aa09dff13041b42148140738e2e291daee37905ba8bb8c47f60c03483e20026b41ea73d4cb03e37b929eee27321acad98c2ffa2c50adbc248a2a24a5739f6e521dd6cfe3b3fe9a1c82e5f115c0d4db7785476736103e5c19c09f4e4a1cb5c91ad98754cd940d12bf369e0708fe2d853bafcfb14621225725b027422c70bd78a9874f8f3fc7186d1c8f13c59c43db01264220648cb14a1fbf82757f6ea9df326fbad873beed605aea965834b2b6e3a6114a7ee2f8e8deb360b376d68b334cee9f6a3286f33b4c925bb698a287bdfa74d5495272b030bde09ceda1ea46490260645a2954e4ed8e19b63d73432d1fea85d46055a27b3337f4da8cf844eb1f8fac625a32194b88f8aab7f73c0a4a0d967dcf5b203777e3376dfe91048c3943118e9093b79821ccbe712e4388f67886da00dc16261742161b952f084ee8e1b1b8791c387dba08f41b46e43d70f1b14da1e30c0dbef54732c7dee4add56ba79627050a46af59f899127ea5a88817043790427e3b0a45f725a3d73a4bb370cfa159ad54200b1358c5eb4d8556bd86d97bef9cf1ca042069f3b8aa2cd80b0b367fcf7301848986460329ad716ca28d885d994d68e3b77f9e96ec09f49bc809c7410bf4639a082657e16498b53f03458d67f6263f805cafc63987d35b6deb66a4cd1e27416b5409b0ea4545e386430ffbda414dbddde8feebe203760414361f46fd365b393e252d4421404f57eb99076af6a6901ecf452756e9db767a10ccade7174f3b317f7f74d7f4ed100cc932c91d029dacd55097fae4d585e9f06ff30326f05c4c63005faa9eeba621e88cb24f2a11c82961fda4d82474d1f71785daf15e1925db1c5ec5932a01d83251ae5b1bd42725b9c3ba9de37b69adcdcd58b57ecc6b0825f930e619df207031d97dae75ec56aefb56250034c2328f73188c57142b0a696041f76d8cd83a60d667366319b109def6e19ae90f256e275e5f743dae389066b08d390d55e7d20f823d0096c207105ad0f648b57a3bfe1ec5aab999fb6221f7a884c1edb4b8946b7207ec9933689f6d5e5b1997e10c9c3476bfcba1f8c3071e4813f8edea54f413120f18d64a3585484e0b7a0c133bceaa3ece196d6216cb0f631df2092c32a4983bfe40f28bbfa749c14d4a2e1d45f66e8abbe2ee2fd80734675e8e72d83e65262102f666245d891411ca2f86d5cf41ecf99b633b3f8d5d1e4d3beaca019a42210cb52ffa181aaba9cd5b570767f08bf03897c71e4903c5aeec30c5829771b3a19dbb2f25f9e9157c07085e2282a8bb525675e69ea51438574374fc48c3d453fb1571afa3a417a7bf3c0e4e3fb4b30f5bfa9783fd415b18dd4dfc09608c75e2a52b07989f7005e4b84df1559d5d0f70fdd6b2079705095ff13e621cc925f0fbbfe1ffb78a9dba7549a952f513bcfbb569d2e52216a58e1651b5dc0c875ab6fa572fc0c3df9c1571e64ea38070a5c322fa2d14d5f018ee6c4b11f94397a9c7eca3feb1d34e8cce54feeb0986696ab0d6f3071e5b1122628742d009bc1cc80f161ee4400c75e98a2a30dd1c2b0caa27202f5a594130cfacb0de4b69f31faef0a1872872b78f7e72fa30990341832170d50664b5629851d23c433f0001ac0cc5e629d8bf6bd73d3ce81867b7b35c5f4094a135435542b4dddadfd5516d9ce569646253e4c83019abb5fda0904f02978b20204f9e8a6b29c7afdaba8f3484d83afb9477946f256c553db5fcdbc8672920650c777f25549dc189b75bb761973e3e8f28d6e30900c988f045404ec877801432a4b113628c198f9d365d373ce815400fba4a1238b399af0470b828bae2f4c1e3114c4a7badc357d5891851c2727d11cc6800caad26a7884fbcc9328a91ca5d79de8e978f0b6e51b4c73cb84eaef3ac65617653928801b5c61db3740907ee37755cfb42fd945309e2c52b5ec134dd5500b710af3d284cfd689dd5e28dddc427aeba164f4eed4b1267ad12ef100fae782f39c7286ae3b5e4ac23a1569ec39ff34c62a5109c780d63ff3eafc4db4f2d1705fea8f88791397671db940b31ae403c057298ba88cc7f64f6dfb4e3fdd624e6f87c59b944fa3e618751bd7b2b9a7f4a09e960b02b056385117adb583f13cab3a0bed40f50a958c276b8792e0d78a8cbe7e83d39a138e3e88f2835275ed89beb5414e2622a0883889fb96109e68dd66c385e973e1235c5567e4234328e5f3b1e4b68e7638838de5af5c857265899d56c35e90af993bcde5f0abe1ba64851841309f63aaf584bbe44af8160ac792d7fead041a97d623bd3288927e13b852745979179ad107415c1627246e703ecf07ccddc85466b77db85cd70e128334d0c577a6854834280359cfa9df1087a2ceb2a86100c79acf6106cd1c37c0add9e3184628b6401ba006b7019c71dc853b37b4b25b9dd75afa15e0ac8c4fe8311c046ca565eab1e3482576e5d3ed455c8acf58769ccc59938287b86cd0fd11dcecb1b4817d24e0fe2e254a17546e80091abcb9bf8533bdd5e848679f82620e25631897c03b2a2e60f7349634b49a456532a089a1923edf85f210e554bcff1a646faeca3de8b090f06803a394b1decdd3cb38dbc9653de120505e8d7537a4790ea03767ca6e2a9bc003b623688f03e98f32abd37dd68ba5cc2650864b7d0926cfb4bc539a2e1ef92bb1de9f6e25db2667ff0522262f75a43c775c3e9fa00d498271abd9510e79fee0919f6631fff62d29471df158bd6640f292fd28c5ebb7a81ad1196455dab64ec6bcaefc444a76d0a78ef068a1e0be603cb6c74a20fd455a6603d502dfbb09cc2ae0fe6db69b969b9c5d00a3f0d1c4d34224e005d5bb1ba327ec0ae57ab5f43e330d8310d3c3e88729e02c6d8f0b8840e2a3886ca78396efb4b7dfe0f6b36168f65a50cf1466a99e397b5ef4e858764b435b354220f5124a3196ee69d1d24647d888eab235688f60d8c3f7ae44ec516bcaa39ec166a235544bd49f432e9c80dbe1b3fc3d9f86448b18b9c4af6dfe5b38ebed8f39ceb9d2debb24313cfec8fd2f0eb3e993f6772c5ac35ff9fceee4944d0de676493983869bfb31242e630b7a59e622f5ac1f789d3450e4d0b02e2e55d830fa7c5a7931047716fede8d7027aa9baab12c997eb9fd38cc6633b454e5a5b958647eec094f20a6c403a430ac1838677100612856d3f745f92f99d3dbd3b1bac1214b3bc3f2919ecc34535c49360771e9fae02b4c15fe2b6efd4e485d986adfe44128d713df2b608cd120541da5da65d809e119dae9b897bbd11d3a64861eefbb6eb10e81388d2cb7b612019f0b98f05b4a4576779ed2eb77fbf6690630a976317e51b22518c5e6c5019f5782b7156b0f5115dca8725865b02e2d554517e74574b45cac17343ce58a43c3024508d5251cf49bf5b9c87555d0daff1b50bf7f3faf4f6b861ed4cecb79e0d019d79981680dc43a2f4c64c9f8c62123cb6fc1386614ae0c666b6cf461a9e426484dd12b5fc075591941d3715826bd5ab6d37c87f03c50c7db56609b4b83d134135fb0fbb1276d5a0e35b9ccdf74c8977ce022cfb17975d0f3542ee451896f86a689594caf1306a35764bb104bf19f138462a58e14e2b2042a0b666fc482580c1862e75368e8e2985931534723777b3c627c169cea3399ebbbe7929284dba900b7f24962b8b8aa982101f45c4d713550d56bf45127f0dc4abfbdb5924da2c7b995d7d78c17775967393b13af08042696256ffb503870d5593bcefe9fafa8b2acb19bbea3443a94c7d5418b9246725bbea9174c7ba4ff4eab74013c596393a8a1780fdfe1eb261a30c3345a664ca5d89c125d8df07fa8a447adfd57db0670e81d7a46f9fbc13e45f0207dd58b7b840cf0e3320a3fd752760a9a02b4c9c2f5b7496e90104c138fc6ed80c78530fd3702edc10d5346ce61a7db76b8b5f8b049de79df952e2f55e8d07d3cc1a2a1a5fea842ab84ee2f062b3d9e2179d2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4cb918e8482a4efd86e99e252d29c2465f7d10c2f63477ed15ee42718f5f829a4a30060dd7575c42fc4271d17e71255ff84a1b5120020512f34b9868fbb75cb19a69a02b0897ec5bd8b9a491701e0a54d2416dd3af945c94d7416328622d2be83177663a412898e88d80cd5ed41f4feb982246361e86914496368ab4cff3e60a1fd6e121d51530155c04bdc0d53715d1a9d4e9ef21e8c86d06820c45d3838f06b05974c950c2632be96c5bd0a41af91e13cdc322761342ecade0acdcdf86e6d5bfd036b6b7663a630636e1ec37269e8d0c67c64002642abb15ceb90a8117f9e0c9f6532f7efb362381bb45b7b0287e9e5ce5e634f138e0195df0c14ac37749efa936bba1afe784801eb08d8f195d64b0c3175feaa905f43b9e3289fcbaefe314711d0e5fba37887c30785b3247e3660ec2c82cbd1adc27afede3683a6c43b2f432bafcf5c1175668eb4c65b676b9ee5781c2fb6d1232feb83d0480e6c762e1bd92f335f13d668a2b8c83b857e6750502e848c84a783d6c3b1665fdc0191ff9ad545a9e360c6bd723177b3ea20e57dd856c8c083f0133f5fbe66963eac018ea1976540c6a75cf16f2bc25297ac6b95d3ec2d32a4ddad4bec70bb8f4cabb8a1b3c970ecfc79eb576521449bbb0b996046330d70106c55154afce7d98dfc4d0baae3187a70a78018ae05d55cb245c61f3d597f717f83802fa93dcaf0ac161eb838d46a081d3dc6185d596ea7fe906491bb2b3a875af654bd58beefdefd9535dd1d2ea5b169429ce8015b1e5e6c776ca6c0f7ec893568bb382c751a3161f4c4bf2c7b74c96cd66a3c258bf524ac6d5ce09e46505612a4c50314a9fe09f7ace93ce3579dee3c6bf9111e93386a81c04685c377328a80a267d1a814c02d22b272cb4ddd02516e3af13e2f8a0228dfaffeef06083ba015628e089f3fd4d58684944f0ac1c6213b224b9347303a794c322a4f144a5c5f44382a4a7db5976acb58f818f69f2b1bf66e90417de516eb4fd0e087fd88c63235f42703fceefd0dbe907b1a40eb712cf803e4d3a712622161b950c36f46359aabbbc1bf226af010c2613e6ff44f07e92a11c8530ec80f8d44259eb4a77509874310f6076bb974774e386a06214a892f29f474b318aa8d090d6310fc74b6a445bb04775abbd10661cc8ea022fdbe3f8c2dcb906c53444d4a197a828630cb6915603bcea414cfd616861a96801d021fa5ef99001cb8aa6be8eaa556eda0742565f2b54ac7f76a9f0325bb1a5028985fc9d8c32ca9f28ae1b38a976aa522f32ac1f5be20ebea84404915d77ee7274169a006128a2a7feb0caec458c34ab74f182fceaa2c2abb803215e4d4d75871ddf72cb4d9c0787c3f487f1cd72057f06fa022ff18a6e269e6f7fb12548479ecceecf3ea1423c4bc46c9d4891246831944f4e99ff9f0d783cf654efe1c56b2bacd08e6a0677d350e2a03026abbb11a1e358288957c649c576c2cb32a2b19fd1d40edbcee502152c616aaa9246380a4b2159e81355fad893ad2a0c1b465e03050f07989ee80f504588dbce16dbaf2038633841178b7e95f3fefe88f3b0e89d9a5b09db98bc46395dd4a7ab4cd488bb408ebed0d6324c4269563abcd87d03e07d7ee10df86090bc2a94a19ff04fbbfb479094309086975c87e3602f11ed06ba3c0814d203fc0a313c8f3bd24983fe2c717137fb79b0690033384688cddd666a44c592a1d1e54b3afec1c188d19ac10c80c55bfdcafc2442ff1078ab86eb871abd917ca51b2d37117f3c24a9070edf7faaefad662d4a14411de393c5cb1b53dcdc0ba8b7a5084c27447c24995bcbdacbcd51b84236202eb7d47bdcba53d47b3f43def0fc228b98f1d3fb7ee9c48eae5e6f5e1115a92a0c0f8134a702a448ac8161a63ffe5f6fd14ebbba98afdab68b9f19855c3a4f062b528aea67b31a8f0c2d78935ce1f42ec6ee304df60540ac94b937faba7b9fb6a2044e68a5981134e1ec93be624df0c8c44c4fabf9c1174f58516077b987e6bb53f72d54021501910acdae55b34691b4eeccac18202b8737dd614087c539dafddc4c27cbf9e1e5f2cc57211ec71cddb082432335baf0a6bef1754d7922c8c58f1a715f07243f479ec08c57083a7b6080c85613069aed13be95eb1b2dcf94d978448227c27b555d9108eb80efbf777450fe88fa472d15471f4f8296a0bb30b87ee54fbcadb8d4f7cfec9e2bccc0fd035fbc6a394428a0c6e6cc72e3b61611532c0f8b67b0eaa8645858e5c157992681905f87b6251fc9d3652665f23dc0680e58a5da5fe29bcd01275e03792ff334d211a90bd1bc04e209f933bc2b1397466e6a5acbb3ad8d10fbd7917995a909dbbc4529a8eb9dc7d06be0c7779fc89bc1617efa7a889196183972d33ae7dbbab99aa05edfc0bac8c23ee1ff2d9e5407be578ce0e79ba017bbbff46656f62e7fac7f53cff5938d406a00d7713c1fd125b292863b7ddc27a9ae782434300acd3b57874da1a3f840199316c4f8c8987f1bd7295ff163dd6686704478bb4f2be7db6520104a4077a3910a99b4dcacc58d4b7007a33b8a320254b544fb1b41f4ea9153478e0f9600c9a506fa21e10c76ce0dc22a315e089d938e18df34a8c7a5d017ec85ec6faa18fec73226d77c4eeec43a2a2da25edecc8861161e8f8ebfa8e1078cfca2c887d5482d59c70979f7a7ddc6ff2a93147fadbfc5c312c013eddc4027753691073417b7d871623f1bf2b8b770c0ab4ba3de61a7a90588ceb90416a5a12fb1c8b1b8965720991bf6310271790ee2010b87dd47b7a0a2734a7ef6afda23487eaeecda08dba2b6bda2510add61393f09e0d0322253df9236d03f9643559476f4ad17ae9f3c20ea00b06839c2be497bf9a9b91621f68f51d1fb53bffa469294c6ccc43d44591a76d521baaf091f8809d820807bb863582cd218e9ff392f9eda1c740882d7199e1fb17c1cc00724c3b70a7a47814d8cb2a6b3f6f9af493db3b345416fd11c83226022a02709f9fcd0fcb40c992314f90e27bf39fbd936e7d6bf0881df3e007121dceac35d8789b83074d8af011ede4a60071917988561ddba1eb0f05b888b3dd900c6ddaab7fd2ea2b38d0d4e04410a064d55791c906c7f7e8c0e807a8a19bfd67b6e5ad6e634e25eb42337c27506d15264e04ff09a5a1418f27bd395b81b7baab6fae7ef73903ee6b100d72c1ba1d0eef6f6398fd0ed2532ed6aec1082e5d9ff32d3c5cc321f5552fa113b33a362202d3f400a2dd4cb2be38510301b418d621d9fd6b34d2f820329beba7382327fa6f47c3c7ae456000f16c7a73f14702f72e2bc68830604852b0e746379034d343e0dfc1330f1558cb375fd4e6d0b9302a9bd0a9166898c96a86972fc789b2b3a94ee34faefa93de5bd8bb489f0dfb6f6ca6ca179ca60466498def0fa7ca1516e2a4f49bc7af32b7c5f0bd38d499ba97042968362b3269c1f8ce71fe1f3e8452fd15ad7373e22398d7f393ca30f99bf619a2bdd082b5c7e8528a042e321067c313a7262e90716a04eafb66d53073a19aefd7b5adc7637144ee148daaef9ba0240aafb44c6a55ef6b5df8e57e8af31d9de6551969ee99c8dc625c703d1c6f0672ffa7255f174f7ffc512979150fad112c0a2a33b781d63a04ac7d05433d380cb6b471d77f4e43db2c3bed375d853324c4d020bfbcbce65194744faf60c2e8fc22fbda0574fb7e9cbf9064b40cc58ef4e26184363be52ed898da2db226c404e8ed020e26c548fcdeef0022a34dee5cdca59411a16bf2c8460b2366345fa9c0f9a1b05185a9f3da79b3627d76deb0bd70c173620bd871103f708a44aa4f8eb73aa3c3e5c937593c47fa769f86e663ea78f6e4fb22f668636911fb23b2e462322f2d3b5ccff6b0bd70e25d4457c57b9728dbc9e36a339381ec6ab22a1ad2b0ff8728e686b37d7fc48832af72c47956f2633c6b6857b7f4ceb54e8754d8809db3a4bb989f47dd634c3b0e8d7a0fb7662f6fd8ef49258cae6864d8695ccfc9c4c46c1300e32a412b951c1f50b68c1fd73518593e8b34618a9a508fc8bdfe15c5b9a0a33c9384cb40e25c0ab77858b30f11c1407427712e1824019668e0b8a34f7d2c7585e3d7ca6880bf5f9822a68ced462b63336eafc831d2d3a50319ff017aaa7b7f0e586c970b52b61ca95adcc4b9d21a98ec07d5dcf8e420ed6d539e96a21dd15d0a871faa103d3d37c8a46dc92272bcfe7c36d29b9743b67fdd86fd6eae41963b1ef608ed621948bf112123e632046042cf41aa800c2c4ca9ae6d9c10e9aa109854aee57f4775ab8f8955c5e85bde541ef9cfab5d9c35f42221dbae18d13cec2e214e1d4b8db087dacea115e604cd5ae45f8533791d2f61643844302c8c11dad25c8c0bd31861e7962d337e857481b60daf58d559594a4c5b7081f31e6782ee9abb40f1fa9ded382b2a7540c209e8f5108df7607b3d1894df0e66cc551e6fffe3cb42a7ee57882c2cba36be0bc128c25bb785d14a1e97c1c53bf1cea6dedb059515d3feee5c79296be79cea32e01746f83fef363625648e8276b2f70615231c33ba54ae688ec67052a300f4945738458bf9c1a39b0472d4e96e600853614e67047ada6c143e26ecc31645b7a355896c65257343af57d14376188082f6950f0bb8bd15afb02f69e1ef5cf5d0040b76aa0d3dff80ace26df1ff0728caf4e1a809770679fd6be58d7f57e040ec6f90e759be0405337884c1993ff3a6be65cb75b5189f677d841a24bac5a6cb31aef14e9976e006451f4643e6c100e68f67394fbf3b7467d0d2bee56933b9cfbb15226a77f5e52941fa9b2bfa5267dc31f8a2537c21803127b16c16432c5986147027f58d6e07899f284ea50f702f8a575d7f16ed2b196da01eb36c7990a79aaa2a4eeee832494e7ce3a69b942c2bc87e59371ca66ba3e052e024f5357df3061447b9f460096bf774811ae2194be4b5ba5879c6b3cfbc036b0c1061b30cf82592c6803a21ad4e9e410cad5c41624e52d9d51ba93ec9e3be9ab052def9d31b2591899699b97533cc584cc62505536854cf346f22977059fbec8c3207f0b798b4a5ce27142a9ecd65a5d4bba5b8374a5e1cb4b366c2f941350cdb7df6a3d87e9be3d49d59c719894bcec66360e1486db4ec4ebfcbe23e8019ab023cb16f3d9138e34b0ac0558507d24e0c95005e5b64c48e8b044e3d1da4af2b7b3965acba098f758a4fe8ccfed1621858aaa98f4388c1ce6d7936d58c655d3055a9d8a96dbc2bfb4cf14683c168eb0e76546d7e8ec4c6ff5a7202776cfb1fc8dc2f6d6895918a0564d13365467d4c340498fc308d89d3b5ce0ccef3a6ea4e7ffcbafd9b5463289ee74c0fb785c12f9028ac090bd4a6b8da3cf034565d684740c412873492b1fe9b0024453e6d59b836cb877aa93659fd8d31105f77e20f67d33e2559bdec18119d9f9d334e26a2fb8b521e13d4d7b605cd73266a4ea151df35c616747ca277f671981339d6b02024b3bd37eb9cbdd8d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h93e674c17f8743b3faf16edb055d9c55960157d71f3ab7534a6620f7abf85e7f1b3e3baf530288381fec316944cbe6c27e400b71988f1fa0a59354729bc2905c52ed7ec3a1e9fbcc3c4d6d6b30e60272c9ea164da903ab1b605a1d1c9f7909b69f756c595f928221e881300064ff0ec5c7a716b2f1ff8cf68c91badda83c4436cf3bfcd8737d305873f0c6ddccf2376ff4508be75e5cd154994e40ef4f691d4e7644f38518e99500b40a27a5956e3806c12cef9e74942044c68c6b7b1cf2a51c11d15e685bd9e1296ae339967f5214c76fb3956a981d0e0b4df0426295bd86ea9d2819e3f47d56711663023fdc403afcf12504201f8aea67d63093f48ede0cc2dcfd4e8cdca2f2b7ff451326802a71752d002b896d82cbbd7fd48ce59c0839a674e9dbbd7de6c93d9b57a1c35ee437d8e57954734f29a13e048f73d1d75d19a72a06a04bf0a6f736e2c43731d984ac3332cc65aecbb569eb455045f966c9a243462c54537c1f1d6ef9583a7776e238dbd33f855d5e71961bfe5297456795c45e4bd2e8bdb1517f5d792aedcae6b785ee6673cac2a82d3b9da6c8ffbb6c6cfc7bf60ec89602103dfcc3fe35185be529f5588a36d56fbbc934082d82da321009f6930b4c4a6a18746f79482765e41e5d724b91f353b657095555c2148b473362cb45cc46cfcf5efa8441994af64e2b96bda01621e06f79c49e5346bb0123eea6e56f74a55f243d27c0bb7ad91947cffee5da4841ec24631cc48627d514e6f69a17b8711c266b3a33b3bd1993cc585153100d6c6b5c84ab6b2e802682e8507a70d50d9b220634aff006e11b4068597b59c7dc0c44d237c8fa02d9f603cf367b1c100b91cfd5fc2dbe6dcbe3b7bf7668622c1e7dc0f7c04e6f13035f7e79d10ad769e8a9f58d6b0f39b6c30423ad3f3239634410f20e422498b1afe4868a3b5459ae765930d535fb6b3d4d0043c04ec6dc0ab1ac230540aa159f8d51dde4864a75728d17304ac8c47a97804ce3a785d9c56555d48755f5d559004207b59be64087f27801771322737c6a0c115fa033fb6be562d373304bedf9e01d65abbd9b7359fd5a086c972c8f355913c56e89085bb01dc40a14ecc73387f58119b82c2ff1a2997a4752badb700b13b5f44a731017d7a2612f77b3cc7e4c49984b5948a529c25fa21fd7e2fca212bb97969f5e4c818a1669c59acc9d908187476f69e6b3fc19e01b87464477d3e576e0abd6b38378eb8f8dfdbc538797f66a42a507bdd573e62672aa60b45c5c8bdd32425d78e11ea0b19e7731f20a02ea995a8818cb9d39df3646f639418bdf051bdb0db11ee88ec16eea9512058083cbcded8649b06e2b18fd4940b7eb54cd9fefb026802d4040a91bd0c6c7c264c4cee3b54d6e885c4d3a526fe6cad86e14110d34acfe62c35a03270d0794e97db3ada59d046c89747da0fa3f107aa3b453c04391898548faa93f325c73483ec941bb47e9b8a9eefac5d1b2f0c73f917a31ce1a5779d4da2a124ee90e556e9934e0969fa7f971de1f473d50241b3b2c05ec66f7daf0f83dbe29b616d8582adfe468bfe838bc9f103674d74baa94567f37f54dc71a9d22161f1823edd0b0812fdbc2eaedfb8061f6029f3749b5adfe0ce376f302403120362320294316a4e58eadc3ede284a32993c668445de624572fdbfdb216660aec7c9303cafab1c978a91cc2f755af5f3f46e121bba540f5cd18e9d01b88eb106f0ce7298f262d2c7d803f7e969799965115c37c1f5dbe1bdbce4de84972f3d82d83dee62ea932ac673d62c7faae0f0da7f79cb7dd2b7db53f03757b61590d9a472ced91d8f0e1485384964585159c6d65ab0ec9b1d4780e2b48cf5c68edd3d1be353b0e78fe669fe93fd94cf173ee1585a5cdd905480cdb3f2c967793e1ab50d36e4143d8a28955547b89320e06b0bde4e06e1623a6c68e3c032c9f69a2fa1a5260609efb59cfaca6620c4ae85c874d0b8081e3147b05fb118de26589b92d647c16206e393cd1e4811be64b0bbe28e6a0bff57ea48f2051e11dfe335396ef1842ba76fdc53ad6b5b55494ae2d9443484b0093e18c271e9bf294f51a94f7dae6b95ba0d861ba4e96ed71bc40450ea12e3bc26ddb28d59d35ba56fcc8f7be516d41000af03c15a77cc738a0c7914aa6d58a7ca961dff3c338c8c52910396a2aaab84fbf9d803abc1c597e83de5ba2546ea8a8bcdda4ce4976b07e47f6441b59d1586c394b21af98e934673d1a07a671334a9198ddefafbd646eacd1cc9e81f95c622d6740d96ba07fbaf1bec86fd955528658ee22225755b94e6f5839cf7db5949137e42fdf7123dbee43e89b4bb5710b5a3b38887bb725c967dd9ed4803a298a493175a3434c3b61f2d1c4ad10f5e8bccce2a5676c8495fe7ecf00c1a716cf0e8a1116b7ea5dcc990852ad8195109f0e2a0bf3316ce703ffa3b7a74e863b4ce3eb79d6f3fc5d885f54bfb15fb3c8c16deb3c9399ff7f1c052d531f2e2a403f84fe3f2bf346a4858558d6e8d31affebf0a455b058f612910f7f4ed481a5057f5951101e198ef567001ffc4a9f6ca1808dad212ac39045e98c2fcee44a341f4a0a18e31eefc98f53ac8d9ace937a7348f1e5ae1b65806e38ccefa422784ea2055f0b27b8dffae41a64eb4348df9b1ee8bd8a3daa8d94fbd8394f2d3eb2b761729a08f8d78c6388b152b37e160b3e111bde42d3da42b0a81a965c3bd249a59fd7335464459755d30944553b19b04ec251ea74065b419bcde49d408af5c5d4e604edd0ac17716aa22b89096b9abb7c722f4fb5d4ded428abb605172329e601c9df9079649f8b6fd4aedfcffd9e433310d239a38b5699e2ab56975d1a3805811e9b07ddb231052497c476b5677f3ea3035236d8d8d68caa004055c80da45c5bc9dc722275a029b2a425617d81d2718dcdec50a07d8c4595241e083f49700d409a672915a1095c1ddf8547afa797955b6064669de30e3c9ee93e710192ff5c6818fbf4de0310a9202e2c8dd300f787f24365fba0b79c622ac50467c6689e134ce040e5b66ea2ed24b1067b64ee43d25e98acc990c4b19d4ee19e3a679c095a851dff265c246fefe23387a00c9b651b3dc0e420cc25f1e04d711ed8f29bf602eb48c9e061291129cbf5ad3cea01b3c3465e1b7979af727679cdfe4aed24023d1ce0ce8691430ec59b5e6ac662110f5f5166ce407f08031ca4dcdec4afd63027953449c804f36a3391d6703c98ee227438ef5c27098f2da23008bacf14405e6ac9aad696e754a8c8a0cefc5dfef8f2cfad323ff9d6a0475412fb1755961f5bd6b673642a71d103cadedb0261e123a5ed3266bfa5602c20cc76173fe0a369f2e77d3abcc2b819e782084d38564d04a21bae4c7a81c59d3a12672cd0916a0241c95a415c1548773d153d88d16c78a100a168ec58327a9741d9c54dfdf3117cfebbda0d28ef293843a7788be7a16ac1080cb5ab2f0ce1d57e69e3181bccd9d5923d2093bd70fbe8b92f29248247197b97b40914044f0c13a808128da56c0421d5993f9a6192b6a15348c81e61feaa2fd1c3fee6fc30e22605b924b5644729a16ce239543df8c72f70d0a19938970e5535c728e587d49c64f1c96915a7fea875e39e9a2164521234a9eb2904b994f41077ca80f604c879e24b4970aae801b4c9963e5e4e6df09199104ce87c51d5752880ae6377194a6867ae2f3c9742acd6606f208fa4f3a423dd66cd39403d060515d232114afec253025a01bb721e4fc97e33852e600a51127d35b39745e1738e58b203653b8af0dafeb50649d38396875b747f8e26b7c131a82e3d903c17147ee8eb1a388eb455137dd922814cb8f418f46f5d16a3b68e72d6c0554f088e38bccb61cd832eefe3ad75cc41d8735a34e57c675a4f0f7e426c18472dd2c4cce7b4cfd37d01bfd19cdbc0cb785aa4b67650b0538c0984b002b561c6224f9abf0ca161e6f095a083510836a8ff53604f31b864496df7cb8de4b82ee0baae1042670484b7e411b36fa4ad734fdc6267933fefa3bb05d83c174dd47dd3b750d6c9827b204c0568ade7cf7b11f11a567d369c27984b8eb4ebc203be66f9efa79989ee3240b858e463d479acce90ea69f8aa0b51c39640800dc34a79991bd90177a2a535290c1c475deee90a2aaf0872a47c586d9892cb945bcf2dd0bf9a0f05ab6e754a4e5c84abdd67864723b18387e4dc593730e399815ab80e73d89b3bdc90fad392d297b58b9f616218e992f11a7776c8607a1af9e668bf4634f11f1770181491ad0fe11c695a42df779a1440887d3898bebcaecbf259e034d7a158074f3021f0270362785ebf75c562a21d1d5d0df5be439da1b63c0dc9fe9a5f65eceb1e5fb3caa8f1b09f03481fa9be51480871b9f1936dcc2073f179563e39f17d79cae3a09eed1fca1c73a6b9232129a1d30e9589e4e8e5ff339f5e527a3ed17896395bedbade46229230976f978ff77a82a2cb0ec07ef4d38e66e75e0a8918b579c1f72f9658a79ba0719562ae6c0b0876b9ec9ca425da976a9a531b02ebf48432ccf81b53fdcc634158a3a81c8a507280ddf2c3db360e5589e8a4d2097141d5de4410fadcc463bce5b8d9943c813e559565e2e82cce498227ad05884aee8e28506da694982515c833eaf52c2fa4f2a8430f0dbf568b02b5c8d0e24e0c5ebd2d607f2119aafbaa1939e261730de71fecea729174292be6f653745def214b441fe4dd00484be26ac4035cb28287b068d7195d828af05a3f10a2f2a95879a6f6029fd040678b1de0dd87d402aae0c1aa684ad22f5cafa91977d0139a22fd602a94ea82376946335dd471bd7f6c01faf15b39c627a80e428a90d722c06472260c47ccbe5a8078d5a344288a152a9444d412bfd435c3a2ee18ada6229066afaada1c86505ab8595f2f8defcf07f78bd0f1781b584b6cf88c07114a70050bdcfbd92de6f9a64e49af8d4bd759be555e0feafe081d23c3c58a5da427f39551658ffffb20802c6033fe60af1c9780c3ae8a26460aacda4868bfc599ded63832f3cbb387b957e89c9a3e4b3e25ef74fd17af614cf46b3e75ca117c104994d60f52a25ae301302ec03db83c66135951a115b0843a81976403d180368bc4d91994cf0be6bfaffc585dfc0edd77c75f3b3848412923b3c9b6ee3225e3b8a22bc964c68e2763d46ebac868137e5a95533dfe54a66f79b010fa4dd23fab06a42407fa14ff7477b7e6397a7a1a2808d6bed1186160501947443005a4bf89861f27e960851271199bf8a10d4e221ee94c00a0e36a922068d98d884e24e3bc2b6b2ba06d8fd7219569d71e57ca0ee01085faf3ad64bc79a70f25fcf6ed54122e0d92a80d5de3be8e411d24b28bffcbd7628444a160c721d86e0cdac172d9819b0b394b152b4e5a6c9618b1fdf6401108e84ed3f7c5c408893a49be7b6aa702e1ddae3c5d6dc34f1306ae59a2b4217a764f79067d9dc8b7c6b916b0238041ca6f78a08eec43d9c44266d1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h643c6057488966618aff0835cd38ec8926763cd10599c990148fb59d71aae673455a2bc895ed6f2864c0f9f2c1c8664d2605bdd7f1d2936d90b099d91dfb139bad832987aaca759bb2e69f0a695be3949bfbebd4c4ca7c3ec9083dd3895b8d68b191ffc54e0781623b8f7a8cc9a65e9aca3a8710ee479935926e4b0c8147b88d62dcd49d9b53da0092298f009dcaeb2dca781a29dc8df2e7573e3657a21b891b544490ddc7aa90aa8410d2c6304bd1bed7f040cf771e22db750a2c1ed6ca7e921aa3bec4ea5bd36ac5152fadf5878770776674ed5183389eb596f1f106bf5145755a25631457458718d29c6dbba563f579b82a482a086bf799f6c89fe47ad69bbb41ecb635cb6f1364c8581bc906816d4f68df6ae86e27400267031b3873faca92e42150fe105ec506cbeae4dfd88700a145a6dac70d734275d5d6c47c057775c2a599e10f8d4036da8bfcfe37f1d7eca1ccc42a63dd083441a09818f66e929c93cd43af8e1dff6fb67d9e058c06f7a30f536c7e1f56f959df8db3b08c22a07e513bfc56db3bb5f23a3a855ab73de9f44408761de69f2d8345e88fb3c579d90e61ab3e90b0526b6d7c17167ab72008f06d36c941817925672e5ce8fd7cb6720e003d3eb6d72367f223fc279e7ebc0276da4482588e6b6da4089f4f9da7d051e5dc6e94dd8e7f456867b617e1402665a28bcd7ece03a977a9a9e33f41ff4ee04efae845963cef86bdfae7e8c190e8faf55d1eda9c9e9c6a18d64ca94c6ea0b7c82db0e2ac21605151d1b8984d9eda3afac1cecd555c74d52c5dbd88d69b65df1b46fa536372088075a6c09012f9fb37ebd0e6580a76ae7bfded99e58f02a343a3547179534a833101766e197eef4376821a229029cb4b1cca51f72ee8670de1e0dbf9f46950f793a043126fd7e7bf080b05f342ae8ec6835694cfd716a35a53118ff86baf33131842777c94f7fb70c0ae0637d76c9857c6698f8b126a70885c86f5c04d5ff69aa5f19675224a43e98c51e768e1831d242e2c1a1e3dcb798461e3cf4945e3701b3a3e0ceed1cd2b66cc6b2922666c6dc7a4ab6953b6aa8bd438b4f20f7f611115d27cd1cf25aeded644865831460c935113a6dccf16566257d205968686886c29eaa7c3550281be4b9158f05ca1dc930239e16a4108a339887635f781c36130e747b0bb14c54667894a4ef29a18b3aaab5b36cba1cef58e0aa8798d5f2b2beb379575fccc74fa2a234c6f63ad7607ee9bbfe3c3b06c4b1858220a26a938566edf1c6b5799957bbd3e25f3188300039f4a92a644078bfccea932724a9a10e3df2ad1bd03ac8aba80564a0161dcb23c1079f67ad37b97d7e10137f2dabf25cfe9a459ebb68d8f962f297ada6811cf1cb11596be07fda4d7427a04000fe482e9bcab5e8cb1191c74d6a8291682038de72b9de87f66cc96e50405d45487c5ccb592721a9761005b722bd5530768b2220985b0158e4e00bb7274f7cbe4ccba593572d14b830b37725971e30661c14f0cd119e600419e86cc08d2d51de24c9d4a22a7252388db636f1cb546371b3afa91dd15be4a55883dc6d8c16bb7481ae3915afd9ca07cad7e93acbdb3c804c5c06046e9fbeb06314bfee33c79aa8df68ed8eb2c5235696eb79ca341d9b8be2eff62d058e0f9e185e96691c9e7c240ddf5fe4f2034eb3c177e2e40c51e8ab309815f1a68d701742af34dd88c8f321243c886e46b781243c67db60af5767a65d90b0d8c09ceb0c68c30973afb5ca234dbab7ed5dddcafbcea6bdc794c663c575e8264ffc84993f6dc6ad9a437d5aff3a8f8bb93ecb24eccee764cb7ae3e2bbad9f667a303b50ab678609b5b4c37df7d215b7ab2f90400e04346c9c97b6e8c207c008d075fe05110d2182962f64808c060e4a1294d48ab5f906f0c96658735b8809eb9258e9e14785e8fdff28cdfdf13772adaa7f2b2c2db23fa1ea97ca68d8f887c474c29d7e9c35b5164c5c7579d75db0fe8451e07d847b8ac317490fb7c002382da8b7b09cf45eb62875330a5ffff847d24f1010f32c313201da18efcb683ce9b0b66499f7bf0b8f599b6e6cdf0d7a5481d6cb584e0a0ae352400ef2e676a401aa830b2b24a160233c388750b97f0c204105b5a4b1489a7a2fc79895da268f1a3a91e08fb16eae65b752ace16256592a846558805bb22766e463e2201b19cd6857fe73dc46f6f978b79eff43315fd8dd4c18bf506ae21acb5182990f640a216bf59d2c905849d47a638a37a5060b26aefd45a5dc69568b121d23a39746f79262f7ea1df7671a0c4cbea7bfd4f7280b1837fcc8bbac80bb0e98c8ab9e507257e8a629a403eb2e0ae640c4ed16d8d3a0971c557b94a223767246fe940de422f3860ac520d0490e072bb347c1dfd5e38bfd2045fcf884b24daa33367ef51f9e828b9cdf8f1c47c84b787bfda2bd6a88457c069045d2d3cd9b077dec21155c011dd7e0e79aa04e9fa7dfae6198e7b60e8822a8a85901465ef00b2e5b29f2114953a3dc9cd87e89f068b6dbb39d8a9d9a35ddc0c7ce283340962a3049de73f5cad466c80bf21d5e868fc65d26fd3123a4473cc4bc0b4c1facdc56e65e06b6f9b1651fc1d9dde057cd7e9835d93ce669c0c20220c44c3218beeb6155b4a408c720a0159a14ecc54af5a440efee2390471caf2dfd9b84cd521e9d8fb712971e4f9cba57df8253de6eb1028dc0f0fe46a42e4cc6435af299ed6bc31e3a4daf8585b9cab4d2400b14e09e51b7b0c0cca4917831b0a0b1c8fde33f883bfa40bf0c8b56e6c9c1169d5f406d50b9f68a9aac9b76b60e9027fae19f55a45a9f2e4823dd5f42f94973e8f0024d33cb6a8bdcb4907880368b5ce2a727613c6e5cae1e9170998e6bed89ce3c7e18ca8a19f0467b51f238480426247aec70945acaaa595be22ff7582857d4153dbf71dcac7ced66c3b777300c0aeed5db35585b6c15e51eabc843ceb9efa5e36700ee9c43b5efe826a8fac2ebf2c09d7237c35edcc46ff9ab05f677832dc7b3b895c342b7c9dd72909147fc60d075e18e2fa7228bee19199fc620f0a530c55efaff59690ce8fc3bc517029c9aae03027764fd813dac59e639b42840725d91541b566598351df46b238e5f1c42de2eabb27ad57061748b2000f7a9d32a6fd209d2a05e18d2ed902d6a879a9743db5052bfa0e2fd7792e9e5996d9424a03b28d58546b2bd391b8fc6f78fe4150e604a01499ca6445d2dd6633b66396cb2756bfa1a47392fe8395de340cd2b03fcecb8d5cc8465c2b8bb3d6c5f022263064f8c1115877651b58cf6673b33b2af2d2bddfa4b003e760967943acbff19071815c1940e9531e046b989fe6a208b98290ac278437fe9873f44ac6c10058967e5db5456c548ac90de1b076a5802919b8e8886de9d6a83d310269e63d9e23b4389aaa64924b3fed94b047aa066f6250b436e6c8cb5fbadfbf5a20352d362fd57bf10e2ff421845cfb97b36416ede63aeb047e594a9dfb831da4d4315f12376c34d19a9e80d7d2bd8e989de8d35eef9274a0dc5161d1a41434b57984dad81e3885a8c6aac2ce225887dda2df461c44495fcae63997ea3a97f69e03f479aa578763a02a8b080ebe80899d0394e6b1d76a27bf6a8a1d1b040ce1337e64131a6c9e15a7bd3547212c6e2a4e81a9ab2dd148db8e2d931419b97492987d1027ed0d3fa713bbdcc36f9aba3610c34b4be1e3c4a0aa5818dc33f4272ce91047c2e4be88c5260e7724df972ed520a7d82c3bb2f72aa7dcce7041fa027eed95b3b997b49cae72195f459b796042ddd8db1e33191bb8f0d071f30e4a2e2274046e6de5d70a5a0fbd337de3d230d82696465b76add489d5f8078236230535579692a455d0df22e520f670e4301d64dd4f10e918f497c15aff3682c3d20f8ecaff34111e059a5804574e15e16225741ddcdb1dd3fd312facafa12c3876bad630822638ef683dead647b0f0e1f6f0058242c0939cc456f27e0b1d91fca5f353a18bc45e6ae22a07206a8fc15a95db5a451eb904ac658b6e2d276b364431bae4428131153f1da5f8563cda3a85fbf876ed379df75ea679c959b677d1156b9911bfa7d081897fc11b5e5457125e07b9a567eae2d8b2a70348b3bcc5dfdecb1c1cae3e3160fbf71034b6cd374d3b0e111f4608d3c313a2a4c0e4d207ca8a0f3b2f2d5aa21db34e3ce6ad0d43a73e730d329d41db475702ed169c8cda0e3465f8b48b5901c9f8481b5a77ce4c07fd7ec4d772307ca3281f0506df1a84f136505f6491d0a439bf07fae51c89c26db7a4210e88c39647477a540a9f11dd5b0c3e6cfd0d305e975eb3a5834effeb998584b3ec687661f05c84ec37501d3eada99b59b6f1dd666fd518010c05da92040cf73219bb333a3da6eec5a70fc78a1dd077593eff93465eb3069f00dd8fd830a073c002961f4cf98cbaa36fe86d0783d56860d0aae60c8515744e4f6d3382d5402cbffb9e6bd5c1c57e68319368a396a78c4502e4a2daca47ae693f3de71b8c13d2d792f9dace51f91042c337cb52ff5e7945027c846a05bb9542a2acbbbfd5a52682cdac5637c05aaba0229e89e94c43e0caf511778d1b484d517bd7ef00cd5a843fb3553db5bcf49b2e0c10659a3c39e563edad2a404ac11d6ece7b011ebbf47a38c4281d9e0e74a9fa7dcafb7c92dbe7119b4f16602eddfe2bd3fbccfc9f0ef7d254ca17d5ef62e2c36b9d974cbbd9cd10ae79ae99340b8b6d91bfc38f2a483771334295d61ce2c5ef8d7385a0fd735590ee78a33a6e8ec3d6d54129da689c078a4afb415e3624b120d8bed588b8632ec8cd37a71117551094ff22b14bd888f663af32bf0440ed921549cb78518115eff39b27babe6efe277138bb8cdd6aac04fc94345ec53d79ceb74251f7e1c83e86459b5d84003e253a738053896eb2a7d68e69ee9b15666e9c5536efe64dd203502eb8b8a65d1ba3746d89f93ea6688780708df75fb782956fa7b5f3cf4ce85eb3ff0cb98378f21454abef03901b110ebf3c4c12e813f062e0c7f5111c967df8f401fd504330b3959a23c6c98a1e3dff760492ae04ba6b0ce7cb9ee6c09410cb2b4edbb2020e7c8d7fbe6492d6f534366f3476bf0882a4b0c48a9b95e5574c5ccfb264c890135530b7c0d96e42238bf0d62872ef27261d1437339520a4dd10871e97f1e686f3c0f0f64e85245d7b468b108a5b6b1055021e590ce9f44a34888d9bc60b1fb52971a86407b57d21aa476cd9eac9922befcd403fb3ee70440f1ea048b6b708e03e5011b48df3a07b07b9aae860378e0e455ce9b3ef9a49ff07773314fb8e343a4c6cf69beaf529420dc3d2015cadaab60327ca34eee1825af337aaf50320055d279d885b131998c418501587914ca3b29c4ffc3c52597ab6d9d9fa02d4a49f396e122593538fd571eff435ae9611c0049d038f6cdaf9c9e4497a1d3e225d763cc5928c38ba53a68a09586beb29ebee38ce0060847ef2960865ffea660e88e03b9a88923b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hfc47ce56ab686707d0960e55fcae7bda2b41e06e274f8079042458b89773a40a240c32da74f2ab1d2037729f801e4dc5798c27acd62edebaa075a05b99996e7490e17b93b75d017ebb368f4939af0515f02e03b8340d0c2953f1605caf64cd030879bf4d28169ebf90728d35a9ba137cfb14a4ef7764638ba82533de523d47ffe664fd475f23b0211469e74ed7600f54b387371a5fdc46fe71d6030bd00b6f8778eaab3575bbdd7b9ca16ceedfeb5da2d2a20d69de8863fb9e3e4a681c74225015880ebfdf7fad5d58b4bf7de2810f5850c8931eb04beed69beff404ec3681a1764fb37659fb8aa7cc34198cf102a450d012165ce5ef309a9b90c190fae11b0893738618bac598a027ea1f9560e294c70f8e204444b6f5394a6436e09492a2a043335702023218d6bcc0f1818287960eafb8701a64708ab022ec18656f87dfe1b9c89ed3ff7ece6d7c652155e27665e4fc822cebfafeeeb024e4a32dd0567fc4a8a6952e8d7220beb9141c1c127edb43253823c7a33ab9381bb4c334123a9bcb733dc8c63b602c46ebac39b02a30148cf47fb8536576010ced8fbb7d526edd691677bbe2582716a5895ac951b066a29bf015defd4cdb7583846c518f0e84735c626b2cef735f42fa0c8fed0649280b388c7553ab868bd896bffa2a133d23abad01bc118853bba25b22856e74b095cf6d6add8cb026b8be5da840fa275ed30a3d571066710a76700414e248fd26d0c097ec045e9b469e96ddcc6e308f06bbdaad576b62351220a799d647f4056e8ea74fc8537fd293f93d9887cfd992038768d378e1ac868af24b00f64754ee77705926a9da5890cd87414c71cc78a4065344c0d6d3b3e7b4f8dfbc957c39cdad77abea8926a44a0b46f567c3bb61c4a413e3acc1a4fb533a4542b2e8f72004113ff212431032e3409968fa1b14e56083218ddb6761533198d4c674774a10ddcccc224f8cbd49e5cb6ed9cb43d4f0580562cdefee5d8d9f3821f00056ce3c9e0fc721a6d7e85f8cb127c590afe4fff989fe16b8d405a288e0e6e5f94c35e0bdb2d33ef0a6a101179c3d9b30e45441733ee828e31a96d0c05477bb21961564f415da86d0af4e14f9c4e54e36658d883a8738cc9ad3518efd5b6454d5b757e82353aeade2a78f433fa9f816f899221b8862b4e27347bb1b11a3d679558cb936a1dda72ada7ebf3184d5ccc9eed5723c192c9324dd8aafc7505c29b1535bc930dfe97fa69800b7bce64fc7115b1620067ee8b224c1ffcb2ec9bfddacb4579e6bdacf6e8e8427b315df7801bab02bf4fdc2af844e62048d7823e28537170b895c7e1b6477673eb5e41638136e13af5f3c7b1da615998df211c70482b0d00ae135b4243a2353108900c42c25bc7f919fc5133952bfa64d96972c4eb43c0e885c77fa55e22fda6e700548e5a1141db328c46b3507fd7d37ace583d035c09847f5d6a50735222e2de10ee9caadf6647604b50e690c5fbfe95b4c4ff22f29faaae63446dd35120ca84d835e2dc5581dfb0643d610d77eea8d3d70de4a04dd2fa044565f2818e2c176271a4d090418e2f31af3d78d9d4c8941c1f9c3e46f115b559b95dd3d7233ad63258b3ddb2d4cf0070ad0bca1ec6dee304c3a42ec24aa6eef3e4423b30d294559b3a4718a31b98233355780527dc91e4a705bbaa9b6c9e5555ab4036e55695df05f8513b0187dfd8ab473ade343dfa404e7eb6c4c38280812910a36a44b9b4ad09ed4004d42ae0d8ed9995b2178f4afd86bbd40f410f58c0466326a873aa9bcd4084b048185bb93460f29dcf0b69e8e16d79c25df6218f8fcda4d73121d31edb2f8d7bd2ee7dd50a69c3a30442832b3e4f8bf50aa09a7975c5098a820a0d1f99a59893659b81fe1eba186c7143ae05a3b72aaa453fbc501e429089106f656083b37df45edb664533d3351dd703c626759dc60c730c281a6220ce992de1245e9a56e451ddfdb0a36eeabd309e611214e6ea2dd60127af766d6d0af04cfd3ddc6948cd5991f4fb529d0a1e885da21d319411e888f036f5ea61a1a55578e4e6831360c9af5835839fb227010c52880e67df12427363baaeb277eab003f8d5bf2c4371bc2ea0446ad4dc64d3c3a66bbcf7c4f9cebbe11e7c81bc9bd8e753983742c4f9e4c520b52f7f85c36087bc4655677659bc1fbe50fd769ba8154b56f22362b8668b1f161f670a0007ac747b2b158a25773db9e8a4c0dad8a5014579566a6fe94cd0d09f3fe589c5ef8f8c1414cc5fdeb34964be2e1e3c1cd9ac557aa25afaf71a8cea09149f254396257499717528e8b83841593770f8231c6579f5cd2fa8d7e552287e92145e158f87acc80532ddf4bfbb1a60abea96a27358c087a3ccb806da2edf010653ede008545cd3904e9fba2db76a4c94d493a849665ceead4fad4aaab24ea24fa70a920bda68cc775ebad0bba6dc78404a5a63ab56efc977a16d090e27853c6a7298f26d75523a25c40265f1a5a894a09c83687baa19b27631595a9d7fa9a1a38a2741cb1d37e846db08fd230f6eb841bed5ebdc32db9693cf59ce29dbdbb4465e07b1783e2f452a947149fdf90a473af3ba901568f87ed544c6bdc2c63bb5a4107bc9bddcf9d9b0fe6eec6c429ed400e021a90b0ee876e878d40d172418aa70dc613be12cdf44a51970ed60432bc15e3a666f5bcb10e8ece46505846a1b866e68c5783ac221e0acb4619b011d97777e779614b577a8085467bf3120db73bd55aed10dc728676769184272e517a0edc5e3e71bc39b230337ad6a5aee3fff2b3062c0aa472f6e88719ddf68cbfcf578a089bb7c566286d85add8342d2cb536ed6a7dc37890fceb845146e4e302aa62c967470f13dd4865b38b264bb544c1d692680c3ab830785969f4bfa3f20cb91c4708a238ada45a156d6a9085d1faa7bdad79676d86e8825604931eccb02f100f9769bc3b34ad596a097976c3853b84357596945d964edb012e6f6fd4fab2527a415a050cf355ba3930e3b582a25e243fddea033a2eac4ca0417905de0f82d4ef5a5b7cf183cd28d189c3f77cb793897eb8cc4e61f3c2e0d5b7e315abd3e9c65c51a3cc21f642f1b584bc2fbcde14e0324293265f13baf8a868f9d405d6ea07fb22da002f5fd9c61a594dfaf30b484118bf9a003a2dcff7fad1d835a9d3f2f557f20c71f94946492adecfa7e5310b721d495c3624522db65f477af17282992608b9fe2a6ae7095869aa9a3269e91e6b015adfeb840a5f80df6a8e0ed4d69e77eef51587d44a9b2f1cab237e56b569c59d046f59c9987b4578bfdf4984b7715b30d0e3ccb945d4ebe9ba72d89f5e665c527d9694213d6257d7f272c82ae5dc2b4f264a467bffb02dd278cd05dd0662a3eb13a95fdfadd8bb821a4f003248b0351f3003317d37a629da0f53e1ba77e753e4242ff08f9b24d1c91e9d142456e143f381e5685676ead41a650fd895c0f3516912f7d44fc4a63a9d1865ea5aa1e2eaca6a62ae452056fe9def62356959d078235c0019222f2902cfe30ab8f269b853330a2bff0a5d2cd9c4ea039d7bb4eb66ef3fd420fb8458b6913be51aa5c68410958a88162968ac84f7274d873fe4406396318ccd0f998ac25e3190150926b1f121fe978352fd5fe1c2f09a82363b16841060af4e3eb7349bb018b3784f07241c0642ef40030c00f0f41ab3a3121a3c73e855078dc5b93e4d0c2bbc1e866fb9279f9832703a9dace37eeb776641ca7a6c3f4bcbee7edb67a53e7516144b3b37e7efbbd6b520b5f7abf082f4bc0048d5b6b6e83ed40f8db216ebfa5fe2a36f1000da12d310d3963cde4ef86e4e8c8c41e56c6248b5ff031f84faa92b1ee39f93f32c767c066ae31ec01be754bf4f5ed5bb4732de7391b005a3aa6f8b1766e2a438301c23fcca71f9019b85769c83345c06e14521efaa09937d54cd5d3848c0024baf3e5c3810b09dc879e6d3c035729296563f33e36fb38848d5909a585565102bef259f9e451c6b5832948fc157b44d29aa6d63257377b52d3b233bf437443769d6df6a2c1e8055ec92a2f4717be9c8483fa9a6e5887352a546a94468052f4ac2fbd8c12fd532de04996fbc44977020f8e4ec86aab63bd1ab7b09946739049557bce95e145400c52ff987b1e5a7c48ffd38c9919bb2f1efbfa48c5a2496be5511dfb07ab6ba680795d4b6d8ea8bd7fbaaf6fbbfd5987b1a652e7062510c77ceb887208b4c1b3fa2733e31e63bf0e16d02bf5d8a1bfc738fab10255131db7490d9714db15693b40fef0ca272c018fa56b3f1096db31b5ff6b74ae1f289e61d19ef1a1b44edb015497d3861fe23dba066b52ba925da024f59bc0a41ff9db592f7f91cacc502f6204f2a2795f75d152bc00d0bcf0030388ea39bb52bac0ac61f7bee31f7c4379edf0749c25b3b3d951510f093d7ea28e985c979897952e9744943e2c043c5762a1f0d06d89a9a2375d6afc2970f3b817965449de2ec11e398760a15e683049a98fdcf4075ae20565303457e6f13edc04064258d161bde4aab77348649ff020985f5cfeaecda91d6cdff008998adcd0ecd3c9878f58a8ee642d5e2454e22a1891b02c72cceed800188fcad81f6ccb0d47974c7c009c20a5c56a20d5ad8593530b3a4e5ef2c72853d8120d0d38fd5b1d18d84542a78c091efa76071ab167c08e552142c80deb9c9e7abf54ab10ce948c88fa47a749234720ffee5450a55140354419e876779538c03566adfab920fc0b6013b8cbae8aa0c08fcbc6d136481717673cb0cb26866f9fb929c848c294a9a446817517e8fdec722e07bfdaad3c1ca96dfebb326694ebc8534f87e7ad9cb9c088f91e242c9d71f70a869a7cd7667d4361474d49f8e24b1af132db7536955762fb6eb0432e5e8664b3fa240e14e83222a6352cd2de99d0a3e28a4bd82382da6e53c0a7a6ab8efdf5222985c7f10b6a72e2ed7c9f5ce15b84a90b4239f04e8b0f8cca82df3d9b40ce105ec1f7fcf1fa340462be4457901404967970d9ee85e193dd5f8de2e2190351ec9f44704e607736ea76198bf9ea0607be2dc663a224d5bb912238ca4b4f60fa21fdd55e4e029594b6aafeb5478422b83f13e9d9e2424eedda6b41b706ce54c86748291eaab6149d3e5e4032f5ba5886f360d775c156a933cbf806820c8c180a26f9fac822290201837454654179ca50dc35b0752d584526fde01f1d37db2a86cdc5d9ce9812993d0ad54ca3495e34c2ad769acc931b2619d3fcce70b9bff86f33fa1b6ed314a73d62be18e62d69dde8caba255cda3f24b1707518dae4496b1a89283d789c20933669c3081149d84a51f90a44fc8a8803bf22246de4ebb7e51b213b1a8ad57342f5d648a4398490d2a513a1d33661c99d21ae94443243b9ba35a674eeeb697474252033f417ef279f9b9013222df52c65c61afcbb486a0d500779da372b40e2555a996fa1335c7c7aa73a2afb96b5c529a21aebebc5329add16f99c3bd59ceeff02139dd9c153ecb30732f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h86ec7873d062ca3663ebf63007f1481e3d608b3a9ccf5649f7365a0ca24c6754cb59d043b3cf5c0ccf67c295608553531816b1fc079101691c942c1bc61618d3286308809712df2af5e4c06dcfe77e17de973af99a401e3625924c294feafe0f5a04e107f19677357734eda0058b845bf76aea69679bc72e37deb93a007b7d71f55ceae2826903f997a5cab16fd173d1b9a6d93130155ff19e43ffc34d8c42706972e164eb21e42ced144b20d98be95fb3550163d869f17edcb95b446c4984d790f84f7f396e284a4c55f3de12a10e464abd65fb1b3ac5cc4307b1d76c4006d1e9a8679d0d9f4827ce4a390bf725cd8ab2b97ba6c08df5322abe00a7ebcf3f33dffc61d51e21b43db9498310388cd15df25970fe2a5ba903021570f2c84608cf4c79ec171ff43a45c4aa4248e868f7bafb2730081b64e425cfb61581b2f9917ace96e01870afac68a4e30b18f0047fdd6c7ff06544b2a14a0a3e59f0470ce356e0f49cc067dd226b5cdd4e938653098cb053d5887cfaba4139472465c501613ed52166062248a44b6e5a792236b7e483541336c968c1f6df06895888c1690bdc2dccb61f76a5dd281a3f4d7940b8485aabe021c2cd4f6c8bfb074856781fbf8cfa9b2ade095fc3f46d09919e716464703fdc02770d5b87aa394d0b8af1720f686db0ee7bfc40a527d2ee7569359ff30def8d5c4d01a8511814c52dc54fc75ecc220cddff9228da4c6fcc4773adb72b3e0c8845ba05f1a0bebf41d7017ed108bd09f490473c0f7b086b0fe3b9fbf435176962e02e4f8ff6632241b5923834a0a1b48594087d59976ab9db24cbd6cb4657a88e2934b2ab8d3417a30af8d4297eeec7cb96d8074d64180dca2fee73882b82c0abf93a6384acee03fe786865fb0fe51b8c635723571051fe0188232a1820508d632302200218071910b9c12549320a2d8c52db1e09f844f65d7d0e6e335a7078301d4e7b373a289b4adfa89d60312f4d5a3c545a41ca309acf6b6344769464cdf25f27650884e3c822433cdcde4a536e57dcae82bcb743b7245378f1e51cd17a2f3c9fc54fcf0b731c48ade0d4ccbc098745fe0577243f9cdadd418361e0c56de5208205913cfd802526f18b4e6d8049d0486353c93272f4493456c1db09a572a8772ef3d2d206b341e2d4a7b70ff4dc06bfbedae7b45f785faf7ece8df03da55d8dd6a67ed824e7ef17b076dc30c50c317a091903127aaa4238971e330d3711f0060ca87b0c19573f9cdf11d92e8522d47fde1dbaafff553479607ed6bad671759dd47373ea7a53fd2f7c15353b3a310cb776ab289433ad36f5dfd81497b2121e81ecd12f9b1874a1900d39cb06f060902b7648acf45dcb626b968abd71ada2a9d16de3aed1aba2d8620cb2ee23e6d8036d7d472e7c80d40d1591d33571043d0b28c148f1ef0160a3a732c39d2a3b7a7402d3ee41ea15e7305c39fca3d308100504fa54f680db3e87a75ff34091365ababfafdc9354134ec62003e4a4a067d852ff22b18e424cc018773a223628d4f811467a2721434c6d21d6c7762dfd263131e1b32f0ebd27a2dca18c521a3794c670364fdc9688932d5a007021a68c14a3acdf862843242e3a13d816c7fd2c2d10226ce6c05536c0eaa3012a3d121556143867e865defb433ac4479595f338952d6e004abd486e4ef5093b1573f29721631cc83a65b67eb95742fa53614b20ea6b535b413532ca7c03e3500a28de17e1e89f241c489fde6e34bb3def1e4106708aa7b3ff749b3fed09b418cf3fede4fd9b877ccb698d5579b197219704f42f5150cbf74be278d1fedf96499890a7c595038d52b9841ecc9145e4e299d49cfad22dc1966973d117a6e71c41aedd582bdea7d261260a5fef986c0f0a87277f9a64fa9c59cef2a1802742e4a8b5f0f3692b40e6c9267d27ebdbb5439b7d1011b9d337c8f3975432d946562797ded026aeddcf57169b253ab7c74a5df9d97a2846fb22d87ae7f584dfc6c2b04e6f54a0c31b9950080b3ef4925667166a25690995a6554df6910f41bb76a23bcc741c6a8aa259743aea9651c4295dfd638d38ddee7bb1daaea5590e6465941be981cd25270995834b1425a22abf76d7a07b74ac6339f3aa7e7674347f577f168430f71f345a94c609cb8d7fca43c1d7498eb6b9334f14ed313bb2148981a7d634b90d31cf35fc13b56fd3be2da00814ca0343784923f85e75b22362db34004bf0d008a2641852ec7c97aceb949211ffbad26bad44b235475e0803ea6d50a70c1f7fa26e6840af9acdc69b47292ed0bedd238deca6f935492b7f530cb5bd2be4dd4572365b9fa3173fca79a64f6299a8be2115cbc781951692b01829a2107683742d44487cc5fb04dcb131db715b28714713c4e22b9a6ebc6afb0ca8b523aeadf94063e9931853aa2cbd2a8f3712daabfc0e6740d73f0754e39ce0cd3b6c56605a753705c3d6f03cb97b0a258e0438d646e2a241837106faead7170bcdc3e26b5f8aac492535e979f32a5c1754bacfaa48aab9b64c89a4aa0010d6235470f46fe6b42b10a9aafd71c3464cf10f5682081ee870bd7c9212578aaaa783bb1756d74dbbbdf97aa91a87bb9b27293e411e272f0c33cf4a4b43606c8850f9235555ec6a65c3fc472d6ae9ad6cdd9a84cd4c7eba5328f63b61fa0f0d5b85564cb17f3a6fb5444bfe47b31e1eca1d8aed9731ec4db23575f93194811db6b79f869fc0dbf0dbdd8f28a2f972bee1a98eb55df1d6ffe5d9f614ba66bdc385781f94ef3822da8a0bc06bd6010ae50d3250fc516ee2d3a2f3562ccd64e386ec37be02fef4b0e12f6c4ed140145d54bc5b4ef796fb439e59985a1cb6ba5f82067b4025736012412e79ed5bbc0bb4e835de5a102898f20fe7a2038c82fabc9a868cd8b7300fc40d5e1e856c9bb20988963f393af41976fdcca02501b3e0becd0d87ee444aef7df99ccb899e1787ea40ba53bca4d4f49139ac97bab8d6eadb1bc2f7a97e12af69708f2d5a894638886f7c0063d78a1764fcd327eb47f162e9565fc7c402aea4c4b8bc59898aebcf37c6bf9702a52e76f9a2517e27f2c1eede2a1f2eba846b4f8eb7f09e011d2d28320d46a8aaffaba37203c1551066bc14c744a82687dde9e88471fbadc885d735b47917750a1bf2db4dadeee6850fc25b814d28831022d0a27ec50ab21d392f1336306531b1d74d084ae34db69230a2cb55a9b536ec85e1eea4ba77b8358d4e9d956bf6e05c6dfa88588a8703ba98e49666de66539f76ca97ab0e357682bb80c467ed8631c07f25d84a993d07eb9a749f980f66bca1c02d0bc0fe4489b058672da4f5ae950959d649d38614d12dcd5f755c892ae1ffab986a5164ccaf474d8994895a722e75414ab76bf18fa45bd532605c7c2d3f02cd2e8ceceebdffb694ec75b0f2763d61047188fb000a822c001359750af968a0343c2aa89fff247b0c7d2900464b7f6406e186d7a5083f37d799609738a18d98d027d7977c1b5b65891f480160c0a02f412082758d88c79fe3b1d2c8e8fc1d8b3c28fe5f594681aca6d3bf0970dd00d6e956e4c2a989802fe7ddb0c75798eb1a1df8ef9f6449b1e6ca1d54bc29108469f38aac63b0ba1ae23f0d28eaa5e914807d09559d28dc9932a34ea49fd682ccad02b5fdae25b6ca2afe86319c86c1de9e7d8637a2daaea3c23abc552a71d49456a704b0c8870608a90792c8f4ed8c72d8534b2533d3fa6e6577f6c4efb5d193c132388e93a4743c69da649cb0da09867e570b4e00c110a4fb3a72df2c306d144aa24fbb9ec0f28eb7dc7578b163711c8b636fef7b6df587bfa8f13aa6b518ca66afd93ba240a7cb530b41a19ff93d645310c8b488318083866fd401f52002d04e7428bbbe106bc794919566560b203b8f811cb77c3878dd849563e7bc8bf488b3c8e9c39123e5a62210a115827df9b7c9d58d1da6e02f68708feead24e709db25ac716753f1b8215b7f809449016330513947d66529b0274346e4b90a5c22a62a6a63502414f5baf8cac99b3134b3130df02d8045e257be1b706658c3fbae1b7fd0777d7fa34afed8cbc0d1daa963ddcf0bb6b01fb088009083c6516205b4f2bce05fe893b5688759829fc86df1bd0ade55d79a6e45fa88087113d2a117d99be6c95b4383437c5db91da34ed9f95c33c1d97f03fcff65a3cef8cfe87db53eda8ad597b8eecc6fd09aa8a015d78206b4f46b98ed675283135743f9a712cc82ae416c36c680acdd0286cdbe84dafa9661081287af079cb4c6b8b845279feef483c2531e28c0fdc5d2ddeaa03fea0682cb6e4055d38db14191602a2cbabb509a556cc8001ee068ee3d4edf92f96ad9589c8c1ff789b3153ae64721880086a7b7e7e3cafe29af3bc8ca5f5c78e0961b47ec7f301fc624b73e76a1c34a26eae1367ee4d40d0ed847990e97193f01174e1a98e0f0f382ce560028b49ae261ba0d2a10fb567e87ec4f5dba83baa3edc1fea4efc97490a72d06e87fa03edece98645f43a28adad9263cdf5467f0b8b631bb1ec2697c56e72410a2a026c1a8fd48a35903a489ef280987337bf8d43e4b721388588990c4c2de4162587bb4d08f7e9985435b803635eb37f318b21a3dfef1a3197a594a22db673e7c35b296def7758e5484fb31dc9e38c7edeff3e91694004bae238f739b47f46781e0dcfaf262963ad3cc7411b8a8796ae51fa941a93d57f162b880b569a32bf758ae2c55ca985ac13364e39fac8b7cd41bf1d6f0b0df58a459b9f6358c112bffaf3e0b3db9fc8dfbcbca150bd45f01adf94d4d3ad8f9bbffeae7df796a01d6dc7481b1d285704397b0426a51e06fdb4d96732a401d677b3ecafd7417fd20924bd249c6a545f20d19855f8f29fe053676f4aacc23b31b3d669c2351bc1e3b1ed3483cd6e61044e85f19ca66262500dedc7b820e03c0d581aa7efbcd493dcce63bb82f84a4ad3b9ccda2332e460fd6ba53dfe76835c43fddf6150e83bdb7796992a892ca58ca09ce55ebae027dac02e49271c18070bc126b706a1e48116f026b91a06d5783093492f64087c018aa9e6785ac7ff4b1b4b7d1d3382ef498291e8ca7eb025d75a877c5bb89e5f2a75ff2cb93d15a8de119975ee50baa28eb3b3b68948555373b80e78adddf2e217db3e3aee790f85ee9bf6aee7d2acd3c96beed2bfb4c6b26d471b1d6105976f05596a6173cd1020cccd9dd282ff2725318cde303f7eb433fa9d7f3de11b78dcae3971cb8a9752d34eed5325f2aca271567841dea755082a8b0ca9a46e85b2af097012830a0c52fd64bcae126cd28ad3157d40c57a055f88051f7da575a63722ec8f6733bf3b16b721a6719189380aeb2e7c6c49ce6f763bf9a396daeabe725beee3f911ce48b536ecba3b5b2fb3c1c73c03c81587dae994aea30be1b01892389dc501e8fb26da8e28e3b211ad89a89464d8ac85b12070a96700509254cbedfb8b8818482d03285ecb9b61c835f921ead125e6efbdd27a8087399;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hec76d733c6afb58b62c9333b1f01e98e9049d3408cc4d12f8c2ae32e56bfaec30969e67f1727a8a154775593566ea1ce6bf5a6c53b7df8ccf08ece31608999379f50045cb3101d6d867838f76f068ab045aa1f7e5e924f815f4ef99d09cc670a65a7604b7da4a6dbcafcc8008e00491c2a27e05f14ad36a7df9381a0cccbf5cb6e117a0702502e61af48702cfe7ced17e8cde4482fdc3db86483933c1d69fbb847f9b1ff697f245b211e6baa5118e0f8f67ff471cf1e5063a34affdea31ae50bbea0b751ad8f08d650d934ae24b25e86ddb0bd5935b947522c6575e9614eb7157c9d9205a1b39470f5fa29b5cb4687c77c1d0afcf015a608ea332290ddcb80e5ca367300b0b5299390a3debb72551634a0341b2b94849b369caacac036af9adbca5ce34363d16a394b564e48aebf432ec9f8f88f98ed039ea9774649442905ecb4ba81ecaf22349583fb994c8bf1090a16490795a4da8fe02af735daa955d86ac8cd6e2fd55d050275ec2ec5aa4dc4b3b43e6d711715ef2535e0347f6976743cd1ae357e8652c56f1dc06639f345c1c2ca90af687cc35662ed70bda5880a6fa1012b819b29fea837888ad5dee31a3ad4fada877c565d09df2c84e7d5f0ca3a0d7cc41aa4d9fef103fe17783f8c07844d0f6e5b0cf3fe1cd98301afa0cd41ad215971a06d42ceceb855580c79977d0cc023f9f12949da13f98752f9c9de5ba5143a1cc43843a756e02a2b2001ac8522bb85710bd40765f01ec5c02a6bbd1a495421690ed2f779b4e8ee7cb9d15a9d57651d6ff0b98f8e16150d8f8fc855efbf90345088c23b0222f94eeaa65fec4ae1ae0df7f419842ce8e3da7d1d4d11f0c00e3556c981ffe74a02ec5ed532d7b2dba57930fde233df846d9ef924d1423526b9e232379fb5af33c21d444656831009cec9d4c6ab6d4419fd0c1ec8669810a1d4e45000e4b98923308cfe1c16b6952a556def5be692aa0e972e0dab4ad73861efc5e1a02af1542cd1fc59b06b619704a5dc710c119d22cb34c545aae88e9628c937d979fc98858515776974499597f755a7d32bf21723bc88050704dea906cdbddb0908be444f5d86d29057a0c2bfe479d2c8ae899d32549e99966da043cb40cef7d69eaad726e89ece1dbf2d006ffc0130ce81b82976c6821e05f5f84b67d288cd1328b440b6f02e99e13a1fd947f7335a51d86b495db534fbc6e1c1120dde022832fbb8c73e13fdc153a728fda9c93800087c8f5e514d0cab7e78e62bd233eca8d9dcdeb4185d4f52ca980324f02ae2d46101ee2f8732fe259da0e4c4b0047349d4cec5ce205f04d666193c9ccd0171e99de2713321cda5d8448c468c5e03ae745e93965ab1ba40ede136e63e89c115ca62760de0ba02c36382f05efd41237b7b3334785740a40ea20fefddcd2ce389e028f6891a93dc03e3f82f3eceaecf991638e4b9ba1a693107f20949796212ddd45de0ff7430d35591c00765f9127466964417b0c16a1b98ac61a65687d943ed9fa3b8cc078cfe0a418c69b75a326128dcd6999767a8b6356345e77f5462393794f1981a4ed6e7a21fbf1430836e3aa11c9a6b7eb5d4c58852f2b4353763c1eac286b2c4586f720c5c1b1f776871f97643b1bf22c760a660537376775d07e170b8e47c0f59abf1aef4680d2a0b6e23c48f765b4598f2a5c9556ff6d01236b4074b29c5f0468e936725d3251121045cad06971a0c25edd7fac289f4ca6c746145de2141a2d8c9e1dfff5a9669462dabfc9cf4d73a997cafbde68ad6cb1a68ad31a41efbd50498371557aa04613e079c1f58a1520cd9cb8f6833929ca7038e9284a92fd1c98403aa636c4c0710aac06981d60ffda9ca8ffcbd26c045b50b4c7329b2eb847fa7c5e07a79e01b3d84f9bb37c49dd74d3e6b712fd64c6f0985fe024b77971f190aeca517d986c0b2d0b6713d181a1a12b16de793bd82577461708bfeb9388717fd90d110fbc3454947a97fed282aa2ebca18f715f084b6ad954c0b5fa2e0cc13c9d5672f8207f1d0db22f920a50b90841a9fc5e55cb36b60d8398f96b5e99ff57ac8db5af2b5062433d3652ee134c44a8ae18c553b54584d27a6d3ea209df65f1eed40b105ccbb1008b7006e9aa4a6b0bb8af7a086521caab2c8140d3d00d14ee7aea8a5f9e2ba9ef0d4b40bef31b71ad587cc8e9502456aa4ed31258891a3f63464f1f2e274c356144aca10a97aacdc1cf3645b0de9cba66b6dbef0b92759c70bd02f7b76673a9dbecbdee1082d59ee52295fa056c969da09a926ea26b5fbe9b7e380b70253c620f72760371f403ede94fe38216297d74f98fe6729c54380635a645512902a764c190c4954c82948c7a7a359afbf76be481c12a108140085e09e10e6d2d9dc47d95b9b13cbce9b9f5f8644647e2047da1f6273e369eb92e85f551f00570e1e4c44e6fdfeac88a6fc50fe7dbff75c642719f06355617197d2af6fad66b29b81841ea63574dea0846d3d5d781f5e8847cc303bd4a6cd6a305a29f211c40e57fb2c554e0b4bd681a3d7ace7ba1e6bb9bc28c04066c8a25a2db5f72625c66269c324ffaa47535f392a4981d972faa95ce2827ea0a7b4f42bc20010cb6585ccffe8237b1ccd7ddb86e34ca4b5106a472849fea5b5f52367fd10c78f0c1bd9285343bb6001e3bf319105b601df2671ac4cad681fc6d76e905cea3f2e5e1f28fe36fd3d3ec063d0fb45b2ca04291897c5230cb64d8100e80cd94b029524ea476220399a4137d2f53d393a5f6837bd5bc9e69dc0a7fc80c57f5301dea42ec4d106842e0898d1074ced483b5e6b5c613b81ac7968d2a82e88d3dcb16abbb47e8e65881d80a69773cf9f28868b32eb67afac7384efb174fc2bfbe7d86c3f32595d5295f97dc1fafc9d9945d199794a9d7828ab724ae9887cf3dedb47c6ae402065817b8b6b884ccef98e4397fd1380b410467d799cf1e17deae3f214e6ded2f78690087ffb3d8699ab3adcd59a547893315b5f83a97764bac75816fe7d97739f56b5df16f6c7a476f3344cad92988380194511dbf5620288e06878e6c2a75c1addc9ba874670795e9b910c72df61bf4d08fe490ba6def350890870d906c6b926ed117972d6897882533e1430f41cfc70d43fd45577452c9c23ab60b559b46c90dfc4013a0f4098e33a490b306e93521c044f089057e0bb613a879ef45635f6a7393b68b223b1043e5569b068ced741e5148f5d2f08efc25d78541ebe88d941619ce02f8b5d6136aa2f918234e22ebb08dcd6e36320483582b72d8c1defaccec336c485683e227ccb983922802bd94121e05aa8af95359a9ee38ea81cc535223c737f8ed81b28ac7314c5459b40ec65308689fc911209b3f9eb73286eaec8810f703c9d621dc1354275870a8f6e137d106a2d747dbbbd0f8817c42464abcef7a4f2870d8fe4b898f1665dfbc7bd814cc6640401b061232d42f16357fba40afd6570dfed5522f870c190429f7142373873c44bacd93246f0666ea0c491d09d06abe764d5fffeaff9be321d50ffa712e78e8e4efbe0f8e3c0c85e3b450ae69fc08aa2e032cc0932ecdb5c796ee9e855e16f589db1e5516e78c32632c29330120ed327dab70b3f552d096a3cc03b81650713a55e2811d18923eff41778058930ca481d331f25e006bcd0ff66455b2da6ad551076c5c893ca1a16cb4db9e5b00f7be18e9f3bccb9788ac0fa3d57e77a428fc048ade1c5c2cafec0ad90d2cd357c89adbb5692db0c7c894fbce6433e119c51612cd1007370c8c256651200d798391676a73bf65cbad02e14d33a4bcc5fc68232e1001b291cb26823f196f98571bae21cfe8e66552e9911ac964b1575e3bc0c063a38540d8ccd9edab806daae1e2dbd54f30e073993b65fbca38449aa357a4f219975172d027b2c78966c3e3f8991ef0a7cfc7ccdee57b30dd7edf0b067d1e7695c68522b1e518196e64c288c7eba29957e4ffe5f148b6c204f2fa6e40857dbce31cc083cac0f98e9265b4e88ef815ef37b37a7a841c713fdd8106892bfb8cc303197cb8285a5c7d415a75faae9f091dbbdcd8e589e403d435b352dc5af90b75eb0903d84bed35679d1e57b2207aa677ceb11b631ef52ca7179ca37417258ac8fc7de5c32ca235c437004b0a3faed58f890af75d8853c78d07276bdd72475c985e04d937bfff302911bb84eee59df889003f52033254752532f20608aa407086b37aca6894d7c12129837e49f01fb6d29c9c4cf476a5fdf47cdb7861aa5505518bb65402c898e97838f20261c1804c523587b5fab1a454c721eaebb6b033a4cd95d69a5ae14fde7965e07f142bda1a1494d4c239103021f38e9e548ff77bd1cb189f2f6b2a712f9677796b9d0cc171c9f7286b32996d35660655daed86ece624a0dc55b5ee889d11f10f53f732cd6c62a27183a24b8b5f82699920b40a4358469b2c27e49fb10c1a7fcc2af806a2e2ba958672e1dfe8c84462235fb87704ad1a9d0354b73c0277390d6eae0856003f34ceb064cb9e92eeb10e0734ee316b91ea1125e5f6eb0a1f3ade11e3793d58101464d0c10f26ca2498103cac60e960c71d133d687ce308d34dd6587946ec812b3c77cd3d6ff53ffb1776cbd43bc1a979ad453029f5876b48ef10f11d13e428b320959c54a0b24e651f36c3b1b70f104cbecd89ca51f17f5c36a3dea38b289e1101071a7ff406d61c24cdc00cd5d4457ebf6c2816357247f2c62e7d293ba788251dee985eee0f2f8dd676f52dd0982feabb20781d8dab35697ee35491bdd04cee507092a356a41349388abc5abbb3d05c5378e6bef05b3f1fca3fe4bd4897b997db8a7037a49c7a0198d0caac14bf799c507b6a07c4f4a07098fbd9f8796eb14e88d908bf4259f94a1c93244bdc4243fb9f1311cb8910c39ca987e8c62c360ea58f3100ba4227cb7477ceb7ce81bc313079352aabdf64fe8cd156c173e2b2407f853e99231ff52146b9eb3907d65ea2b464f96dbe4edce2e0cfaf87ccfcff68c905c7d71812d640f5c309ee36cb57ae03a65bb7864e206285396306760e494b3e6f539b5fd595c9564ea7b4f470fbd53799514defa12ca8b778052ab5c739e0780bb87fbc6ebc96faa7764b61cda2ecc3a1c460ed70a76cbb1f1cee91807c435e29564cb4e89ce1c67870dec34b88121b4e021fd0230be2977fb67e8979d6011ac26f0bfa1b8be9cf9274a012cd212685e9575fa7b79461ceec141ef93e53921bbde3242351641216ad1ca0acd8f573169373c39d9bb1ada3e59d4909d65b2f6e85c63b1eed92de2a2344017536cc6a2be46c6dde791c59100d4be1d1e0cfa8daf5f87094b7e5e5aa43851edb11b8192e0e6050f0e1d67715e84818a5ec410d61c4dc9d2324d8cc39d05440d79e30276b0d63fece63f57740cd2b94f9c38df34e93018d7374bdb4823be3e17a211ec6c5c39c00dc8f34dfc95bf71c9133b0c9e63803e38c69557de2008f2ac951b752928af4bf2fe6314dab06758dd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h49a522c6cf2b9df8410e954632abef40f13b12c97495175c364b851173d5928e500745e039ed8b1ea0fb0c023b4f190e9508f2160d2ce427c6acc6e1610ec21a43fc51adc06aa809b06081e899b1baa024e3e6345b1b3d5ae9a784d67abc3d2d285323d2698764aaeb770949bb8ef4082b7a85ab6f77b6212e9c4d38657691b1edde98fd41d0fbc192d8b444e3da04697cb9861e571863c22c20d7a9c0ac465b58c941a21616f3aeeb427337477cd60bcefe29458d16c834ac7f8146ff3b5d55846131e1558efa1f6433662ab16f8adc8b5b9af857d8c5055dff4c9db6270e99a959ad507fdc49a435b87617303900059e9e6bc3cf2870616570eea40fe36f4a92cafe4b40f5ee7647eaf0691f2d0d2a12826b62c693f58eb95cb775c2b35e44dfef0be8b3881a0f465ec58e98d5eabe6bf3a269a589ebe486e2c6998fe2f79ca22b45554c086ea37f94e08aa2034ebcccf0ac37d70fa2888f4112aa0eb415af13000151834a067dc41ea07a6014ce282bd80f52ecf61691834f5f5843371431e13990f978a782b36e3e36cebd858a001d12dea68a5efd2adad5d2af67f03303e383d1b24beeacd8dbf76da01a22c8852273b9a70507b020649b695c3efb9e9ecfcfc30e4451246c511ef88e05bbe2dab7011715c4521214448dff010f241bcb58fd42698552d636aff7dfaf89c80a56a1cb3dbb711650f141d64e7ec61f11ea83188709964810335213632602075e6b5933c08538c724c2064a805079f5021a492105f2552120fccf5a8e628f64c06bf620c3887637cbb2f84a1cb6c2df4f9b855118a63a20b7c71dc4657ce28efb2c4abc443c0eadd8a993c9b803e43278cfb412fdf92e285d498cf080cb3e33e110551bc2f2d8cad84e354dd747c8b3bbcd75b8f14e5eaa1908b394a9718193e312667cab3e03b381f41e2f1502b2842f627563484636024439a8b13a0091b0e55e66f3e337f0c53133fe2dc6e7a19a1f927c17cdfccd51a5d0b9cdd5e7899dc504c6125e97368d697af92f424c85551fc1c4a54082e2fd4651dfd9941ff1264857f0a4731f99df0470fd888f5e7368f4911e7e820b1e9078ec0a4ad0079714666cdb77957b4b02009b3d435ac5259d2a58567d4fff4a7c5c6310430bb6338d1accdf090c3fc16a2ff323861366cadd8e534df1c85c89157e8ecd580dcb63ea87d7320368208ee41a649288e08b32d5202f4c8f8624a6d7f5f99019a107de95656d5108658165ebbcc4f8009a217a82f6067d886dca1d27dfaa7324fb49b746610db783d7c3be118171585eaa200e9146e3878f005d84da5985a60f066427dcbd7c2c76c21843be4ac409931f6f17911cb0ca529879bca2bec18df59b52ca65dd429b90ee1e6fe7ff054b6b4abf9cba6e28c4308de8d32426393f0b35ec537f4d40ec325d47f7675246f93406cbafee8f4a9088f9df62678ef5f67730afd2fa49b389f6eff0dab31b2f9a746eee1262c7e32ea1f27c01585a7e4f36f7ff137532791ca34d9b3eab6cc58e01a92bbd9579f74c0fa92f564bc22b3c43b905e01b0c8b9862e25b56f4fa8108fa42d71be53a3c4dca5e8453966dec0d4d1494e459b135b26a1fc444a97900cbc01f37f25e9469d25c01cde284f5330d4ae6a5cc7fc9f1fb3851679f572351a37c84cd65338d551f698707bad076564d61f2115d3ea55ae905cc8cefbda460fc5be0883c891880fb0fb430fa8fdd7fa3e96a2e757111acfc56317db2a638db8fd87797bb292ceada7a3fe121c22f958a443e92c6a5e5fe02075d2fb950f50ee4b71e135c0ad9ce6d3006931410c7d456852145f0cb6b8158079fc4734ce461906b819977b891033f32045539781cc4dc88b57ee2ede99d448b9bb0c98ca9145b0a1ca19c1231ebca3f8302b5ce094064a8a277053ebae3d9f91bd90dd7ae077a445e49161ffcf071ab23a57cf843dc226ce4df8281417cc5c907f0fa3c17b6033591791dabc7b96a22509db24cbf026d610d68d67bb2b9936df33b7bc1eb698159597fdb060b622b260719ba9bd471728cc8d2d16cb86f54e9effd494e17c5b5e251620fd0b30f158a66710dc65181c409dc1aa7ba939be1e9ce7aaaa32eda4ee54bb2ced2a72b3c91ac9bab603ce870c83aa9486fa5d6cc8e95ec8e8603b7347ce40cf317260feb18cdf1825155695650bb36d6d4088cee2bb68bca55326a6aca9b36aab48f319d73bfa98162307a8721b8721881dca5431c87fd8845f9dce430780b49a74b5afc2c9c46204fe99257ecad405995b00a79f18b0be0d1a5c4da60617c400bd9686b522a2b201e3bd535883519204a31abbd9227317b8f9df2d15facda198d9ca66d26128e94e89d48e609999ddc57d6076e844f752a664f327391321837703e7a95e3fa6c436c1011d08f9ffdbb91f1023d4461c7967154c48aaccf293edd1713772364dc428081a0af548f853ed70fda6237d9dffc6369e42d877dfee5dbf5639df2c0e060b29c07ca7177f03e84825f73a48c0b38c839f40c048937738c6259c90f10f06ba2eee22b671be9de9dfd203f5059f844ece9f808560089c8562d61e7e4b97a17459c3b9319a02dd8ef7b9545cd892742d69c3c5eaabf540a67b41a904af122349875ef70a6051143d0e2ed13d0508051a5f18ac908c0b7e939747aa93b77bf15b24080d5e1ec2854777f2032d3f96cbb5a0a9638b09fd3637190782e59da8dcccbdf17372638e9035ce9bf1570d855b1736cd7e492ad2ed1d1afdb78d606184a68e7c6252a2b0cb1ede679365be8c393487bca3d46e05da5c1f0e8d3f5c3996e576558c7aa2b1194074b324b8c45b93975fdcf2bdff7481ec3d6187ba40adb89e0ef567083d3bf7bbc869164f0c57b083e9db84124a8656fce0465a2dc4cb06625eadad96cdc34dd3cb5957198839166f498dcfc6bb86eaf8ecfa3ec5e4aad060d0770ba5d3cf74331fe3b2a1b00e0625fa99ed6cfa0b6b69908e37c36affc2ba23a5c2ca6458c7eaf40e387611d583858ea8e1b9f587ce66a32d1520f616f0bc3c6222e788d6e89be0cfdd17bf7de5576f867dd7857563db0787d1988fa79c87e93553f46ef46359160e7898e1e7a2d39f093877363f00b701da93d0f01ebb7eb2ee197c376347c54e1bd51e43f7ec531a271a276383275dcef1bc69ba7f4fad009978b3bf6a645fe146e6dfd5f4364dffc6ba7dd7cb5a5d285063b5eb250fd6e247fd01fe58184eea8a029fe179d09bd2e8415cf09dc863dfd3ecd87af19faf5d09eff543516b16cb3cad72895b539ae623be6f3175d85c19f820daaa70c89c4800a89a8443455f4996a8211b5395c501179c7be6212f35abb9823a07dfd177a0800ef78dbb1523bd620eb66899899cc1c281d70b87b89bdb2c84849589c3e7b76cd8e5e875144b0c20ca2472eefe31cdeb7409f8a65a1ee44964de81919ef0422d377100d343e4c7d92696726e011c7ac67556b0284605a8050ed3c2808d706440542882b3ca945da125a348439fb42ef542c305c1289974a9009c43b539ff9e38c64c59c989974315ce9614dc5fc03efe16bc9c1ca477ad29826959276bedb230a26eace97a2d0d7a786cfd823f3ead2bcdb73e323b69b79b40538c91d14f5fc368f3d831c523e31882fe83e981b5af6dada62ad4100135aa5d89de4346dba2878ef3e7506e1ffcc65a01e4984ab65f83f6459c82be768e446148312c2c723baab05d3633ea19f34639c908b16f2293819ac674d9db908dc2a66a49b8a4efece2e586077674b79811d79ae65508ebb5b7df70c7d4d689022ccf066d1e6fbd104415fe6d2b7a6e74beec0f18b36b43c03d94f2229667e73c3c5df84747ab047ba25b49ea63eb8bb7d1a260c95e0343170cbeac3e93a5388c7cca96e880dfd7a056372b241d8f13af36a9232dee3e9ee1ae81971389f83e53e7412acc7793f840a4cb72bf972cb53df3bddcc5699f7424daba9e4d40a4f4a7a0dd4a7f8a8dc7e1b3628bdd4869b39b719a9ff2617c73b64e3cd20a64afd595e5bf32a4bc8331e3b89d90224f4eb1ea70476d9edc25c55b622394876629fc1d979387d9cb20933da2b34deeef32c9e2ab8f66ad6409a7f4b9ffb134c03385b6d6c036e58b9aef9816b295be88a3fb790c4769b97ec5dc515f0d91a9bbc52d53085a629202793ebff9fd8247bc20d3f260b75786f41adcb8ef269a7b0e5cb35b0ca6a77795d57ea273fe49bda066b2cc9ec9aec0af922886a8580f3f695eb1df085e55c5f4732ccd0d6090a0e4586b2feea45d39fa0061266ae1a16e7bac2c58dad6e0776e6b7bc1cb807059610d4cdb0d6d2b4156757cfc6c91b1a71bd65151dca5bef20768a6415e68f20f7d30cd18fad5c73bcf47cc34b33217bfdfd5769882873d6977f0a6d64d81804021f4f53f3a9b82ad79cec666ed8f730b0cb325537a7eb267d9c3b49ef8536f07a5869afee83831c7a9c3a44204690208a68f6a85a0e535cc9c263de8d268981938b1ac5f9c155cee1fe22bf33668577f4c338c5168f60d26c5396abea7133ae0d77676ccfbb0ff889b2971188fc4f707502413bf1798034f67bae8092506ef2b2086832a178ae75df0ed58e6fff8dd2e3dcc4d3192b2a44c5a9ff132b3908196a3ecdb8707d71fe2e7322631ab4ce5220451668ef04cda97aadf95e392ac7488c1a25b3f5cdef3acf35c38f26ed36b5ef57bf83527ee22a792a8f71718cde1e35718bb62194561e0b97e736bbc99a7a07f3db9a7e95440b41ccc351165a598a3e0c8767a5b91da6e360d66d5dde730e1e7d9cd5fc6b44654706b216d103f09383b73bba74d2918c0a8f17de174df3fa74341853ada6a47ae842cb8d1ebe888f885bb8f330a26494ff00328766b7432278106754583d5e3d85b54ef86026b6375e438dee87f4df45cccbaa8d7ba222f57a11b747d9e2e630bccf3ee85966de78a4ccb26d9ac4c0eeaea1ffded623a3b679dc9bfb3d460d59178fac27eae921843afd2cffe6e9b0078e4e7393cd3b0c7d78e449faa7539148c03a2974351a237b138ea14ba585af80eb647f3cf6103ff67eae639b2bd89ffa262b8d4dc8cfbe9b8f431dc84725cf78acd1a7b371e34b14cde3981266864150735a8f4020a2b454c68af370ad4c0585d3282a6844a15e03e0b166e5f638d8e873f018fd3e0011026574abb1543e7e9fac496f532f975855e3e7bf2dba0df2217a93686cfa9b1ec65991eb6515482b6c2e278b89d6b65a3b44129a9bb6d04bd5f44d96ec42b10a124d5279feb7b889db185998025775e91080f72bc74f3800204ad1ee7e03fecbe6e2d5f5773030211487c7f0202372af72aceb2a3eb2b689c5966217b1221f5cba279171fb819f0c0a96a40f39d67fbf2f381858694d78e96333f0cae2f17aa2fba2ac3a8005ddfffa84b4df376edfa481af2ec4bbc097f0c8772c71dd4266a35a7c9873702de456d2475e58af3ac082576364f71862fc841ca3867fcad6bfe78d73974e1b7461;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h9c06522ffb1aaba97687ff2a1b7f01be2bf28566344f809c514f078db769ee55aeff4ab0fc03b743814b3c38f1024cbf562b0bc0dd2c5f1b9888ea89a8210a6644221088f4b6b34cc8882693bc09fa99bcc65424f8dc312a3dfaa62d30a270855b0ed6b9cd1f2c4b7c312ac74b144a6ecd037d0c84ae0b56e5d5cc20052f07d1e150ad0833e43f78e46f67a1075ee9471dcd7e2cc6764b20a2feb3cf4ea0551d2b29ca7b28c83c0b1af3ffcc93110bc77dceedaef504897d19de0d0d1deb959059f2a3bb2e8f247eff6493679d2694978881e0b1a7f5de51854aaac05e4ab8b9793c23e8436f21adb136a04d0c70fcb06276b6cccc2c36e7c503da7a7bcb77391dd3db1f31859cccd946c44b6e8897b08ec469d9483c6dd77f08024906ede69457adfb42e31c94055de7bacc0136f9e59fc4b74e5a92633c2039924cfe00f8cd03e382976ccd2020e68dba2fe48f53c4ec4f348e8823e2b9be2d2ed0ad4f008c93b39972e643e91ad06998ab52da9022b464012dd842b0229cb9c3833b3509bf24e021e67cdc61b21b7137dcea1a707af0ec43348c6ae0f928ee99241bdf8e0d19b9953c1235777eb5a9822cfc8e33aff746079c4dc60bd3a5e5c4b6f3b71464f75f14dd71ba3bb105f332467013af9a3f20c8023a7cf0f2722f4c4a22b2e1dfabf39ef55d1005609807db012e678af0553c169f70acb6dadd1ea6e619f68eb9828bcfd595053fcf8076cc7d2f4cec2807314e860b38ac105213b5b52de3370b867bf334583e4bb98279a64623306545bfc932959a0d5588c6d9986930e56e22181bb04fb02faf0614e1036a9e0718a99ff88336ac1c8199fc5b9d3995489ecc457af1ffb40342f48ce007ff730c15a7aa48a57441590f491af5231fc9c3ff877a7f7b62016e77c6c0ef4a207353e1440638ffacd04c26927cc5ac3f3493acc29fa2b978bdd0dacb043b93279f6d6137c3b74fc3f7c9693477999fd85dd13b0e0254904636f707c68f606ca10a11fedee40634f5ae19ec48baf95c271b26a5b6570b2fbbcea39c94cf757f3d4e9cea8d9f5445667d056d5704e1ab12c9b621fc3d1056223b9706fd0eace0c224dd2da85edf167dfeae458da48e601b879eddddafc4255ecaabb2b032074002f3f0d6a71865c55dab521e4137d1a42320dbafbbf7612199faf724f618279d75de90bf52be46d7f0e0aee54d8c65a18791b7eb61c534b28fd4dc7f6f55c7164901f771fd6b3cfbc4c0a05474d5a4793142ef3612184cf2087c53b01d7479477645260d8e8e5f1b628b5e622c94d5439d9ed14fc8d3ff2a419e2941e99c786ded2b190dabbbe5943477b71b5e12ae939a2c935d750a3224400f4afe8351b8793863a14657627e26453787f86ff2a1dfdab5d95669c71076cab279beb59b20c0b0fa79c4bc27f4e0d85821333af00da384a1d059b53dcdd4d74cb6c58e55d574490cd7ed83bd75873834a94a5e0d083b9cbff6b6c0990c421ca36163dab52376af2e4da0e7bc2e907672f656080f841d6f029cbd22586184485f08eb71c0b80b24a849ab1bd909365865a5cec2105e802202457b19a08c44eea0eff81e631a623230e686d43a9c7dd1f7563d0a0b4b3d1d224dd090b834c5b431e8cddfc7285622fdb55f3ecc1fc4f6f84ddeaeb13cd779def55e5cbc59ed4f4bef1b26bd4a491978864ba0482e7da89a7ce89fd57d40ec0d02a59a5b2048aa147462cda29fd5a295d25c735e0d38196a7a49deabbe7b201b0dbaf381a3034178cbd0e5481ae027cae0d4312006a85fcaafc664f9d608c5897a938a4bc48f8a1fa7b847689e02e85666a3ac4c1a732f093f0ffd11e509abc8bbcde8fc28490f2e8f7fbb2d56cb658472e9378f19e9b0721960202a2d489b6c6fa766367d78fddc6035e5f1483588e6a81385f6125c4fe8fb3a26de8a014c47843d49a0c35eff55acea305bc7f834643474a25ceaa4bd56137d61c6a9af6de34fdf9b33c69caa40c980ee5623623472e045dea46f6f2d2b47df611a75b5c2bb3df9367ad87c5577a4d375e1f731a65931e759a0c31962d67a98435e1c8a9b16c536d32f3306c0e87838a6dcea014892b6bd76abddc29bc3c54efcf67b7c84faedbdf9d148d298915c968cb16382d3635ed0ca34c1956072aebaff9be2e5ff963cb976655bf032e88be98848473632c3ab00febf73746026391e0b152cbc5c634d482c151b35f328b63d72f4cda737ad9f9f3e18f1b9202a7c38f1b13ec53173a57fc0ba4e20b2c150cd5f13ff5c9f24756cf31bc9d1d64bbd93f968ad6f9b316b0d5c8519f761fdfd1e39a2d076d17beb21b51a3bcaf9bae0d453867b9d8814500f781dcb472d107a8ac43647a3c6bc7f8a698d38b1f49f1296f7c5ae2b674875a93a8c1ba99a9f471564ab762cf25de1632de0f15bf73c082803c4301b56334a4f14957320651ca141d3e34f8e0706c9cc424d9cac115bd4e23bf5e69055106896b38bc0d0d312f992ee0d92ec30fe0b9e80d3c0bac26a220eaeaf7a8c5952ea9270948388de568775b93978642321a22fc7687bb94f9688e7b8c995fa9bc170fe7ec05ffdbacd166415c11d67cf2a40cdf70d8f7533e37c9cc4676c4d25f8a95f520b52e12cd3daebc5571ad4ddc53c9858775fcfdc278f2a1e377837e0e23786c7a58ef3c2961fb4c7ed02836fd968a1118bc855209b0843a1ec9ac93189008121f03121f1d92836313875da7db925560f943ec625277cbd1a58d7fcc1222c80fff4a7258be4dacc54716033680ea17621dbe1ff31e5d1c628f21558bc32b7f49876fe6713ea5aaf794a8754ee6ca19f1c8c735088ac70e616de034e06978924e62ca14f6409e7de71cadb2beb2be5a3b2f791f726535988a83da9543b1bdb77efcd16172cae0f8674cb5bcbafbc4243806da67cbcece2fbfb446ac683959a2d5cdc983ba2891c86a9f7a968ee0aadd3c7dc86c15957d231cceed95edbf5a193a74a46979bcb78897873f99eb33e27a2f4ecdb0218dde6be21c4e50678870301d854a120f8f8e072e97e3ee61b4616b414d0f2631e2f254c36d802a8ce26b2da24d07e57039e4257f591bb65585e64bc30f0c18d141bd524e0541a54481907f4514499a2b5bc91a6edda638c19f51d3ff48979cdf8249c069dd627684d8ea905d2258ccc989dc7804f7cccbc46f1b7e4271569a13887b8a8e589a25c76225a2d0544726e472efd8e81e90d1ba9edf9caedbdaa71ac47acc6b03b956b8a4f2faaf4df2e6b26ceda07dc26779146ed4d0a475ad1e42223fdbeebed2fdc65a7e22a99755d68fb94625f20240746d4a06d131d4ee61dc2709538ff82879b170bc09532d0adf72ffcb3efc5bd7faea4ae8260ee5970433eec53410e2703143268d11858ff36c5e48224430f6b411c858e764f9bf0b0e6d359805b6ba6eed5e24f7217c70e51e1021e44cce9960daa763d78b6e816535dcaee670a52005a5721cff7807d16cb1f36a51dc0bcaacbc4cbd0fa9565852958e1c867f3c755ea949cbeac95f8aab1eb1972c32850970fccc302212d449506d130aa34f8f77388158804aaaf6ff2e2d325752471fb28630f0590ee2f0d6c837d0b560def64dc8df6c1112b622796d81c5210461efd2f5f6c9716d76c333cad6f1e8a9d4fc5e9723de57b35516e063f445c70ac4458d78cf029ec1e4d1de93b807d12e4b155e26536c603977ea34a63c5d17a25840601b3eaf0ccf2f2eb4305ac9717cab484c9105a618acfd72a2b6a3bc0455c54ce84612890724bb9b07f55589fbb5588c65dd7a43431ebccf5641d661bc22257a221ed6f3f4fd29bd571c4a8a0d998b208696bea658268671df8b6ba2d81ec01574e4213c410b7d91b2e85068a67df34da3740b217daa57658d1fbc15450337151015cce9e21ce4661f16f46597f2f067470f81d64c97b6c0e94f5427e8686d74ac4bad18ad128b980c6adffcd924a2e24a0b5772f33b8f1ac7d083f5044a378b081f91d3d5cce3afbf37d636e65950efc30a545546c935d19594d44e82492c3d8e8297e42a839f1cefd80c0f2d5ae006d983943e6ded761631b33f006f54d95247bb4bab157235ddb99b3afa0ccc21d2d8bbb1ae8cead1fcbaa0e3b1bddc6132342a976001f473bb11aa57e3af9dab1014b5c8371ec89ff7b8554bdfc69953d3274276768f2dceb60f58aed35012dc5fe3cfcb2d2cd2a4115881742c2a2bd62e428869ffcad3819ec7b4da215749585cc2c74ee7f9b63db7b1c9c06d601e5c0ca93c14eab633c79ba850900b9e021ad414ea7b36b9ddd389b98397cd56da6cce24cb9e30410fcd935b17d30421956d08825612b997fdbb140dbe362a8d7117d696369b52c84b787abf0acf483874ef0ba9365fc61acc3a1daf9f171b5f1b8495b98f8326aa77694629bff3109d022b30b4bce7248ef70f98f3dcef631a6210ba742cff92f69531e6f2f8e7f8b4b33cbef7179ea08cd862ff34e90a5e23acaeeae1876a82a1755ddc8096bb7069a666972a181b94797ab761109500078e3714f02a427d05cc02bb87ce42b104a13319b61c220b3af70714763608e15343d368bc91486b7593f01e66dbf30825e4a12ab64a9959368b1fbc4dfbf1db8831432fb39def73a88130e7b0a3be2369f606ee6010f31666716936943fe55a9b6fc9b0931ada649789aaac6bd077eca06f23ea9c4dbb4cd5f73818e828588b10bc9d05f1011d695c1b48753a29e28b8816272fb8115261df9315e89d709c48337c98006dd03dd2f7857aff87a4e152240212210c8963a6ca70f9d140eac486b2359e1541de0084ae2800efd3fb2b20792ca0dca604f0bff3940b3fa1f7239ecfbbe711a4c8c28972c3ebeea5717d667f10bba90eac5ee36fc35d749c3f05038a06403cc45a2e183a969938bc56ab8ef71fe0ee9e79800f3f26cc619297adbac444368ee7ee2b1fad5755faacc479e2bf82153cfacbc48264348e3b7fc0b1f03c6de7c867e01164a4075b5afddf11a516b17ad26934995f7fe5148e5feda381b8aa0a839ced4ce01ba96cd80b150eced09896dd518ccbe6d29db847aa86261a557c352bfc7f96bc44494e95e94276c2e0646497bfbb5ccb958f4d53439bf7e7990881a0601c7d32a0d04b78de0b541b52f54626afad7a56e8fce3594df3eb933cf168883668f72e5da8156f751a2b42accaeff2f9d401c084cb99fda1e9bd09b2c3ce278ded182bdb87ca496e2adcdd4f5fd7851e6ffe706c4345613b92bf32e920ffd51d7089fbf39515a895294751baf3d014c6f2b722194ca2387f8cd54122d9a559729d0760712725a29bb85255d6ecb1b8d7f6b567a027a26a1ac1596927198a8899e73e46a9dd550cb35e35e86079f33b4fa44913b38c6fb09c11444ebffde28418d9a7166422c1bd91ad630fd25c6bfd1f314b950ac231a1985320e39ae6561497b0cc01ad32a6fb9b90f035dd43fdfb85779144640127d52a6f656043d4e5f9939d252e514cc71fd7f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h169d0303f2fd86b773edac76585d5bc18549903db2d6d43b6ab1a5db59c96316a3485c8fbc2bd011afb8b86e6277c32162ee8632deb805dfb3bd281f52dc0cd06e207078e4deae3db785c4418feeea42aebc763c89929a247b658a842a8a3ed7f4fb35d6ac7d712bd3bd2d6b30135839aa8f413a5eb256c885a5cd369cb93673075f550ebd98808b960d61c5f2f9c340af7f86ac34931be08d0004452308656658512a32e9d8b6ee734f614a42c72ce94c8ac3c94c36aacc6d36acbcc6dee9a07dae99ce174764cf4fc48036b09e438b6a1daf8063347af701ebebab83fe7164552c29d30b7a5c262dc4e9f01a6dd649a52df3687172454fe77d7962f204a42a11d42e7861eb5b57ce3b19e0139a193f249778652f1ea6b111c0844615ecee5f6100e5ae2fd4df4daf8de8b1913f673c350d92f1e2bd0b24832a1683d62ab153e540245b2e455a3610d9a7cb8dba1128757b1e060bf26a33457986e5d68924a75003f74bf7bf0c5b9168f733bf66006240ea64f04f95f7d76d2b5b8d1abee65edc4b26926f7efe53fe2033b31fb6a20c0ced4f2d785adf3d9ea5d9b66fef84d53ade4ca1091a02e2b6692b39edadc062449ec59c0032a4d2bdc51e50869d94a86a47d35c1c7301467e6d25055e716ba3b932eebabfe7581581ba89509c5e31e2c5c0dbdb34e1117b1a8b46f69d3f81d4698f1c1b9c062c897af07ca2d77e301ae9089aea694234faec5ca9fcd551456ae00be3861897dee9e3fe2c4ad969dfb912ef3745c56cc4cb0c6ad45a4283eb61eb2e58b1e4207ae5805c36c48eaed20f0f32e7b10b72dd5e56ca6f1c9bce24266434a6094e2e8cd64486c22ab547d73df2f83f30e685de10981fdf040d633e7e3fabec32c9ed97563a5946c2b145a59d9103ccc7769cde20f2b22265a40aec949cfbb71cbc230600935325a982dd426597cb024a745b83260d3036b61139624a189cdfe41c1f4b15e57e401118a7e7b37e9fba2216723b7e1084f8f01812cf5dda404e7fe97fa6382a32173cf4e1138fb21439f61d477266896c6f9af237f57c26a70dc3b274232ea5aa5660aaba47c31fe384eebb798bf036b637f6eed8c30277dfdd2c5beeb13b230a85699bc5a96ebedbbe93c698cb9184e1425beb64801fee46b2c501c52e1f7973010dae43826f310318ddc4def9385aa43e3e39bbfc15b8c5ffce2a37d3354ccef57e812b84bc77c67b738cd178d5046f9b406fda4b1eff0a2f2ddeea0fc6908eb495571ce6497ff8bb6d6db09499b79e2b7bef1b5946d0d75929bdc5b395197d7ac12ddbe7ef454b5822fabee92305a58421aa745915136dd004704d6de15dc2e47125619ad015988c0bb425cfce5d91e7906fddfb3bd84649e3070b2f5937e60dcb3e68c52b2ee17b7fee68604ef6ae2f181941ae4399c518daf61e4708ae0d61d81648d008dd93e54a297bcb38fa2ebd65d43ff4bcbbcc893be9ae40347ff2802f7300dd64eaa6b16fb20dd46d741e886defc507437a50531060b8e382eb7cd5028eb2f95a1f4788036ce628272525e90807f672472ab763527c7e24cc06108ed0a14e4c8fc51d9b1457a00050721cf3eedb918f80b88ab31b51de51849d050dbcbb6e2e1e88ca908e38e81feff78ca6711eb57926e58c20e8b4fdebcd47e0cbec09214fa6d3daac978729b4d7a134be4afed8f5b604872eae0feed965f0ef0eaf65ca64710a5ac8f19461bc34e313f6bc10c3349cca3f48dc3cc349662f57d15ebd33afc3d73006b8f7515f5cc472b465ac7d579acab747d811dc43cf53309db869add31b50d39a65975e3743085054a118dad533ea33063ae9f86a0a650d1d2b291b4d1f816d609456e4130c23cbf3a044dbe200ff4cef3b6c60955d5d2fa6c208c796839a77f44f4f6103f5616a4703e23a2f72efd1921ce06703ba47bf03b2d17afd6955279f1d6a04ae323424259337d0e82f8a3b89b67c172b87e88ed62180d9d70f659500d3f3562635bdfd85f2aff9a8d7eb19eb529b778c4a8d293857c8c26a590ab15c1457a86b0c36ecc1f9e22ceca104f7422c323b53277b1a61b335ef6febcef35b4c4c49fd1ed80459110af32b14efbbe21d99470f19b58fae41827d659519cb1b24fdc9bce1497aeafacaa3187815186db65ef7030fc53345bbcd2f8f5ea7c2093b0705dc6558ea41be09851d2f683172cf449bca6d3661132f1f3e89cb6da42ddbd87aea057ec4b8ac97863d7e4849a367d3db18b926f0051764fc475b22ff8c5711cc64a986430d7defb902f24befdb4259130842cfbb075010841f3a0cdb686e44c9bc95bb728401b68141b8480f502fba12e3d058ac43f297a31ffb6e27bf88082764d447ebba5db2a98b58c35df27e6f85538895bb42252eee3317e1155cd97f0467812c24782ca760d728d42a7db7dc39227952a6096ccbe21430c3c0cf504c4652ef7bf66b373939ba58024ad30c3cba362a51ca71c5264e675ca7711d6c7d1be4b8e24e41577721c6260ee9ea814519dd2f8322f7d48574262e8d0ed63c7e3d7e235672e85338d16d291646b9353178847b99a387247b01a4a78fed275db12bf7d3fa266e65b75a633c85cace4a6cdd2ea45dc0824d0bfae1582313b8df912db4633d4f4829f263957378752360881d0c03b7c32cad92dba4eba0bed416c920916460b16454fdca745214581e5abe3b284d6792105b917973913f7556501f8812f3f21d249ea78378657edd83ba4b93cec5cbe7e89d99a763ac822a7500bce4d821f0f70a3350c757a6e5983cc2a644573ba358656576e2222504819edf81d6a273ac0112b15b86b5c52c50d2902c6a6d977c4c2214d615896c2357b4bf04b86d4c299cab4527b9b04449da86569955708bef62d9465e8061b0ad66355fd5be5a8d894db2101ed74c22bab80d811ae78ce742f623cb737b11287dc06bfc34e789b2c0a5188bbb5dc0b778bb9432e88c1770e1cbb96a078f7b836d99989b494f324cab55359abe8b615c96db31c9ed8dcdc5708ba61ee7b9ac42fe9b9f4bb2f102da406b31671c39557f5aba62821fced48a7aab980f168b20091b1c24664566bf1b685dd3c3c08a7ffae171eea7c21148d2ff5bb8b17e7e7a221e09e1423faf1111bb86f3f9c57b6c9e79fd5a54d5b707b8166867b74b296da50a483abbe9bca57283a40a8e8475606b9cac7db955c09a26e953dc974204dff33faf3b7083dc93c34aea178d45525f949979829bf22624717738b63f05b9fbace979db915e5c8882283a1b091206ecb24771f0ccb4457198161d01a9e94b17a9090ddd9a3497c77f3b39a24654d6dd382cdc506e2fa48d47663b38c53276f450a162fe46572cdf3741060da17a9b704eb1196c475477f78efd15a16abe2f0358f33af7d986fcde20ffee613e94bbf25da7ae5ba449ff89b4cf6b317446dff6adb60b4bb43621b398816210843e8479fea6bb710b4fdc5855f109131241e06903e7feccaea1e9dad5924e9dcb076397d2b8a80570e8212472e329774bff68d79256f6c807525fc656b88b67a12e8521df9115bdb98017e9e00442aada160b383b345bf90c33d9ba127e6114f1ee7dc38e806d4e23e66025641639c72928e72441b50d0432a4307f695f68ecdf34ef01fec092c1398b93b4777599f178722c456ec09ae21809e84f6c0d3a5d032369f7dc961d49139b14c536d91a433337cb4da7e48febfb88aec719794d149b3808842d846d191fec768c59fdb467630b9ff05d0ffafad560ccc6cb42a7b6a3404bfeba54e3898ca07b4ac0f1737d620dac114675c70e21e9b219d6a32111b98429d9bc819f59b5f9d848b73ca3804d70c48cdacdd696e4fb1302a1d16f6b0548c545fd5cdfebe8a88183e3ebdc8585e6637187f23b48501da5465182ca853b20b1b8632e6ef2b5f508bc1496e11f6c4cda966ba8a20c553d8af47b78529e5b2c989cd6a0a333f0c984eeb86d05cc10cd57288904c4a6d95138978a4c80e82839f439c084edce5e374037a536483ef881f7d5e1f02397999f1a3c77555713cb8a0280667fd94b23aadf3e831b1e495ca2b3ac27b072c77b507a6780f6db77a42a22d7979dc8a7a9e4ed62ee94d7f6de4b8c33b07206970a78f68e632db37d7fdbd95c76aba2ce716b7450c5cfddb55b6bd874870063edfd5e7fcff61a1ddb50fc406d92ab0e0aa06fb429768d4eb48dc0245e688ce8d55e98b97e10ec59d4b606fa412fe37826236232137058d863b504124787122aa364d33a3c36ffb52939f8b83366a2ae375021e96ccff85937c6aa0456bbba74210d5b980da612d0decf7d9cf4b3905aeb2c2822c3a5fbe6d00306a0a8118ab1bc5d63ef3e24f6514d7a52fdeaa3e1f2d4f82dc232c19f9189e6fe3f54a1a6bff62d2bd283041ec7a6817d678a513aae84f5a41a91f562e08f3b0552c45494cc50298c552a11d3172306976b5804dba3d00e22b2b3f2f04e9f1f58cba86f1637f914080600ea617ce6015b573a9b388f65d73f83cfdb761f746992226728e5666ffcb57ad862b9b5b622d95f62ac1cb352d3afb2bbd1b7ca2c35d3334e88fb3acb79c08a439a488861611847e0717695f84061c878dcbae9692e3aa0a760dffefb708804f46568ea3d56467671e15e1caaad0d50e010b10e0ca53c35e2355e4bf8072bc4f6d93063c11eab968ece70b2162278a0887650ef1d51117c2d5a95b8034cd9196573215c8cdc8a636c791212b506f37c34385ecd9f5632407dda5d0fa876175df821b102b03a2a03deabc4e84b2f6dee80ddeaaf84bb6c191e9babfbfe4f2da24c88272d4653a0777deb71436e55954be85cfc0fb6680e8ff5058488e04ae9a863cf41ddec9cc471c57c2021e2da56727acee5ac019ca5238957cdbb361ad9aa18183e9ddd040d26b48533390b0b58f34a812c4b2f809ae432f616db7f95269930d4be7ca7d499fff7a412132312fb40cac5686d821dff48701674d64c625347835c8ad525088d6b6e40571b78fe2f35f248db32100a39434f731741b5c5e8624e8bee2d3b9a4bc86fc0a23350395049f7b725c50c7e67b4b201c2537fa05570b3567bacba91e2f4e3039d3c72afa633dde0f2482e7dd98468937c4ee7b1e0217866bd1f01a0a05e34d7c55794ac730b6e6ebea2efb7dcd56ee2f59ea293292d8241bfe9ae925876c7e726a27447dc33f2a03fd7eeffac4d258389f09d7eafe66ec3916aaa6a95dae5299e7c76d8c0797d1b3ab5e126e02b2838e00492356c12b0b82626ef3bfae79ac6051bf7b127f589279bd39791fda27c6202c28d7921cbc7e03d2ab8986f366071f5386e7c0b6d1d25c1b09124096f8849aa622ad4929379f0d5b39cbb705425829e709966e2069fa57e5c898779b6aff29c6c38a66f3b8bc0fff98649627d4491766919c32ef5a586a323046246b2f57687f3ec9198cb0d2c46ca2bdf3f9058d0b12f6928499cda271b759edd4fef0ad3f8f86c539f66251d8e3df6c866ad23cd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hb41d4b55ac58ea2b594ab0ec864626d6303ac97ad8535bf636c3d1b8c2bb247ee7a675e0cf4caeab0793233c9b2347265a3872cc79c86ba25e92fe7d19c33a106b1f3ccd5c3725171764e18c2296fc4e7f67652e6b17fd8023232f3a07f9d1d0c9b2873e8d561eabd0db6721ee974d2c6525a669258c96b340306decf6a8eeec54bcacdb2f64855a73456865ad34fad12455b070e689174f86c329bcb13d1fd9d8e08dfcc87c30163f7de90d6cd3970f835645e113aa1b4cc089cc56dee112c285e98940579fea147f8a5aa56a46a9c41fb3c4b079985df726b34a97779ffbdf23857b051ae3c88474dbcf5749e6526e38fca769d77c4007e4aaa330dcdcfe1e470ab7837c5f6ec9ef9c03758f3ebb816ff19fb65d62db427a4722468214475874f31b7db79c4c84099ab24679a1e7ffc3f2ac495d88c444c8de277f33db3aec024650e2cc821456995e98fb41f2e327b0349c9a55add3290b39dd0d304b29ef129bcf4442e58f04ca91dc4eebc22f01c599efe97a2e72254fb398205357d1720bed412cd84081484fb341e57460c6e3f32dce7078a407710877ed4fe8edea9135a81d7ea9dabc4387f93735caa1d205e7caa3a277225e72e4b88263cabdc7da00d1582f9e2c0d137641769c2775d548cf095ac8b6e5410832392d3bc5626ec0b1effd99f15dc527415d70286c57dab9440a721ae71af14e14d11d3e86facafd3078558a57338101149c938c54441226cc93c725c16ca3a2468385e627082cc0d85f2cf96b727c074f9581cc62942924df5d8e1dc097f3773b2b7cc43409e79bd71e068240aafc5cfc9d0bc43aaa1afcc23ea8f17dd00f1ac35bc61cfc3d7c046e08d5c789cad14df321f07289e4a8e1ec2309d84e91fa6adc523548fa1c03fee0c5865c66ac704b264b6b96041fb0c361ab4c77e1c14d1c4fe88aa0f6ce7c222bb94cd469713a2d23431b436d6c282de7a44ef396f63bb7bf1108c5dfd08f3b3cb1a872d5f4d4ca56f65fd6e990588862038ae06274ddf40de4e2d79f3dfa8f6dc457c4af8c77e7b9166562a1c9cea8f8a32eea7eb0d522a25462e4e7eb2acb2c80274062ac6d8d6fff8e5abe09a4d00b68708031ad90da6a50e9e235ad522883d7162d025f3641c56dceb9833c29e3eda8ad1c2e5f6f5790470ada1ab85836891728b7acac8f2ccd506bfbf36c9fd4f30fbde6a1f509f482217569fddd328e39753660cecd86cd403952185783161b07acc7a0b36d34ab3d1799e2230c383c190b9c34e8d7c0ae7a922ee7693c3a50280041b8a55a504cd9889935fcbe7f6f1102af17113bb2bc8918ab9583489445c13307a91a658d8cf3a88ac844dec951880fb085e8696e6cb8e893c039f15e581bf09956226efb9d0fb6f8ba68ec3e6f70d0559d80c3de92fc1ea1478848ac0e8f5bd4fee112d6b7dbcd88a2a7c747a39f4ae2d255f5c005decfe9c059f6aba0de4e127e15786fe8f3a754ced757c55c22e7381eb400385da3f13a8d4f0105740866f89a98106526bba4fd4b180a79e42c01e8d141eb6e5f59638a2e00bb550ad84609e5add6bbaf1a859cac528773e6e3c358da0d0979da56f38bd682b18bdb65fd7360238cf0e118545a368ca51e499fb5802e700c943f398cb909fb54e93d400e2c29a9fcd75b6b0788c2cb56b867c4fb568f1c6837fa746858d51db8b69a07e71e0407993be5ecd0d5c2c944f2aa79fbc8a0c5470f23d4ff3a1922cbb09898a62cfff9fce0500f68a2699462d5a5f37936c7f466b9def01da49ba61afcf390300bad08a74bd70a7b9db58e5db31583b5b661f12edf8307dff61d38aac0336e285567270a2a178758340ad55c72abf41fcfd65b14546b59c6d1f69722f24ae14bc3e33f04904f453cafdeeb57adf8840f3c3c9269189c9aa19634375d0502497dfd1814b0c0843d92a25d77c4f37751bc851c3ebf309fe461048fef069dbb2422c697d527093a3e670cc01361ae640ac4faf767e70ed13f6d3047ed03d9508e96e5f58eefa09aa55718fa3219ce9926c44af99c207451e714b1ef93f9499b38c6c2804b66657bc2891281dadf90aa8c83dc8e9c5e0209866b17d8b3f2e05046432790e4c76bf8c79500851413ef74c7cf9cd23e6184d41670526c90153e297af533a635b2aab926fc4bcb1aa0868adcf7bf9e2d77a5d8bc68e530c5089efee6af6fd77e1770f2a9a9c873499d7c7963bc0b4a38bd4816817c185dc610f6d945431769833484c9cca94d478e8ea7eee3aadc3cef7f5ae228148f4e025e527f58571c88d0c0d46d5cd3195725abb4821abc9260692b8a7f4116d610fd21c54d888812339327a35e373623999adff58d035af341719fe6d8bf0cbe489d5b7cb1741526ab6ebe2613f17ae9c7e425ac5add744e01eebdec3bcf038f677a43e4ac0d6cf8fa745a382b9a2f625d7c4051c7a3f8fd66c763365e10a020dfab6ee25e2112cff827ee896126d5f09b9d7c4952dccf34f74025212f7dacd4a0e5272ac13f5b86e8e0c27bb7d12bc3691ae1387f108031d09118410fd0429fead58c588ab48491c7fe57f6a66a58fa678d8b1b8c905be8d72291a0cb1f681b7ae810e4fcea84c5d90d04884ed512e5772ddaf9acfa8cc33d27e96efe9d878c328c2ee16345624344ca6ee0988188cd7b51d0e82ed86ed424c880483376aa4809e08d573c23345c1fb23b71637eccf648dae92b83225327136b7aee2a5deedc67f5bbc8eba6ef588c88ff20312088d1f1835489fc9269560cb31f7619b236566774b38be1302fc0af72a856786ef17a5367a5fc09404a9247c1643166568c4ae9def2d71c28975ddd35a05d19402646f5b4b310da57f7ca3d98091316124788504e21052ae050ba03238e51a09a1a57640118433a89a63293fd042cf3fa6116066ef17a49d0d75ce7824642fdb45219ead074b07382f759934720106bebbbd22bce013e3bd30be08733b6d8bfe4bd5b3c17d1e26df352c7dd9a8d79076308acad4ce68ac7338d3741b94d8a021d4d467bbd03a49c27337d5dafdcc42147aefdb93dc15749ba492cb948d629bb8963122e190428f1a30e921c0cbbb898be4b73fe0d0324a166d66ca7e8cf4688b44046feb49c287657e5df1f61c4a809b34ebfd1ea3e6f595ed4061b5f5c922b8d5131471a2bc8fa933eadd286ecd641ab37c25679bff89b2ba57767efa0a56370e526255712b5d8ebfb06117ada8d6ef143aa7dd1a51496d91c553e15131acf9b438f8194b572289873785c30e17eda162eff7cbcc6138dca05c78a2235e0642e7ba169acee8adac84f1e83cf45b4983d20f98cf3faf72a1e95cd8ae842827e8e060df4bf139068d1ca4876e16ec5fa1b508401d008c6a99a4d4a413d92cd2b2cbb911e5ebf574a50bae5d80293a218368aa675199137616f5471ec309017858c90e22821a95b8388514fbb1eba73821f2f7817990fd4dd17321829410f696323fe95f3e646575cb4e07f65bf9174c3afc635b502a0bbc176e739481828b55f667dc05d543268bc324c20b379cf4132309dcc018065d267b13860100612e464de3f3cb40e6fd3800909765246537b311de659c94ce4036d4e850d0b0e5b98d683a98ae079cceb12be5ef5ccc1588ef8cd932d3c97cf0985ae562f72e2b0a32422a5b46315bc33e142ef6426fd4bddb7ba41de0076ddb675727c4801220b01bba9ad400be4c2e0415d4d90ac7c752b00f0807752bc9c25c6e6a3b4198ac1c812fb4fec29b7e60f077bce96d751312fac122fa3b0e50ea5c8257349ac24fcaca74e492982b9907d6c4cf5933f3877753dc98130cce462613b142a0b4ff2d8aff309deaac397db75e7ff1f978448876efd67366096ccec92779dd85359365ef8e87dab6bfed52b473c57033e261e1b8dd99b7d7a4417e8200cd9ed7810713cbc343983636e4f3dc4b75b3233ff4a2ee6ccaa87ac778567d1c1ed3c7980921342e25b19e590a81962b05aa0e5fa4ef46b94d6a4815f4dc873369ddd9eeb45865653c9b711834ab046a9569494bff825202818f70395d3c5e8f7375a199fc60510bee62664222d73a9fe163446e2a4ca6ba3e9687f39f1d6a7c02cb9dc2c7c627ce954715b5acbdb25cc84ae723ce0f12ab451589025592dcd922fa78fce1ea08135c2dbdb7fa3eaf847916977eb264ab4d1c06b335b5f6ae1f338793d859ac1d3a2ee3046a2931a53fe826c5c67f1cf754828c83fd7354d47366f7a7a5643062e81cae4c30ae54d7f62f3b3b8fbe855602b129f08bedf69fac6b0febd50b63b02980155f20d59f980528834efeed1544675abed54938ff7fd675ef8a77c9e9420aae80513a0b341ca3f55b3518bf1d6182ffd20b4100b5c66d50371ba55648a1b06ab7333309b5ba6094214ccc26908ec8956a8dd4054e8c8c7b6ad07712b8d834490a7da82e55402e461b7ce635f9bf51eeb90bc764911d775bc0c13b021b1a79510e72f056742c2316252ad3d50579216e2bd03bade194123fe0b2b10b78120b26e06e89ce945d005c01d3f670939971ac03b5833c6ae9f944b4720a62962c8423a2791835e628afac50af968bdc70e079870ff0467659f0d7ee384beea63e23c275685965a0740adb2c9c894e1f7496d4b2fe75db4ea1204bf1244041e7a66438fcc3d12d0c205e9ff366c04d5dfa1e576f54768fb0a16a296035f342e00d9059f2f8a2dcbde461fb69012d23f1f07b04c1d87403dcf7133c2028535e0ccb9a1e88ec6443441e2675061248fbb7ef5e2029a7119fa100f89cf2411e4c68ec75ce7d38ff93cf7012091cf989a98daddf216292c53a01e96b4a8bbe0b2932e23884d7333b2dab544c806b092a6b1b1b9ce295663108bc9a9a92114ad5292d497c394ac027f5da05ebd86467c625caff8c0f5a4463a67de57376a2cc8e35e285d14c460e2f3822124c04d8dff98eeac94f2f6dbe34f9527297d38af7cc7e9b1fe129c24d4a20e5653ab390137f8cc3502c005f8416467ce3958617f39278d9936801eaab366e1bd6d8d3fccfd22221b91d79fec9142c39c1703f1ebf7b6d63c398b09a8a32787fc6e332309b24b9ac87eba78b08986c4d8040db4375a0f276ab6c8c30d6fd4fc405216cb3acbd14cd875669bd783d0dea4cd7f48f3bbc77d51e14f9524f6babca2934d0d219ba972d6f6bdff3198d25dc856cd7d636e7b2daa4c2d9af7125de4bba53b2d63aa0d93315ffcebd804130d702ab268929825f8c135be332344d8af14158a46188a2e5044f2f850755f3d457ee264623d7dee4743ad177a0776789560902e22cb1c53bedf3999c1c28b4c0652aa998e4294e20709d8e580c6d1e7b77e1637b33e597222208634ac0d69c89e8f88dbf18aa729a0acba4263c8090f9e42a185a3f37fc6265f3564882db1309e35752fce8bf7a4cbf8310f9155121869ef65e4dc2d853f0b3437c5dbf01b6e1cafb8b677a9564d7f3f0202f5915d1ebd82754aa07b29b79daf334f97d0ea86d79d25f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1486c22b8fc409091c1284d787d6740f4e28642ebf7a3f7619383e1727c43d675f2efb0f4819b54142d211bba6b731748fb3a4a8a3cffae41c167dec1a64919658dc0093548c638bc7d29f9c1418344c8150d24e4cf3437f0ae781ecacc6bbf5c36c8416c0b20b98d6aeb32004bca495cc038ab2f898cab5c98dff9cec4ee526b58a9043c7ea7ac2134e12d6666d93a31fbee228aee351671e21b55dc2d70bdebf673d170af6f4b5b45017a8881605ac537654b40a83e2bb8354a59257401530a1ad86e77ca526eec82bd6b603d7173e4f2de27883397a6c64aab205b1df42bc230e297fc6a63dd1d3829d0644526f963e0ba1ed82c28f8ff77932c8a18495f4081a93eeddf8829470925cc4bc763cb2976f63001614d65ba3108896b88b2af931bcb8ed1a070d82a93361cd34b808cec1204ca42900cadfc7e822f71e673ea44c25ae8cbb1b532b7f23f344ad9352bd94c1ef2f9445d316fe0255d6a28b27feb0fca1c0cfc3d2dab133929e1e004c3c6972e0c63240175f6f53d56a4fb18f678074e4d718f3c6eb81297787b368fe73997cc12ce27bc8692b2927bd19f2367ecd0d86a38297decfc5b9d692b5b0a1a00c7237a35b3c1b5cc1b7d9f6b8329f34ab0fb016b31257079c47dfb46d64cecf90f8dac9b31acc1b0de54b6e82e357101ec46a049056191b7588b5b16ea8b6662f32b01b96a4dbffc8f1d3eacb915bd43c3461cf4a9d5fc6e12ea48d4622121a9cc2cda6b3557f00bd846162cbeab1365d483426226ae382a2b874d2279b0307d67e6f748558edc1a7141ebc2469ab8589078e195fca58e446593df4dcd45ae0f08ed0e8757d8545916e606bfa3400dcd6eb402276cac59103a16a06e9482781a14d6a32b43be77eec12dc9634193678d553e8b08791f09765e59d49ab3a212e022eb819b90b3fc5ddd836d084e2b7b40f5ab35736b15860cae35bc82cb29e6876fc3e50d55cf550d18c5b5b59e4c7527eb44ca6762b2724f920e230fcac18e53c51e08d5b0498fde1589e6808c577aeb2c06edf092b554c246a641bf419edb2b9d34c667e90cdf742014b216207bd431c61397709bbe788addcd830a21e969ebdc2f892368ae6e6c9479d637521b81c59c1b696f67f63b2ac7ada6415972c02c1c2c044e21d5daeefe0c7c9b5c7a1e1184d3dd5a3f0055ee36938434235c587a36d3c31d2c4f62176570b18c14ba34df5ad0415d3e9e173599c6948fa086b409c87ab3ad7876df384042f241bb4c5ff9763c7e574974284f2b78928bce98573aeb90dcfbda0d44b5b965de0b36b9119e1a6173e0f7cfdb282e05fe992b729d8566b1592f29d2b6e53f6e62bc0923dc4849e9998962f185e85627e53a058ee0f3b5665c5cea9d6dc3694c811905a7b56b55945439ec814b7bcbc5855b7798758a86489f953eba69fc5d12d3eb65e3ab9f4898d37d39e4a604f4fc27cf002e6c8528257f599a62bec2511d08997354b70f1af3ed6f9fae7883a7547c5f8b8088070d654c1f06ee2ca89779e36b459f828f643e0eb4dea95d2bbe5c6114f58f2e81c7629c0d27362f858113186b534f6b8aac3448f61cc2c09f7346a6f0c90db94f92aea7b0162e45cc308b0c8c5079781b4027eca69639d6cba90ea8c5afa9e030d4fbae5bef30914d302993468ffbc6eaa0fcb14b6d4f859a4922fe24ce403a063ffe5294a26711df614ad9a2688c028efc2ad4ee0e22e9a7f2296b987c334a16694517afcedda7735695c6f04b671447477e152f4afebcd0f0dd00d0b6013a92ac3bffa000037e40f1e400517abe59a678d69890e78ed9b0fa1a548322883936dd259532fcbee31992691e77a917117cbd1364978a4eff58528b8f63531f5f1818ac64a58e025ea8b551f223bb5a64eb00900e2e6a547deafecaecf924efa769c73c5b23670af2d9616ba9a2dbb9d82e4950279b5d5e3873524f2f165ffc9967f58d55b0d8dbb2e7088701e7195884ad3899b84f09dc9d2e72a24ae24137fb196624abc6bf1c727e28cb2526cd2f2fe24a1eb109cc6ce62357cec68fa56b019d8f3b8e75a0afa7459f03dd3bcbc424b8024758a1904ddbd03ea0d9097d3d7b81d2f28977e3eb5e8519e03fc8ce79c27881a9a71bd37fa2056d59779b7b0c4b4b67a8d1c4e09959aae7d89b6f43fdc335ee69d5becb317a7eefe5d258ba8b5aa1985f5dab791c9fb43729885c75c88a3b26b7b0b334b59b54645ed7a01e515559a94c57b48c78ff7af000bbee82c17995b52273e7f6c0d20d592037de8befd5ec297a5c214dc3b5cbf199c875e5c818df537d418e994aaa155b71c90b705c20792ee231af0a0d4397ea1e80eb4c62417aec5ce878d428fcd84c0c7f932aa715dd2dae3b6c6a80c43c29bb68f47ac71a7cc2f0301b9a1b2233ee1f7f0809a0cb542cc8d0c0da58ad137ebf93b6877e96fa28214b1a69f151d19bd03ae6589a914dec2f8b520e2c66c666aabd4137bdf070199dbe0c403403ec57d11556cf075ff861daac85193a0fd74b097a80566ea1058652f1ca06db133f185e189075e5305262669241e30b48ebbf09065ec4d3ec0aff4702c6ddf40cfad1292891b3c586fcb58b864d8b74e4c0d663ce27fce9945dd8118301a8f985cf50697e5dedb10e533ffe63807e3079ded3220faa5bbfa703a95e63ea4267daaef9b8ac3d3181700cb31b13ea59d07edae038a9344214cc87ac3c193e2c6a517b2ebc880f1d5797cba62b0ffd74f72386c49892807b4f5c9e87f449a1f5d0ce49309fadc402f5e56ed3b587b222934e6d7e1a884b89d4d7d68032e7d045705fc0fb26b5f8c9ac7dbd66d8c053572f02f4d6756e3f5ba05d57bf02e3231840b0efd138b9ae68189641d9e0b44de6be20d4d534d34844f6c84671058e2b761744bdd49cb6bb3f89e844963347750f870f3a9e776282d7425e8bc061e922e7ed803524da3c8527b81998b40ade70521ea398e7c39404c62b87959564c876bd38b3be5a5106415837f21b8cf182766db75031b6e92fffae578fa9a5189de78428960091255ef8aaaef2ae012c25b76eb94ac1532c8018d4908b88be016c3771d2a6d876ca0e6d517bd87f65d8d6de88ebd53d89c3bff205072bf70e39f9bf85db928f869f706a0acd510d1f3145ce93b691b87c6a8556f86c0602bb8313a9ee59451177582578bfa7bd0546c8a0827d2075b466ddb6d02e34ef001b83304d59d5b0e1637e74f9237d3ec45c813692d31b7ede9757e6a1bde139060e027cfeaa7e499381454049f842cfe32a926853828e25f95b7715c1f8086db5361ad0ca9077b72893be72ab49b847f659797469e74f26d6e9fbc1deb89a4a9a42a0ad510569d7e9a20d9d025df56e44997c9b188151a212d2337a4f52d82d1e35fa022b3e63f97f7d1d7d5aa0a3397bbc7d3b544a48bc039a0b1a157cec1c4fa63fa884c7ccae04db211af04963ce4e7abf6c3949fee9ba45a341baffad96ee3d363e099f2f72f96e2bfcbd639a84c924373dbaf5fe3443cc0028e919476fb924e5c8608c6c3d06916ae8920de45d5941d2ae633e230964f800c713beb04b5c0d68f8c461a341deb8826f0a9ee1f36a279ece5916ce3119732c4fe869609e19357efbc04c7be34bcb47ed14a569021d12625d54a261312e369768ff651f02f82dff932fe2efe57587c9de72f3986e7cae273a39a0db06be3b746fcd7c76b033cbd7fea9b2ca0f088563deca9320ca4ccf5e3f4099c7426601bf545aade8a6fece7bec34a1b3a4bc60b46086d2318ce0ea8d173b5e973943d02d758310fab3ad9ec085b64081585138a2466694bffee824d6884408abe8459f844ba4837e81af260b539b66a565b754a916824f5b87bd721b43cfe5c87c991ff1620eac5100b93585d4af6b0c802c7efdd56c0d5c81d23461d639a1404c24d09365021f8d0556838a7ac361af485d8b5edc034007ee0f3928190dcb1147a4fb942529a4be73d0900a107cb62d873982baeec40b96de1952bf1ca69bf5b1ff8b9663be6b6c8b37d20d78a22329bdecb1a9a359b1d730e5242d2e8bcbfde4c8549f51cde7fb82e9dde23a352b5898d78afad0fc712604cd6575d155dc07719b5528623c14f4bcb7331e451bf9567a5c2e72ac58ffd7ae776721e4d41b0ee9a7fbef7e1ecab4b55cbeb6031ea6e5eb7062b5c99b1862c492fd3fcf7f08759f266cb118103449b4df6ee2385d7b5fde926adf25b0bd9143f1906e51ce9cc830deb4bb34fe868f2e7a8faa6a20df2115972055f7dda2c683bad0e2096ed8bedddd285095ee3dc5b0da885909003e761fcfbd7746b39351077dfc864eb6aea0ba1b5a00a91e4ac5503ee7c033d128bc8a6d5af70dc335c3365c4dea0c661b9a2de9d37ff54f4380c92cabddacb41b131906bfcec33dfdb10642705a9d24334a7d44854b8e6dc1b0a57e4980588e9ba6b1b0d79743f8b43c11839899a5d87d07157391183ae389e6d727444e13191d68c282b0dd8bcbef03a7b478c2b08de484c1174c72358ba0a8f4d3bb199708dc6ce70dbdfa6d3aae4a0925b01780d6d3706a6fecdef605861e54ae12cb902cded907bc60a9e983e3bd8d2c1cd7ebcab9dcda926bff6817a6e78848e52d7639e36e3edb61e9cd36d0ca5359b3569617fa48118dac79c939e95cf4a7cd9392173312d47e117630ac52f37c5c91b7834cc4f832a6882a9bfa02ec7701c87ea7822de9d267cbfd9b5ef0a5db53ab96c8f02320ed39813a11c57643b889617293da68cfffce709367652fe7b211cfeac36ab920cffb7b2d9270eef334f156ebb5adbca3bf272fd2d0b07740783e070b0d25a4fb6c40ab08aafda9ea54daaf1aa3abe8099d94a203f11e8a0cf5f03b8a1c2b09954675a6c181f8527f69c54ab23195e1cfc61ee7f68c5b6e6ac8c6dd420b3301bcf1b8daa9fa80f37b551492c3a892ca5c0d04e339cba0fa2dfaefc28dca005be9b8572652abebec5e4a63e6b5f66b9373bebc336d124ce355c5234f7632b0832dff36bdf93ae7edf9f5f273c0d7096e24ee509463cd56d089d370376b590baca57a2921f579a4b4cd0e0ad296529edd47976b1bd6d7d61f8d4bbeb962e8535ceacb78b5225bc4c572fce6f9442665fd22b8b423c7c154f23c897a88600662822981e8e7c2670e3594bb9cb0d28ff8277894f41db51adda40e1bc41f6bf2ad0e151dfac53782acd65ca7b45ee74dfefc690995d0bfaedfce15b7cd89c75903d34a5ca669950b3ce2192784bf76392a1306bd22377ba350322c5f6fc332b01752360f5ddc930ece14b6aeba9ee3225523a4808b7832d9f308a68411f0ad87eac54d2ea45c953f4209a59672eeace492ee0a92dc2ed75371fcb36f382463d637e3b2ea4e6515cc54d459166d5351f8517bec115b39627ec6382f292dacb97827c11a21263985793a2270306be847c5c2fbe8ccf074bf1eb35fc85800659ba27d14d9783e37e388bbe13fecdaaa0ea42c5101e44f1de85dfbca7f0e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h54b761692b50ada6bb9cb46762d122bd651f61b453432fd3abbc8e2312cc9a492f176ff932435e8cbfb5907145a0c72e39c47fe59563ce9fbf3255aab6c0b31e958bde14730562eb90ec0e6b4f8107220ca16050a652e2e3181e9ab25a58dd0a52e850396e5870075629e89b8168b285317a1e67f8f24bc47ad3228d54fedd0e381a9e7e3d2f66410708ef143c6c28d6ee0f2d03f68c2c73fbadf6edfb50e723fe76b04e7bcdb0ed31739943d32843611112904b81c61e287ac85599150250997f04fe494f248a55f9c7801c408009bdb2cb5267a8ae2480fafdcc23f8c7ba425b014b38530178f18408d924b94cb90c1b627dfac2914f751ce21c481f93bd773cb55c92475456595de5ab72666c071ed2bf4eb2402f2e27f6fa343dc7862b336adf5eebc00d0ad2c32d6c768579f643fc87d393c8e6bc377d1589c6388c512df958c15690dc300172a040535feddf2cf8a60e3bbe7798b4ed04e1c8cd2592108020f607f0156e622de4666aa42b5978ab9ea79529e92be6c15fb0c3aa2c51292b0395da683897e62c0eba6faf35b845258752e0e6667966282450f0ca3b2d4473580ee3fcbf85f4ebd76e1c0785a8a5c5f315a0712786e6740ff5215a929f9cb72f359dee8092a0a7a1f48a98c492389120b87682990b58668c3450e42e6e91ca36ce8835ff9bd892d7069e9aae2ca12c3dd58c0b3ba47a8a2b0d09a5691c4456b3e09182ebbff0d184d4a5ad91c7c0e75fd6036ce61f78cf84e109ce6bfde0f6f0641029ed3b74904ddb2038ed668c4722ab49364a5849c1915fd0c7fbac81fb8808f03b651400f8016134d14df8c4e7b4a85772be0cf8819de2d6734976b78a3e39cafbd246b944370cb49cfce0ed9809748bdfe81f189f7ea6d3e2677345f70df0135ecd5bf4df9dc359d0994924a99717bfdde01e9da2dee1308a48c41f8b16e5e6c7f631b8b560791a9c47d31eebe96ff369a38bba79c6f8612e7cce518825f6bb09667736c0705423958f3d636da0197a08b397023d07a1d7de28648f5e7cb94a57449d034736d4d7633f7aa3d1cb8b12b21b6784199c0223c72c82a36cfd1886c13ea9f10dd62834f36e2ac72f6f6ae0ecc11c0e4d6f134d4c5f6562baa352ba2989baa95a202b2ef4ebd2e90547880b95f37839ddba252490aa9dde0369c1dd596f4c67673a5f42602e8c13a60e47e274111e72a35d5b2b0eec19f7e4fb3f655f055636440d3b5a5bd6c84aaeb9981494b41eab0931cd0cfbb91ed73395baa5dc282d263d48180067b167d9065e2c17d0ff651fd739358c2745dcfb7e2eddcb4e5237b63c7ef43c28d867a92b36b0e53385f8aaee3781aae58317bd1514938f5df476774444268fc7efffc9cdd0f950288fafa4d7bda36f50eb9782d599caf8b6c7353544aa098a20dfe42b2283fcec6b7dadc86d98515c10d2241075311ed0daf82df47b0858263c15447cabd1fd22a1ba5140236902942a11f26d517061bed959d962d2f5162c6ecdac1e400f104125695217e3b29695e84039e6d5be6ffc05f24fa1547f776412a5ad0c958778cdf5b3f3e3f1460fdbca1467ac475cccd2bd70f94387c9bd426c65000c98cac0b7f11e33508b900bbdd40d4cd7d3a4089ab1b42c474a3ae53429088d10a07d093ab0f9c284910d6a31a20d0948506478bae736032d767877c00b052adf8a1d88893de8e8c0bf227bc4fc203bfefbb9b05406b3b6d7c875909edd8df10f3fe4509b144e70471cefd8b22055e2fa1042b8a0cc2a9d4cada2d949bb46a0bceb16d1832cd7d54cf0bef042c219919609197757c5e01a2fe0b8fa10c07aa6caab6ef4e47eff8d0580c15f98c4b22c717e0ab7e29a415e80e00b87c6e3c6fa52a7f58bdaf552816131f1b860e95dbd7f023f36c43815e80aadf8b53bfb17b930856c74363ad0ddff708da5096eaaa5aafa4d41d9b906061762afdf5bdce4f6fd5e615a2c896eb35947aebfc54fe7e628c2b37aa5f4a207fcd260ba13e02815c8f4856f8753987c9d882707b2396f6d580c533a5696fe404e398a2c7fafd77dcbbba06633d4d7b9b18e1c21e45ec2db63ba38077583c267ed3318a4026a03a663914d9c5eae50ddd3661d518709782899a1fd1081f9a4414ba7b51a0a6022a153648d82bd04d6feabb3b52c86b791519d7da9b5c7f732b572e1ce43130495e11928b86fc1ecf438ad941836fc718dd68ff3e13145e3ba9d75bc76db58a193d2b74ff9cac2c47ca6a0bb04d94cf17edcd810efe75ff73e151d36945391bb8f94cc470484f22eb4033d909f3ccd948bb9dd6fd5825ec247ac61c1bbcf58227787449f2716dbfc358c23fd97b03ded15ba14dd1f1e13a28beea040a49b1c308a332cca3b3b9813611dcc2b926741f63f9a14e79819c9a7c9120ff566449623fe549a83914689203627e9c7fbdc333e2b2148d3d9f5cc30766fbfff2dd49d260f41fee5e6c9a990b5832ccc24ae92c4b55254c40dfa2eca4f35af8b7a1c6a71033408e4e77c6a33fe3f8680fce297a594875475811ced051de3e2bdbbd3692a2ec3370c6ea08f435313d1e4c5ee1de15e8b148c8b3f480742e2049b55e3665e8642d1fc21d4270217cb98226c6ec74530c1ba33e224eb8c94c1ef6b2b3386f7969a90a8f9659c6f3317a58bb6ddc4f1dd7f091166ee0a2abacf3ad8e8529aa09055db940effd644349264c2f26bf258bcdeaf8d634141d8733528a271ec11384fc67004d5888430af041230c2adac7c9698f0ff1849ac2b3a3cccc9253b88fbe0ba88aa84908d479684c1646b04f183f63dd443c060eddb51ff707d822274ac95f8e9c407c210aacb6de0f57d37411a316ad50ebc06f6bdca457d85e707c41a6edf0fc5ab3c87ae8c1ff7b3363fc28f47ac3b9219df720ef0427e29c655541f7d643d28d3b76c3fedb2ee4c8d93ba0df2ca3a2fd1f47a0f6ddb78a066ff0f2da2e200d844ab7aeb1117606b0d43d6d26e6210850d8d2b9e02f50b9acf8dd4c69640cb761a9996390e17b518543b72d6dd1dd7a45190ee10cb8f0417275a8e45389d5274ff138334d1d0a5187ccaae620f6e5e0d606ccceccc3ae01ed8526f519007bb7068cfaf6080b2285b475b5f5088f33b0a8499b9fc62475dfe44125c7bef8e21448bc859f02d59e2dd39ba5abd09b86f672f59fe0491229c6b7142bbccb0a8d571c0c1d51f0f6ba3fd775ef59ca8c07862ac1aa587e1b6fa2b649b16cab8d7dff7e80cf4eaa3c336fb5e7b747e729f9fcf492e1d90768ede34af1c740bfc363d9d879e2f0bd06c10af8d963c38bf38b96d8ab641171aa832b0d7158ac0f2f32d2db0157ab641810a94bab997424002feef83340e85c2810378a0cccfda8db36fdee1482edba91a6136712464c1ae2da7fd04124be7b1aef194c78c4e4c57428b427e9d7393e8bd756e7e8a842473b5773b791d5ae5114640cdc54ac3db65fd163922e06f452aa13e9fcb563e3d983bb77cea1cd872c4b5ae35c9ebc380914b0dc5ad5279fe46ed303aa2177f2e7b8dee13e8808cb98719a03499d12280ea419b22793999a693c2f9dd7bc6ff87bb72bb1b3c85b4b5458aec949a1c65c3464743590665da7d90413dcf9e3294101b4d9d4126114676b63210357b4b5bf8525c8776d97e77b467947baf5ed63dee6612b4a46f4fa1d31dc1596f61cb12335b927eaaa2a6608aa09fcf5f395b645138405ff5c598c9bdda9b9516fc5d38407246dde2cec256c2692fedc979a69215080fbe73fd18472733c76894d02783c07d66ed41ca13679d95bd1bfc6b91ccb66977d33cf4d4cf6dca18372099ac9a1092abdcac4c455ca3ec627ccdce41f54af795747a87bb489e7e1b6f5edf693af2cccb5fc49f77f1e1b25459469a22751644a658efaadfb86c0fecf3d440e7fe36c10b8e98588808567a90d9b7c044e8ec82a1a4ad18326aaf39de419d90d3d40ad8f12d83be91063120b739d4aca4225a860cf8f070fab4447269423f5e7b6b0e8caccb7f5172f5dd51f6d9dca58acacddee1b3e3008810b00920d6fb81dd5f539f4db1d19ff76e297a7d4acdf2bb57b8acf73691c9b34e6577efe2756a868807d537df1b77cc6243915f2555e83c7576984d99602fb2e0f62734b07ce07d0917cad1090815bbcdfe0be94a9ceb93d32f507481257118077f3aaa9cbc549653dcdd2ad9a55b53acbfc0053bbd0d651639b7577d061847b34478bdde9ad22d6eca71552b1f0e842b2f94f24bd9b3504679a9d494a4d55a6c87f70b02a85440383bb74443b37bb64a4aaa868b09353983f058b1b3fd4d7fe8923193700ad2079daab694882ec0d3712b4a7201799b2d820670066d94c6d38a42f6d2c967c0604ca592c58d096a7a896e6210adda0d6415f9f003d292fad38a419614b9f5ace88b3b14a3258e1dec19398aaf87fed9855c83eff0b18761b91ad4b9f172447a34eea143f43cdfdd445420b0c8149230c99da699c155e934122d6e028669ac84aea463b29a62070d35bcd8b769a9c6289fec43acd4d194a9bd13d622c75749999aa1e7df6dacecef4022ede23db47b6696acd3cd1d794550c1c76f62c7b09b75cc342b48c7b0f3cdc9cd726dda96f30bf66ba2ef01c66347918168ceaf990144cea2f05272c675c1e141e40546c43638a8fa5c48a47d05d06daac37e565b6fc9665c12a1d39879cfdd8d07a40ab8090c0507c19358909e2f9a53e854931cdf9627e3622e1a3a830008e480100905e7f3eb9e4ce1bf8cb7d0843dda014752ebc2915f2e903b333ac4f126b80b77dbb10faebec4e955507ae1d5c8a607b13cee45f022f930235891f2f4e86a322c32ea4b61327bf2638f0b98766eeeec61c79e5d1083978549cf3bd7ee45fa3d85c7bdc43153fe4d047fab22df19eceb5c4642eb8a9f5aa23d8eb4866289cf0e856a9b2ff07aa964ac0924435cb233a172fb7a8a4115a7e1fb737b80dd6ee56fc2d5c418b247bb33c2b32a22376d3c61a8b1b85f9a5cf81c1d0133b73176077952557245d6402eb4199adaa28419b36372b23ed87aa879cfacb6e0723e3df07eaaa5dca2a8ec1e99ce99d0d387ac9b37a68ce4e826de23cc1a981e5d423ba92ffbd34c2107b290e03c1a8d5205a3335cde8db0e8268f6f03418c7a1ef752276ec36c728543d12ed1c68588a92acec1c7ed3c65773ed899ed15bd86b75057ac0557a31d6fb3e154575583ffa8186e7ad86bc3b9fe47e887f4ba65b37f0ae9636075c5c4dc1c06818c6cd8b1bca138b747aa3bff4d4244ea54d61020253b550525f024149dc677506fbed19d959c91df75bb2f848f1f888c0e60267683177ad5bf1492806b800971df78f8be733c58a712cba80635edb8e6ae69662ea4baedf8de586c893bb07df3e4f70cde2b9e5c52666ad0fd7893b1208268b59ddfdff63272e0465d740151d5cebf04c1638e1f3ab8287666690ca166d0a5d964ce192bec072cc38a763603b965a1ae0d370aee01d575baac04a35d6646d2ec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h53d9ebd796cc50a74642859ab7c66046f3477171f6236829a5bc6906e4948c2bae23c3e1eb0b841367e3bd23fe8c684403c237f4099a1235233187d79b3217653a0e4f07bb6eee103178d62212be075bbd504a87f0f8b5bc1253915f910e216103b971dceaeab535e0e2363c9ab5367d1e1b2ed18a25eb22dbdc59d0631a49a104736a5b91cc5956df6d2c1755578920ec1aa1bb634a5d9367470d4e21911ab6b48990359cd6606f7b6dd1a25d67d625c14f85c2dfc2ad64c180eb95da6de861266225c73de6be7ba807868d6b84e6c27df4e5478d802caba3555c73d165607f429015a08db8b595e92efdb293544dc95e89e628e916a02e4c120c24a820ab4ffd1224cb135f0873ac16d3142bec7008fbcb1f07ed90a2e2157f1cd9c98fb900f39897aa7514e006fd13a2be45679db952ffff223e5ac96f235f535a01dec623a3716b41d224019df02aff4aa435768aaa1e14232d3d539b743fbe3b9e09894079a047d7e3e3d82595272ed9ef67e9efe92f5a013a33f468b03f789fe0e47ce7425267b9e753d407acf62e6aa09ff7b9381ca3b7653f619d88d22cc8f3ec62f70fae070dc90b48772de06cdfeef8da0ef5912e404bdb0dca8da54b6e9ec43389da67e4ef545e01156397fee6335c412ab6e46d8c0cc6c872149962cdf62b2cc68d331ace4da7037cfab41e4e2823a2e40689f5775e3ca64b7dc1160f0a10f7c583e0c08e20b1077571fd748e71dd48d518a5cd2e65ed5e70f4b208cdb678d196d7bcd0b38fe13fd9c685bed4d2478f6c95465ae3f018386c1a5c9c830707b27f7c65ddaefbcf613f607285a9fe27a3b3cad8d142de68ed22b005d4e9b1035f127c614ba18006a9a9f3ffc4221467132ebe7edcd5b4b119e62223f8cb98f6aade0d43bc536b960942602b1247af04b573c351e62db618dc442076fa1f4c6148b2ee33984b54973fbfb4babcd72304924154eb363a5617d098c7a17a20fae68b1283018230bfc999fcc59dd133c67c93dc3606e157bff3ea15b2f50e776ce4e50c2b01596e30419b844e24bee55920c9e485134311bd8461429d6967560cd7d058df19f3abb1fc8eb95c15e62b750a2ccf1d8a03b72fdd1ee900f9da8e288c291398975e7d114f70ebf8453c169da13e26f8f383ddc4f853bbf088a90f190fc0851093a56d46a334e90df18aa1921d0f91a0d77ac81a657df212c0e924a1aa5c65ee7bcbd5b807a9015682ed8ee3ca7c403e01f8083493a0ef2f79304da68c4bc0de87e42d16323788b3684bdc192ce9a7392ff53504b1d6384667429801df9a4cfb5f360d33a5eef4ebfed120a96ea0c854335ac91573d6b0c9f784a5ed88b2e1e0fc0c5c49f0c6265be27dd88ea0d0326d9b4ab54da0a55a5727e9801db44b72e204676022ff7b4f28073fd3fb8baa28fb25e9d4def42a14d9c213ba896dd6bf6b4995d1666d5b45ec8bec0d2cf767fb0bd5708ef13e11dc2189e5055c2337d76941f733ff1e88a173c7253ef01e20eec63b29b996cc81034da7cf3ce8a253f6b29cb41a6ea51efb0df213a3ce955d206020e685c781258b90f154761a620d2ab0b54fccb93100012ed958b47e4d21058283c35a9c98b3848bb923551b9fb7493376aba4315055cdc678fefa44e841a3f53ba968be3a82c0c09c3ebc33421390d0c85b5733ef68a67813ec03ca95da66b24e86d8de654e61574f6bd3f026bfa3c7b3fbb4139780c9d6f9f0f300ee6dc75c0be46948351fca0beebb0f43adcee012cd1a55b0d3dcc4d7257342cd8b6cd19160865b1dfc9b8e8f726b6995c1625903db8124b9412f8f82999e66dc80af62216ec2b35ef316979428ff40601eddc4b5ca3ea512962af6b0cc53795a897bfdc90116b84edda90faeaf152e6761b227b640a525bb72cddaba50717fe9d1056962fb4142bbbd1ab539c7f65c0534a370b99ee2b7b407af99c1f6d38100a9420a2016da127ad099bf79d9a8f7f04afbd551d67432838ca3745f207544030795c286e097a7411db1a9155c862ab4a34a0579f724827bfb3a0e204d1bd27240f77efdbe359d16f54cc91bf8d37c96c1d5157fbbf5d704d70c1935ecc1c8f4fe833a4607adba70321550e1411c4abd5b396fef6aba07b73ff607b6e428789b90f97e6a1a7e2176a0b5b9acbdfe32d39aed199518693439cb372754dddb3e975a3ed55b5482c07464e21986d4121aee8d5998a40ec92cb1d12c79a84f3cdc35bb5deee99fcae1345766ffe0fd610fa176ed6d077c86576735a76ea589b7a0d98d638feb68baf2a339470cdd60b84bd2c7d797029bdef3bc840a3dc039329d8f95a11645943ee1f47f0befe4522c058b08a6ff08bbb2bb058523b6d0ccb89918deb71a02c277c00c067adfa13a27e192846b6661e285db0daecb6722f89307c7e333efbea989bb0df2fc8eb5c2a5cf17954481535f8675418c938c86276060417c0fa26cb1798e1ecc425e37400c4d82ccf6da81cdb77fb01e46ffc3c4025d5b32dec9f282865e217ac99047b83e7795ca894789ff4858410d9e9ac55fb4da402dd6b5482313d8de92c0d09fa41d16083eeca5ff5f9b707e3f4453fbef4e75841e6c0d2073c6fba05425d71eb259626e255a90fec310239d4dd3d10ca235c9acdc32126b6309b61ad83a231e7b9259f9674fd1ba1c972fa0eba3a7b331eb554aeac509a645f50881043e6b7425a283a229ebdb222a156daf354a7a24d05a8d9ff16f1d92f4c70a6cdbbfb6f7f762a0f406f24028ede16cc8142ce1cb5db8926a343c47fda8d06e0baaf2b9366d01f9d611149248d165129afb92bee07fa3d4e16fd0f4cc9f57df9453eb271b9a38a8189ed1e331925214193a542645b44cf916545b198b46c749db43520a37b681a4fda1c662706eb18ece506768a7a6fae3d1f74fbc07ba71a9b5346f15001d79cfed16dffdb9c3b5bc8cc558f0abd47ef2c0dc5c1ff5e284d371015cb8fd3146f1750cc918de525a1f58d244141d29d2730edc752104153f383d058ffea34c67fba8bfa8f03019c436de10f307f7efcf282c764cce2620325c59c5a3aabe8477a67ded6ee55e09053003618c557bc0c77f04c2f4c102d4e5319039f36acb05570b51c813904fec635019cdec2a09c61270c1ed5504f6426cb4771981585405d4cb70217fadae9b343e6a031ed7b86c4e751472c1fe0d78e22ed22884947c3fac56204cc2c905575c59d785a047cae330698d03e050600c8c537594592f14bd43a26623a1e5dc46318284133ca76b110773d8023b07d261df0253ce038febe387f3bfb02fdcbfb228b65e4a2bf1d6882bc8df32b7fd47524f8785826f6b4d225c85c96bc9527359e63cde5d97670886905867c3f2e187f0437846a030a7b4a75e1e2018226e938ef83860dacbe473497b63bb5835c3865173ba3fc52f6c9045bd7733720f6e64ee2c3b7d149e648840daa313db0a6ffb43906a08f5b23dedb789cf8e6e8744369bc39d1721254e0a04b235094a4d32f73d4ed7d9a89e2b9e5989338a264a13536a019c8de8bfc7b7f3c10254bba19949c53015af531f3c22a78799c8136e62c6a6a0929ec67a5ea64950ec617366d3de5f2ce4a0525f96357cb14df463432418e73c095c7de6111c8bc1d903a49bf0f298107326141d6109d5f0071a5d35e6733b5cf96257755d1a33152a3fdce4032c374dcf547d547f367b490e576b784a9a786222245cbe28f429aebcdee642ef32257ecd33b8518ee6f79594e7b6e302e4f50d75deaea9b8dd18a49583e630f536d7c3f4c67acc42e6fb047597b07a589a06b21e4c4862cf1dc495b0b95145c55a10e4d08fb19ea8517c3a17a998cfc3477519ccb61533201b38f480ac9be8fca34123e75aabc14a13d158207c11f83b172cd5dc71750e714ed893662ef647564b179c03f8ca9e05dbefc7a1d4d4b92bb4bc8bbe61cbd2f7dec651e3a9a72a1454e14e69dfe2caa9eb75c67da62df75a526200f4da4ecb8e1fb65b99717e9593f6f68358dd6f3341f0124685c3a9576085187e7b4233df4e58a9202c363aa0c94e15b4fa4dd11178747290b2f04f09cdea37ace841e50392068db999fd517fa1e20a6f099b664c06ad722b518b45ab31166b9292b6166f29596b19b19ab86f0bea087f830c88f7b2424db7a78cc71266af404aad603e06aee61382246d7ab45de1d147c0869b18c1182c3078e4066c45d196d1724ce1b4e8577cc005d7b441c90c07a307bf20b10bb24e299b7c2a04e0d876658284f84b13d17ea373f3274e9d6c0010696db5cbddaf64de588049ece4d88f2b1748751f1ff3d41b8ae57ed7627b167270aca85e49b83e599465e7318fd8738273104944c02cad5bea56efb7a096c4727b06b3047eb178d2f98b31978a37935cfaf515374f504cdb54db8f311b166e4cebb083ac0cda08595615574dd40ad3bfd077d05d7d1d09c4f92438c19918b04c777fe170e6823f38566cf33eb2cc5d9f2f539e105366b32e4d664fe5f3a9b1dd559e7445587d22a01b2331fe7539c3232f0e5f8e3a34ab64188631ad7f2ccc84ca7c13a13aa97a128037b576d6da8b56828b4ceef8fccef0dbb5f8ea3c325943fa3426933e2e07941cb8ba84ae9b7b3fb26767f8b8355653113d0e8be63f5444bced55c53e8c455b0347a14d65c941be83f02cd573435742b66669e111f90a1e9e35b981f9759bb838585cb8edd7b2d92aa77f813ee24466062fd4f1ce5a104e5961e57ea1c34a9e15f4bc0732677098a13167fc8a8dfd3d3a6a5a94ec34d16a6de1c318650d6a4595065219f045f5c547c8e7605c56604f2cbb91b65f402ec46d5c9b3c0e502693709f967cc444c6b2445fbd425493c636583ec3a99aa27c48f38a2afcbffd23238c3d8174ff6c73a5741af09857eaf94c176ea1e38ca495cf02b1ac13423f099a4fdadf7492c57ae59fbf9de3043d7c195e0c50638cd6051c8faac138d89e64d330203765c9888f89f119f9a9330d591cf2499d521352a359a1c789d565cdc3fcc50dc0deb0b4c99ce51bd70dcdbcdf6632d413855562292da6e6ff5b0664bc0f169723b4ff0f5a6a82e6ec0ff1bc80c5b63927f649a2e8270db303299782faaef218cdf6fa457fd7f5914c936229ae57c682e3864b2ab9a8d353b31e71b312490d180b077220ba81136c813958c2edd00ae67442a1757391ca226fdbbdd8fe63b1e6a4f633fcaa1554839b3e99700744fd90f0c81cf6b8e6c9be4e5752e66fe4aec042e09ff312ba749aae5f4f8dc3d5cb3f185c2f5d288c365a0a1f6c8efca28e8a0142782a10dfdf05f1b7dc81fdfc046ed7a58fed9a87723198df84225597d97ed45472b9665efc619708bfd6234698e0a0cb2f5fb917fd6d8f8b5628100012bd8109a218b96852c26c4420b55a06ee30d85b0d66f9737fd87a91ba9f8ba14183150878454667bd5e05b9ea2389506a393d0a82fa41dd2fd33ee4587834d4c6283ed58f735ef9c681f3dd912c17484c0c04ad74;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he8492a2d208cd332b352b57c38eaac38d1de6e9412e7dee7d582c8a7946c6501783f7d8b0dd37be699d5f90d0306058f9f5c08732ac5f61cf6d44f7c2fc85cf5d359ebace2bc68aae80f8d42864074bcec299c4d5b2dab6f06c1634cc576cae0cfc29c322baa3f663dcf89863121b239d26e16c540bf68d5cf34b9230f59c88831490ae802d05f328758932e2183a859bba5f928b95370595a41d7ff327e25f012b8f220f5c4b9caa8a771564d5427af679f2992727b2e4740ced918cc4c04217e0df5b08ab05f99d55509f3ef8d5b2a4f3cec6c18750698c324a850fe9cc258b4d700e095028f842e4851688ac9bc111433bc9291f24f2adb8e0b8583ceaafecd0b0f93fc84dfdb303d25537a56efecfb36f3f13a7cf2e880b8bbf3eba0942ab3e895d3ba7a7b5f0f4400f20683f458fd3456ecc6b2bc127e4d3197ee1f72f88b99327dc4c26cdfcaa60ba4d43547e729a0da886bb4b6dd1cb1225b0965cd936084696a47f4ddd0342a10652ce19cf1dd6ddbb1d93d341e9358048141ca11f9669a3142ffe591054e40669fdd48970c846ce45da49f933c5b1ad3671ff9161bd49fe4dbadc69a6e638baa100fca89369a234bf90d9de2c1859645e248fa25482e5383db610c22386561fc7252c062efe03c02bef0987eb28e1830842cfd870dea1fc029e38afc4bece00e5617e2e5caaff4703cec9f595743985fea86db963dc49b441b22f0e9ad9177f3f2039b7ad89b5abadfd7c04de4310218039aee38c9d356dfdccd38932cab57f3df3e6bbf3d8b7312e59bafe9d0f42ea833672ef64f6e132a2f788a161d30c0ed0cd67457212c92f7520ee1e0c6cd724695c42fe290aa9ba552015ae08539a8d2fa34cc4576403c0527e948f20a29bf5006b84a3db11f46f22f730025aa66d84b14ae180c80ea1a88c5871db982085ec65ff7333e77e606a32cf044f39771e9d163bef77a047d5da3a15829a27a59f0dd51519f85d5c8730ea58c9727f740886ce26234fba802134610f1cd59f66e3dc2de933f0c359d42ad8a4fc29c4ad08b7bbe01398b2ea3ed7bdf0528571f7c64ef70bc8fefe706ca0debd883fcd05bc23e4611f5be2072d32c97caf8f90abdef5b78fd65aceb12ef411fe8fa24cd47a0e74565fa7c5dd4f663e17a28cbc57b9768dd3b84de71b2ecc6924edef4cc5dbf5f9b17e65b010c45481b2ff9af8ce6d1938d154d4e5507bb4d4ecb214883689fea31e69edc6648a83634251f89e2e4a4ccb6321af2680d8800daeb564249eced716c781da2a17fe54ad78977044e234eb57abf7a0b286b6350ba7b98b59254b4ec8f631395205f822f96448a44cc84dbbc425dfc40e2d01a48f3d07de8964a5d0665595c52d8a3820f20d2ab8e1552e308951461f9fbb7960e6a6877b575906ef208ebdd0a5cbd3b9e7edc899a9bcd10992efe3feffb5d3b664e9fb603af1cae56fb04b62afc916adfe9c7f3b41308ab222a17cfd166ad8788c9332ac982117647fd456a18f7508115aa538ebd391575121f17ba585cbacaad88b39af33bb3f65f8eabc2609b6d4005f383fa14e5dfefd6832f92c9c8d8b9d858e1804e37467ef615f8889840b2615763f778a2d87afff02596d3aa06e5feebd527afa2b5f0a7b8f27e0d965372b4e36295afe536c061dc54f12abedea3e40045776c2e6ea8eed1d68627db35989c2f6e83acbd455b0f373ff1e48716912516df9f76368c201dce45201bce81b4affc811872656392445b5d7ea55233eb82979792c3fa277a315e9a49105569575b3bc76463578ebfa2460e80b91892d78b18b0cb660b242bbf948ef931d51431b0b8e8bd94b9d946a87daa0d56aa9ad477bed521ed8ef24ccf6f59e6a0ee68e1f9cff183efcdcdf1edb5be79394db294dded5819abe288309b5c6af5995451b04b7eb8bea49b80b9bd601fcc822ee5f6740f9f677332e499d35668e14115a7589f4a2668959d6cd3e5bcfdad4387b6992f8af977068c646bcc6dfd212ee586646bf9adbeddf339892ecdbff8395a0e476662ccede67087c538400a0d8238d4ff253b0ac4e6282545081578cc795a50a6b3c894ed15c342f80b470bf29e3b8ded94fbab3889985dc2fad13cf55d164dd30d06347a8d73c9c46f6fe922e81537372edcad70450d761c4a9697fe6e14f4f03903cba488d4b800bbc7d3282a347416029ac9def04b4297b3ac79f5b69511d2163cd97e6a22c597ac3fb213cf41f3489b3c551d59a095dabd275ea66e2e10b08c4193e26a80d2cbdf05b591857bb24bb6fda7762faf8c9baa570fa0d0c7fd87a1f78fe7e16d1d182a44162815bf430c4d5b3c2ef98f5c8fd8a979d3f0e332d6dfc6ae9651060b67362f545fc6e3ba7ee507929f65a66ef4c2667658b0ab7559bf4ffba232debb06f26c489de0a629889df889aba2d5dbc0457f36fbc12351d2426694ca3b8e117c0279e9df21ddfefcd4a4152064b13e0eee549090451a8e7df694060eb6073ee4a8224dcd4fb7a8c6289d7e7fee0e50002734454d5fff811372606755325e87e3db02895a21b0097ebb5ca3eacca654a013d5b79fc77b6773ef714ec8b5067ccbd4469e207fe14bb840cf69b204cdfef433cbb2003e61d71c18f0da0c705775e9704ef306889597a052ac1a14828649de527676981504c84644cc060bb651ea771e4eb5abf3bf05f431b874fc0411e6a6f50e793d230ce508ed55b5b1ce04e6e5b7488085aac6e8e838be7e0d8d907f3b23681d2c24919a948fe889f08414dcf9659b07e555065bd865c50dca76f0930b08a3027dc80807ae3d008f9655005ef5cf4677273567fb5d9341122beb8100e6d104e1d48463c5221c00d48d7b1fe3c44b19dba061c6db2d614c811f9ccf37e7f55be039a8b7b26f1557966e66f38cd0add2e70b8de277995da1be093faa04ae569d8613ac9fc320a8679cb67e860557afd2eb9569ec833ee11bb0cc7c3a0994da38b95fe373d8dce66daa7ddd90d5bedeea3b729c13c8aceae685a23fc53c246b77dfec2a98d69d96ffaa1f192a24b41f422a97391db1be86492031f84b86422a0fa3ab73e095514feed2e850475ba771e38c5942ae02b509d4a93a5fbf8a8282d565479e2d3082aad49c525c3c288f58cfa3d03fe5f898ff3c9af12653be12a8a530dd8f86af943b5e38930b53890d4c4788778eef8892a7286638610ae6975ab9414084e663eddbbe1beac03dcb8eb76f61c65286591f198d6a788c6654bb792571fb485e06d60f2cd396da0aefea72466dd07e86e23e3b4b610969a23786760284fd353f28580fa9b6dfd52a4cdb44c503d698786fb16b649e3eed640fbbde9c954000b0790597a4bffe125e95d93e79be956a12866b8aa4cb1cbabb34e92238e13d145721adfe4eec313733bd17d3dce3bf7db2c00445ed8a2d0cca23df5d6a3d8d6d09310e02c9a9f4547e3db404ccea6b3d561a22ffc442a2b369c8d5d9a8cc273efcb91767ecb80e3b0e4e0115e33502a18495fd8d393f80ccbce4683296b582b6038c7819b97864b15ddb8e9237738fec4ed1e55521aced45c624576abdb9be3d93cec7f250345aad910695524cb2d35b1eb758142d2760270489c4fac755afcb6d181688aba91cf585d2cc214398ac275f5287adb6bdb5692672e51ac89b1140b0104c8cc1c9c8174f0fa0b89b1848cddc6770b196cbef8aad28f556e1db2be3d83d47d1e81ff9e0c3d7907afefe58c4401839eab72392408f5f6319e54b52f42a69a5f8f10fc714969cd16ecbaa62ac80a429d10a3331bed3833db046eeaca333190c9256898e7568f440a241d8d0a644b6a03f86e92e731c810554c4bf102d20653e5916e87ade0edd36d054c6950f02899882cecb4bbc650d0084cf0c3a4e8682c043dce82f223bd925fa82955e9743e62afbe8a9e78501b051b1762144b9e4963d235dcaadae7ce3855d895f62af77b61417535597928acff88d99d8edbaecc40b0fdbc8b4faeb5b2af432f19e5167606f59b94be8624e4a2e46afbb4eb97ef00473fde5391ed0b5522d43d5acafd1877ecac23561d5e2b3acf1fee8de5b08ee2f1124a6e8bcaddb9a6c8734363bbe8f5072243b7845d3d38d319041c13604b4f5dd4344982b3a913b8e89e1783b09073e3c159c5d4c958a58b8e25a9f0efe20017e807c69af587ea454f2ca77af4010581d06b944e85b4e5b37c49162d20c158dd0d9377e09d8cc803cc2e251c9593ca637760953a5803afd08dcdab8dc8cc4ef83f93e1b23d299e961dbcc93dc3ef6e93bce5fa1a7cd00b6dac1da8b75baa743681b0a5786e4deef3f4b7471713ea1b3cef3f5fe8c5e5c0b3445458e492c02224a8be248343f0a26e456572ec7cde8af458142dd3c25884c49e0416b2bc7b9f0af0dd333ba879221fa18ed81029fce010bf6783e2e507e414e81fc8e9934278b54ae80d4cf521975e1535ee671d5705b7cccfebd2c2df71b6cd79edebcc267d45f877cbeb94309406bb318e39bb79d805b5317ad634f81d4a588c93e25c0cfcb7f7def4599cf69ad7dce5ea03ba3b43b5ce8007b4ad6a956ff4160b396cb5c307cd12651bbf81395ab2ea72ed68bf3087063160a6957f7c67c67b7219c89d171b48149e8088a1304c1580652cd74c6bb38499db0ab1842cf098d4e112c9fb28fe011d037ede7d4420e440a1d050ba8b1f88afbe08b8e6c7342eab037f3f5d1b3fe0f494bf2c1c8156526eca2f4d2976511adc43aa5f9fd34ed2f6b5e803f05a889bcdd0fe89a12dc48fe9aca04080242b1c29071ae535108e0f909c6abc2d8322a6a29fd572235f62b4db30e58a8673895587a30bbe75ffdd087cf3bac1994c96c2fc053bc7c55b199e34044660845920752e5f4cb3608cc3a476a6b450b51f22bed97a1827f45cac4d1ea12a687320ea6e5f91017d3c3c54b7f70040a7cfd100b2331a4f528546b7dbc12b07a33b6f18c189fde942ac91d5a3ef643d2dce3402f626f61ac36e05ec9eea9761b9c546c684a11f982569aceaa9bbdecf3a07043f6244557f8dfb1d8398f5560584ee89b9e9ac19c4b281322ccf75e90209503d0dd0ce0a9d7d26788bb95c092ed14267b434dd23d0a96dbfaf4e9e579874d18614b92dc165962b0fad62ed9d7011286ef4b4cf9a91f4f4a8d928b194e7f2ef0f2f535c0b744e4f136003187e18692af62424f5500385d2300e97880a2fb0b74bca25952fa9ba050e15d45316d462802fe1d08fdc26855350325fd9d706d7d7b947376c0a8536f64b5c31f7585dfd409f91e9a342e53e6db949653ca423f321eeaa95886d5c8d02f0083d33b7aceed109dffdcd01d2c0798170a6b880cc729b0f23acdb1874f64b9481955ae857881ebb3e500fe2c85da4ccb0603b5575e1a28ee3d2bd742e94d93597aa06bb73a624833ed207a1610110a3ccbe1eef39648edfe52255ce8554262b6e366798c50e1569bde04fe4674088bfb4176d1e5c7796e90a5f7010830f9da16ef7299dcbd7c17;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h216c9bd0cefd31a260144de1400d30229e02900c63d8aaefbcfaeacd3e5636c1c18a4a5484b247fe9c1054941969b017abfc4a86118aa0ff560abbb144cb436f4bd24efc96f7c5b02e4d0508a9c964feabb43f4d1e7c53e0f6c8d38a4f00128cc8a6ec28d981d2fa638e1c6b6cf6e3aa2782cecf9b8964d903701b2f363831fef00bb66f6ee02619b1532e106b5435291c3142334faa0829176269580480336c28edce4ee40f56669ad5c70e1d6afbfb2a078c058e7c2abd93cae0a1d4ab52ecb1950ac73c8f2e4c1b66188eaad38c7729b74f807d01d8069fe1740cbd51bf5d42b4fd4029c9b80abddf6aa393e1e7134265512c13645b74b848efd445f0efe5b1e13c30a7a554368e9d6136a60417a7fd0b8b700db49b5ffdc0ad201459948446c0641897008722935223b86251bce56d9705d3053178d196b843046a030d96c929fbca986b8484346e8596e9dff4e8f02f6a5cc09af87303c7a567ae564cab48a01a079d9efc104b1c9f66e2416b387af0aafe443525040b39f8341a65999aea6db0de411b1ef01866f81acf5b7efbdb2ae71fa835a380bd9cc176a287402f919cbd30ecf0c807b1bdc2beca3198caaf3ce4c67d56f308b5dfa42d0815db228c5dade758f4bd078ceda0a266726a4ef57dcf29c36f82565f13ae908f3086ae873a6137046cb0f0194e206b168d932f74548d1751a1a7f952109d08d8e5ea74d3e2d8b5b7ba024d3b6c783f908ad12c64328e2ef149f0ae9402226b2f467701ad00ce1f7216cee17b92697974d5bd66d2554393e062dce74f4dc58b9399f3c564e4c7de93b73eb19c4a87b5a191bed0085a145b26794a3d1a96da5ccf98c331978771eaf7c9d3b92629e2fc8db7fb62a0553aa089f647b13ef306d29c8ce134aca9fb91d2674ac94272f55e4041bbe8e71e7bab4a3ff6cebfc6406998b8f307864a04f50a9ad9b68f9f1606ac9b53bf9b157305e76f83d431d8a4eabd14725358e06562bb7a5dc471874cb722e92c218dae7bfc7f0c0b79fa9a71746d85ad5860e3d545d0f1c9339ff73c00e29af9972b90a0febf76ca2b5efd777f3ee7a36c7bb6e1e7c716dc89526aedffc01f82160f1d195a6c27ccefdeb2c4846589dfd53a3c5c44ab7e40fdc547a4312488fed76956ca7d56e508e03610f6aa2d72561cdf24cf8573aee99068ee8b77edc0d4525165224784182c67b74b32d8746edace93792e3ea6207344a0ad99ccea600827eadea97c84c942023fc4ba8268ae4b724ccad2f8b618c1af859297e92fce216139b5d4d9bb55154e9fa03b7e962ad6ecfdf5accb6b4d163a62673f1f0320d73394637fa86371b62f45074c02f20c6e5eacaf9e3681ea4b5e110f49ec37281951594c40276f35d9b106433fd5c60869bc464af48da403a83fc3305d5168d4d92514220ac4facc7689df1a3f503a794053df44647773caadd5ab8d06d98ca29ff38e9dd1c6bc1daf56c77cc4646d2ac96819c6d980faf88b668ee6363cb478957b0cbc856e5031d185e0f4e2d4125d9469f42853b00bec11b74e3f26e0b81d1abec566fc40fe9c6092967e360a6b585ee9b294d324cc29fd00f43c3615dc62f42ca5d8575160540286b166b9487980c950611d1ecf6f1db88567e5b1b50568ae2f843718f4a034c071cd90d6adc8c8f34e50ab56ef54f2443c536d940a6de443e15de15aad23354b57ad354fb2d8c29f236f52b491665c1e5d73a02a1d7d92d35ba88dd9b5f9798a05b560c443ce0e8be1398970a7288d1d7c6d943b6afb62d21c30789049a401e7eb8c136808c61ad589d11fdf53439675fc379a174cdf20f39d7349e85d60ef40274dde232170a77b20870353ff5d9f3c640208d45ad03e9dfd3395cfa3b921533e86e9320a01c888e462c7da973de9d7399709462251b718b4da3772d46e3b0d6dd922fe953190cfdac6aa33e423c892c786bc21021b973fc4fd65375f8e1ce41a682475af2806f5b6cfb037bc4c04912a117921874da17dd123f61f499d99fa3f9c45b7a25773ec72fc471c0863c4366fe8b057734d120ef06656241b3ee34a7e9b1f38665b86099d8a6c1b4e51e4c00d0d86c9c79a5acbc90d718eb144cbe87041507c4f9dcfa7185c9f49263e2fc935af14cbd8e8534bab286e5b3e93a05dc5bebcafd66dd5ba6fc6f7780063f87fcdf337cf1f3e5ae788f96ed4af4dd8f9aa7fdf5d49382f7677f46208859ef1a25eaf9820af3ab3f0aa9654742937b017ee1bb79bd99fab3e5e0514008ac1a59b0052327e617fa8a484ed59d71b5bb599cd1c7efe60c85ee9fb76f27f53af9b2c647c36dc7f55b0b8a34d12600b2eb34c426a93bf8aa78e7bd67bac0bb11b656377fbd39dac31e571fb9abc40ebb7e7ceb4ae3c82e46023d66267a0e26e8c1c4a0985cd6e11720d3e5be0f612c18fd8c61a68a5030f5be675d2d7c09c9e712af213e9d936ecfbb8d4bf70c4ce23f3788cbae6c4bdea271a974977283c495dc86dbcccf41d3ed6e1d9cbf737a71000373f2c08bfac8a0357074e27b5830e488eb04ba71b0ed1190f39bbf0e67108ef0c1f9577dd204f97fd2c57d3c1284a25dbbb96fba2d20b4801c1a37191e81ccaf26891cd4d4c34f3d8a2c678a3d16980678b8ae6da2b47b3bb7f783f9f4f955b6db12c965c8aacc32d32d02246b33730eab3c84e9fafd4b688c3ce28ec890be955bd9bc1e8fa52670ec282ffb546cac871c9f96506ed4ceba73c00e606176d4071ad642cb207358a50fbec99fe80f3ff497fa09f13ac4d80b9eab35fcafe5d8b4579e073ff7846237a20f7a10e16be3ca7358153cf59368da37033768d819665ed2d0d6869a4aece9a60380747bcb4339508aa68ee639d994960f07e0c2724cf739ac30b99556d02126ce639aaa4aa623c680adf9b4f1e1b46fb2d783e92d22fcadcb43a1a7d123924668554bacfd2707862dbf3cc3e0fcb86f4e2433c5f2a98b6b492e4d0c552b1a1de20a0c47349c21d43d65a47677843321e19b6ab2f94b13dd27566436110950354b0357a65643e89b49ddc894db24fe4e251bbedd26d46a768724d19453b7ab2198ae54bb81e0b2fc53a9cfe037374f22b3be6e358111a9bb7a2074b35b68bdff323022e3e426593ead78b9f5a209068c0be9f49c00541a96330d0c5b891dd7bcb3d8762dc0367dac7e92f6140a8a10aeff3b30d3486753c441498cf94a579d412d942820542c718a4e6ce6b527e26e8d4df3e869047c34f9b0b44e38752d40fc15e6a89a277c955f82c4a66e4e60814f7c8340e0be0a76439b18d25b55f1073e9c26d6437c4716c896372eba8945b9386414e8e6e1ab5b2eba8856bcbf8759bdc858d4e2cd6dec59a2d854ee22421444f2d094260fbe374855109d758f81b3c075c5de7dea57df4814e0f342d29336a59a8e5891ca4e8790be50de2f23a10a729fbb873e71e656436fd6541234000472cd0441a5f2085f5690f1ee7b4a8bb2f5d481fab5508015dcd673c16ecaddff6d21f3a2fad94e35543affeb599cee94eb2f3524d8cc1fadf7a5a25fc4311d95a550330530759a561a1ed4c24fc2ca35a59de3f33769aa0b212f993449b5f4327b692adbdeb7c4ef069817a9ed343fc81de154678e77fa527d306671fd24638220fb504ea606849604fd71623eeb89e708c3f9765a175f765752f3b396f4dd752a70396461f2a2ff2ed47258300e701d3bc8a03183c55fe0daa28857435411908d2eaa1cf92964f9e9a4438d36b34a05ec037f417cf4d1a591fe17d541bc5c3ee660f1a2732aacd9706da09f48e2feace85857da5b504ea41b947472d2967ebdceb530dd831f870cbdd4fc0bef61a3df368dd744e3dbecf804eefb9e31a9f484f3e1913321707433d36d4591989ffbeabe851e4d5f06af80861cbc6008e4d5bfcb6e2284aaf6e7075cabdf14dbec6dcdb3e45db755bb32c9870ca737074d3dfe81a228d78357ce75ff8041353478041ac2094fd67f6dbe0bff090dc5af89fb9402029abf4b4ce468e5ea3cd500cb74ec8d2f6d5c89bb3d224f81da8a4bbe0abaf2062d42a71a2813e1f9a7e805e604179ff6d92596965391ebaeb5de0168eaac4fc9b0fb8251868e6e10e51393e639913059ce126a13206bb05e0e474db63d895c108596fd23feef0008ea5db1ff8f1599185cb210f8f72f74c49214ff54ddca69c389f79055810f1c06c14f305a2c83619bd65bf03342605eb4acbda893036f780c4272044d837aa39a463be18d477708ba6fb3add61ce475deb1681944801aa557232b9b264e77c1b35ba7206827f9b8530ef5c6d1058abca0ea8a3a5ccbd988592eda0c8ae14f94a75adea11f181f79c9fa9fe578f2c75ba45df7de981bfca422c2c7df1c9bd47bbcc9c16cc91b1dcd71f077515803b9df151f244fefca8ef66e47ba6b70b7d4979fbee82112a38165ece27f0e3a7ba0e2a3e5cf8e420a3124c6509101a6e4811bc715a05cac0a6c41de1d9c18b285ab82a68ca06b3c82938e22713c7b371e77a4fb561e60c0e6081b8c9d881db0f8b840c1e869c19fd6a2fe7fcef0806682f52cbf5537b56da8a2332ffbe24101ab34e0774f00f0c2e6b7422117b7e3415207a68c228a01cb3f54cd35017ee78f8d2462840c8bf1dc8e11c813b1e8d5cf19ea852746a495838ca3722397c1e443aeaf5303718ad880c163483987cedc4d4fd05853d59bf0cc83ff4b2c74edbd7779be72f3bdeb418dee71f79642b06b18494222e01b6e04f078ac7fc9767186bf70c23dc845d025667e0b0231e474b91749fb9f14a83e7e576314aa12509663b7a6aa3649f208b6f656c7ac6351f6b8b8bd236797247734c44878f535b2519e9e5c990e2b37d40b5faa6c443a25c966641780240b38df08b24b393ea735ed8139b9aa9aa9bb02e985864ef3977663f53284781210fd4c734ab24e18f4cdff7db71b4792a39727436edf0819c3a7bf986565c65027e65dfacf7b3eb2ef618e411bc4afb72bb33f4ccebc866fd2b68d96d1ec77470dd70fc84e8a551081e17a24e066ce55542fce03d93df526017f34fba3b71f07eeddcaf365de61540d515fc819e3d68946868d2e4bca6c874af5a70e1aebb7bb8791d9465d68f09f20553a3d0b2b98888fa159a748a15f383646c4fa8b54ed1481d234f9fc2c1c7b618281b2daa20839f274821ca4ba10158393d8b89f04dcd2d6bb2092b82501ddf0a17085989afa865b7d7e4e516649e1c0e7957ae820fbde5a0fd057434b0a1ff08ccbac8470512b8c98fae1286de4f515fed2401190e25e4d2c9fa26890de497b0a08ad522036663f0fb4b72a04345d7b2af52979a8e5620fdf85b7d1131ea464f0559dba4146df847e990089416d69482e491c69d5dfc9227016af5c6140d33b46f0e31f96dd2b5e22b9012402568d691f7ec7633441ac24b1de60127895c3af89a8ba4ae567338f94d5ba4c860e19bc118b2812e80fce2c5df2e4a6c9db8512b951a7d614ce0d7c17f438a46a57f0a68;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha543ac14f5dc41895e4cfa89f65f3bc27397ff32d8d91a6bb7e91e0ab54cb0050942ec85541cada3d479200fd6b03a552d9eefc12143af26f11b00418c63ad265d69476a288dfcaef47608cca733149f7d6a587ec9ce751a36d13a7194f0e650189c055f5067b21a01e100e1a81604b1785b4137980375f0a21f6483c3afa650490e98296c256ddf218775d98f6d8398f90d5f6140429d7dad8fa8c849a4b2d86a3ad1c89bf4dd00a1915230d187858da3da31064966a90b506b582299f74fb9061c932a56b510f40a0ad7bfc7c28df6bf005ff125a16d744010e8c2fac5ee7e393dc63b348a094dae2169fcea9da895db617a1fe9e8cb19ca0eba38b32e65d1edde4c5cf2bc49dcb920e7a9c2f73594ca635d6d2526b0644c18a52312cdc5e22325402f5ef7bd566e645fbae6ceebcc484073ff5e3d9a1fb62e86e6b2102dd1b12b2e8d1cb35b312875b485dc81f1475a2402734ebc6c9c9bc83e5af3224686ca368e8585f6d22523af5f289de4c66e1964f53de8485f033836d9ca3b95658510231c74452e5aaf2cb80c67720b49d4e0f4fcf174b51498873a4108f9a6d394c86cae519fdeb4f44aa9e6514bb491fb4e3a1aa57f623520812635cc3071d1055750fc0797d7f2ac07b12e63d8201e3b608e8d1e7ff648b2ba9f9d840e11976ba21fcb7fda5717f5fcfd3516af58355e2d5fc7ac95472966585e205ee9333b46cab2000ffd727dda80291fb8ac60d2027760e478372ec867cd68f8b3cca85673bf53a4c07bcface26232cb95489199bc62759fd9cf23b0c185e606a375b6f16aae46e2c5a14dc9e6a9c2ba96c2db8e96a14109ea8228a1deccf2400274d7532c79a8b787741c68d37b8ea467bbdb664b9834571304962f9f0a79b8be462737899888a741c030d23ecbaa8028cc6ec61d4c240fe40b0913998319a93f0629f061add0e9fb420df5da11b5c99c57e5743d6aac72522fdc91f7d0cf5c5d8e285fa43e5527f014a38fcf878f7526181b002ffdad1b1931a7cb71b560e425f8e19c4197d4e24018efa802670ac5230aafa1f71d3b6b7eea6e91cf57cf8a1c686d39bdc4b551308310c57907a67be50baa8bce9630b9c0a4acd0f7a789f10dff25f237f9444876867cd0637b32ee3285e53756d9335e71117e5f3c8de6fc2d5339868bb8f645321fec2fb16cd3b132b536003469fb7f093ddfe92b0ffe76938bcbadfbec38ed186e2180d41fbd734713b823a6a3cc96d7cf4fcc64bdd7388daeb8dd1332e2134075dcceb93fa7761a6f4c473ed11992696ae1684e0b90066217f5fa5e0b5768ac435d7236aed07e6879f84bca47b8594f63754e50ce6969dd5f002c4a600b5bfb18d904a3e83a64db23e0ddeed5bc1ef2c52978055a5c3c482d97b232614a41845abd9c9705ef379f050ce1dda1e781c90ac84a408f5d6f9f7360d4b40c395f4e33f692a1b6bf4932b23b494efd91bd05327b2378428e3b1fea0d206ee3359ebe27b5ae156461777988b724356d3d66b64019b04413176c87e65c9cbde71df5f635c40b1e3a8e897454e72b87741fb9891c4351cf3b981c5339072b453b2327cb797dccdfac2f7793b7dd24e0426459185e204367c9bb1ee6b0adbb13baf91eb3fd67cc6b43d99ca3d06eea767bfa56efc3dd71af56917713683401c037c2f3a84b79b9e884ce7d39152acb31b74e071c4bf21f1a007f1f210ae9931142ca65d67ae0a906c5e734fb0fdccf02d944098a6ada8143cd6aca236193ce5c847329191614d541b2bb443e95ee78df47be85225b2e46ac7468b0d170bcca4c95f6ada583d140d68b221d66b5ab2a3ccbc527f2b06599b52cbea8866e17ac444c9388769ec2fbd92f09b5711853957e32129e665756c8d4077127891a7756eed40d02dad67c64d6977fa36828fe413face13157cfa691aed52138466207c0ad853705a6a2df3a9490d104b79e1bc1ab561ad0443afe4f97b2e2010079e7a6e170485a5afa291d0b422c439bd91596cb48a8c17cc20f28e600081fbe35e13fd94ba810dcfeddf24ce5657e337a7444d3f3e1d57f92644e588d29af434b4e1a35601f13c1a5b40cfd2e01076c3fe72c2cf533ddac56a2d6934f49c60cc8d28db016bf647e1704b545faa6c6e49485de9fbc7401a57609dc227ce2e85bda803ddab58cb1d1fb7d0c91dbbe51fb79226cc713640bcef4e3bdceaa7398c5d7d792d5c90ed83e63dedb16ca6377877b2ffc838ef1d7154127b462e1ab42fb45d42dcf3e6feca2aa5041d5c10730b1a13792752e753fdb1e05e00dab54266f3b03cac77a9b60a52595d15799451a5360e9d96a8ee2abe44e0a38b0c73d8196f4e0a1c9d0124a207fe1db21650262e0d6026b9f7b0946809d128917d314d9d06b5411942a24c32014858d8fc651967ab2e8c0b46a64d382c253bf00f5fe0599f3a89959d2f8f6e4b957eed87591c271d71a973255eebd5b4a82db85f5ab1d8f9f87160c2486a0a5a866a46b0bb61312ddcdbbe5dfd8e191c403c3296b4453d028edecd383ae5073ff4668503c826effbdc0ef286608e8de217501027a99d5aebe97e6873738a0230134b3b8507400fc29e045ddcab47d75ac28c80ad55293246af05f515e32a90f07d490d76e5126a6b3c397c5e6c409de91ed21e70cd20b5849180aa9124c8d4388434e90089c5e6d54bba92fc0aa2ab2477ad9b5287dc52f2241c3286d3251dea884c993938b57e863590676a86f98e9bf513855847520466b3421a42f18e7342c1b1165db274d224ffa314f615297fdc7942310b1295282c3afce9856565625adc6c2edc66ac0b9c45a29042032ca81d2f5c7195ce044c52cd6d749eecccf5b38965f622800204460a77b236b8478ffd303274941af15056fe2b80319729e24c37aa7191e4f894cd790f234250730d885756cd76191ed3f93956469c1bca87e0755b7bc97576364bdb61ba5681a2f23880f20c9f9ccf5157f59d317a197fa890f30ca5b80eddbb3788911788945744063148e78e00805e6e5c312e9280799b3897593bfa65cb62ae9f7659f3ecda8d8fc578685a92755a3fc8756c5a14b44be7d6edb93cb87cc89b1cab692ec85c01fb918fce5626bf2c0ae65d2ba0eba2cf1580691a85646715fdba525777cc115516941386cc9ea39dd37c201d66343cedc7e139a7755c2b8494d21c622294b4e7c6f576f5f93d68e601484fef00f56ea3fef8e08f0534c7695d0b5d06a77c1862da05617422619e90cec1d2c9605f1468c403bbd00757667f8a939bf61297706a7ff7234496b60bf4470043a0924efa247870f6b3a0dfc4ff45fad5fe29aaf3b93518aa1468782017ef6ba89aa9877acd713d5d67732752837b8153f3cf665377d32e9cc39af44733b88c1f886d94cbf580b68f99927859473b8d8476e011beb1bf11eac27be1bfae9874947d81d2a7d3d17653b4a4d64b80e05f947cfd4558d1e029c075fbc51bc30c20a23ab3431491eae3ccc8b5cfb5e468168b253b064e49b95bebc4503a001672574f01c584bf23190e490f2dfeb024fd4807dc889ffed241f0f57737cc067b63fc5983379a97fe1284415a86bb80b925f82e22a813be2d184e2ce1cda9a9f63ff45171cedc0f2c21a84659da7968efdd10d3ba540357560e8c65b595d177455f2e47a66646156ecda9c4d718d1d7d2de548bddbe4c7f5c3129ff896fba49b37361178519e689e669a01bbae971949381b09d94fcec07f8c5f928cc3b0280238cdf690536ed7173c7c03b9add26f2d467077bf28ae102642017b24620a554db3c341fb77e4e72916ecc1de75d5e4388dd1ca2f99708e1d1d50f802334013db2b5ef415e9acc65a6c722f49aeb7908983ceb09c41ae8aa06d51d989f6a5656846d4532519830d5b95d6d07ed5e5a66cd4d13187ae6b1c652dd2549d32f07abe3a61970c5ff8331ec5c15b814e88a779ab1663a510c26852e0220a62a563284264f7f9931befcc3efe4a51d25d3d0b08ec397d495a034fbfac13129f0f592ce9f755dd7eae0cd3be0d18e1ca63b3e70e529056ed1b71c58ee3ca3b3c443d646c44d4ad426c23a7b5b5264b0d582166fdb4c6cd3dba67683c86a41b7bd913b78be3036a3e9af7585f14fb37f4ab779af7733321856b0d4a9891cc5b119d9df559b3da4843a6fddcf48951c0a4725b0d862bc26158280eb244e490a16628afe92b22d42b0c32f4fd56fa4b8605e323b33d1ed0863fe7a28047dfb151acd7e2d7e592f064d2d1bb52bee6a31d577a9150280b48930526b60738b541db6d41159f91933411f531e90e1fee1a91ad14a1535565946198ddd7000c4debba74fbbb26e78d0eb3d7ae447cc2b5441cef3c54bd5b41c59a5409249fc9ac50e3294caf87174986c85695ac2b96400889b7f8dafef0109f58b31e50497883c3b029a2103296a5398e62a8ceea2b6245b2450420573eb8021b3e1c168ab27ce2d2b484e216c27e814c225c6f4fab2064bd73093c5ce83c859129f1f67d15fe19f0ab22e6641aa4ccaead03c7496d1141a9bff86ebb7e9beb5a68aee570b3f8dd83bd6c3ac3c946eb09351bc3be9d2563a7a44f6103dcd8e8579a1640adca4acbb9d5910a8cb0af3def126ce46e5af662e36b877fc86690a4018e1ae7f0a89712c865305a88d28247d58c2647c2033e6ef88f6ae5794edf9b8a54edff66d7b874fa7b0d6114d2647cb094483dac062dac104e4262229b311b155663dd5d13f4d85fda2b7abdd1c2901d7295859f638311f9087c13f772fdc90e4bdb55aec3266e1901e63d8420b6e8412550629acf03cdc87aab943f6b44bfb478f7e58e7f464a08ecf6a9c6dd6782f1d017f49dbd4657d9a04e29652d5074c84faaf2f1e6a0d24c20cb810df6a1fb1a64cc82b3dc4b80325f1fe16ff8af8c7a377ba045b2aeca530639a3bf7bd5ebb2c1d0c998d0b4153690c1bc98da7aa160e4c94f431482a97eec39f7524a8a16c060f17918ed9b2fe0f541e9818bc4b46757093930fb77c39408dac191937b9d3e8fd8466e903914ce6c1ba94c0bf33ccce134685a4ce1bd1a95e934134f8412ee6c6fecbb50ea20a770dc5ab80fa96f577b222b0a9e3e63f90e09810a7e43ffd42266dfcdcc4e16dc0a95827cc16d7a84d346a1c4c14c619ac6eb4ae121e4416ba6e0b55f9380a297f09a6b8c7e0e7142146a5ba80e6bd4c3468c4169b1b17ca91a8b1851a9b36486642097a3d5c196a28026ce26e48ea107ac92fdaa482c68e8d446c1f5d8a217cefb1f2b0979e0cf1859c3cf68e0d5a2f0a28a24a9f8b24639be5341bfb7a389898062710b714ca13c188fe4304b9b79be4f6910d8dfa1fec340d3ce427e3a288d59b8ab0e9b49e5c2a2a24f6d553d6954525528ca44be4e21ca917f0fbb5211bc556234af75b1df12a95f8941de5913b7e1a18f5193401d0c9236801f8a5ba85a147fde1686bc3442177f0dcbdeba04b6e417fca9217f69fe50b56323f134381ae1ae71d232bb82cd5715;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h2550896ba6417d793700db74827895c3d70c453b76e81673439d9db4bd62a2fa7f934d9295024f908bbba62711333c2feebf60ec05864d2e96bbd0748f0bae9b37e925148888feafa7b00ff6214a9fe84789c3e246a7235eb204513caee2af1a5d0dcd150b073743562971305abc805ffddb6e675c1a74f454814b3bfe4461132ea90e8f89f43dcb8ec93ef85da31898981572b8c51c8011d59c1a30fc970ac47b277f4cf9fb74559eaacc1dd0b9ffc41e7c14030cfbc6705e648b79bdf69450cb9f7ef62489ec6f84561300f4b0a931d421d2508fe004f63ca8c27ed25533afdc4423627b2fb7bc4df68ffb07f97dc9945e56bae0682098262c540153585e23dad987e8f9605379be8e1a43646b04ac59325420cc35da4747444c9e7df1f471ac0a177379f03a2c71be30bd08fa845909daaf2029001ed0d6c4c65fc395636bc4e5e1fce0bd687b6e418d5e1ebcc2fc3a3eebe0dd12b6d2aecf12155aebef852691668143c038812ee36ba49f9ee8cfb9fa2f97b560e4fe11b59123d991c855c2fa1f1a38068a9fa3cc893d13cdd1cd2ae07cfa1123a11ddb9d3017a4f16f02337c6722b406068550ff78f2bcfb23c4c0478c64ad781b2ed0b8c3d7a11ed1d0897ea88026d89b4975ce11c37adf681f956f86e1e17c34294e97117fab71e204134638fafadb2868d522ac73a9f4d7dc82683e6cad27a9fc75c4b06c68fab32be6104291f9f780fedbd6de4cb43276fce829d0aa97b55ca9eeef77c38b31043651df9388f2886d86ac59250c8793e70ae57ffcdf23740bae470319813cf096ebc7dbe20eb1ef353a34a5f47191fe3e4bf47e4013f163945983576735e17002c694a32687e14497e311ac11359eb302264e437e5d4141d8c9a871404ec11b18f39a706374426e9a8c79a36d01375d8429481e7090844528e38e81163258af32970f7bd1c47a7acfd2bc19446c537b77deb7da3a4bdcf9d492e7dd3f77ff894aeb51d196e6e72c4ba7ea05075e08e343c78c5a9402a5383f259bc07e104901dc14cde666abc2a6d0237b8f8bb640b31703d73ea415c5aa42fc71f98f0203b3f83f9c7ef2d32c646aa30177a579c7c2e73a856da5c6f01f00f761be9aa005a30d17dd51a8356808e3cf9a5796d9501110ff0ecd4381be84df3c96b97366333234c0e4caec93175e3a169d247c3646b9aace6478318de179d9dcab39a9cc59a0dd80610b11a4c03354c9f56788331a4098775bc754a14151fecf611b829ce674056e33ef30fd3ba5b999a01989c72037c005f73a144261ac7304713d5a13af7ee8ef61119718d3c87c814ee887a9de8f29a41683a522cbe8325847ee24057495279049d09a43fd76141021f0e7e131ddf4ac8ef570830bd98ec54a701cef894f337533626879bf621b084b9078878295a6653a7e0bf6ed96d469fb65ee387bf93ca3cfd9143c4f9e451c4f3f0cd0da116fe36af0733118066bb4b898efbb68753a1f900bcaad767b545fabc6fcf703290d275a83c5dfae700a56a4814804813ed6aa5a304dd9975c79969d0d79085010753841f47f17d78e93f79e8d50d441cb00547db3527ad1188a58d24d96a7b3d3a659131f8b841f7b82b75a037708c4bd9cd3058156e6d5e7c6810a7c6e6f3d4a1b88db663af8dfdcc7d51bebe5e427392e6cbdb89f2279c23f41705f622058ca32fcce9562a29b86a27f8c2631f1ec50a741713c53bbcb3e59998b0cf8ddf66904879249fee7a115bafdd455c51dd17ccda5d3a154a619ac9dbf3312b80624572a495dfda213164e6b39af58efc5dfd829bc64e02c6023dc9dd1501a1825356531448d3267556b8ddd59df4e546d40eb426e154d253e5331ed027973b6dafe1cf8628d23ba73fd8f94afecfc2141788a9ee92aa575b5807a3211acab976912d8a296283cac5c68f5c132bf4161638040824400157d719edd87a2c1d5e936b703623cbcdd0f1c28ab8274b2e2e65e97ae174526e6ad9e7dec0a4748a05452d759ad680ca67de84b2d1ebe5e8b363106e7d2f45bd68ddbb1969f0de821f4e6e14f2772f76afc8eaff4ce59e68b77bb310824333b4e60d00f72abe497e97dfc454b46adfe927f497bf5bf0d9ba73902fe21389177e1b98937a2dbe7b4659daf17f193b04c44625141af73ceff2d6f96f72c014422c6e5f94665e60176af019fc6c5993cec8b3b3ecc98af005f8526b58108b1ddece2bb9210f45895741bb5e9e57b7dba67a2b578eda87f6a7382714efd000a8a0d3dc7b72528e306d846b9cb491b666fe48788ebd86ea7c13a3ceed3977462612277920590a32f0b117d1520d0d6dd880853c70a0f5b9467607b9a850ecafde3d4e1ede6d58850b97af1313dfde11d5b04e5d694dd310f1d5dcb793a3846e9609ea6523287be668206b74340f35a3d5404119d41988e7cf8e76b38027799f35ca5ac1e2eaad6fc11b30a34d78d8d069fd1b997b5c494b79cbfa4d057eb759ec3c9926482a4d7758c9929c1307779efaa931d3d588d035940238b6c631764440342413a2cefdaf6349eec6abbe877a618f1ad5c160018800e0cfb031afd0c0ea7075684179a2dee1ae6961eeb1691cb345c32b206545fd793fa7d7a01fa2414b54afb87fbaf910fa5b9e6a392ca43ee697a168affb386c7f7a32aec609ae290649c55ac4f7fd502a62e9009ccba00474bef3ecfdd85f918d05e801bbb758ed1479bdf82a2bd391b43adb41bc29de1e711155b645f62cd2e1862d5ff2d051c15b6c677073f3870e7313a7b81ab46e4ff71376af135a2a0e35f7d208c2fe16c1388c41093b8f7c09b7ad260a288d2b1bc37d46608938e29dc2d559e7d049fc8311ee6c0ac2572911d25c48e0c8965faa676e6f232f46dde854e9173fbeb8021aba130829a118e1aaccd20197e4bfae958e3079c6adfe72f55e64fdc24b33e0a1874428472b22c9a631b96fb1ce84e6af0ac60c9895d837a97f08f09de6929774e9b4c048a6b21644fe0f0d002697afae9f6d104a0eebc4001e7477827f4ab0a397998d0620a6e127f551ea0821501a6e2aed4390f9bff4c0a45162678467253a9636c4719e326c13ad7a8b8ee37b83afb29fcfd25ad88b5673d5a813435d7ccf176e8172e515112b97216589ff8fe0c0a3d7fbdf14412a6f11e4be3a67b3c9708392c18af63bb072a2c2cce6d053cc510e480a550efe8a14a895f3136b63a74bfe775e86d33d47038491eb2dfaba3b90fbbf364ed0115c2befd0256f169e1d7b74b49f37f19ea66a33fa7e8c043a29ce4b74845a90fed5cde6682a0fc992ffb70c08b942fc96012acd2824c6312ec514d3b2f5348de8536d3ca943fc7cb38885586a7effc9af3d75261bb7e1339fa53ba72066ce1d1091c6fb5e03e651fdb5b3a71ce44ef2879678c19878d01ba3686e19094f37ee70425ea4356e8da218e64a53ff4f74a17a2fbd4e904a7cb1ee7adc2fdd41eee5e7235550c17b9e9977e7ec23a91b9f0bf191251e668fa0ee5baa1a691ad12064a65f5492d2fba925e1a989fe8a39ef22e0dacd9f0e7c8d7eacc526db6b84a0e1c4cfe005ad3c38ebfaf1ecb37853554dd668171669c4f9d09c28c327f1ab2476af22f28810a760f008d728201886ef45541881d006a8b18144bac34a0c6870d0189e650bedc6ae2888a86bab90d66bbb1b2a87afc9cbb331e6131c7e5d29ff5ef17d1743bf6485f833c7dff86d8616a7a1031ddf50a1efe43735b34846bbda43585310546e6306f722d47c2af9cb645840cd3afc2fbfee36daa9da96320d564115fe3cf9cafa0701c8c42607a83a2a59a9fc5b6ded058d2d4b5f97b8995929072e653663714368f0b089956a8bb09d2ad3c82edd3d31777b304b7dcbcacda3d251fb723103c387a293190b652ec3b402270601f836eac86e95d9514fee456030b6c5ea2c12337dab31a56f6c1ceb63022e908dbfb7b005ec94b1330c631529a96535195b42786b3e563ec2a62868615e6dff5b638b3eaef791d02667c46afca1f71eca89d5c517cf615de9ca946787bbd09beef09bdebc912b8ae397f99e3278c72f63460372ac8dc65d68e1c59ed1f6a809d6df9f0b7a805746d340d9d876c3f2d7c8d22e1e15d099eb51ebda5d4853e2ba60cf2a58e8c73ac3caa7547e45612596d6db2ed9291f9059819b7a92e2b1cfbef90a3147c25323fb92c2322d1aab904518c8f7ac4e58061006feb73e30111ca317047416936c62ffefa7e5d0bca6aa17af002a59fdfb95f0089a858a516a5dc070fb8141bd9dc02466a7d4ca1bff542b4be857611ac993795d562f89e97e3d38aa2b32a93eb48887ef8c3b9170cb0f0ba75ef2ffb504e3a1337b13f12dc82b43f056c410cb2c362ce8da75d56c69aec0838c1aa005ec30d72f1bc4891a6ebf4dd99f0baf4dd081eeb940744f0b3b528e5f1b6369cd5947b01ec14fac422a2d24f5b24d1186d12ed1e6c78b67c9e0250cbf6576a596308eaeaaf4dae4731036548af88601da54ed0ebf1e560b0bfa710241d89655fb4e62e3adef1f7b0daa6c5dce97ea11acb03ea898ad65f4d8f0951477bcad6d1abf5d43814ea0612e3828a0e8f5e5c3fa4720764ded8ebeb555c2e4346dab4fbaabf4feca51f9e0a93b4c2eaba55f5d8846269f5fdb0376e863298e60d7675d8a162c4cc9dc1c8f7b12c70436011a2e7f3c7e420a40f799b49dd018b5988574ff4c039847ec3a5cdc15aa2af13200cb31a84f6e41d9605f6cfbfe77ef6b2a2a058a012666bafc06b2394ce913c532bcaa71a95f31b5428339370958c1b4471ea76b0cc05c23a5416b31d88f11084e0c239495501c58fc16c3439e7ac64640cf873cb4a81d930b8e0f5e860d7942c5a1602938899fe67a480e2e07b560dbe85ebd7ce74a0bcb75e94a0e4946e2c1d84bc18f067fa4b145a7db045321b73ea958d3acfe8d871c6fa4f8631dc13d085abdd56734caf49b100914e96ea595b423943a29241967f2c4e20447cdb3164934a6b1f7d40b992dd2b9755ed9000345e964afacbd188e5906e7660e4a05b92cd3bdafbe64272c9c30ca97dde7520ba1ba167a09c1af41007f885848372eabf7b8e2b5014a0806208896f7c7b1ee3ab64e570536690e8e93f4dab98f7ee2d83866e48a1bde19ad9beacce24b99dbc32f01fdeb1af9f682d5d337e7d53cc1f539cf9a0615f6b2bc44c1ae82bfaa5ff261cf45001cea6b806629b18de7b267872969def3da88d4100cb3dd1fdb893b7b742fd4373400f69caabf89631cdb00b9cec07751e8b954d76d6b50b88591e027637e9f102f2ccbb0f08682c509623b79a47f35260c132d35589f3228552b95970be8df736e9fbec37386e940deba64d7ac6b803130ea100804fa4d46eff0f30d6dc81430823d13a76ce030b3f36f0bb0f6186e9964f0000545ac8b03440d23699a713603121c03008abdc0803b13cbe7ef596dd73005ec120d12703a6697cf5c9c724a22d823175900722819a1e5fee527a38e27a2370501a2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hca0e0b52159e46cb576e4de48f0e5e1bccdac58a5a731dddcbbb213c7b8c7a7c4da75ab7d1a39d9736dd21a5ee545319166a8b1353b392487f3abfdccfdfd9eb7f6fb63880841ac287f618abe590db6d8d404420b0923b3f6bd3f013232502f3d9de4d00d5632ae7edae6f1d55ac03f6cadd19db0753424b47378c1b28868833863b508f299584338c7d79ab58b1f0f633e9b9401bcb2e2eceb58104e89491602be407fd4c92ac433b5ce1a99330668083fd8cee2c6073aa9c9fb3c2f914791a85c8617d08d32efd597b51db6fdaeb41ab443831ac2046dc0bcf5ea35ae0455a89f5983dc3e315919573f5d81d3e3b1b0bc958937f83046715ffbb13f478e0fe43a211034678ac5c981a73e9f5873ee6f0d467866c4fb04ae75fb949493b4f9095694185559cb1122912acc0c726eb312a271247c29fa6a11b396deae4639e2935cacd591e7d3595b019653532d353c1ed57f0c898782ca30100b98693445f6bc2799afa97f6958dc6ce296b27f827a0eb07c002d6cb7aed0c3877639cb0d54eff621bb4479b9d0cf2902af135d9a2a518781cb784aecfdbf1f7ea77b5fbc28b0860e1aa32574c4879e15c01dcaf2b19c71e45e7e831ec1575cee0a86b593b45e0454b1a769441987906d814b80262feb590634a73996e41d2e9a56ffed99aeacb111b8e9af92412c57217ea6c492ed581f5cede7be0798d2b2bc3da4f52f65cd2db1b9cd69a1356a44c67978d86795810702e89b4d37782cf1330282f71194ca8dab06e5f53a32a52266589fcbe31dd25ab6a879888b857a59b8c0a2ee9888b3363e1a022e2f661d08684d8299a23f4febb90bee1e4fd8258382570f2677935c85a0b2766536e9ea1b6350aaa951205589b53480f30b4a50d2dbe3505bb976b72415b4921f96d5ec4961b9e335715dcb613ff2f4c65452eda94b53c3160537e0e1f5616f8fcbccbca1eac80ddcfc4da1bddd8b35a45fcfaaefbe22c73faaa283537eaa7432d6fee2295de74bd2c661b20170b682d5b77d5fd372bd0defacdb79600c886bb7e8ff36196c88feef8641ebfc9d36207aae170cc12a879d9b2fb42bdad1658ddebcecccffbd648104b4f4173a725085d6de5af66aef2df61da2d0f559e84fa440321e1ab329827f5c7c0b7998cf7ba5ed0df4a0e7cdeb92de0739f088b2cdcba2cb26fb01475ec571c686b0814252e86bd548e26f72f7fa7986e8dd97b032a93b6ab13e7fe5efda9186ef326fd1173eed64e417720e7585240a21444ae48d762f2e301498a82bd1d640dd8c0d8b00cbe1681b127dfb766281643c61c4bc82477901597595c665ea830854ae2dc4f99f173fec665ec73282055f7a73e014bdb939b668e7ab28625dcc086fdc937e55927f14d1aee14540947c65e3ff7767c22a1e4c88d129128560419865d639965a1173ec6067a0d2012a39e0fae4a2ea33d1a505c5284c990f17200acb02e15b889747e1bdbcc7cae4bbd65af775c1d450b649e587bf96b66eb6b4845a4e80efb120a428da2917dae44f995d48679aa7740310d7b76c1229cef21b21fa7c3e3b1a868392daab56b058a5a65b99e342de2187b233fa65d39bfdc831ea9998906b70dda8523c295d737aa91b82875525c719622f0150f524f457bbd27b678739095454b575bb5cff01d170e78a597b19d5c5fb59f291a6fcd7a45a6ad6aa19cc18e8c162cec1c4f0e22c6cba1a41a3cd49d06c3e7217ebe30cf2c677994652c35f5e5e0a22f330d7e2c9c6cc92d53e1160390b0a0c3c75ce8892915adeb5e445d109d2b62351067d383f0371cf68d45db87bb17a1bb17dd04ef8c2d85af69a6708c9504f31a6fd766b06ebf507d2083d033973817a9a48ab42e5ff2535e010a432c894256738ded2b9551b756b768f03f670821da38d9236df343d90122ad56e5eef27e32c47110312407b647dce3dec58e7e18f57ed562cffaf0060d63d790def14aa43719c59542468cecb96c9dd835a422c1ab472df89e9ab7400a23925b35b14bb3a493fadb75cefe1a1ce0f4b8eb12a3a77f3e1d7ab446d7469528d2863590a0e99aa434e8d2bbdf5cbe46386ff73d6588280946e80644c6ba106c562f8dbfa257750ada31503c5d2315484e17e992419d1661abafe932107118cf29fdb211935eaf6dab96cdbbbd7dca88dbb8e36045780fa6f9c9b90f6901ef700840034d464f372aacd27cc2f83e5081103706269a05246df648b33aee50c369714469b3158b2ae674913dc20f3b7a78812ef658170118f4b2d674f7ab9a463e20880bfa49baccd26cbfdc520e1e2a495c9f4cfe30f2a5b7c80b37344cc479937114be9de3a8885fa154a39a03ad3160ec0ed9558a96acd692314f0912017e19e4111f670fae4eb6ae05eac6088c77e91b6616bde4f1ed3346026df2f2fa28a16efb358164bc6cb88e870aca06d44ad5d910d19773f37d0f8e360ae8d77634cabeb05e2a3ed74f1f13b85603b6f6ab0922d80aa1b8e0a3805e35ed5e4dd6aabd3f98e46f9d6b6c3409f1e75b65dee793f116b12f1c5eb0c57915bbf09ed9c27c5ed6e124aa4756542fded8c3fcae077bc5b778f4d67a1353f3bfcb2363bc48422ca515a0c235a819c6b957c9cb57d23a01e7337ddf99e9117267fe7faf608f23a7b518e00e86c3120da636f112dffd08df92a8482635b14181a2bfacf9ec6e426451192f4e5cd1fb3f028ecbd918b3ecd8174793ace7b06249d448b46de9b85b3fffb0b9c08efe6d6588b91f01d3e8ef91718c4cf88f8a01e07227ad43c55f83cc48d64bc8ce3175c91dd07e6ec8a579e72bff37ff727c735bcb8b135a6854511130fd9ec99f4d6e162cfa700a0217a6ae8c1c561f34c825cd489b3a1649992f98c3cfb71266cec3295abb4034219dfb33e48de8beb7ba288972788e34534370c856e38dd01bff7fc8541ede97656bf39f2fab85c4792bc904b74e250c4f47dbd9e93a25651ebffc609ffa413b6db8dc7dc4cf38a8189f89c049b44a88aba77d4bd3eb8383221b7a175adf07764dbc12814fd2b529a2247be7d272ebfe1b6ef8242ae3a477f38d677760201ef083f544850b8f8b061b48e132cb9c69a482a3d09e171ee904006a7414ef4dcdd3b66f7dc9f9d51b042f6838699a886a112170b06e8441a5b1b25dbf005dc1b20111ae58279d028b602a4be04dc6581d4db8d65adfbc08bea1efb53ad7b733a2241a68612276edb1781aa89088ac1eb21b6ec130d498d17d01ce485304fe87934b12f2d06dfb3812f44cfa04188bae53d68f55110584f1843415a80a8f6d7466d4578179dcbbf8453ffd8f205f21488c1567ddfb40e8af4176ee78e0a6433cc4a5f98dcdd5cd8c90695f3071484a959306a6a40de952b0f4c0e3c914a516ed7fdf47eb002cb835041a5e9afafba09f5a5f35676233b542380044f5b325e88d38654cd2ff9061f1865b3219356cd58628fb1cb817de2f17568d847aed73fbb3cabad855fa7b0c2d10ebf91ac73735d5b281de34f866153d154a9fb55767f842432014e4331865286f7509bc06eb328820a2b0d4ca594d100bb9cf9625263441d52faeb01d8fd53bd96dc52564d89cbe7991b2d075c272bbe2d1db8aeb84df9da0de7de766369f918f8b31dd24859ddd3dfcd6c5bdded33b1a15deacb08d2f508e44a0109bce0d3f5dac641c6e6a52d92fbd3f42b69acdf01d3d35cb93d3c76e0779891072b498cd6594eda5909ad3f44960436cebf3577b536d4740e429d4684160b6ed984cf0b9d1d1cca7d8a2e6497a3c3731113bd1c88f42114513f19a11097410b06ba41a8944111024454be9560a0954a50de79ec9613c5005b76eb864cb6b85f85d42622bd9c0308c877f1f8f3267865f9470217f14c1e0164729e5904ae6ad05c0f53081e4743c103d1ad77164962e842947cd65649b04176b4275736e1ee39b45de31d53df4975d4be29c0aea6a49b255071d52be3ea8a99ffe95d5d844ca6239b801877b24bc89d861a39f1819d345372944b01bfc912f428bbba1ccbacb3c6bec7529843fd5db0845327d3eaa395d67d7fb331fe8718678568a613fd5a8cf4a7a6d742b1a48c00a3ceef96ce4023b2a273d5be7f1a26ee04c108a223fbca58e67320c118aba69ee4b3ff5c2af6629dd3131070c7d209a81dd6b4046d53f09419ce83265f3dc87c7625d92bf0f1c7042b7501289c7f6d5564ef5a62857b966a265212c957bfcc069cc223b5cab600e19307976cd7b2810c6b943d48ac5d9a8b59f15ea16041423f526256e347c55280d95d39a5339e5355883c1232c0e1ac688fc3fad345ef4a8d21c6aa6fe8804b3fdcbddb44ca4746321587da91686f63aabc9f9c23340cbcd970f2ced409f90b7e01bfbedb9e9dedf2f84a0bdb1b0d51cd8e88052e2fe3e2341d43b8be93f5871f013f820bfb2a0f7c0a73d803877929182e3fc614e46e70cc4f6466da547440c025debfea8271047f8dca025445355d894577d84251612f4884e01db2136abe1e14f56c727b2e117439a178f6fb12a492fa531d04b3a16dc5b2a950865917e17dce0e1bc713d436dd7a26834680ee97a4d0da3f0bbbdfe72ffdc44ced836b76210abe87696c3355c9ddf11821cad307da61ce810966afbc4c466eed782764453955be5d5e6cde57f38cd407b8ebfb5f4c88f74754b0ca1617bb7f9dc10f2a4be590b21ce8601b61261f8e0c3b1d5ee24e281029e1f2e3d5a40858f4a084dcbbc36281166b9fd7c5af16dd1c5a6d882173ac6975890f0ff747c7db4e52078a6e6b3a2433d8dd53dd09e7fa441bcebc56da7ec6e7e86d2c1ca58aa1464d09ccb068b2eaeb4fdd5664c7f4ca90b91f5eb7b764fe8fcaa457dfb94a66b25306afb35b7682eae6caa00d06182fbf28c2b8641e6bcc0e46debff835909fc69dcada1a5c8806c2b424c7aeab978afef24cbe8b7a8bfbab76155941dddf5cefa0a7dc7644eacfbf62595144efffa42db6e5b5affd4f096db76e3cd3037ecb91ecc6a915817195a6e61a4be9b030ae6f4baf43b27dc66c400214232b0c144e7581d0ecd997dd855ae209de4f9a90107a34cdf2ed265e800a0eb3cb2b984eb356aaf25ccf5e5d8a75614adc17ff8936accc44f4f02bc88f49418a948c2fea16aa80631da1ee23615ec159411829310d1f25b8c6745e1f042ed400db49e2799c3b2b4aea4d68ffdeef3ff20f007eecab1bcc051cb857281a1ff2f419e8e89c3f6443d0fc6afa4e68cfbeba7d1b2c8bbc6fd3e10a563b3fb4f63a4a563978d87e0477a645d75eb518f74e142c20ce05839323cd8770cde841d21c69a505d9c984a10e90d6e3622693c84a96826a571f33b4aa4d385edf49e146299e1138c7d76bddc8367fec50e07e96a641e4c797f971691993981f1a7dedc2b121904b0bd74b586213b407a25359c06e2e3ce2319137f2b1187b4cd787b1bc94c6be4836e648202f499ab2a03be0d94d7984c8bd6f19a9c9c7bfdd731a2ac0356a9f6680a23b41f0a7bc2449b48;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'haef488f777c4147fac58db364a1ce1e0b2ca53fe48689284255b6b16479c7f4babd9435200731ceb949b374912facacbd8a5c0b80edb50a73ac257fccaca6299b94b3e6655c8300846155d12b8b1d0a24be8c7c31775b721788b1ed6647506d2691748a5c3b5b9b43e9df805aaff1d5a570d50045de65316c243e1e39c73032257216b4198f620dd889b81e02c8de279a9e0a1b50e1d6b2be2bba6ef9b8be78894dc4bf447ae69dac553932ffb4f043248ebeecf9e36b840f71ffed582eea8595adbc8b8a5bd6838ac07e22b861809254eea3395c3e89b6fa2e665f59b55140508cb5dbfa24531a469866a3564776e84d3128326b50a4b7f3aaf55270d3a51d716a392d205caa5b7b118f0deba76a0db53074e6414b78514d6f4709ce88c2b64ce2047c6bfd4b6d0e971caa614672ae7916d01e8ab6d6379e2bab42712a429612988c8180e394a182c9a5f3b6f8538daabbb7ab118e060dbe5745d3786a652f44d3d304e0945dbb88720e808f6e89e6ab01d178243cc12ead570c26f607d190caf7a4f29702845206848ae2fde19146a5ebf248f8ce4b8b1c1032255199c6fc894fe8742039d258722dccf9d52f03c93c6f342ac2086fb9e9fdc7cadd3c5b3964a2fd21ab637614d5c1d90ba4ffc3a744f0b3eec7d3b26f2559d59deba188d7f6937ee6ea97808a6dd71a794502d9c63509b056595c29d7e683a87717bab457a8da2d7a3e4dfed41d1045a5d8f42c65bb2cad04c50a6622e363932ccbfd3b03bbec94407d2b60bf187b20368ad101926f893bbe14c224e840045339130b7ffb857441ed3bfb7244db18d225eb683efe3276925f5406300f0aa721dcfc22a72b40d6ec33c35918c2e8f012d4617a80db4041e5d04f3bf83df8d5da6f7df8e61d7015fb8cdaf4dd35f695c9f46173f55231b5b07ead7c41b479441b7cb9b90040ed5408b3296ed661eb91f65d280f7602543f3427762ddf6f2d800cc0863909a11938f99f9cffc0087644a55eb89e2d3cbdb170a0eace7c80d1afc776a49bcdcfff59078fe1cd024e045776a263158a00620f020b3135232dfd8d0b4f21d40d617cef0e0ae09e18179f612cb3f1349f12dac2975456bf9250e7113d4495062720edb5d651f4e74ce1a1b0c5a89634d63ba0753a89d5198191fe198f737d00bb342958b374a0713e3e77ef90a379142fa4aa74299c421dc16afc67fe717f6dbab2dfc296a1dd94f84e6c59e6dd983a9956fbbfc591468b7327e0474a1cd719f74108a3dc0b8a5434bf3f6de35fe7ad4bcd4580842718211e11df9b7fd9945cce8cdc03664dcf20e47238fc792cd3bfd3cf6d9349e42436de5fbf3d99db15dbe344ec28242e1bd4b7d471501f8e916da3b1f2db516efbc98d93f73374518a1d142447c13844f3221ea82df74389e592bafdcbaf5d59168f7f2bc1a66bcdc14c648f223d6c52736c696ee334afd64b874961bce6abd11c496262cfc6e0328f87dd77f4534fa4581320e5285aef49efaa44ad0c75551bd5360855725ac73465118846743586ddb5e070a69e20b6b5ea4f9057c7154183658f359f0b457503aed6874f16217d1486be89a26908fb0bbbfeed8d8c5cf6856854c9672df4cc04feb82fe4e96e428ae6126452dc9c6c7b2bbcc6d8b7f84e5cf25338f8bb1acf1c0aeda573ea9b94b029c13e8f14869ff156e02c2259b33b4b9e1e20c07b4eceb427f7172b4dd66061df577176374cff9f0d4130253fc5865ca8293dad59f45716924129162c605e45eadac81f85fc017f27cf626fcaaa3d94022bdfadad819f2984b7f1715cca1b01f22d00317d8bc1b105492b192fab8e0b1fbbd8387d9e47e62e31857f289b06f31b5228d26188529b0d70e90e76db5d8ba6b58f088c1e1f54d190d32045a810bbeccd0536bbc3145946c45d8cab2811b727726ec9bca5102e09db0cd1bc84a275b3a3c7d235af3d5c31e6ce6fa292a8492dce4c699c6a1efc684aab331f01d08363a0e21577390be58e5f1fcecfae0add425ce28389457589cb1db4758d9ffacb0bad9481ff2c3ff35de338912e1a5fd4fcb989f68d02adb282bf40a22b3f73316d0738b118483776f24e8e44152c0ebb5f962bddf0a85c22953794ad41cffbd1fed4a19ef1152dc2173099dba61f04c62490e5ad02b204386bf08ac1dcaba60b91b81d0fad518ae64cb7e9efb2ba3f07a75c46dea2fb272e05a5de747d6d09b0f8a1c94c514efbdd2904c781eeb8dd2ef86e73a92c0f2891b02904ce94ae262c3adbef72201ba76c6d9339f2f65e6b38f3bbbf97ec685fc2b9e6f2998b40bfdbf83188731e67ff358eaf200278a6a86d8e9a2bf47d5a1bcf69b96a87750a4e797de4383cf81a95af808d47041115ba1764d3add337fef9184a45f7ff4294ce0666852ee5b338e7dbdc5b71e2bba1a58e6655812cccc170fa3637c3baed38933c97830f757826f7ff1750733aeb968a089a59987b9ca708c01fafe81034ebd67ebb7ce8d3f74f29f2bf6588efe757c89c90ad820889ac72dad3e2b7969a67b516a8648250e07ae4465f5b71cbabf316a05978e1462f74f408862bada505a3f016dc121964239723d7bf6b1f3eda24ac930b4519db6678863a67cab81520ffeabac9b3bb6e1ebd5d5df4858e3924a994e48c946da3d6914107987a8c2907b3c690efba4c9f50308414a5aa8426f751135187858c52794173c06d5fd2bfe7b1fd083deee9fba9e54f1e12df316b8af2caf52502e27fcf669839f2e269fa37222bf35d8282c35f3a7b2b70a4630cf8676d11a99d9baadd413d079aefa444ef0ed6414b0b2160c53bff42a1ec43228879751c65778945c6d536c4ecf4ea0b38a19371bec312e78e8892dcb592a86cbd4efda8fd52efc0070df7302f531130540820414ec989cca73beccb943b2fd51c4511caf83966f4ed4d98b23af17dcefbe0f555c2f9f77035c25a09f66f9d6459adc14d80ae0ec68f8e6e1facd66a051a31cf912814bc9d93fd2909ec3dc6059cc305bdd617caa9896ed73dec2dc9063a5596caa614dfc2c3c63a5144edaa8ad6c9f57040510795c3673878cd9ea2fc7122e5d421624701fb1cc740124aff82214d3903c44db5a682a4ac07ed08dd21ea88d83713466efb4d4934429eb27d2bd12b1207c117b5ef3b9eb64c564d668121e2e99927a9dadd35647e4ff2864aede710520c15240e0b92594c93431adde0ab03bb0a3d1f3ab83517462e833d4c46ff75775e2faa63cb3f657ce1eec21e02f93215670a74786eae6c51b1e0e6b3329ce46378b1cf06d1794085cb215a9fb6eb7915037d9046577f390f93fea6cd251dbeae0d29d509e90619718ee5b487cd8b0ce576d0c9e4c41375b0beb37d0573a258837fd15aee0141a65c395a02ad130ce6924256aa2f73d43d747688a12f125f16ec588a517c41909fc8a7d240d6842e2418b0afc57826969aaf435a36b336f4b3c0787f2b92adf57d3cb7cdc662a7b2bfee90fc13e296ea381718e99e37e1de9a3fbe51b980108c69a700b6b79d01acd40f12b6fc92212fda44dcea11bd7a267c0197df55d8d05c7f31e5d3873f3d4cde7a20840f076306ed79443d1732fbd11d216d4ca8efd11f9f1e7787a3d39a6ab31c0aeaf75d4c1f8e7ab0eab3cbece5d99149a7ec84bdc055ea84f635bbc3a22d77e4c7b5283130467ba59029610ad505a5d7fc2468cc9259c49e5fa86db2d6ca7e0ff8ee1012678f83e7eacd6c76fdd13900cb71af56b0290321b8359cc30fc8db5037ff1eb07f49a74be56921c0cdcfd323e2ddc2f90d962d9b6ec399717a061f1e20c188f583b314ec7a9d716ef4625eeabd2ee5c09977a425d0c75f8c0651489e43911712f3510ef5dcb0c9c5bee55a45374ed9b792cc31f05c4d99bb3e756ef82762f11260738cf143ea58961b6fd3e15f4dff89f58e3a6a8e7ff09a840693528b244c78845b5c1e25f01be6532c37c6f816d5eb4a249318400282043763b12095b6b22027ac195a57878547f2af754c597dea2974d954dc83cd6fa34a52cfc49fa2d1bf2d57fd2d0a1d9fcfbb8c5066dbb6547f95c0d044837514cd77d52c32dc47af2b40548a5bc68edd181169a9a1f38bd91582828bcf76778ce6c7ff7e112112c2e2220beab89788d209ef55ca206760f891b5c43b7eecf9a7f72321ee8a3cc6bd6d711944c9beeff6c8c451639af28e6e59201b443e0d6173e9326d17175ae06815110f9c921ab9817452325ab363b702399a7fc90352a18b330b093db030c024e2f26393b8a558089d3dd6c45d82ea9b0ee8dddb271b0984ee2d019baf2b70f39564c21e909088512941bdf022a82025308a7e4db5e83f1158f65fcb2a7db859795d5351849129041ee5bb2e86ff56afc86d188a86612e77e949b87dcc8c37d4e67d900a4e18cd2279f1a4a1c4ef8e623ccb47ba53244bfe1402cc2150cc01b511212cdd4e15c967d6fecf5b22713b537cc4e8ac7b7cf007f8c7e7d61cd84fe3a437ae55746f437a11368351cf02f9886ed34fd3c04e1e0e98a2bdcd0f8e8a8c66ae7819b81da8c9bb227c304f1a468c4cc95a79dd462c704a0ec63a6b5e29f940f016fe2d49092920d89defb8f3c29182b9e6321b3a36b0897d3c0d933abd5fa6a032c774ad8e08fe1b2bfc6a426b433a85bd070e560be6bb2496f2614021b1cb4ddd9907a69f4551ea2d70d02388d2ba5b5c7b7a4dabe0ca011254eba09f3265195218455fb20899891ee69437016b00c55add7607cfe4b53b2c0c37764e864bba2922f0484f22bada20aaa4d2251088dcb6d73bb9fe2232b97de01a2343bd58daf8acc044f0a544aed700f383c563ee973f1904f94b8e39cb33c79d890d5de1a733645573f88900c6fb0528b691f738480aa50ae35754bd7407e76e90d1a694dc9df29cf87e4471a6b15c1f41edf13250a698ef9a12d3dd6a38085defb0fe4a6963e16375ca9f5f10f836c7939e709e208a706470219b2aa44258f178249659170ec933dd0182044934dfd3a6e033c8b1e8ef35ea940a9efbe018b33ba57f55b6a985b3c9816a1358cbc737ce6e030237ad97cecf9283f6296cab5a552b9ea93ad08c5730554cf40f1f33a4c51957cc037c0ff744f918aee57c1c0b23f84e7c6282128a5ff63da134d8aa7da715faf25c6c783524764191fdca7ee050a3a7dcc877451142c7211950e01e3b0fc89b63def56d47bb16762f6ffb55ed9252b3666a83927d1eb26c133c02032ce2138a52bb982ab77d4bd7fe8fca7b2e430c5c3aba829b97d67c286f37b2d68d1ed447ecc008c0ef75a2d689143e40e8aa0cec20700eb3698a9732ff6a44bc66a81574a45888942c0cd72ed20f03a494bd72a1808527df1b946af207d9d8d5685149081da909ea1d48297c376a59af9882d33ba27f521f97ec1f7a59d15ad4df600ab4ebb5c0d345156805c01e170da636bd07585f14bd255abefd21c24c0a94fba1819024a388a19661c923206cf0e962dcc0baaa238e7db986b9576;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4c7c5a4e2fb76c937ebfa03c5099d8566ce6b6a9b59fe2f8831edba4a7baba9739b676cb6f265a234c96d9e767cf383b2c9ee8789e120528bb27df4413c2f847ef5bd9b64869cb1717535884a6677e1cd5b32813b24131e86dae0d2f747ada9bb0c1d58e0649944afbb2428cf76c5f13ecb4ab588d2c0233417e5b7f8c83b09a77512030a7686be9ae121ab90b6b72eaa5b3758e1dbb268b3088fe9e98c7b1ba60fd8fa6b008dbc9a17ab64cfa2336c0d8e963ee24d8e241dd926b292af59b955b1cc048838649de28f8a5adc5f1a97cc55e9e2954a782f05e6a8b143a31f83d375b50e88d375756f5f5e12b7c6298f7b66e55d4e7f9c399dfb5f5852aa7345674ad3a7dfaf899c6bca75f0389f9035819f7f5adff2396e2b1033601778d61f6c5d4bbe3633e2fd34e9b4794c5b1a4a03273d7e56858d97cdccaafb913a3eace1d45014f30150b3189f39e48ae3d6e0964bacdd592d6d51d6b6c6ce039a63ceda3776906e099bbb3636ed0c6ca4f29b8a16dd88b68c08579e4527f60e1943468149ccad939b9b283b11e029c77683c7722bf92cc16ca215933f561561d3a865bba11a46fa6f323dee6362ac9826dff80be5870431ebf22a332c69a8979e42f25db6d9309f49ea4d4f0600906f230c74727ebb176ccc32262b550bb931ff4e883c60ea27ad3f1cf5ee77ad581fec61856463d311ed680f47bdfc8cc83f0864cd6cb0eff21d3bba85b1afb2d4cb13502a303aad81e5d2e38bc25c005f0610979e028d2a00c0c16cb2e173a8acf3899076b55d4d6314411a13cec8f81486f4e9ec4ad07aef9cc389f7b3c4b3444c265976b2b41f78bad41563fd82147b5bf98bc97905ec6f27feec8876758406ab1234e98557cbdd46d6658afd00ebba9eece289173911daa459588447747acdabd6ca63926946ebf50a0d216980c0ac6baaff5944080c4bf34e93e8edc92cc9c2c0787eb6f0adc8e55a4eb9f8c854deba3af9c808d924ecb901014ef4feaaf466bb70489bc83e85d51a94b1c63826976088b67fb34010be7a59ea94b39648f6ca9af507446cf32712e7564a79a9ed4fd237ad23702c8b6666be79bfc889ade1ef7fa0a23a83d9c281317f9054eccf5132c6990097a6677e4bb9ca32a400e504c365840f8872555ee8e20abe2042713a6b434764d26f599c7e665c0bad20d9a3b579fb4747daac6d743a5f15dce86ca8e44bccf6f43af36ac5e01ea01ec4a711258cc08b46f32e315a33f0783958da190cdadcd1101686d9f599079307a5fd06e4d85b6f8c2f8a54aa3532629d52a6ea0ab1b348e5139ec1cc466300e7250ed6039464788bf9ae2954f48bc2672b93a15711adfa2ee2864003aa4c9e2da447eb02923bf0a97fdbe145565db5f549507317f198973bc32092daceaaa8f121976075ad73665e4aa989e6ea89bf099d6208e19c1b8d924156e0b8b6e1a5aeb88e1a8a698f2ee466599cc0f46020609f443d3a2ac1c611ed1c50676c081b278e8f46eb1cedfa36ec6c9e54f89dc33dddc8c8f20ba8bc2185d30568901c50add264038c0d18326a1ce9d983e3b5e4831b28466de4f456bd7a319049b4f416a0beaa0df210fc032eba9571c04df162630e56155218a35cba4b1b42059776cbb593e6c134d7932e7d2838b8f1476945f86ed9fddba99a301a90ee0640b6f0d0384aafbfc057b9c03480405919314559569de78b4e38bd41c46cb303715bb0b2b702de50c8ce8727e885c64859ad534f424e754cd3a2d8135f447bff37465a71538d136df864da14199da9a935d17056060c34eef382442c3296f9efb12c29cde179cb4ec15a1245f130e6ca8bf08b78144fff7c9331e010767049af852ecb059fe3177798bc5d1782e0e945ad7cc7824308836c3f6ae1a72d0ac9aea5cacd137bcc5196c94197d4b695736c8ed714ad27d9b919a78e5ba9e8e5e04aa683a9b6ac2f967217492db9ced06593e15a8c0ddfcafed478aa1af39fbf5aef21fcb2ec3420f91eca786f7ff0649af00fa8634347aee8a971c2d6944b58bc0009394be1250f2bd99d8162f61cedd21e2a664be82951b4fac27587e20e9d688a1572a90c2e3af9e2b2e9d4456b79f204c1982e768d4b570037ff4b7bc5468d4367aec7781299a487d74fb981f59690a08d8bcf470c2d4e5b08327bd7946c6fd0dae5e9ba5f92c7688a01e8d690129f0d129f5067500ae1a35a421f970182654041578cfe90a84a7b53972ad56a8a89e325d74b2636b9e9faf029ed6a205f1c711111deb8428dad41a452cae49644194da4f90dd2c30a379d1962f8f6c710f288de54acb5a5cee4e8f31ec3c402d1a4b459d536d94bf6dafd81d830ba82226fcc3806dba98a31564eea33418c3c7e6c0e69f7e8bac4fe999bb093beaa04c8931742fd0a9bcd5ddf8e430ba17c51f4492d77296ef1f3c36f964b58c7607b8a26f6c026e3da093250b133873505a8bbbdc0113c0ae7ad2da93aa492f719fe92dba5a5035b9896b37e6895b02452dfce6fadb7d40f1230fe4d420c4b6c9f747d33c343c03f55416d1f2d86115d9616757e2daa292daa139b2540eb1d4535169a0eeeb02c6cdf9a3369803397a9007326d707b744827dcd80478d93d84e7002596eb06e1cd407f7f7e4421083c9e440cbb186cdaf7918be2dc176a55123eb495eeb1116232bf2fdc549eb2a375990b0fbac425224c8304e7a8fe2423eb68eccdeca3b6fdf274a4494fcc19299259a2a42838701888966401a474020557f5db29f9ee52964a5af11ce3322fdfd500be6a6e14da5a08e2179dfd97cf208cb045c2abf5a17722e7d712cf353e88cee1877990825b57e92992f19ba821b6418cc0f32b62908200d96e16498b1b2020c15a0ebd4941dbbb1028ca98068339753c2fc414841ac2ce90c00ded17eab45eb15466e8194e42b3e5b9385af277be4e914d7d5d1306373d6cb05bc18e3d9da54ff30fb9745bf974c63ad449b88b4e07576265267503962950f07576fa4c426c6ac739ceebba37f6e35a946effb97c54fc234795deb55710ba34ffbfb72fe11117aec9981f9697f0a5a2600e0effd34d882acb52966ea26482fb57e0da029d46d934820cea4d352252d6757af3ee0dd571cfdef86eb61a50023c67abece5dd39f8638d89584b4efbe96a01391bcea6d018461f7977c4643b8af660a34d1ddbe38f0ab0ff19d099ad9b7646b357b1fc8d8fb5a22ba3d4af36b9eb8ae41fd7806af4ef04d7e98653474668728fe2ca08a5c3d80e40a308a52a2f4a2aaf3734197e3309f33bc0c53ff9e03706efba6a6ce3c1c3506b00d9a8b6b69a93f3d9084e809b7c2bd91f32f5bc6bc2b9f7fad1792f71b8c0c9a7fc63ac2252406ffc99f63cf99945314a83e77799c12732a2436bf87f6644d32e1b970124d7b11034e99ef1a088b6ad536aa96d9b6394c9bbe412a48c82b1d7a4fc1de9b832c0ec96fb8ec5ba2733f9c9a845df4d12ea3b02b6f9c6318a59c0a24d98ba1b91df70f7fcaf73942c2e75441aff6679f7b7754538e6db28a7ae46271706006a4f539ac2c15a97a99475e43b629276c36609dfadff58a9ec4683064361807dbb604f8d8d9714511cf05552cd997b20b1444e7be8b295e6a9bc587a71d21bd811c86770837fb8ac902dc1bdfc4fb4ba105ed7443ccacf94882afcfe3f66bfa88e0c9c753f682b75ec767a8383de8c90e5e72bf1080f420c16c84afe87e137868635d3f7aed287f5babe67670cf6e3aa5f9658e4b687c1ce31601a81358d65c39ae5309fdb4743bf841ecb5dbabb7585e8eeaef85d1f3832dcb738220432f0331127706f559d6ac2402edca9f0c1520e327fbae21711f9d4bc79fdb0653725703f40911a91d2e2293255cf7a1608524c8c9c47e4bbbfd6d53078a6d3a909f88f94f3ae3d558e3d9d639a6951365dcaa763094a1e7f121fd463e234ffa7b53538250b06920728b046401ffd9991b8e25ebc18b37fc08e9750d16038374c52e6a994c122e64a5d44ee66b1fd1c93d3fa7276606097846920e903286da2150961ff948eb71c46ae0c0e022480825ef2d82b90bf5b676e540174f7dc2bce42ec4215e53409e557cf997249098e1cdd3027bf52fc21477b91d87dc549a52139bffec5f20581e1110d21d0f0ed3b0c33cb448491694bc69d72ad03cb7ea1e928a6fb76277ccd47092c458682b6f967da1509520e12a95c59869b1b2ed66694100c83989b363e9e8ca2bbfa176c0f4d13e99357c0d4947f5eae831cff3fd0b190718cffe1e26362ccce09b5541bd69ba18c3188b09f87353242fd12626e932e8924f3557573d001b3dc387fd57b9e92ca7c27ac94ac336018f769a94779333195f15d9df9dbe78d24da3f87dcc6a402f1145dbf4672371bc512ae2e24036d51a708e4fc0e6bd8bc6b9674bbafca726b088faa2fae291be3b329006b68db48567b61c874a889412e2d21bbba41396c6ce36e1538d838beac787c4340ee7bdb9b913ff07d60006330a909050389c112e30d1c5bfd9ded76ef69a705f18da73d47d4139263d3633e63a2b1942264bd0b706dac6478e731fb62af025cf2a2845ec73c6e6b489f2b3b4e81f817b251f82d502ea7321a84b5fe99d0a32444bdb6c86cc82f70a114ad250feafad8c4c222e66b1437a4c72bf28dcb6d616a8a6d8efe8926a6f7c12b1a6f988dfba9a4b76ec04b884ec1519c6f36187eb297b2e2069ff4e0e4857b78a80ea766a410b799ffdfb0d527251be80374813a3bef8719271ddbf7a34b04ca34890fea7eb28aaf250d73edd6c05d8d4a1f1d6479e3a8633b2b45f9e6c045d27b7062fbfd8e7926bf833ecda1f068d0cc70daa0a8389b2a2350b09cc22bd8c59120408712234a5077746a9534b57ea3b0adc70145c0f9f63db7b71cff4dc15e5ea77107e2f1d6a4d116bdba64fb5e05aa76fc711a80ae1f57c5eac7077289fc0fd695e1994c36515ad3ad65d6a1ce11358c59e242eed1f9b6d5321d3bc85cac0f2578978a99de84c143c5a0078d637450d1126e7f3ee19dcb46dff631d3b32b7d71c199a31bb6e008fd1af073fad9bd6bb95bab9418839ccabec2285ad6423a238a30bd263b237fadfc38b8b79f54249ccaa93bc90d8a110d660290af80354a4ae4acf290f54b61c8235e2559089d0398d3f25e8ccfa799e5e50cdfe67474a91d37f80ddcf6ed2c4a0e66c92d3d9e4b4673fa5c2ae0eb444051100d1f57ab029bd274d515f4630beddb2e167e4a916744a7345513b825a32999601a53fcf2b07cfae8a8e4a275c3d566553236d828b111a0d93fd9888570318e44977a41a35083de2a52c51ac57d1b123172b2b4b7ed57d39902866ff28f767d2b7919ef7e94676d61875608d10585089828a3313192713b95b4faf5c9d6c80e51f702b1928ab45fe22df958b082e828655b114edbd8057b361394e858a77062458cf646c147b1b1b723de5698c522c262762bd550d6e0d98f4c70eab2762fd378b4708e7a0bd29f7d646eab69e747;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hbc9c2f0f9111df1383a464d735e91332dfdcba32dada35f97dd6b67182459459e4467fc2de6ded2459e9e22435ee2871200d5586a27c062bfe07fd08ed8656014a5d22ab602da40aae4c25fcf9f0b6e48fc6a15c2f27c601204ac5f45aef4a1f3b99bdde01845aec4844fc929897ef2cfc9d52079e35ff3d7487cb9af853ca61bbec5e8a9c45b52b00da4a4e82dee7dc68b45825c90a2c7ce856a8d15ffc2baff5c4d3deb799097831a514823bfb48a8a6040e78a07a0a1f4e09b36938ba63c5087df3b54facc53c6c23d6401f93a92d64d85314daa3e8720d11bfdd3da9e923811b0972d1e72367cfc925128bc2e166ccb78daa4fedfcdceb28c12a256fff70a17a8798339521d5fe4fc11df1ea67bfe1cc118479744bffb95427aaa0468837f954ad63cc28b15f789813bc910c1f5487eda133507e0e4ebce40733741ceedf1c5107457208d9e305fc1be201cb966cf6daa7577fed6dd334f2bf92e21c61d7181e5d5f8301daf3e634680d77f31ce7ec610012ce003204f1b14dd4197ebdc3b938d434b8273c1c4b78df6f3104599183e40eea817c14a8b92c98f9927e23410fbb327cfe7e46ebe0d2a00e42519c5c4fc702d731dc0019fd70469b0f83f82d2762ab04579f3a24a757464878732aef41baeaade555290e2caf083664fa4bfc3c06870d270b4154a5348d0e990ca26738adb807b9e216da368aee184e6fd78b4660c8df2ae1f85e259ea76fba6610ace6d9e962999868e3222ea60e4cdf02650de929a9a60576934d7cb92600429669246bbd069b5e29b8a9c969780f64fc4939728588f54c82912e4e78af8d7e834a383f254954dea15aee76bf5fa49bbd3953d4aa2a8dc58e9ab0a4434d32da845f73029d059256c96f5e5d8ac5a7473f138503c83230fb679e83dcd4ab0abde4f2848b1d19aab9e44ace6d7b1bebee9ba993297c4db85fc1f34c67cd6c8141e486006b6f8d594cc77a993aff86c8ba62b34abd8f94f8dd9eb1966203da993fc83500301340e5a11d1f6721141c520cb2917507b10ad4a2e88fa5701b48a6bf4f897fa3f1e04ec9c9dc7bbb3b8880733e4db5c31e9a456c56d4ece649ef085d0cb300a60a97ddabf80d70d3e9ea751b26463c127ec2328dd8141c5957d1262e9f62cdfb746d243d3fddc660f943ef5b753c5bbd1b27d55db083a11edb3d5cb13cfadd5c24f33d21aa424ef474a63b91502ebaaf5ce445a1fdb8c1cb4cbf8d4450f300a9d19e723e1f04a5d22f99221cd54535185580a2ba0162eed83463ba26faa029afb2c610d1c614953ea30dc9ee90baa6aceab6afc8ad9f4f2c4a26831413ee5b2927b0e0bf348f2314d8a6421b43229b4e316002ac848631229f2de8b319ccfc6be1f1f31950798021ef52d46013905d0800a5299058c441c202e0e88652b7d016fdfa87e12d9e3cc8b19d1f4425295f8899439eafc1c2b73adb915b0d5ea93e0a5485f6e772f8ba85bae810f1d9168d89da6ccf2646274884763151e067bd1b79aa9ad891188bc0000f612645d066f0feaaebea1a97db0fd21b9205a44c5964268f48a583d6378ffe59833d6af5c6e3f9c1c8aef09d87f10590f81c421c98a9faa051a34a27b12400a6e9fcb5e210542a7dd4199cbdfa9242d508235d39ef3e3c61fc4417746e52648d6f8c945e24826da6bd151ea3a29bb48328cb0246b4530dd76a46386cf3b2dda7dc548b0636377151ad87dbecfd63f4a852d94c001b68e31702ab8cca5a8557295a9f044c9dec1e667dbeae8d82cf839f0fdd96b95fe6fe9c8c97cceef9ff1260b557db5e3a2e27c83d14fed1eecb9cfd829ada7847c807b5055670f3d50373bdbaaf7e2e1b4e89f32ac6253fde93734c2405cd7866ff5b6e1bea8512b7719db7d1b19803c6b2bbb3e0da6dd6d7cdb9be80f896f60a74125c2784c3541c160c802b4344fb5a51e15e0409b3023a23c0d499a04ea4f13daa447ca9759c1de6081601a2f400056eeecd0bc2b2866b278adac856c9cfcea7ad3dbe31ebb7e3a8ae2c12c6decba4f6eef88171b17739fb6abd30c7b89144b873d348ceb6e5616521b98c80b211a2500d54add6db5e0c332cbc36ee7c44778471d6d6f67b746a9d96bc0113ed77c09836d94dff18815bc12bcef3f3d03de1111f6031189f44693886cbd6404ff90516e5fbc33f9d2a90b27cfcfd1d7ee45c427af2dff3dfc176717291f2e6cf0aa2bd83cf678fdfea0badae785ab87ad58385147432634853e8a3d137dda142288957d53be76c8266979123fa3783a8c40c4dadba15fb6d5fc854f9fd5c752a368e907d62f6aa5677f63e8e9956e7523677c86a34170d2618f9aa7e9a07a9dcde9497dd1fba92f337b853c4e5145ebaf21be56299e57da6d0c7cc6641422d7d7b0fd173d5759db874e3cedda7b5d7b894d5d7d392c621f6085cc7dad142fd1c160bfb9bf139422c9bf25c0a85eb2da4882ee21e1c1cc7c574dc71c4119da5e28f0e5c367597d5705e78a7ca4cf6a8e5228e4bba1a28a9607d2181efc5bb05a0e8efbf1a41cc3ece24359c3d65baad4a91cf41f1500213f71c0f7e51276e56d5abfa57e830ad4c803bd6cfaf30bb2b02e5200fb235566f17a5368834b1bdf091ce325e5cc6bc4251ace394e92a12d81857a0e1ed3b15938375277fdeeb96f40d067195f32ff0c34f03e9815e9c4ea6f10bed6bcf3bf184a74f242973a3763320b7b919e283218cd6e2758b7051a8ed6274d57b4a251ff2818f397230fa05fe96c6b72a610e557d485ed4102b42b2de50737a719abb04b29fb04f4aacc6ce0f1968427f93b0720107fc47e81d16fa4818fc749603421042919867c045a6a0879095fc137b0c565f922217fb1952d4123b74a0e138d2ee3ab9c4a48b29f78f00f11ddbdc4486d776c1755da2a892311e3d3cd4df7806e8dcb230730905ca496145fbd64738ad3aec0968c0f2d45d6809aa377722fc32ad3c70a5d58574d232443b0a31d51185ddb0bc432a5bf76578d56b8fd9b82b28e93a998d145309461bc7e74f07887296e29085017ff4833da0283486caed8686356041f5b5e8d88a5ebb956bd683f3adc11f24c06712ca8c17a5b4b3538f15cd80041b942ff688b2d369573b14ce217501e941e26771658b08b29e881b0d3f0529d0f38d0478ac36f7b8abcb55f93d92541926cf95a55bc46aa59c0521ae71627e40dedc78765c8ba3a0228f3f7760cf57c58c7a96ebfc57773519827e700c68000393dd61ca0d0a02b4c48ee25af9149252afbe8981f2e6fb15e89d8a8b5fbb61c1f804d55346b9eb90c83516b51d766bbc963ccf213a7f611c6f97c060ee938a27575b19ed9776d00f79470c98888375ecaba797fe3a568ff232868a08ce5642f32a7f48895a8f027f2ff223c0408e2fc52eee393bddc3208ee22f81528eab5a86d37f3e97426879913a2da8539526bf5882e16c95bfc1a010e65ad48c2b672ced477dc2670a337329a4693f63ebbb375d9fc00c5f930fd0fad0953a44db99a7fff7b326f3ee1a54755657443c8511c60a06772f59464fd7aae717a25d58a6e14463c558d5774e179cdc34c7a869bc112b83019dd5ea553aa6f894fc8531b3511ae548e2695a044f3980f159f5057107f56d4be819132852515e9e8f94d13a6aaeb357a1b55e81be76710041986772fd924ce34a366f234522ea4f0a7eee229907d5d142347b40593d7ce4e88d4308ab21a2bb1ac013d7d260cd04f608c49f42678bfdb618479582dbe405bf3e38a7a8e41c158f21a32a9416b9f3333d1a547ea4708070dc28d5104f99f0539cb15713e0eec784b5e8d68248ecaad592cc83ea839097a0d95853376379a6b58348c8a3478421e71a6e25658b7a5f2b904752e32bb473174adc2ed17ee2bb5759773049c0d605ec888f1545a1b6730027844dfaf5181a61fc2257ce4b9b9e62790665b96455f8c8de284ce058368a27615ab4163b6c26ca66e50fc55f92e257fb197570e0368f56f1ed9159cdf68a1483374f7a032a22c4cf85e31e1207cc4550faaabfbeff902a2f7fbe188646029ccf1f87a72d67a80ab77cbd2dc42f739cb0c59792d62c9a7b2e3a0b70567172214161432763446b08806cdc57152e97450bf66a8f236423136a454d7eae6fb7843b386b1cdee50f2e5d653b0cbcedeace84897f70dfa833880201b9b799172fc6101d70db8fb6ee7b23185d027bcafdaf74029a006810bd83d70c229ec3f79dd5a5d88441bae87dc165376eabe1dc858015c8980797d97cc7195b1ddc40ec06b5777331a2428c28913a77936cdb98b8071b6863c41360ccb2d189038a21f591599b959b74b014cde41658724cb235fc746b6682486ba1c4ea7fd7fb04219f220ffdeb6333f33293f30eb51773b17399499fcecedad4ab26ec3505eeef4e7891b95a36b18d1521d483c1731d1c5bcd90024a6403484f2d3ae3dd6c933ccf25648e0b255f1c018e198857d4712074d941834425772faac5cb2f5aafda55c6dfc638e9897f14226cd876fd92a3b3a18682db0eace8dabd8a704115841151bc48d6028e611f360c9bf25b48e610f74b20de0be668475c923bb454c12e4424be30715a5f8b74a4c1115d12664b76fa06de159bcdccac04bee92d4a94dca7c98d3f5f019eda312a1a86fa95dcfb6bbbe789e1995cab92b2274c4a9eb540186b01740762eff140e6cd8a162630d254a0e81e4f0a06398810bd1190eadc2722ef24bcd3190d6b1cfb5625d565463fcf007ab813df16f6bc82bc26c86101a62dbedea0f44fb2fcf63c5fd2a6a30a95cfcaf1bc404b28a46b4d2ed8867980aec91f9f05ab97ec9506cbd1feba85a78418d03bf42e867be04fc4e81dee3b95581c73752df312e1aaeb6f4359bbedd30b6648fa58433d8e15ee03a7b66d3bbb4f80503492bc0506627efe1ca99f6b1a1a413605c4d89cf82b185db132cc7664e7224191f52872d0d99d4859c6822ede741c85676ed01130df177f43205944f83a63db4d3ea5f7715003cd1151e44bf6b798085a878d6189c26c7ba9bc400d7afdf1ff6232341f2e6ed3faeecd5e7d873ca2492a193a587508a2cb8b07228b9e1391868190bd57fcfce892a9a5dd64de1af389677e707d20adc98fb079b1ea0b5fd64d0bf886fc46e94d710c70ee0758eb18e421beaee4a44717470e17ad8a4081d2c153009cba16d1ad0b778bb98a286f8831c3d68e9078b437d0c590277c532781ff559855d8e107438906f9a36230bfbf1e05b45d1bb3ad533b4d66ece2917efc7d88780596189d0eba45009ae29c854b0b127efd775a7fb2765e2dbc0cfb1d73f11300a7d344e82e5453041d6ce1083402417829cbcaa6d7818602dd1808124217a815a78f51c395713e801402a7007ef95d6aaf327213de74f5f63deec30edad07460a5ee6da99a70d9bffb29e0cb258bb973404c29e090379d1e850548b9560b08f2bd866f46148449c957c818e789bee912935e869a180c831da80ca621a24e9a6db611;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h6f78545ab052673d64436701f6faf2d774486a759f0e64d8e0c22d831520a4e964e4dc09521e73576320c96ba7686fee69c15b68a60bbbdc6cc1f5cf96ba30ce069a7d58581e31bc74c6a328b04a0ea131b53451df09dcf193bc62bd717673ea3317695ea385130f6eca5839211ad2434cdb90b5c39c5a2c834bf332f0bafa315ff251f1bd514ef3133cfc3f778f6692eba358d3b5908ed52fae3542874b79fb30965e952bee29074f3a2da985bd9364134c1997cae1958236814596233ce499c4e8066114c38bec7e7c8026d3fc42ffae0c28881c372668e88c648cf6841dfd6e12c0009be4f2031060506b142d44e4c7c3eb3e40410e49402f54b72d4162ed16732c1a0e7e1b04204cb8d49a0a6c4f74c6ab686de9a1f8c0f67d29a061c8c6633bf29a760dab19032ed63d68ea60a63958f9adeaa13d946ce4d48b2428425f8dcbfb064e508045ff5c134448e51bd86b88060bd7d620348ca16aca045fb6056be32a7c34820c2d737efbf2464d0515839565d946111f1a603d52b764b8034fe0443535bd3a3155cd3620d31074cf0857ac5a6035021b998aa4faf0a851f98bc876942354e341445ba7c6a23bdee3d7f49c2a73dad651b1aaa148612e1dac3ae736b5e26aa8cb06e9e36dcaaefa1bdf4469d01c53c01870e4e64ac86b70a5f18529c18ba5500b6130049f77a043228dc7381186e2a26ec7f5077c34f60ddc1edb31c2df7fd6267959aafbbeedadb7ef7841e2ad82afb894b4a6243e442012d799cd8ed5bfdab2b91caca9db63bb768bf8a78dffa7e0dab9b2bd76a49ca2e8be309e9799c54f849cf23318c07caddb3491584e00fce2e8ff18417ee45bea4d19e559d739fa1fab7474c024a658709c13c3353e1628c9fb45d39e99ba29389635d79741c4a774c401a752ab87982aad886a691bbde4262376c38eb929268149c0751de625277c21448da2483510df5a52bcb9cc317b9bca7b5a1f4631d2a052aca321c86279f3a309e7c054799c022f694c2657697b3538eba35c540aa52e31de80e872f7c459209cac8f5f7dad9963bcab72b6bfac5ad1749734e4d1a3fe912c1c87d898975d848ec3f7680de4903cb91df820c8ca0cd514d94c5170b2f239f5b51eada9006c65e555af6bfdb5b9da8c74b65499f0e7ff15d978da985de22e3bcf21032e3263a1f370acf116a59819e2490161db70e848e2bcc1e6e435c2dbadc55ad646ca6d83a76eab3c4c1c3ed802e10cc622eed692eaae3354b46448b7c16c2623a0eea851ddcd87d663ec3abe9161e8c806a2d51973a3a77d98142c797f0e7a4bf0d74db2dd831c0b10d68560269a86c9acc0afe543df65bae6e9e5edf0d499df1dad2e085fcff2ef4980642458f0f1da94b8316a6444608fe883e08867f9c02949d6d092ad6d4a951a9df32f6dd8791029f7dbc2c6ee723a7b4ed8fc8be36a12ff5030cfaa0ecf1157f072b2d0f22586ec4a0f947397e830946bd78773998c124d03260182e655cda3cac22dcad99d3f3c21c6240844dcece9ee2b82e1de8b8539d0432b3cc6a50b00e0b0820ead876284d835c5ec7f102d6efb87f731f35b6982c2d765639b767f1f8f2c105a76a7ac5b4276fba9b521242b109bb37ffc1c00b35c2f010b1c50b868192435c38ca0b8ec47c093c1986094354025e712d61d9de5e9d7d664507e155bcd4cb80ecf8a4baab760ba8c1638964849007c65c8b3fdc2490838a153bac2238b67e07c450fc55ff7ed1b2108d33d8f5c6a4944eb7920575def1113b08319216970884c946393eff05bb8de8a76e34abb1ad22fbe699271923b37f31d6fe978d1ab2380bb0378d754e704cc8a0da12153d2aacaa32fe23d97ecf277115c435f5b072e66245e59aadf625603bddf7bdd39f40fe94a3e97e0801957868af652c7227cf365c78b54bc302bb561a7bf58eba25fd2d99b7ce7356bce704a9286c942ed56f4051f09d72c4031b649adddac284070beadf80b46412259a47de5d94e2a7ce2b2fcdb9945c9b12db1de7c89c2afd8d1827616e3bcc2361fbc4dbb31cbb803857d697278c791a784b6344361adfc8c3da00efc05283ea7c5d87323c6b65656ea4a0fcea5d3ed58e27cd2454073da065a9a2f34b410fb312d366d913a58e96d3af63e1350e059d476a65f827a78b84712e930006d5813d7dd6759e159b0067ca3c6e24384740bb08715aa2021824fe1b7907902f6c7e92f7b82427f5837ba6b04e934e6603bccd2fe476385fa0786b5c457fe885d427ae3efa4afd805081d65461e41eb4be80fc611e4527305126b963fdeadc88cf8e608353e1df85aba7515d4c07c1154745b0b2552349f2463aa414566bd9e83765ba9f974f05e1add056524196615cdf828a4c539e7157c5cc3aaeae5525f5c2b0a3dd4b4ec761ff4eedb562b1e02221b4956446c79e5eb77fed52e11a11bc7ac1e83f1efedc3e19d7a35389e0e676d9863503577ed1ba6270e76449dba527476a4523bd71b570bf42a84d9ad4309b0aa2b17204f0fac33c021efccd4e2bfb624c72493e6c779264bab9053d7201f02baf1c3f9aea7e59d6ab42b5ef891eb83e3e8264d927cff24beaf3d3bbdc04b161c78ee3fbc0a5cf53a1f2a6f834680b7226c6947fa8041fd920cd364e4f834bb893fcd64a16622b9294ff1302d4a166fdf2999851d8158a4ec5b0237c9a9a2e3ef8ffa2c1212871ae7c374930ba43e4a318fb6b918162aa4a3ddf2b3cc444d23e80a798c9ce6f45185279f18b2e103dbc39dd077aa0cad759af48e0d4510c6e5cdcc680bc94dd101b0e285c7f8fedaf923961c599c29b29438141f45c63db070beadbc3b9dacdd98c59b27506126a1059ac3879cbeef1a680d4e98e120e913614dce4152abf14d057572b3b9842660c04e0b1615596659935cea44fcb0139fef79dcbed7e9411d3f9121258472ce7ea60881f550dc25c4d1d18abfeacee44e18f4b3ebfb9bafe1175410b301cb3024ae96b098ff6d6f8046ecfe05faac7e49e0ac09d3e8001abd7bc38821d0c887b9fe35a85267e43e495dfbd3b3ac582da37f1ebba78778ea0662f98ca4abcf1e89fbfe6e1a7a24e9e1d824e662c77fce2e9eb4c444e2fcda23e498744008cb671187f1f48285e04070759fb7230f8e730a3d1f62fa426f0d9c76add05eb827ca3885a8c751328fa3ddf769a184b42ac48f75794afcb4fd39a13b207247029cf6ee98cd9a222288a6f6f14f4c724b1a26419823ccd3c2537cda4d5a86c8a7606b97f6a13f3a7c2d73503512f9f8e6123e77a142f1b52ba8d7cb347bbeaeb6bd580681460166816058eb7cf2640adf59bf3cb7634150d088c005b0d07ecc8a5e0b4cc1ed623201772c07de1e4113d79d294ccc87ea770d16ecb32816971b82f40d75788c3be47cde60f84cd23a214183c9818ed8266d0d64d344c6613b4544942eb15c223f11e6e4a82c9797827229519a3276846cf42f5ad36160782f6d247a78af6667aecd37853b0ff80358c16125394974f7d000fcd5ddb62b4c0fc15b3fe1dd42b3e90cbacf80b14063f20bade4de4068f7f0f07443f5addc2e09d4b644d1b7ad65d0e1d47ae330d511a2b4cd111131c41dbb2955fa833c51cd3f3ee5a6553dba7ddaea5f3ff4bfa394eff8393c48531e85416d9071e1b520f6241e053507edc73a51843e006a4974240be28b38cd84b24af0a053190a4871c0ea53d1c4f7c7eb44ff0d42ffd10293240830b6a944c7a305d62e91f5730120a0e4174537566aa30f7462e62685a7b184d49c92a76910e76d68f439eaa8535ea1bb0c79e06d34a65948e9eaba4b36354d4b2599c7d00a6c5bf9998daa82847d2b30028d4108d1bef6fe573ccb528ae3583223f1a3c1fda17620624c056a711093d50d555cdfc023edb6bacddacdf8424c42c3d4f071095fa484b3048cd80cf6399b11f52c7c9bae0add279e28a3583cfda8b518a7e929c02ac7ad8a53d3192da5fa1f7f00ef19c1a378f4aee03837463be46e06adeff0e1093ae9862f75843bb6a9cc07e6a8935ed230835de50ec9142af46a485b2b28f6fec4767b8c86473ed85819379a430b7e9a46f33cd319b097ed583c0ddd69d42645c596b30894e4dd03981b3b227dee09101354bbe68fd87dcf0b6033961ec02f1fddadf8c8ec7ba691f5b897f39c00219b6d1ddee0577fed1f227cb742aeb2c4bf768a0c58132415058ad1ed194ac6baec0b967b9f6a583bcf8aa8fe2ddeb08d3be9479750d91b2d6ac851d397486a0cac44045943875ec43ca3cebed951ce78b095b82865a37689fb750f8b833f3900c241861781dcbb75495f70c62e9f3b56df3a264d57812a38596da92329df040ea11593f41b30746f41319fabaf34d88a50131fda50d395234852daefc8176c17e0ea894da7fbe47e57df5e02334c9000ee6c3c96e0d0c008b354f7d30da36ea33b455430d9af59c654fb5ea8955e9a8c54e6554f246dbe699491baa02c8609861c7e249f5a3699e6cec243bbb3ce1b0efc303ea7746d8ef1e81e42b5655861086f93bfbae743723f319b22a257bee122e11cfd0ef758c1affb06543dfa064d3a5046ce453ac4461552657e76a211c04f7ea005cdac576d4fcee08df66d423ac1d7a7c991e33b134c3dd1430b9a7e350892c5169c65c038ffd6fea0e2d061f781198d857b363035c71dbde6edda95dbf2a67a35477aec85242a59be11ca4929aa004d644c3eba03eec13d810c1430d33b5b9e39d3b8e514c1b9494c4147c95583bf851e551f45dd6e7f9a25c05b9062c6ce488e383a2b6a8a3e52fb77b06658b49933e7021476a4f0aeb71a5278e0d1244c47e4385da0c377d8f931447a823c924c51f68654162200d8ca02017e33da0e52c203c952bc23cd3a141d730a7b7668b1834e36049900ceeb73f9b97b328d50a772b44814212814c6df86270432caffbb71006d14383060e3a2c2910158d0ff1fe44bcbc2de06c727b1b42fd191d346959837f0afac30ec1a4478bb61b93495fe81c506bfac6a198acb1cde9b4d1d1aa4a878f3ca5ce08bd79248f56395a5de8ad514bea9ed7b459f65dcd941cb6f087a6a9c44df14559edf58590cc7ec31550e01b2c8b6e5469f95af4fb4b5e7db8facf1d15c700bfc4436559bc54d173497fc3b3a6c259b2da7a3c72589ac52caa562f434d515b7eba4f23237b7263bac159837ea8ba7883dcb622b72a2f6d1c69e07ef30bbdd855128b1c884b8c5cc86127b9b4d8d304f7db390f8da0b7accd8c78d94605975cd0729cd3f7fd33e39c329a04237318bf47c45aaa5f9f74af04f5c7b4e2985abe75214c00c7852fc132dbb01cdc429564a7d9e4507410d35eaf1861dcf1c6d228a22ae867658017e650002cb52fa65180c3e7ae4372706d3cc5663605a405f4faf369d03737987e5412a073d7a9a1f790dd74ec3c2f043a31cf57ef4f0771c70895aed3337a42f91db7b17307895e28e3fe85391e97e65cb25058943574ba08e258d70c74469e6d4b3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hdf5fb92c1eff8a41d5c69601d12cdbb2424f048f5ccc411567bd15dfa68652a27801859ce7b186ff94c99ddb83dc109722f97d506953ae472103f1095142bba04d1dbb8ca507d9fbbcc5eda6dbe73df03db621131a041a6a77aee6eecbec0f23abbc9c238c4e4ad768000bc9856556f52cb8a621542f1eabca88c5e312d38ab0a0b4afbf5e634b6284f0a3d57d97d68a4423c624a4783381d9c33ce8ccf43c87e99ae16c1afa79a28c1cfcbb5e112ced365cab498d8d3255bdf9b6a44a3b9d9ca78a104755e2def05739071521b261c0efe0ae9879086c2d3e6e3f052edf7a462d8e9ba8153590ec0b9fda7c5cf4b1d9116f6b5b68ff412a74bd41ce26ae3e34f9bf2c60600456d8ab8f5f99338fd1ab620345121f41dfc7901e933714e289fde1f0df0e623c769ec6b34e47b79f403a2c85b16161fb55206f835114e8deac4a818eb0b28ef61ffb6756002371e1ba3b0873eb8902cc85a461577a92f020faacced3a1de5616308bebb872f17b3eab4a23845933ea07fe27757e8f4ddab99a1c73d954124169be480d737c40a7a0b9730e8a8feb0e845c19944a720f5c7736e1d548540c9fd467483e69ddf06c1337f53b8f57042126957dd64e0ebd4dd62fd27374e9d205b67316d27293e280ebaf4d2f847cffb0777494fa82f18950edf27d360e36d245b9ee9b48a6316325a06a05942fb3c73a9b8e78afd8e8e36629fe048aaa7e3be992cd9864424f4b72cb7414a965ca6d8d06412f88a526b93890e871dc1e99b498030ae72d7c8a628a9a9c2e5e79684aa38d2f299144bc1757083d189f883ff7043f0888fe02b2b6d498c864ca38a8c1af29f17653c5c6c13e034c5812f6f706520da3462927a82f610df0ac28c48941273836f30cc572475167dfe42cc2cb0689506deba7ed3cccaa9036f131b3cd462272e7a6fb6aa219d4a2c1fbc87c0277961263aa9b75f8f433f6d261ad1a3b588155c1d2836e4fc71103dfa5d3760f97081a6a9c40bdb8106c3423827706d3ef28b6e2b87040fc25966fc5ae04cee7c0782d1340d538e9b144b9668833262f603609484e1cbdd9f05f61db225f32ba56599dd9135b633b7f3507ff98b77b7060026e7490df2da27e41de56cd5d9992b6f3bbc9b0e9ac82969448d3f6e9c35540f9870c7ddb30f847f59c8b0bf259a16d9af4d6bca52fc9df145ee4242a8e569ca67ead6d39a1bff2aabdafddd9a11a8142dc0fb0f9d3b4eaed2b9f762fe221906a2885adb9bd6c73ddb16a1c3d48db8165e6b724865c733aaf6b9454dde77bd27f11faeb335902933a85ce8b24bdd3aa026d47ea85c2056522577bee72c0802821326d39ffe8e509a220474f96953872e0871628128663c500cd0015555ad39dbbc69e892cd7f6a57a9e969b20ae44a9f2060553b79961a6fbb41421c8e1c3b2c562015d27503dd4beec32b997e461474e13b975fc033c906123452d03e65acf1236a4a04d371f667634bde06b93f6f1faa08de772cb845d4d65250f19d4ea4c12310d3a3372abc7fc5bac5540fbd927871c5710620ad604ba61eb29eb5a67b730b70644b9068ddbc33a40b6eae407b9cd75f801579f5f1e7371b61b645388deec58211a6db2993bcae9134f8935f5fbd81e87fcf445911fae18cf397a22f7a305819d4cb00486c5119d9c4fec64a403844b72d6b869e20a31a8e804c406c5b54340ebaa95001aef2fbb8cb2456378d04a1296c2b55cbdd57a87c8aa44bc7611e8ce6d8364af9a5e57ec71bf25369832484693a2931e90d679d1d8ebf68078c66ed2abf5c49ba109b2f4d4d8aa91a8abf353d09a9b68c65ddf2dc64a8844fa57ea5792713c134c2d5edea24a69e2db428ea37656eaca939c319733dd876ac25252522c37572f55a9f0ad7126d6b215441d0d6c578a71fcb761abaf5a847c73b539a3bb63a3df7e59ab0384d1f6721c1fbc00617dd1a77dcfdfc414d922b101c1f1b00bbbf00201de798eda8c890c262245ac5209e827d3869ea8ce2a1382362fb10e3ba815967b61206e571fccb573f87b25106f2a62f57da0318df09a6041f85379f73178da31ef43a8a73c8274d7c7edbeb7428eaa4d307609d089f881686a3cbc7684c068088ec8531f50f8fcca052d48fd3e4aad1c65c88389f8f261e1d700b462d6ccf250e8764037242204be81c16847439f351a360a81a1471eb87bc8b3310c3637aea2c19796df6428eb8baa6a498bf764803cb64ff8ce4e04ff8d1411208213a2fb737efb09018e12eb9d4a84bb963228b9e9a0286cf99f5cf556acd70b7cfa848a6d4ac09ac3eef8bdd697798a745c1a1f82ba0f206cc54538730235260a26605ad5d118f79991c4c7a35f540edead4614a8476e582b3dfeb964a510cbd85280159e7f3cbb0af24c88798a7fd9564c03b29a6a27b84c58634600ae1b4993214aae66985411f57ec2f56e24cd4aeb64e714da9771c80fa36ded45b251c1d97a5dfe6b3a03619da0b4b045c0812490d48553fa42c64580f73dc36e85d4bf440c323fc0f868cff48135db05d2b8d88eea08c9e6e98dc942cfb4be095b9ebcbd3fe954272c16091d12b093ae71b3b94baa60c9e5bfac7aaa76e403c5449e2004730fa88f0352fca738ee3acda302c044481d454a72ce8310821303c99b4fa1e4bce4e7c13b576e9cf7e7dc2c667e2f673a2546458384d1907467c946f593343ca0db45e3dd279aba97975e0f0db939895d137c41a87a342b38c21c89267e65e366a191aac38416496c77fc757b03e22a596c6bc680bf096cdac75d2fd8ee07e6f07d7e0b627773354488af01f70fd8cde63cb349c0775e3119d29f5cca853dc007156ce1e555a22ae58e692f5fd52a44eea0b3f4bc327ac4fda51835579f2126844219e1e72e28540d148449572d0cb5056c30a0f7157d8a60ddbaa9eab369e1da9cd76777660287ea1bd641dc597904082acdb85bce3f2290a62be129ce195b70cadf0c4b059a9b822c1e5071cd4371525599093acfd849161619f3b7b2bb64e35ba2ec237daa671f972318e28429c046b6152ef8c0d7998518a6931a32c5f202ec60dee49f9ab9b5fd50fc6028a992a812f36a5f2c01b5a6719e34712b0f2f33ce3a070aed8dbaf839fe64ae4af6ef7ead83e677c5d6e226a8b94db4fe27db0038893b11b060a948993a02d5c56aaa0525132e97552a0b3e58995135bbf8901234762db9a6c73bde5184446da97227f5d007c3f052817bd1c0234dc0b00ab63c7fa19f3aea3edb28058a49bcca0a9cd779b2421e4c34596d28ec83e4f44a96ee5f7c6e5bbf988e79819e2f1c7c479ac41252c9315d7d779b1013f1f1c709ffe238d17767fc57b2caf6a48cf67f7833f8514bfc991b365f92c5e07585a3e00235e2eb6ce8ec035ae3fcf03c8c731fd25ea8e2e30b02fe40c9686ea035309756a3d4a07e1c894c6eec579be49be28a59302c0e0dedab9cdc9fca29846b49bf67006c45a56e6c5aa52d088173c756d66a8e24dc9f4808ada548de788a77912d5e7fed7bacbab47fdde66e562b2c33d338598160383348d388585ec24ee527705e5eff79f0e1955f9718aa4c6685140845a8d32c91fe7ec9e1f39fedb4f21daa8af94d89124a1d1d3f1c9fb9d91f3c0fe2ce5c2e802aaf3725492d2f218a28c3dc9eaf6133fb3c55379493b63d629aa8adb3a3760785fa45d78bab9cae5a54d57dc7b3e5a7d11bedc094f452f80d41fc957621a220f3b13d605fc71a354072653cb60b1c9eff40d7928dd29db3eda2b6edaac626187ea1a65a5363730382348439a933321f650ef3eb15edf97f2d341e8ee2308cc95cd92a87e8ec524e4bbaf2782bceec4d2a2cc277288556c283eb1dac684d7a69b93d3f80b646e4486d758abe4512172226706b417a732ba1af7fc8fcccfe3e5897a8271b7d03256441679f208e58c6c61a285b77bc78b50ae6a063303ad9db830014b3048628a1f29785d26d8212de72499e587022802f8de81026da850d5d18a91e0c2eb3ddfc772e7143aa39fa9ceacdfe90e74ee71091149fbb8dd319978422afb4281127b4ad3e9f7283644ed1594c0b4991180799dedc10e6305b4f826516f03f9cf59f7cfb49b5404b170d69c0feb30f109dd73aa1b7dd3cc84fd5699ceee7e9993d97f6e5d724d89342c2737d84e96005a703c373410ec5b5c97402942059d12feb96c3beb72d5559fd6cb1a4ec87af8b0a3e397abe6eb42b97bcd2a1d32b800d276102492d336bff34f46fc30af056a4243f505520ee9808c6304be04527c4240309d87c0068123c687903fe339080f93f0814960b387819ba3ef69f8d17b197699a83570180c980f71100c8416109a8ff41f4e6e73b229de1600022bf7c9a99236dccc47f72720c24e05ab0bbf4784e5989e67d6d72fb84849bd6e811ddcec76948f5b9c6f777b9102583a7ec6dd1ee449d9b7ac7b5f76cf4e534c721de4308d5f1084b166ce7c1e7b2722c8447611268c61b240d84f8e35b054353e8a8b7451b56ce16dc36abbd2b2c8a9075933b7fd34360c94f6a8f5b2cce2ddad71eb9fd7149dabb2c7eece3be3a2fad887c24956710dc59b8909a60159cc0d1e10ae098a1b07c42c962b2c3cf0792d394344186f3bb749e300cf3a3b2c745e88482c2f2f5a65a37d0b2331f139c36c466d651d758e85f41556d1728cbb85f7838d4ff61ab50e7afa19e8b504a94add6c50b29349e034b95c3821182ab041749e99f4d66dcacb7e990152fe7d7ef98e7af8403119fa41826636ac2b758ff8624f64a4141a58d710f5a654c7f41b74f758571ce7fbcc4caef73ddfa7d1728dd3c586ab16a48b47e996a4787217105d93aaa02a5bd60343dca6556def06b89d94f522382cddeacba360c253cdd4ab34dea08aa2f45f3c8ccc5050fb8701c7682aefba7bed5a0b07a6ddfe565929a5ceb74e6b82e749c0e2a9f20be922e7fbc8710a17e9f82c3bfa641576eb6cd98a7470b28224e61042f5e7d777d770a02d4942bb2d41e8a386d49a300d190f3f18ebfc852ed9decfcd28f2e23fe822e9c883feeca5adbbe753cb5526bb44d1716921ba4d8630ae3fe550c92b60e44960d10e4cd27153b4b8599a483b0c757af28226bb9cbe69b30e18df4277511bca20597355313d17f6144e4e2ef4df17fb6efdbed08660eebd8bbca45f47ca166e0c462d04b5dca137e15652f2e41a82eaa3c12c091b1a963b752b343f91ead30e312060a453429bbe5ddf87615972789b82aca050400063a4f5e68e40dd7bf11d5db8b3ebbce2b419cd435532173a54737b18a0a55717d3c25d171d4b5f4870375976bd0bf320eb504c7f55349adfe5f64debeeee3a4bb2f1d8a00c3d001ac1952e8e7eb32715eb99e074e2445713de198acb433554aa4b4e47ed6e352632b4cb21c9b455b55aecb5d1122880853ff47302ac8a55e865118f1ffc0deeb39c357d1c9d4ef8a136e41b8099e5e0d8aed3f6dd304ef31e80fa06c0ce9b66c86bce0731b8e12fde251966c63;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1df065ff32eb9f2a824c5a5944db518874589d4cfbf636ce36ff2142c029c46c3ef54d3649f81c9d66a9f94edf0f189987ff6f33c961a4d3a05fd3423e63bfe2d1914738e1236eb2ee380d20b2052bd6fafb59bb6e2e0a2de5649849bd0758c7afd90feb1febbb5c65126915e4d26ee7feb6557ee622e5892f51b46b0e096f64f46a8843b63f73d08f21637dc2b7e87e6ccde260166a6037fe513501c2be553a78022d0820d1ce50bab84b75edcbde1c96833c878eaa094afa0f9a83af7f58c2832734542483774194c26c27ec6cb2e7f7f3616c0f579a4959b92f9284b06baaafe6658f3e61b5474e1388e7b09277ef2a33ffa9788db26e7cab8809d6234576fd9f8872009657b14c354ba4950ac9a74abeebf46890b95a8b404e917968827a892e3837ce69a715c6146c58305340822150c1fc3560347dbb09ca83e15eec7120e046b3563d3762c50834159e54f6bb33e64afa7c7969e04c2831d60dcf767209e85830e7c94dd1b40a57180d70bb4777972cbb9cfefc30f1a6c7d46261081da9212f550da1b9fcdcd3e48ea484ae5563c176355d7aa798de4e0f2ca5697560735c7db70889c22d6d8e38de192ea07849b137630f0d83fc50310e3cadc81311c1fb3e9e4516e3c7ea83eb19c0e09c7038f501e6d7df570794ea4eabdca67934fa2f8c98f91e09f6946b26727a5f4cea1bb89309e8387f7b441171a84486f560910f48055dd315d3b083a4b5588b287c1f7231c9afc243ee8dbe2ebef67d2dc0ca99e2d7205a955564076fd17cdafb992c8e6a84b85a613d514ef8104766d7e86ea309fa4f5f2ee8889279c8bff3c6d4da81aa7a5dca96fb65eb99eb162f3ca945aa60a87ca63af540f35dd3e701228eeadad8b9b50b8880456023d28f9fb18f698e4a9ae0bf668f5b8fe5f84e5a576ea00464d7290e1fe9aa189464bdc4b6a34efc5db8e1e554e228e6bc21a0994333bb240199dab4e2d30a29fd401c0417b0a2afa98e080377f7d4952c8596a9e65bba37951de2465f005e750196134d846797e68faff72c519b042ffc0ae0d7c07e225e31537de568a8b9a79638904a5e43fc8aebf554da5ba9398d91ab70324560bde7ee8066f0067c4395efcd8642bc3a1d865114c4c1a52ffb083b38ac7312e1f16873a9f4f801a2f4099f2ae6493225daf7a8f116f6a897ca83c1c158fe0bb50ec337e4ecca2aed42a93b83795efab288fb04134db3ff071a0c8cbbbf375ee900601e91ac1da5368e33705911e616c77e59316ee8107521652e3b943175c31f0e9fbb05224c9e9989c88231c8923f20f59855b6edae1bc3129c3b96ba7426150ad1953e0b50ecc76e557f00fa0042f8ec31877b06e14daa0690318ea342508aec9cfbf901b4692a44aa9f3856a286a727300c3c7db706cb0196ec56421f9ecbd4317790e11241e3d0c00acaa5df17474a37987b1d1295ae16ad6dab5e9ea1ee333a813d965a32246f3ab405bcd39af502714e4b6eb36eaa8d391ac61fe8a56f61d0b8f93b82a2bb4d967976a04f0cf544f4e2e7b246b7e0731a2b633cafb6dace81edc5988dcea1450ebeb91afd252a1fbc500c823eb58fe1e79eac8bed20dbe862d2b1d6a314223eac3f77b02f1bc9e0126f08014d60cbac7a69cf6606b0b1c6ae3a03408d64e0c1b06506dd270c00b323bd4116c3cd4973eb774a9893592d0d61e4f36a615935a2e7e05f764242b0763c08dd068e365d9e4d32dfe1395cb5beeacff4addd8e3940a9e5399b09f2d83e483f27560ea67ded308b390732172cf041b3f9fdd535178f1decf3bfb5c27f967f10f20fd318fc3d23a0ac8c2e33d1fb894aea11a81f9c30887803a54ecbfd7e6cd68d7ddf814c03e9b08d2d432bfb9801136a5d08598fc56d9efa65cbf9b7cb739c7d2a0a545e786537de1767d9cd44e399d52a10d62fab07bd999880ce69b5cf801b4b69790973e33dfe6758abf303325e0bec1dd410fd6ee6a210b7d74b279498e7e30e804db481cdf4dea79476d4a0b27b2af22803e4b138e64541c72f8b82be5795f38d94825137b97e19959ffb782a88494b03c8ee09982ba5d0cb8196a1c60bee9a83cf2d79c58cd6666f3f98d7d99a252070f1346cb7b0a96b2c75d4c245d519be29e62a1286ef46bd2eb239c6b1972d456fd9a79d73a68c71b492ea00a6c9153f3b00984c4070e2df9c8383cf87448bad73f112b61c47eb41639edc6b064e715a868f79c0e61db5027f3ff687d43eec672f2878e6d0b9f8089580e85b22daaf572572702b01a4a62166c520473cc7b6fc5ff4360e620d5e769113898e797c2e530ea8e7f55e8d26823bca073162e22cc19d3bbe1c6e0ef69b9a735d0c3c535d9e79079b9088ebbb36d901714da578d82b1a22c0d6f51890cff4cf8baf1177a3581dc509ffe26ca81faeb7e9772d5ab36aa3b51dd60567c2e28ff32614a729e21cffdb43d8cce76ac9e5c9f53b74ead7f88931bccaf6194d47669672361954a7c613fe76720aefa26f6d07c93b53f7f3261ea4250ad7b590ed8a3213b82179002db21c7c33a9d402b9aa2da0e57e6e5a7a71bb8aa659535c34b88c988cbaed1e0e0ba4e3b188a73b80793646c0dc5ae4e18fd93fb2ce00cd645e50c2147e07e9a94fc0c9b2f010b814b45099c0a251391267732e964d6423405a4831f98e8762d1e9e45263c95a002770d37190b8bc8ce37d2e74a2929a9c3ffbeb999dbb7a88aca7fc2cc0dc5db9b18fc883c77c9d1b2711eae25cba5a3b41d24705e2296395f8c522073f45a3c79c65a494068f235745d6e833b52a9571134478d7d696aa8e28a734a3499c7343b5e83315b31e387c74259d3d3c8e2dab4e4bb9a837817364c3c657cd86ad268ed172d6ba1d2302d82ad2c3c91a5d21b6d3355d4508cc8317aff29864d65571c4e7ab129ca3c66a2c7e5f86cb36cbbec082c135341d6a12e5ce2fa045849261559a8d8b682fe988e9915bf1d8b019dbd5d2363daf3146583cb70d0220a604fe5fb204eaf64324df156aa64f122b98dfe3a4c3e4ae1bee6091820b142eab995f4ee9d94dda8b9fc0c6a16b061ca91e0e96b371ebd1beeba7aad1422040a96dbeeb33c41d7dfa9882222dfa431d2ac2fec4893586a12aac338bef82b76f9b1615aafeb22c112832968914798e3770065752ba9c7b50acb39e9a22ff25baf1c5bf72c8f6d2abd4de969ff830d38768fe94ca66f7d4690e792df142f105fd5bf136682587025c436644569500af93c3ac4128cad78cd9b7b1bf182baaf7be4650193b6d9a8cabe7231e80a5a60b2d0ad7df1064cd9bf77e2fab8743cb07f6bf370cd8c00a137eca1f7c955584e52acc4f87c37551951801d049604e7209c5c13d2c39a49de30aa0e78ecacba7393ef4ee63e4afad205da424405e464cf12e816491f05d5094ca9dca9121087188387b143b769e1193f94696c4bea034fc21534f39aeabd2956f438e80f5161211113bdcb8d5284127f1b8b8b1a6956adb14d1f5cec12a853152c9d79e222b9e591b461be75a086f92f33d3b3906827bb2b13cf7a65678363119c9c7a77136d5e767f95cd1473765d8739fc7b4dd3459a3e59d86ea0439b775263bc765909b8929fae76e98e1a42c6524cc66684567a41904cfd2b9c099d2b3259d1059ed85f88c66a31fc2b97dab7c089fc4d2c752d0b9046f19db0e04c9c6cebced410395e85c5ca99f7479a808cbdfe05b32c0c77e2c4622e739636a137fa4af664d94c5aa85ce86129bf5ee6452a15def176e826b328b63c5a3f53c074c2ff38388e526b6abd5920495f3de6d3cf6821ebbb7981cdf5145394e284f168bed4d5c2c5cd0d55e0abe6a9bcea79a16b6e398c6858d3db15d8e52cc314c890f62cf2f31c68086c5a4fb8573c251cecd1a2886f2345a3f43bccb572c0f21956d0fc4159ef03fcdfee4c425834e294b739c20e1c143093f31ab9a3115de9af124651eb2a947c18d8e7e9e946086d20554ff2d990c96f09f9d50a586408e439e23c4e8762d09b861b864bbe34750194441f23f019aa625d26a5a2053574eea01b03925b08dd1bca716c296cc74fe8857ad08ae6481350cb649f44e69aa4d62831c9c5c04b786e08fa38be933603ab0c63a73b517a6499fdb945423f7be11482654e196ff593fd90dbcfc1abc4e51de228cf104239f8dc748c7ccbe558e067a3fa90a8e6680955467d13e304aba9c0b76fcf77a9d321147272ecb84c6fab9caa270ca280a77f42dafceedca23d91b8980d0f914a63fba6a33dd0c50ecbdb61987d3d039f4dd77948d05efb92419751cc1977a859d8bfff2bbe98f57ccca35ef59dfba9fffb742b292797efc6d79987d24e4eda64d5a1973f0e5ab1bed527b555abea29ac16dd9937054af64eb580c43a63cb7cf23879879f4c34c41799cfee2d53b825f3b130b8d39fb57aa15ef255ba94d910345ef4812b415a8de80926b92a955a4f09ac077898d0607f6f983e7431ab2047668064a589cd73d5b557c61a8a05c07d92a92be11245e9a23c4a58b45d6801c082440c83c8e5889f58183fc0f3c2c00aaf3b7b739dbb389b24ef75a627df34a607664fae2e22dcbe583fcdae8f88b7eb184bc3b4070a18c48b23ce2d6e502bcfc13c51d7d809f93babefe0090a32ed17157f70be24e1cac258a68fa44b989ffd642d6bea24810db13490915695cab91893083831e9a2f1bc2682eaf29393621b14b70541b43c8464ada42a82dd9bf02fe2ab37c3b7cd04b9c04595b3f833f46b0bb1b16e584139e3a483bf42bdc8b978eb3bcdb5f37535f3a5e90105bf7e08b4f01a5915536b2249fd8d67d67f18db1679a4327a931a382fd912181d17fea5f0cecd58debe0da83cdd2bab789dbe4be297fa8dac1cc5c7b4162d8ac7c455bd82676fd217f40f728a50f0c28eb6cb688422cfed827e91f04fdb63752b3b76aa2c24bdee7bc9fb68b34dbb0aa556e651f2574bd4275cf46d9345e65ec6e3fbfffed20766e552541234782ca2b41ab0bb92f1b8b5052983acbc29b38da3df0b46e7f85568c19e764f7735d06be27ef6ad05b498c25229e01517894420192166c002ba140dcefefe337230cfd119292e8a39f340c56d18e9d7081b505075e0dd54730425454c68909e7af43762ef4c82e59fd2568782ad9c6ff804a6d2b7d3391de248dafbc404b800bf261fbbee5e342b272d9b14e70ad6fe41ce30740d5016f4e017c67f8348b47daaf0e4451b65cbac4bfb7cf382dd299924af07c770841eb4ac91d42c340e6711b5b5d0b6be98cee69e073a9f6d56afa406995d77571abd8e25695adf92ad3ef7095a0be325c72d8228d09760fedecbbeb8c7bfcba7262769b17efac04a3f0e2b7e48eb7847c68c6fc8f0b3da9f008345653122e9b13e75c7bfa4fa2d6d75acdb1b139be899d62981192cd0621118fced1c182ef58a2de2ba8e427d53f50988106005db55c5e2cd616893ba9e5f167f4080ee7d0e2c1d8659396126ad423368236a18b123f2df0b8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h93dc879e7cea5e3fcf6fae77a6366aaa6befcb4b6735dcb72b859ea6a16a110134ef2a78121920d5e13cf3f93ff9bd867c21851846a9a5f55b08ff7bd46f703918c5a27c19679203ca8e53177e088adf8c320bd504eb398c90c2106a9653e62af9a26c3e86ee5c412a505c932beb75f58a15fe9b7f683cf7b4ce0af93859526394e018baf9f3839ba66eadd39865f2a867faef53e24d057401bef2663b27e991475515a49f9571a9ff9e15e10cc1210af16f757ffcfd0536a2b3cc2f6c242428a72d3e68c84507da8037cd2eee41ff8973456cec8e04e5fb413baee32045d00983a4d22bd380970081c6a79f2187823afffc887092ebf0b9030494686da18f0cb0752b00f1a6798fbdf0870f4ef9274989ee32cc854c9e3ce8ca4560ff1daeb016152271fbf8dc2964e6cb6aa6e946624dfb3edc762e06beb516dd1d794cc8c0f5bba3060cd33a939624f69d8fd02e02fffc498d2523778f1c3e3d57bcc0678323f8954e9f1f7c860919fa89986ee9b2b4b04847866255b87f6e430ca0d6b25e450e3a46177921840a664ad42baa736d5738a582e1cc88e114070d79cce56e8ef2b8895a13b99fc803ed8bbef8e66cd298544c1b2a17202b1b83e59f3ce1d7e47b676be21a7df7db50af410acf9f6d29fcbe77a3b0b3253f05e9a3ae71d80ac4a6b9ad5c4c2af09678b755f2271a0b337c0b1055764cb4de1e06a390a5b5b5ee27d4943a732c16b9f5ca4fc33eb8f68f4fa89223551d18f781212b36664cf606bd8ba017a45b42e9271114b7538f5ed4171d08913cd0f08404687a7d0d85e5ae003292ff048f2ce3fe21b05b7281cdfd8cea7abf98ef3721d06e475443751cc503b76e5046dfbb75e0f0044d979dfd3fa281c8071e3d8b0dd6013f31080c089285c456e00d4dab0711a12e18b72d8264bce91dd30bb8703a3cbc5ca299fecbeb3940c47c69a94418d431a4a2372591e27e3f36f2d05dc1cb40eb5c4eb7386616efa10bf45f344bcbee76067430bf89b33a03ab3ccf3d070c4133db373f33dc96231c6847bafeab6cd1c377bdc51ca55f31508eec8709418f30b134326239a68ad0139d44def29be1dce225a66fe2ba5da964594cc0893f919e057effed723221e2a6c0b2b0e9bdd10747a424b8b89167809f60907091cc5c9386f5b057cccf3068ba4fde0a9e377b8f99d7d11abbb8a7ff2692fc6f82260c82c9f9384da1e59cb6b7443811fac214bc40af6272f25b70da09092f780abb77b04465681d5992f717e46245048d5242cef3ece1e50afed4bf17ac3ae6c712e209101e66dec7075e25055b5dcd5dc5eb177d9c97923364ea4af2687e3245a820fecb4fc1e097c307f01409a69e7bb08fbec1cf8516d9c362b7c4b695d654ee85faeb4c2db145bdacf3c6f0b255d91c2bdd1564133a32a35172d8ee1ec86d87d7df3a9acec4727e33f14fe6379020254c0b748196fb3a99ec28d46fc13d948665e1b1fdb6a418a51f9b3b54be6970845150a85a12bac4ce5d40de8aec517ff400d6ec5494ad7de9f3924da4cba8398700e49561400bc762c0014082fb7cb5c0648d2418205019000e905146ac99cb6ba6bc68d587964ac72c2dec9f852ffcb69c14c766f4c015e27b58b4e25b5bc179bf4659643c7aafb8f0106531d599ae1a4571e8817b0150d3aec94393d43f8ee4309cd38731dfb1dcaff8213da5cf0c746e2c814e2c7a5ae9bc2987c1204bb8f053b38102a0f60b2f03946398597faccb42f740d34bc360cc17a605590d006c1743298a7002a581aaa440735cce26f311f41e2c86d7babcb3bf17a6ed57440a7011a7ec77148e256584bb03a326f35bda07aecca15754f9b1ffd923b457c9edeb583a6ed6030d9f3ccf9fdf9e8d36b2620aa17b84deebf9dced59c0ad25046d109bdeab785b5c4183492bbd3a3ebdbdfb7137c0d5c428e766e8b3547e9ede4678fadd82942a67ff066cdafa2db4aff70a81ae1cfd86d65ad7267a8fb16b588e7f36fc9a4b2f144cc757ee65ceeec981a70e246460aa55396fd4e410f7ab93b44ce2f7b3ed0fe64dad8c216857009cc5178907aed21afe5f1ca2ea7f77a5351cb26fdea06c8359e1c37c473e6334f37c2399c74949928a06f77713c694ab603eacba66a98a50577d36f13fccfb78d03a90d7f11b2f77f96285ea257e716ee7aaa04150ffe529414153c6e5c681c78d723c9c25baff7734f70e0a7c0a047f2aa7e453ff9e14c8d542186f625d77c01821cbb57e56f745cdf6ce7c47edbc2afaf865be97bda48a52d08b4fd502eafd537229defce7b20a55bd1127cbb5091a4a8a078ccecf93558f4c4d87c3d6b8b29489d352b6c90bc66e8276fc8f49fd0c076403b88ff7377b247ce46ece231a5c57fa1394d412cb088d47602f1ed3312a2c7d1d348ec62e518c7be11a4b4e943af9d11a5ede6cc7177f3cf33f43e676759a31d77ec81caeba8936b53a379a7df234d2123686d2a455e1e80e058740bac74c9285bbdbcf4972f4d4e799986ead6e51b80916558b105e5e00621fa631087285126a0af5f22a171b32671e4adfd137cc747ff9a93e21937ee3316a58812a8fb2de8aa0154ba5e82b770d576332cb5517b01d7215e4f60e48d899146fb61dcebff9d4f2864ac5e98e188c77816db56b410735f15c2d457fe296db469a2f1a2a96b596faccdfce39722c250cd5aeca5c876ddc5b5e9435976a7a51d28c7b6faf98c3ad1cd2ec0db5655f504b18121fff5fe52592bfd0fcda7d2dd968cc09c29d9be2042d9e515ce74f48e04b4a39479f1764752642ecdc7334884f4f6bc34ecc01f513fcac45279aa03a26be399ed27afa121a1ded01fbc01cf545a16c9bb13fab5223cb0c13da3f79903fb6e9ccd7c5dcbfb38e3c335da6f63079641c82171229451269554460a9cfc1e022e763f31679e3d5e487fc6046b57a668427c82ea655334a8c80c670752b15b170f1b74a837c4261576b683a30374821a8b1e9d965fe4c183588b79ce3be8464dc4ee88e6d91ad4efba94630bc59cc69f4772d14a3d3bc2fbf00a1ee0e49f4078b48b63838c2b6fb736c4e439a1a1fb315864c86a848541e7519e0fc270fa17c9ed79831abda2de80714eb7847b3a07b592d4afb2ee63730d01dd476d2074bce27e440f94d5cad1b0760eee28f67dc5270f12e6279d270c8c9e7e5bd218b29c47687932a821876a855b99d57eb123228bcd3629c7f63396452d09f708adec2cef53394bfc61348c276d270c7b4838964fb4c3949d902d280d2ed9782c721f28796ab137f253a04da96d26b9265b283ddaaf90eabbd6c37f0d07f1ad5bb5f44eaaf034b095e8194b07c922800b91e733459a032b77eb1c7cb434277b0d9fc5fe94fac61f2b5986e3ff21fe8dc4f1cfede6d6c5ca8acd6c0a48704170d82b33b1f934836b79c3ee0872cabe862cf97298a90795bbd23ef5a2ef85f48af2b96ffa50fe7fbe3bcc9fa567ff73342b94763d345c540ffca20569fc53e6b82598338dae4cee7f43ac949fca7f978fb104056a26ac3b54f19ea5c4ffbac7f770683185a6b9f376b01ec1e85f1a83a9aba29eb06a22ce5c489eae304a569fb1568161ef5e30080984a5739230c30ebd5959a6399b9fbab7904ef328d166bed1feeeb8f682a79af86005c678d044891dbf4182c918fe99c15d0ca22dd8c3b7d2140c9b8c61fed1463c4ae118f8b7401997c2b12fc16d89d1580bb4b1fd0a48183e5d11312be7b6a927551f8cc76d6c86461708bcc9918e6ef0492a80a0b5b9a014dd679aa8e8b66e46831d8966c12068a8888553c22072f0f8a688d77655d08fa30284c73f85a2afe1d411d0fb53fba4b653d2734a261050fefc0d84c2c0dff4ac2fe3685ee715ead3ce14e4e8cbc8f26bf96704603d9f8fc2a1465f4221ae6c4c755b15af620633ddd324d241050ee04df1a78cf62a79d91132edfda4b5857f0ae98f8783d06f4b246e1cc7c38a5798b79815e3317d237dfc0d98800183b8d21b87bf53206edd6ece314773c8f31663aff13b6480501e95f4f7480bc3d8800ceeacda7381e5224d4272cacb0226cd6712e313ede5f3e7e87759bb480c6757f181896bd66a6e46255026abc000a8d8d82bcf703717834a011904eaeda7e61766c98a624cba053962f812a2394f7bc0da8d8416fb09f490180ebbbeb9784bee5d8ccc1fdc257b482c311151286292acd99c2d85de1545a83758c21859db56e0942eb78a2c5f51052089f21e2f1637ac626b652aaa03dcfc02f68d07da020c8ab818f69d13fd226627734e0ca0fd01b980a0a86251ecf19652d0076420d065e51e6183d22b08ed371db49ad736843fd3fa406b997b198711f7aa38f9c70deafca83dbe40fd2641de4266b89fb578a1abfdb6b0ce5e80c85fe54ed1d6efd184781ef32c8b17694e6d680c059492a660d05f74f5d5b9f4b89e3822e6065a06a7d2c1e2767b5c34241c8eaa15a26fc74c7bce48ab95410e16108db08c751796002fbf15bfcdbef4fdb5b6cdf47952c9fe870f57556a24a7531445334d7865fb6177e3f0091eaf48107442f3840b77d87bdd4700d1403abbbb444a6b8309a3d4f70871078fb9101ad2fd006401d1488bb18bfd1aa85ed7b0aaa9c4ba64e93a95fe99fcf261aa88dfd6affa2f6a893069de1b028d78df3af514bef5decd2040fad473ccf453906f65d392cf031973b241ab4fadb43649b9fa914f725be133763a7ef19c78486935db158d843d353d5784d4efa93477dcca393d21556a8eeab0b3f8d553527aeb7ee5b140a6486073eb6203319c3d33641085f24d22ae518647bf93173dec86ba68aa0a0c4ff48ad9a8d9e4b6e80e3e5f20050b96ac591c7c9e0dfdaa8a21a7cc27f62d995e1416fbbf6911c72e02fc7ec344cd20bf252db49bcd841ed99babdb1bef031e49189b44a0d81dc929dc273a1376016c58365738793cc426007d4ed75a895d8913d5f849a45ff53c85931183d587e2f4d62be12b425feb1bccc770941167ff1d4d64b9c1d62194ce9976f299c03a661cf964b969978baf66445d139bf0d03288f816456eb3974ef5067898d40b593f5ac4ccc6ed1795f633d68add71e653bbc8ff611fb794ba0fd7475a95b8cfa376e6d395fd096f0dcc53422f70a0cd33d24098221cfb8bd14ea629487cb79be04f3f176fee25376f83a3640db5248fabe6d3534aac8d09524e4c4e75e349bebd6411cf02edf82aa774ec8cef3ba83411d89b9f50a43431c162c7d1b45adec709137da99a3081c5ba79f213c82d74d72de0630981d5c43b786360e41d05d6fc4bce54c8a482bf0b012e203479b24e9bbba9389a985000e41e9815225cae5f0bd7e865eb1aa3b51ed93a54b4ca145c5765eafaa2fb0b8cc7352aeaa80f47b6d0c9d43b33b039e745d67db1cc7ec431cef2ed3afa451ffc6cfda3f31e249184ad4c0f45989c98047da636baaf3534a2d29dbce06f3724a2c90c8569c3d5f72534009e76aead8de49755de1a5da9e4c703e3a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4e8f4f4b56f9275d66b63e01e21fb0cb6143a105c528cbef7a143d28a8ba5343e2e015996c4e091475b0926524632324804b0c99f2acfee921fe3750206e21b0afb370953304d82402b1cdf2e53a2e67247dc726c7dde9d02aaaea4cac9c91972188b0c1a73243c6a797d3d6cc0ebde05af5cd2c08277d8a39e04430d26dc98842e949d06385853d7ee439e3f70bc8400e4eb6b631f6be82f244a2a8acdc9e4ed7eef68921bdee358fd79909bdf008cf83511a0d39ef6e594be95f341065681189ed28f6783546e2e0229de92453c0938953b089ec3a7e86e243918ac600dbc93361870a80e5347a46f1d397490148a25b0e2bade148540b6270ffb5e4e5afdfda7cfed064ef7fad68d59e9869104c3979cc12cc5bd2fafca23cc859e1640b77985992ce92a9d927209418e6f3e4d3cfdee1a6407d0db3e83d43ef8053d5cdf65739656af7ca1801798c5f3698e557af79090a614e34e549f45b87a2bdd5dece38a1f4986c29fadf157c365470bbdafe80e90cd85b3a8674d6cc2ad3cecda011023d2cfd2460a9ff9c5e4629d99654354c88850cf18ff7ddcbca1e14b0901bf3926fa56b2f07761342c2b76d975100bc472e86961983970d3a0da9ced25042018b920eef4e0c942d8e10632d6fc89df11c5f2a27b5ba7a3cecdaff1e603a6fa9211b728887923fcecf2e36d2680ed5abecba208ceae9c0babe6d2e2facfd51f049c8735f91580e55ca22c4a9c12384db5fc52bed165a18d512932adaec68ff6ffc2d2b033d51d8ca9990040ceb70715db82bd011dd42c2bb95fd098242e7ba6a209262f70ab776dd120cbdda757ef282386cafb2b96410110d9b89f4c4a9c71c16a38db4ec838a50a28d988c350c4f2c6d078add528a819114f3bca80fd1c5c172ca991266efa31925707fe40ad386361200598454ce1938890b0cbf0df6902a71ac1758ed7c58b6ae9e1b9e08492d57a6618b0452d0037491952e83d07c9e86f3aed0e908387c5e7b86396fa306f49886d2995dccfbaef48d6e60098a0acbf69ca900a882bb52f25668488249a588e768ced0cc909377e6521b6a3864fff37ef2589f5031c188dc8f77d24ea4d9620118daecd80227357003ed6de89a54bf3a0c8d014370075c8230b3df6601a374e92a8c54772c99b4715d253d588187ebf36905f6757228820d52892df341e10dceb166ee555d6e22ccac840e6cb1bcb078ccd7a36c6fbeb1a1719117d9824d577aeb78a598a908ccd57686db2d74e4323fc3afd8a9ce14f544b33ac4bbd77ae843dfc4d5eb0aed5481fb0f52f38e2c27703bdc817f6753f4586686214e5daa0da9c45ce0b447f84faf0844cb55d03c9d89d3eb9850997fb68ad2212f5d3beb4c6bd20ae5820020e791c327e2574dd84e84cf0adba1ea1f12f1df551424efa5d7e14982e6c6bb2428d8801f778660eb14617b752d21b39efcd59bf98f4ae2cb3a0e8ed32c02dd9394c31569c10f697cde5e461a49e1aab7b6d34a1a179b1cee93538df3c18b9846199b0d1a59843aaa4e81ee8845117369962ac9f5c64dae9243cfb754babcb88419d259a714581b4d435b93d700c62930f612a10348e4bf6a055fc4fa14437e8d804563251a66bde8a088d8dac615107510248729626d66e7879a69b31c0a08d201a8eacafd936c8aac1d40a8aff9f1c9166fcdb58c2f0d55bafa69a17b11d7a3602c41cea42e1ac37888b3e6e150d6fd5ef26c5119ea4555c9427a8c4fe8cb16f7053f467befac58629aca0227acdd7585d93bdc44c5ac4ac56c3caf4c093b4d66d2d9a529c3d2db9b7a194424f576ae057e0a936ac44ccfbbdda520ad34dd79d264080f29839de31f4f0a50efce316443d2d50af72b9ee369a0fc55adcb689032f77184487f1149bca36d04b298fdf889e8ed379778a4ca6d2ded56270e1dbd4827670460bd10dd1d06bc70739762c20e4723911f1f0d325dde7b13e5213b307283b946af042478b9a04c8f82e4e9d62da483f09dd9bca433850c5366efea9b1947a2dedc3aedf7039adfbaf0c550eab8dffb2707c6c46ac96663bfb9b5cd22caef1be63c6ca11312beb711883deadc8a2b7790a3d0910166aa14bf9f922da27125a76467f9c3518ad560c7314008aa39977c450c1e7bdf3a24716c6390fba32425a1531bc2862fc121ebd4ab697a1cbf094cb62dcef40751756dfa505e68297c578be65f892914761ebcf5c470260a8d2f7ef6d05948906854fdb7b987e11e422070ce097d2df9ee6ceb7ce9954f74a9dd01c19be8617ab485ecd19a7e05475dc974fed22a2bca7790d72bb2f7441abf7e2e2dd1c74dd7b17bae3af361e56230ba288b86c27007e9894c0aab5cbf20d531b4c66a660fa974940f65d65e12a87b6aaa21a08b89c5b1835b73c5c8ceb36182fbf0f637ae1483b0607dea5aa9fe7b0bfe9e0e2084a091269afb5d6617e05c18e7cf9fd5b181b6212a470c8baa9bbdda4106f2f9df437f0b572103aae24ac9aaa5f94f73e3b1bfd40d74622db7bd828fb315a16e1e131960209299b506a3dfd115192f7c2b5a50f67fcc838f37822b4fe6f61e72aaac69753cc2ff352f0ee26c990ece00bb4634479435fc6ab0a67195725a914b3dfeb9e298aaad0d0a6e926e26ba0cfa09524bbd4cebdc4d356a3e1adbf45ef51e18eeea7c0b7884c8c794fd689ba6f304b7ba527f947450399c2f9a050ce0f895ed6176a6606c31e6465934103042823d45f8e43324f7897d7ef01c9a88751d375fed8190235e5ce697305891ec50ca915fa711f5d326a2f7d281bc75f59c56d8f53b62a6d58e22d6897a4269a53bc6df067c8e07dc3042caf56784fdf2e606b9251fb4160f100ff7b783b90ddc68a3ddcd4938ef3e4c3b9edd17f3efc196107a7558e813ac7a34719347f477ca726f4b70376ac6e0a06ac13b375708314eece56db1bffa15814f17d76a344057db8019803a4a9211045b25082fa026055cb4b6b21264e7d6562687176d0f50ee637c40df89388f0df882c0011b9d41c6b1ace13939ae66abfe58420cdb912ec4b9d3f4083df2e084c6b943752e2ab85accfe305a7fadcf2308b76fcb59cb5a72d6d85dcc62bef64a1e02a5b08de37268a347328befcd51350868fee9b55ba70397089589bcf34592d7498f3ae4ee6ba368f75dfefc7496c7c62a37a6127f5b2fcec88e3729c1e6bc5208c5a9b737ee0d291130de99289b28afb3aad8d10aa970925d9ff337479a0276af8e7ebf606072f4f037e99693f0b93fc2c477963939f39242beb721d41c7199fe82cc39bfa9f698ad1a45b507a2228d3882be634822e5427350630ffad342a88a5f4640f551e6799b17138db919ff746315ec81cdacae4c0efbaf1c1472889abade6d033acd12ad05c27a02af425846480cbd907c057be1e5dc04edfaf9f4f80f4385cc9c6563fbcddf6d0c841217d8cd02c7c7ea65c26c2261e4d30ade360fd0a628b4b85f15c0b140fa97d8c09b948b4f2bb301abf27b8d16bd6b1da64da6236fbb8abe08cc2c925c7be4f4a5009220aa3338b31859b66f2c12b94b23104b1f795b2395f38d5e7505a28cac18252141fc8dc5935d84ca036780f9e901f635ad1fdec191720761effe1b8745ee9851ed816755c46afda2d1c5323ec90e694001682b1babb243df9300808276098ef4280751db110ec6b0e70b77674901c9009f85040ca624ee83751546607ceda3753dc9d0231cf7c16eccf4b39c77afe566c9d974f1d35b4a75092dbddcc95ea354e107921a9a97202e2a076365ae97fd6ace5a1ba27ba77d212ea07b6c40f27242830e1f35221a0c407d50b96b05d364cc2ead05a25be93c250778e58f16bee71457c0c7a1b88c23398131f1f1c5447f53ebf12bcaeb39ba067e62c9bff8dc7f65eca56cf52ab7b957d7720a88108f8dbcc78d929e6076eb6d62e329b23722a2a253084f680eb13d128ae49645b6bd138c53fd56527c6722b4212d2b69ad66032be3ef56406d840e82539438b5d164a655eaf01c1ce6bb48335251dcf7eba6487c6fc87c8e8acb94990207dc4eb8137419f2e850047ed17862c955ad84532b2a58fca74b21daccd51386cf9895c79a9a8b6e91a00bb2b0b81e417be60a3a202abd80d30843cd797fed214db6e435ba998c5c19831dc50d8f16a2d880f689f8d21bcdae9e5565c2633566c957b844b7af00cb05089cef0e3a9bb7fb6a2ee3515ef75b53e9d7c4ac48cf6935f943c7cd6ea7d55c15b95d30f60afa5a6cec18d7e9311912800c33c343c97ee7ee4b8cad3a940cac7d35299652c6f2d30cff38c31f7e5c9e1cb88bffbbae549812ad54eeb489080397d9a67e285544acdac24492e9b0a1731d8aef2e2e52e3af66b4086239ecef727ab652b7963d0571430e4fb3a2e98df3c8e8251da5fe886f95a89aff361d93efd011c076ed3e96445c71ace219598223c52b2870fe7e4911969ddbdaa6d9b7db73327c5171fd29856d634fcb617b5f9ab98b01a947b654dc2a32161e0304156d46fb8ed42db51aab8391415f3ed0e8e117bffbbdac41f3fbbbbe798ac5074c3393fcb0d7626ba866b59ab57da1790e1ff937195f46518c4d93fd99d65f7a2e3006a41da4e20207881c50e508c60b67f39e90529d16f63eb9e5a7521ee6c0f140b3b4c4f548ff9aaad3af9ffb70fa43b6727072787c969235730a69e7b8d8e3a86abc79a85322eee51b473e8be469d0b49dd8fcb9a5da75d46e1027996e10b16119412db8e5c00daaaf86fb627cd7f0a2f13887dfd381f1a095896188f5ad2273da5c9d6615486f676e7c8ddd7cbb254c6b542fda6b90bfa0e1abb088b5d553202e7b26e82d5bfa929877895bd177b0cf114971ee0c6c2d5089834dafb3f3001023e579062b8a2ed5953ce3f8c940e469813959ebd2764706bf7ae5b27ed4330401d836222569c702d1dd1e2b73adc8c6ce3d2af9c41617acd60270f6d402447d7132866c76df3644f9502da4f16e4a433f8d3222142983b99a7234a4448ae40f125306a3b69a1f7f0b08807a91b9f407c6c1c98a17a8104a9206e7825ceabea560219d433e53c71dd3f71e306cd882c44a99135c9687147560a3e2b70ff12ea295b16fa0ed4f900a28ce7a6de4c53e89fc63bfc083df6b7a72d08c13ff7f8d5ce21e467f0c570eb7d1975f01e160ae4d2e2037c26fd69cf85cc200f5a9174711fcd62d2327388e3a8d70518ae2f5bd082b914a392c2e6c0b55eda418bf821299b6a7d1f694d4da94742e51a9cd426b37e5dfad5f182ed32953e390d70843274ebd45f754b06b622c5cf82e7e1dfcaceab692a645c1f94f0ee11899dd82eb1d7f5ab771de8d0321fb7f1a1e51dfc0ee787a8fd3216ff6afef4705e46b777362236dab19764b6bed8defe27fa8bf9b63dcf8f4ac37c195ed5c41d6a97fa3c178e258278671494c24c797674eecea53ca5b102a95a8068e9a9ff61666c2586e665d5eb1457c8c0ed1eaf5f1ce91d871c67a9f082ec3084dacd1c87d6a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hcd495816d35b846ba875a78615c7345701be71c21268c5559ba1ba7dd78f0effb99e0fe50b873982e67cf5d3f877a06be5f118d11fbbf3f7d7868b0a4f8341c774c6b9e4b26484165f57653f74206cd51d914786ed2117303914a66ab1702a1f97245cdb2b3c1f89330712d1a29524982d67cec0dcb0b57d0e82cb9c5a1b9de83b939b5b472a44af40d162337ca26a8bfc08931191757f454fa50b4e8335ccd83fea24bbac2ab37b4183f87ee846aae76703d1517d4faaed6be4315daa5de50bcccda4f3039002ba57c83a251926986efb2a5b8cc50c1553845c3047bbee7077412efbed47492a77c2ccef6867afcdcc1be852aedab07113ea68631416841be5eae3772a1815784d7eed50fa5122a005d750c4a103cf82e2e9b4b8c730cde7a1053713e88a4ceabc3b3604ae58ff34e0b8da3aea07f429e75bda3e44f8ee0e6050e624eec3e0ab722fd7de3a546dcfc02d66e5832fa1e140a468eb5792d55daf8ae9a9c4adc7f5fda693942a036dfbb9642b8c9c38f5cb3ccceb0081738162f9aede581972c966266afad7d6d6183969f6db430d325fa73221c9bc355d806598b82237b38063a79e4593370a873836665d5ffbf53f46fa37988078d7d15a8c7f4f3dff7139b6a8e27038b0624b6b61cd50199bfaef6ec5b303b7f252600291a7ac5d80585374501b6b603803b0abe35c34a86d5cb6ad216e3256d04b21a9db08627d13beaaad6900ff2662d62541899f1be1250c0d2a00b9405cd896714a30d9d78f0af4de5de64b07e61a4f178a3b59489d62a17992fd162bc823addad640d2cc0e54a2b8ddb5ed1f3c5dc97035648a2efe14c9a7fd66b410b68135b60f387293db78780a7f139b1bb0210da4b338d34bdefa6ddc215b09f4f8a166a3690df17dc78e822b572ea2711e1deed20ff95bdfaae32d9a43dc03a34db05abe9bfd253ee8bc2eed97f9dc1238f92c2616b32001b09e5bf9fe98283f9951aab53923598a8ff620afe6fcc2f7f832a7413cfea579e834b166546a62581f4d45780c51aeaf2c6aa09af57094347bc87ef3f3d86213cb53bcea5350997d68eb25e022949fc7cc4e0eea1c384d9749416d5a13dd5c26dc5b30791a1d8cd04329c43f9b5a58b6259d610b66a4edaabc8cd88a349c9074a0e6316da4fae08f7dcb4b14d8e2de417257adb495692561c3e7bdebb7c6102b68c2215ba9bf3a1b595d809f1e79279cbbb5d0282c5fc9c66bd1c2d81f1fa6f0b21933581cf9636fd6bd99c6dddf93763de046725548de733b8c176067e703e4e2da512e9f0f2765d3f0a62244846d690444f376e51821a522468c84d8486eb3289cc48636da781bf35f777a5eaf3751f5fa719a98df43b20f24f200b5c1d99ad2ec3c2fbebaf7e934f63cb09e06aa864644e0fad48324c400cfb42210917d66fd21ab3675d45079d3681cae31f3651dd89de8d8c4a5fb135067df4135b68f5f7f6d7be4941e1321e35132a902a15ba63b19cdce773ff9bcc6487ddade737cd2f8e931a54eb6d5ab7c843062731e6b883e5ed95e8470b78f436f92cc0ebae4a50c9d80b50eafa8ce17066722d68d6f49768c371840f10b9a8a8ae8ac4329f73f34be52717a99f237f96e897db99d3360f48c5908bb373499cf1fa9c6a0969567be59a2eb7f5f0b9a9d1ab66c4b5460979564f547d217f436739e640633b0e281aa1b9d9ebf0e754c58cfa781c69b22f24a3d352437377c3b49d721c4e88d1806f9776025a902db04ed6b12686c932b337c15fb64ba211b595819d10fa6d9b03d3e76411da7d832ee2f2d18a89f3b6eb4b5184fdfef0552a3428165d3b3428cee890ad39ee1ea44d1de3e5953ae94ad5d6849a4e5a429b79f9c976ea38fc8e0c6721253f50a813e8da8630819989b3327b1278366515333adb2803b6087f779770c780c0a512bbf3a36f624ef21f1f6459e1329b61b93826491ca6512693eb28fa9c90c0c314b05c7194a59c332f884d85055abc9baa66c567bb8531d1f658cb13e5bde252088b3f1a53f2f5a6f305e06f6192bf7ce6750d7a76597626d7a04ef73c9de9061a401a692308f0971db6af69c94605970e7abac1b9dfa62ab6b10829a4a8bd5a1c8678c5dd81fe2acf0fce02ebc0689696ea5e0474214f600015ae9bbb5c1e102e1b3a5e05d750cd0e58564c4d2701f15df3b1f1504bd13227f6f10ae519216af9ceebdff9739cee5dc4ae1c1d5a9a025355b6cbe2b46a7e39ffd71b9bee94bc5ec26dc3b4283d0678e10ff52cb9fa3bfad7bffbd2caf3adde2cc05f5f724f258b17fd637e795d949a93842ca3d476b1fd541bbe9fd6b253913c39d4409de6b2fef4cb15fdc25d573710fa8b61e66365261db802ae179de01c51239489787af95516e1e5745756bb9d421227ff4ec0542d3725f3dcd94ae7cd2d93b13b4f32763cb156890c7de2393ccd19c419e9d65278b0c031f819396442455831a56878495f3be611d5fe54187929824d130fe178c431db7ae2d37ac16c1ad16719e156b0575f92d0f5a007a0ee84cb8f524b9d9da4e2f27e77b180cf9a3b9153ceef4d4a6cf8cd938f6aa4461ce01683f51edc47c36d673505ef1786f2450e6c41a1de9f2692ac281538c3fe32d97f31225554cb273acd46d34782c08364e2cb2dbbc5d52f7715b40f6ee0f3ab80a97240b1f6b6e25b6d6a6527503f9aa219306a94b440f021e06440c834d6efce8c45980550ceb9d8041fb9cfcffafb372456c4264dfb204154187a53f3f99153f6e34ca0922b6681dfe6727057085e4ca1a8cbe10389db87009996aa5a6a730363baca49d02be0bf48936267101c4af498549a4fd41e10a91786d85bee7fa85d2df608fe40e4a2affe80f9bc837e2a96399c9773edf88348827fd086a37040edea2809d3719fcd50f727945391d1116099dc3de0e11f77ad6f052e7eaab6b521f77368db1e220576ce4811dd7d919a20022257f240ea7922d606bf8b5983f85dcf7c159789547e775218c0f2a66e60115f8bc3718dc262dbc37a871365095e6fc83e2f7b1a83aa962cb8d3ca002139bc524dee6009211ea14fad4a687d18ee8e77ec3c8a15caefef7e513a3d4b32dec9d7488e1f81e737fbe0eab8c512dcd2eb8cfe756242d242ae9b8a53491b10766e394d019fa40589c1b38f08b59645fef8f5a25ff01a1d40d5d88da9716d0d9c5666093afbee088e379e10f86a3283b19a86b0b8cdcf8d6749e16629f46860e7ca0aaddad309085741978a800de076844268eecf675d3b1e54773561e31567816a7a64490f124f70b3e1969b2f70ac3dc3dcaf13329171d590542a31813680bde2ee2a513c88b7bee9bcfe5f273b8acc9c21ff854e4faae0fd6b33f653da74e9b2d52308e1c0a5fe2eda9e18cd080ec67192b13adeec886dbfaf7aabb7222e1f679f967bd8b78caa2c2537aaea49b522fd6ea2aa8a45af54764af6cd367edc6a961398f5f8ea62b71b6b131b81a6a3124dd941c804c69969ef71630842241a425c375b3a9a029eaf8fbbf1bd4a2474763ecbc725835ca4bbb2598ce04c8b11107e60ef6a754a2e2f0b13ae51c9b99926d51122498c17a3c48fd41c1e60be864f0916ebbdd163f368b50604afe3f2b52619696290116a9c15f15eaa68a6392b01bf337e575f8763def617d539dbae78793b697a42dcca26dfe2164cb5f8bbe0f06f197a93c6755ce509f5f772617ab07d6a9391e1044954e3eb0376a3d08828b05a1a79547c13a8507b5983be93d01b534eb94fe54c33e151ba6723b9aafa700b49e4d188a048d616b2f0f23de747d50801af1262b60ef123aaf837455c5f76207f3253c64a87dd318e2bf4c6bcd39dc7e67d8e5184d3459296a3e9931879d3b025c6107e4f728c243995eacc216d469cb448055be8d8523067194840e8aaad1d5ba60827c311b97a5b19cb5de6b0bb70efae3066462eafe444c31759a815b2421c4e3c0528ae1bb35fb4c636848022e0bf3ad07a1e92f50ae3bd073a7794bc95435c4703d963d2ee0a80a059529dcbb55734372be4af0d8a89cfe86f65016e357874bc47224a9ad595c7a387ac51e77a512bcf7ba65092693e0abaf05fb53e4f31022725ab8853371ffe8e94fd8e66772e9ef6cd9dbff867ad666dd1f30b7cbde8ea8c4f7b144b6690ce29e645bb676c851bf75e95d1615cc8a08e5af45bf3666496ad7c0786a92b8d2fd64689503fbc1301a681948806744aed5dd3524424b7a6f5dd0b380b72307637a0ec85c19ba3fba8fab128d4ebe29f58d452d4365d8a21447dfa5af74371b49d499de5e972b7548af32b6f1b7d1312ba8f3960f611e9834bc3be8f6117d1d0fcbe2cbdd81909352cacac1ced234900dd1e85b77c0d65ce50152b74a31ca9f2e62a437c062d6889c54a4606cc0e4bd8f42274affef21ef0cde185a1531cc273fbd0eb064dc5cd0ac8f3b6941b29896ec0c8a729f9919033dc6f9363905ec325fc2927c63b9d234d79fd5be1b547ae2f477a4c8aa0d3312231b54ba6ce0b6348e44299bb79698ac565ce354ef4b01a7a0d820bdecd8f77c7f727aa29abc05c689b4932ddde6686c5653b72433215a0a98f9e79cb25d5bcbfebd2bb254202508e80483597afbf6acb1d5679867ebfc361600d52ac48bd352e585948404cea23dd64b2e0f12f6ec0466bacbf626f5844e15c05df7cab1b919a4709aac2e60f3df0cc011266fc05f6e6e10fea13ccb9a3acb48abbf15dd2bc25dc5486875e215c847cf28b7b2fb689c769461728ed88948e2bf423c144969657b28b721ed347a63e65eb16f26e475aa131110e8366eb1d4478ad4a7c854957e57aab1b5fa0302246422f1cc8fa3d9fb172b7676b5ccc6d81529550daeca57f7d6eedefc6cf26cc58de462780ccc4cb6802a53ca6df5dbbd5f7b9497f03b0bc7c8ac7fde029cc9d90a00b44b8f6b252f14085af920091093847d635d8eed56d408a77672c185f4414b2ef92b7b1acfca2f1b76952442c643d45bdfca5da52010b2cc676c7d76949451181922894f612a8811013eeed0ce6e9705a653794feb8bda67a0828993e1df90f2047296c80c1cccb277d0ef0c29e64ff2c45ab48c2259d667d95cca189757285c56ce37ef7f5c2e6302e47d2ed61667186e727e62b69ebed6ed8d5f0ab9e121628f55d63603aed20e0298da50b46bcf70a5c53dc0c6c921c9bb713e444da4ea9d24f1c208b899917652d74f57a46990d470d71f2a9c79fc79bad64babea06517faf7ddf7a61c41cab8765ffe2cdfc3f072819a461e8f0e631782ebd184f15992f15f6a28df8a5a71778ca485c11062a212a679cbaac8cacc52108cf33f939603b8540d29d45fd3996ae295ee0b18802afdfc3c173928f1168adebe814cad8af0209cf7e4dd6634c607b332de74ba3c9b02fe755982a3cb781bd1894ddd2b7e04e74b2f6111b01b9f93d7d3520ff83b5d34c2f2241d615269641eafa14b363a909d643b5f1e86ba00899113324b5f6dfb6fabc87b71e0ae0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1bd7e2fe5721362800d4a44b4fdcc5851d8e89dbc714b5f691c8c1bc68157374b4b83169fa966505e4c3d5df8da2efb2336618703e49eabab8622b568d84bb48ff8c28bc7736f112f92c6b4cca08688312e22562218a8c0a8aaae7c37ca38c1334ca0c55f2d0d206e884078531e0ba609966285cc4fde2092dc97bb7509b6d50d855c4debb610bce494f86c6e8bc202d56dda7a331a3947d624ba52a2fa2b6ec6c73a4df61cbeb847901ed774f4217d4cf8bde55ae5710fa0b2212f5e0d3cca75692ccd92a919d803fb3619161ed57e63aa5d4a6016d46d15eb99f24a934226a028482ab09fc64d3de63a750735459004e94baff1b12d18838153ebb30fff7734258e5b5df5f9cb0362fb6b75bfc39ea82838ade5fd4baf120a16e297556fb38cdc9083e04924683cbeabe0209094307518b4ba6d202a8c6fbcd987e81555c8bec59cd0b53e4dae5951d15e98d98687794941b68b40ac6db3e56b0801f743ec1f7d887039128b7417bd248cb5ec9f213a6b69892aa180ea0d66099ff1cf4744f329d2e27e4adf60ecfbffd5d80de21a82085c03ecf740d0eea02b885cf119ab3e0169f1c4ef78090f856e97959a1fb7f91a0eaeee4fbb4481bd0b4f6a958cbf89c67f411365a9b242e0c470985f69c1582d4850ba4913dcae88d65b57e37fce0f138c255251a838fdcd91c4573191caa07e4aa73f4ecdf54be998e92567056459f9f2e1e29880873cd6840482816e3c853db7391c608ca0a767c90580775d7c2ad4edfc927b4de925f8263828fae962725cf7f4bae9265e71752c27408c16ebcb90950995d5a33d4612699172009be64d5c9c8dc246bb7f65f1100bb8e5e94f7a8c897878a4be160ea31dbe1ce988e4b318ac440aaaddc9ab406a1b4dd41f6e235d0c16c01a39e385876f5fc3db453d5c31feda61ca0946737bb3a0f924ad4e63b6d640f24d8e10bad8ea19398f76b79b99573193065a6841c1b41f4f85b8eec7463a3db6971c33cf034b7f7313f1e30572b6eb989c7f38dca6a9b333e457eab2e81f2e5e3d7a9681e7a09f6203658d58d40dc532b7cf4ff4a0a760fd54956e7b50dc3ce652ea384f0cd371191ad2d1484fa1cca53edf184806c525afc9ef1d719ded2a6ba618ef6fb8863c36b3efee4703b493c451767b2797c810327cf26ec4660748e3ca43a4d6ae27ecba6f5fda139bd5e3a63ee3d7f03fc8be85b62ece96173efb60bd7cf08bf5ba36eb13d854befc979812ac88bc56d719cb917e75b27e89e41d4c02c24b637577e2e078d049fd8b06305dfdad202b95fd8ea6ef29209ff9f3ea41b639a89e5c82766e6195a0670dfb175e3e48cb55f23f11d6e443ae86ed77a2580c93ef98dbcd63fa1cc6852e9b7d900141fcabd89ca178ea3fb8dbc6f1d0b1996da74b830c0d96fafe940e2a972e1c97204319715798b45b1975fce0411506aea27824ac75d59462a6d4fca44e996be1bd1d44cf24cd42d8279659397dae506089f28456dea117dde101cf373f4314a0fc4d8b6e3c6e6b90ef16a6b501ad3b6747825d454f8c858ddc74a93da33de6fdd52b53be3807125028e2049ea167b4827086b92f6855320de6efde5f150758f2b72513ddbfdcc577ea240c865236072c0031e63c022d987105bfe3da65ae7a726d8fc18c0bb4d77d7b24a408b831f6b23c5d1a79c99f57b8a1c7d0af05950bf234b7df1edfcc840f9fdc34ff7d9f7e28caf8481c8cab7f6a88cda5a445a23e483f1d0d63a9d3b3e7ac3346c9e79cfe080ef850769489e0f2a96dbd7a70c35e710e8dd9bef831113d4aa0292c651e36fcd7f00e33ca5e40e3c5018b4ebe7eb2e3d5657f54db66d7275c90f41921f36a0271207b50b04b05c1a25398a2ef2c90c1bbf4bc4324378d6c09d8d2fb941125f0702cd4a9f5c457df52abad9d6a7754f2ab78133012afa48582a855517b3fd28db60b462a5b7daca41ef29a38f2d9714133e7a0c04bc0d609048a7134e016fa15a3486a59d0da93e7be89fa58cbeeee4774b81dd5b6664aaace68b7582f6cedc8e7e5a398b2b641ef77ab1a0b923c7ebf442418ff5c5451419f4cdca230fa38dccd69f46abf71d1f17f3e4856e226a45d002f7b64679eeed9da204833889ab7ec02e3114c2f593c06ac46949634152c36e23988343e493ef941055a33b818125721f9ea3c9fd2e4770f8c7ff75df24e108b527be6c23b04dc8b77dfb9fb71b68f1d5ddf1ec1cfeedf4c6e8e110119c71787ced8bf483ec46272517792404af23d263282aaeb4a031292b701a36ae5b5638c9b96b1277e99ba77322507a009e8cd723f1b079f8c29660ed5557541a5975682d1f17dbe32d8202ebdcac6e67eb9276715bcc400dbda5adc922730abd91cd0ee2cd649d975781aded237110c9681edb983bb0d9479b3386f271ffc18f28c7122f9cd0f002a2ab96f080c8ee0c225ec4ad7b5fb9ae2ee9460a42c328cec3bc1d28e1d6955efe9b7a559a11af9c9f73eb1a5edb8fb61812b4a48d82c117622f9174031e0c7b99ec5fb96dcf7020b6767fc81803fa39e1b444e8e2e4dbe65ee1e7622791b7878766260b2c3bfa0762425a89edc08c164c27b5b52b8b141997f7de1b6d242596be8de38886fdf095dffe3309fa168d8b57a098ff19eae100445dbe1ac8525e6fce824fe97dfe988e432f008591f7e1b8d788b00ce54f966aa4663e4cceec3e9d55a4620c84868b81321f5d5a37770f8c11d980f4c6070ba5d1759ddc84ac963f5af834a05c627474a680046810e6534d3cef934ee8c1f175a1a9a78f87e79ccd019485ec514c7f201949374ccc7099227f0998a09ac3a2216723516578dbd47ffb0ca774d6b4c7a4174504354f410d2af3ded10ba40a0e5aeb0dda5330e8a3dbf72fc4847a8fc99815230f01006bd920bca076e90fa7b3852c631162e0e619bb21c4d98b60b944b85d695ec6e0f71b7e7d2f54f5489ef5fde55c12bce351f387f2c8ce57da26e3d4bb87380760b4142f09ed19fbdd1b62bd429d215375a162e29eec3e7d3e99223874fb5ea7837ccafefae5f2b8c2ef7785a4c86c3bfcd33a7a62e3716e984f23551f8924031f8c1b0dd4da3fcb79f7db772ef77acd1d7418cb95420b64ecee5b21dd7016fa1f8ac12f463742e111a9f7e64fc958eb90c347b426eb9b2271a02c4ed049a221e8f9dfe3028f754c4c0664889f01973cf93c9ec394ce66168ce92985178f682a312c49eb44fc7b5ef1614e2575c397ddbecc6ddf3adca913b753f90778938103c8ad8ef7a0ebb97dd0739781b192f36bc331b31249f5aefef8370d9c92af06ced6c8cdff76427ef386fb68aab137ec657112d994b11ebdb55432fddd1672b2bcc6a9098d9c531c442daa53f3d52151c06e2a1ff2b9f0b9db226c54e2e56f0b2250fb217d70975b13edd95473bf5d5c4dc7abb03fffd60e20f5cc515ade236de01f713793fbf891a0336e20b6f8187a8f70525d5c251afcf156709708d31bbad3355853142b6b5f160f868a23b6f76694e90e62b47a22f1470dbf26caada17bf5747b6da81175aa87cea85a036ce1a1f8c0c1c6a95df2b113f358ce025fd61e2bf6dfebfce5e16030a32d4d82c182448627aaecc81841afdaff8b53f3da8be7eb3580236caea0818cd2c163cee08c4980ba3cb992c22dd2a81b54d455bfc9cea5c35f173795590788503f0d955fd50e9f91ab1a4e465d1d0bf276bc849b9763035e89efcd668b7da168dbf1c58fa8024496b7dfd0b9e1b5d3b49dfd1c21d6ee4d786041a28fe382062b524cd6d219f1e17d854df63116b0117e3af4b28123e1f5f2d8836517fbede7afb33630c0831daa6bcdf544521d9f73a4273019c27aa7ef162886eba6405f07c1b5d0b279d340e47483dfdf3262a9b95f6dd69bce19c94f5e642392e47c72356529bc710583df98f9da6cfa43df2a0e8201474f2e5d45adb95cff32422b94cd90db59b0e8c82db1c9318be6a9de2c19045c54e06576412e72d1972250d8c1dd6bc77c243bc62249f6523c8db4203999b9faaf939eba932fa1f76583d5c46bef147469dccd5f04f5658b1f73e6f72a592344cb259e3ed77268eb4c430f039a72d9d77fb2b685b69226de5a83a867c8de7b10f7c687cb33e69864a955c9f7fc54520969898111cf9c46f762191e8eee008937f6bfc1868863bcb184f2c56901bf6fbecb88a3a5fe24cec2661ef2136729d54c4eff1e8068da01562fdcb03026e653af6fd16de95cd10e1ffdff043788bd9163097747683318286e3b48e03c1aa1237f9dd306342ab103efa73343db4cff6165c6f1f79673ab1782730fae91ee2a28067c935c3e145de223f585822f0854fcc33d7a6e41aca325eb208768994d136ece67849e81a38d07304229c2a3e4760f94fe722e4d2956ac18a9e54f1d77956defdadf56cd83514f645823279d12c87281a78fa4eea126b5be1470f074ae345e716ef2edba500959c8a986dbdc02737e945219df0537d49f3d61ff023bf59b11ed0618237920f0fcbc9dfc333291f0dd493c806a09894c78159a79216cdb1eac3998ce75d31f268d6bc71db8e2e831fb5e95c174ac45fe7797b7b818aafea6e88364bcaef8d90a2af861e874ce57a152f0fada446db8555f682d7d80fbae44baece57c9beaeef9358321373e7afb4fa576acb39039fd55cfa1ecbf2dbd7de5bd745abb8168480cf3c13b3a4875d395e8d93dd8feb3c61b5fd90812cd25b5b2b65c22b53a0c7810a903cea77ab4de9d3bb788f06d80f40672e48549d72cd76574efd3db88768e33332517fde6b61ad6dc7da1d7932ce04c517765585eb3acb1399e9bae8417ee667b2768c8a78e366740c05a47c843bff014111057c444fb32c176bc7493b28823e019f914aeb23033129509f015d03b0cabcbc04b3a620675f2ced711d22934a56f7dc196052d60965a1250734779014c0892df56ce62e0f8071e68556bd49c9a22c07d21aef8beaf1103041d6f2b391dd2d34d86452d187e02909e1d375f7fdccc60e2cc53d1402eebcf00549eabf06df79cce199b35b2d37426b03836919c7910dbf533adf2ec2d75aef7a151b8f6ecdde12bd11c970c94a6b018bc6fbaeaa23c3ba007f27c4b1cd35fff9c02e37900b6bacf4b588fa7dfbf8f13573e8efaac2c3f1fba47edca3647c3671f46974e54b8f78de2fae8a3bdf33b702d06d9fe65b02637d05d4c12678f5b46e0e25200fc48798237a344f1b04f4bd69b0885fdad8e7f82d71119aed4f857aa0d49b3a4240b78482457d2195ef1bf8d59e069e009329aae096c0fa9bfde83b240853b419657e45084862c1a95064444f3f5c6e25dd8fb30ebe6f91a4fb5eee332fd61e8e10b790a23db28b622b24871544176d18534248ec143bc14ae11c6dbab6c7b12ba0c66d615c71d33f9ffcf1c90b954d3d48c09dd94bf0930708c29eb7fe59ec6cef712eecd58fb113925db96961a56e811b8cda25bfaa5c59c6d83ed086130a0e8610225e2ca9e04a7f92b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc5cea3000c07bf226fbac0eb0af02c9ccea3b8a844113bd4a6b80ff08a023ea3272438abfbfd085af36f482f02581a4f0c4fc4672c57b51f534020ae543c0faf338d2c09551c2544128be50fe9905a4d1026cbec8c91362b3746baee67dc58650370228ce942e1240a99b57b3bf5c77ff8a44b27058e3b972762cb1f2ff699d6853712de1a653a0b2e7b313a89fe0c9237f110716e9e73a03c590481df39a803a372d2ea0508f50c2361852adc6a788d680d2d9f36c848afea5b1b58785845859126fca92635c570e6666298d04c927635e1009af492623b486141e46d9f7b1b367469c2361a64e6403ea94f603357046c19811c4ae9b3e0cb3323e80fd658a9a95528c5a59ab9c6ef807984ad95ce573cfccd22850bf6349a299bc37d0c07804a45b4f31a371fd72d4206fa3e5ba62e8d5c4cb3069557afed3235b6fbab62c8017d322dbb4e52b9fc2b4358235ec367cc6c78f479f8cb653e3f624a9e3f812950a8d4e7360aa5d1c62320abc363fbcd5d3b40b0e36d758c21e9c201833fdc219c0a336315e4051647005ac626eaf95023f1b49f03b67d0bb5f6c0bbbf3c984a3405a9578cd1e12749a66da641a7bed8fb9c33f0dbf862246380ae555f353e820a11fd7b0cc931e57d6f7d39683fa4c9f54141888ffea8b76e2e5bd83437de5e8dca6420639fc2d7c0ed0ab655379c4c6f2030ea78ab2c911d96f0f43afcd9e5b6db684bb8ab41255b3a7ff392f0253845c5a9a51393bb90fe889216156f602ece0047f3dffa4ac213d0eca55f962bf69cbce158820ddc48bff29574b2c3d1ddb6ec4fcf23db55492491a02d31a9f1f99eda10ebf5dee6c8017d6a60404be61e1648feb7b650bf57b745e2c9aec8b8f05a34f23d91aae310809b5c0348fc613b20d2b4f39c7a88c059df14be487456b0ee8b71d5f77bae1f0368b992a83fd0e794bfb8edd994a32498241a79ca4200ff7b0e4a3d03510c8563d46f0e4f07905bbb46efd8ec8f3a95463d4e12d6063cf4b1d84f8c35e85c9f1d55f80c2f16d2daf3752308ab76e0c735b6230b807b02d8da4b86d74863317519092f4f39cbe71f0a1a5f40add8b3de48625a9f8ded3f1b9d6c97eecf33965b69b66c4dca8b091ea6f06e9abb0b5a0d0fd47de1ce6062a1832bf2f016437aedd43ad234a541e5d1037d67ca0d7eaa3fdd00d3bf9c229ac3ff512f70af95137aacb5fe92a1df5e7e81fc4d0597bb1a7a47f7df11a3c277f6cebfc691f1594ce958cb4aac23a2c17997d6a9f9712b185a5fdb7150dba1e3d41fea59ef3f67b55c6203c9517415ddce9131a2212215d18aeb4dd5d2b1ed6db30c3712bb5313cd8d2d3be4c019179ea360cf13132139cb5cd528217d2926dcaec030a284b1cf37acb7b53eb2e47a60934e2717065f34f660004c049a6ece601a958dafc4fd17f18466e4613aa88136eacafd48fec87687f5de9c27072606f71af5a31598437295d11a8dd2a1bfcd9491dd9eb06a25a6c5bb50cffd00d169011ec06445bb2456f7edaed339d47ac3b3b0c4e84a179e5731878d333c69dcc58e741e85af64f3be1743250de90c7cd6fbdb8e1cbe1bd58431f2cfbefe89eb551529891ce59cfdf10bd7725dcb3d3ec21d06ae308ded13021bd9ef174379734be24bd8a4b370fe2bb006a23a7f3c566e400c1ab8c0c10d0c0f2e1752407b77d04458b4cd5e22d9cdd167480b2cf97777ea6be1526e82e76d5756255281518a33220afc2a7990ef2d67db03487908adc699b1ee9310beff65f7ab667c2bf6f156cce02d57d9dadafc64e14ec13c69bc14df6be7f76601b60f092e71d1f3af0d5d5c39c55e50f049a64be3288aed2b8838ad0c46b09104397be8f3eff15c5737c4d6eb80cff30d35652e56d67b2818d03f71ebb26f3745cd67feb121bf7acd8228dfb7c738ea18a2ce9a09ac5025bd73435a2664eb7f72915bd5fb775c95cd61251d6bce4e5a3320d743947ae5557f393b8f1d9e46f3f0c8e6128049b6fec09d1e6ac7913f4991ac32aeacfc297ab6ddc05a60821d2e9f6137915788b9b78a891cf8a1a2a813eb8d094d93e84627e06d76d2f4ebaf9faa17b4357f1a853c4dbebd1a3685c14403774c56d8b3ace193768d9adf7c9355da653e560dde701fb6021b164747f24d9afa1e8ddb815c23225c1b5bd5f9621ad51df191ebe2e51481606620a74161d81ec561d1c01de31ee9146bf888a0c9379124577de1fda09cc120c77639b83dccff113985095d660d4c5e4f20bd68b09fdb291ef62da47be2040ce90725839768f304390cea07ff550777a4dac9d6a0370e85df7a87a7af5a0897bc4c7a96a62ef3dbd8bb8e487cb587f96c98c2ca05c11ac506aad87ec6faa5bb210668d514287f88262cc87e0a4cf5d413682a1edd512f4f46bbce31703b4aa879e8f08185a0367d6a3e82d9b8195484218adc7d39baa60f274edb70716dcaaf763487424bb01935060bf5417c4ddf1652fa6204d2fcdb34df28710882714dbf63e6bf4ecf1bc5f4e3f1311481786def97615be111281a9034e9493445746de5fafdce307cfa996a5a33594d3f454bad1d58f0df8880d2d1f9a21549e6df163b7fac2f19dbbd71d8ed7b5bc964b6cb5c567f4d483913bf0479ba833a04cc9402fa29b3f88ec521da02c7ef584b2a90e3b95838184c8d085299db0d3273a939fecd008bc36102cc66acdc311d2af745624e01a16137572f5b772d6a002b7dc7285f55be62f7e75bd9c881a9696bde8d774fe936f89f11cafd4564872df0b1f16c11c2e3df7c662bee71c91f4c1ff513a6091698adba1c8d13cb55c51f533b9d91d7d796e8c2aba70a3bd1d64422252ea7f1cbdf437918edfda27b951c46ba80f1e25c792c43832fce5d592c7f1ab5b54da8755f494c46db8b550d434c32621b5e8b6dc5656302ff819e49e59129c60187733ff3cd1178d7f5f874d21a392c9ca5b8539b23ef245b10f354d0604b63792ee702755d52a3b3c96a79216fe4a414c3d442c1446cdd77f06c397b05d86dc9a3adbfc0c60ad4a74595154f82d6504b9d71f439a2f57b36e2950081c46ef16e7610411cf4afcbfc9c4a6cf890b31225081fdd5f7746c6e4f6c497de7f4cf5e0102721b80e71765bdd3da40c8727fe01f6318f0e02700ee88ce50d89332628a94e24721245083e0f0cdece1a23e8f9a5cbee79b12881269dc41204e0cfbe0d718da67808ac4d342a45613de4d91039da0f6dc6564c6e34c8cdfee58cfbb96ca8ca036533f2a8fdc3f3d45c66c3dae56cf3bbe57bce29bfcf0a4fb9e953a9b90849c769e9ef182e8c86e62cee30bfd34c08b3d73bf883600c3ca5422141257bdbfeb641a73927700c7566e893703065e02c4c7230c48f133cc7c7f706c45fd49d20d3ca0227b69441a7e9f8d01b6b951ab202de3022ce4e75336099219f882608d3e5ff04b112d3a043aaface2038b55390aa14aa477cdfeb47feaffb555f649687b761692b80ca29b98027729c819d804339dd9c57277954a16c32fbceb95c73f8547b0a01b9f6024e2d3398cca4de59dc1588012e0e086b72085033dcadf3eeddfc7caa2c62d63eca01507ba63110227ff63258a81b6a52fd6cda9009ee0cd46cbf7eb4a5400455f55cd821a8dfddc854e151e85b2cb5cbabf215d80c1d7122e1b0f21fe74cc9f4f760d7e0e383db63cb7a21d71d81d41929824f3e494b1c44c18cc160e23d11d96d1c2e06ba19b0d9bd746a11699cade1fc8c13bae0614c76e096b7d2e632b1c6b850c28153a4dc865776dbf6f86472791660b2a108775a62ba36ccc75108e432b95ce60d4288b677bb53f44d529f9220e7f71fb1403950bb3e90bbe255b7731b59456687fd28cf1d424ccad8a38ffe07ffba9a942a45cec34e9562b7ece4694aeef82bfce82fdf0b2e2fae1e64faa28d313b4e8744f4c36429513fc8b8bd52aa8bd62e1bb780a37560f2190a0025baa25aeb4647c5c2592de04bce685ef8925ea97e28dbdf133991945c1f5a7bc400e0a353503bc05d52897727662a6d86365854226a73737d1dc62fdcb7459afa2869c40c5dbcb91cb92d6a7007034b081952cbf7fc7707b12e3926728edfb1c0ff7ed333aa0917d58fa930faba27ecf0b066868258a1701bc9e9fb73bf29f0cdc1282695450ceb3f8706f860fd9c58b426bdeca82189dc31bc53396a5087ddf88e6d2085915cd91a49d476cee9530293f705faef9771de67f196c160f628ab465ef7b01ec944f36638379eb1ad45ffe86b586a0eb92b760dce614da81b7037310795d9a3b62787faf2cea67a06261a6c73615640fb8386c280f5ac798d30a45a1002d17459fb7cfef22e81cd853bb2bff624a92e8fdd10a40e7e0db8a1bec5ecb16babc9fa9aa2c6d56f672441936576c6852792b16ca0abbbc54eeda07d7273a8f3fdb75888632a9e336df1ea8e53b920cd5d6a616a9226a670c5825cb9283370c82f37283452590407899f2ff37041a1e0c8ddfb598f26093d095576e61b26d4969b1520e73ea81e2be9eec1c590977476723322ecb42a9f10c374c07a35e50bec93ad44b9de0f9afa78a6b2a9f1569d47d9e36a443c455fadb1e1bad35b6826a4e788af584fd2f287f0b7d7739cdfbe1385298cd58f482efc3ab2ad897cd411383a3b097131acbf3fd6ec95b9019212473fd31bfe52566b12518d6e2dca2596a397475900ff20f5f40ca8383596a45d7f9504494577a475edf696d212518bee822a3992fd7dbe7526b2309e24ed39d518c8e856f0869fcd222e65d4188870825f6516836312330c5604f34b57fc3a2b31846d35da21c65593057f9b89605a327c84be14da3ef2b475f2830f897b47b1d22fe1ae3afbfe8dd9debc2e73681953f681421bf758e4d05ea171a694281e6aa6947db7af097b3715753da3f308e0802292ba0e55b93bfe9f7c365be287c0dc912c131aa32e2cddd4f6170baf9b3465195091c1de9a01041c0f6ca00b7b5c80cb6b43afa7ada617f1ff4d16f9b6eb987a0985cdc9281301c91be3323f6a44614fad8bcf110cedf59ba5c604017a5717a319e253d6110a8cc3ca31e9916058758e626e1a72d9aeac3fb9ea5937c7d70e59d5dead81bc09056ec5a2b0419820f4c228c87f1aac152b1b4607b8dcad8848a566cab2d9c7b7b4bcfd7185d12e88b8dec75c292abb92c5c1854a06ad0d1873ea329e2a9b095afc5c233beb7bfe8d542a7f94f6e225636cc528a8a61117fcd19859411e43dfa87cdd288dc2f4cfe3173ac2b9cbe5d02e55f80a38f37e23bfcb855e297ff8ffc8e29d188c6ece87ad6f98ee1ee69cb0f7eeae54fef902f71f7dd5c55729a19d9948a81f26c5927fab78dac17e0bb61fdbb4cd28e490946e468a8a7d54bdc16a8712a75bdb3b305b1cfd6685514bf016ef814f0e90247ce23b0119a9d5a0a2590544372ab558962f7d18f4efbb94f034afadec18af3445b3f1747b3335baf4d11dad84d3ed32710ed6b65a497ba59fa98b87b9506cfb3d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd7be1b9974c90bad3fd15cd9728851525f83109540948ff4e915590572ad7ac90c8463323cee15d9c893de382e73fafb1acbd17f4916b033c147c0ea06f2590b75ec56d2ff747156970293de00b8783ace4a9c54e071c26c8b05f10a027f21dca24cd3c1dacbc776edf3ef9d9b17137292616027a7958d46ab21152266ab1c1b1aa7c2a7a8f2ef62b35b6b8429ea85bb04015a10cec242c35a1f9d1a5903ac961249bf2090c72c060d55e3d1eba08a52d01d97fe27ebf55c8d1c911da2336a91c9bdfc55b86b7dab9cf64892a1cacb8943e0953af2b8e99394c282ad3728350c0984b83e84827fcf635678286bd024f7d9eb81acdd158fc9a8141544f391cb1e03a0ed1b5441a3fedf0d511d5fd570b8c71835a0118e60ba991e5ea2db8fc3c243040c460d4c8aae2cb469bcb7386379b1c717c4caa0e4a8efe6723e9ade4f8f804f80795c41e7b527f0be9047b07f190423e4c3b77f6a03fdcf1a3bc7877389ad6327123d40e18d9c2b78647d20242e17952853c9430f0c73a502c151250bcf962f44cd28a9a84e7038e575fe3e94df76976a706d73c46126505e580dbda7656dad953c780be6428b1712fe64db833878a8080af1b6e2fda8689582f8da16ad34d209c1fdfdcce0b8fa2d3a3eb992127f2df5484fd0f2623f998b146b348fcf3d89797d725e188022072097190112c4d05bbfdaa17ae79fd092d9452db2c38eb1af918e866976813e38a130820e8b6274046b74b174bd4ba63a54b096dce64325c4a7fc0fa3a15a1dfaaf600ae44d1a6b2baaca52ace8cb88b402764314d7ed89f4842fbe3b59c17632facec48eff88f38122aec1e02ad66b507ab31a36f9e4edfdd1a7f9f39a5ebd3d59da4ee96327ee93308df4fe559b95c1b2387e332b17d9e0c38ae35b6098f0a74c01ff14efc41dd732c321e639d3a237a619fb8e959aaca0faff63b36c6eb74e1c2351b1d5cfcdde3cba08f44556b6b70748b2224c553cda744241b69d9bcf04e1ddb157a5d80e8d0a08e732884445c7e0a331358f0b59d9db55e620ecd372aa7c70c5b4c50c8490be0fc01f7fcebb5e8ff5c81c79585bec56ab3e23e3121ed6435c372e55382a94c490e76ff4bb71e3ac54b8c63d23bc03c8aa9c72fcbb2fef45fb1867f53cb63e1d868e2166ab6e2274be56e2ca93328429b7db5dc1a8237b77cd9be197c56cddf05df467a4f82a53e80fe70e8c797845cf5ebbd334d7604969b6efd18d7f086c90b616fee8a56040e3edeaea13a24a9b33138f87fe956d70d2f38d2c2b57de54c1b54368544ca338b67b4a5fa78a28bcfadb238d3d8f4eb839a594ff5fdcccef5541b395d3ef9a1d9fd594386f2a01bf051f6e62e8afc07c8d6d792775af046029c4fceedfba78f4737d12a5cbf4332fb2e84950a1d639b2e96de6e97be842cf3ded0537c4e3bcabfc2cdae90db387268ff9bab0fbaa5a8dcf34bb11c4ab9cf8f287a2686d6aa4446a55fa74171bd9d96e380de293675454cfeea3134076ede08907559cd7f3cca017938efc4907c8f6af4cf69229350a988fddfd9f438d76791e07c45f1cee2b8e2c91d3d3aaf03488ee79bd448501b851b693f6667ededf948f4ad9c73b7631253a78bbc097844aab93c53dfc9d399c6ccc1d717e35b86e9c4678669d1840a809dafc56ffa2cbd7f9b30e10491dd992968951043a3e9be1fec5ee52c5dc3e07e674bd43508a031b6a699dcb863e3c81735bb2aaa137fa26d200e46e2f5a4cc8efe35870432f671009ad7b25f6a206535739e1aa111b2984fe89d4a2322975fb4e4c5acf4542f566db8acf5f22838831421410b977608be135c205f2aa9cb6148159b9afa0c3843672800243c0eb479aaa51570defd62a3f884ca2208449ab36d03f59a2fd5aaa912e41c4ca1f8d8722087f7e829457c853727a069e046b8c64130726188ac4c32288024f0ba644fc39e582c28ee95a3464352e9426d8b28b92c6e59427d49b3478bf436dfa8acfb53082775699f51e0ed2acd4d944361b45d8628260c319829111f511661e6cc7082dc4b93bb159860f54f52ce8943a3fa858697f37a5ab81f59d4fdd0aad53e3397e8cd9ff15bf3758e28a4c5ae8d0065e303e592619b3a4a54675dccd408b78abec37a9c5f039056fdad3225d42d7f64e0be942f601763acb185908ca0255a457e945e69b7d9661bd69cfc90a530d3e9b84d6f2492f90ccbc7a8718f6c42aafc5a63d0263341108a82c92cc971e28f7ee41a150ef1d734e2098a3b2f02ff31ec4a69ae554d5d36dfa90eb35243170c052b2691f5992abdfab36eae5132bc61723dd04c70f4981aa9db69f04b89fe24079d123442dbaf9829df01ebd91ac33ad215f5d5a8a875a3a7ab3ba9398b7cfa43c0acbf5d47987efe620b2fedd622710a8a01d8ee538513f5c23e78e47094e33458b51d560c9b48c5371c4143cf2640b72264aa3b228da6da09b86b28bad72385673e739ffee99915e47ba14e68041e5bc4bb7745e14c89c4ed2708d88ec3474aa6fe5497fea1de2f07a973970bd14026f8f7e21ee7cccbad197f97e76bc29da1b243fef505f1b93f971487bead8bb4b2bd741ec07dcd58b332e24c5bb9adaa4b344ff7228465e37813ae265f6e38fbb520c76d777f710ab581bedf0edda9b9d4d20cc877c6b074965c4bfeefe184613dee3cf209f68f1780d2a4514fb07f50ae1db52daf4e847017a8d836f4701bffe75a228d85d1986b4b8b1ee6c7cddef257f03801e6d60dff0e51e08da157ad8d9359b00b2309a43d071f1305b61e48690d594b5ee83e3d57d78fd6aee7e893aa8da5c84b9ab31cdf803ce47a999272c5084961e36ffcd1a8d68a16d912f474c3085dd7325fcf7035fb24f919814f76b6b9b348655112699002e330b19f91383d7c86c7f652adf7312d57d757ec84b753a340b5352f01d2e62a064f616455bf9100f2a7ce157669feabd40f23b64bbbbd9b9a0209320f58a40d0be64d909efa8a098613a647a91a3ba7d3d9aeb788103fc401cdf63feffcafaf12451f8519865509b1e210c86ced0a9aa03943ce91fde0ab48d9081c5da4a328b3aae3235eb329a132694722afcb252656e06b6e364f2a067ed35cecbac6b938c0e9161d09642d5bc289861bc91db51f134a56d7333b62c1199f73457c115c30f1f74673fcf26fede618a21956e8d47ce51f6e015396b216f913d5ddb1cecbcaa6496cdeaa817d0e17bc28f559362d4433e31ecfe3d8448e213ae6dc90f12bb5092d892222dd5bfa96d2d7f5bbac97f32e4f0d73b88e60986accbb22944b5f7f080ed0ca22eb8ffe78f59d6da3def9d1a916efde47ec9c60bf8904bf85087ff02ac1e14f12f481f4338ea4b2d7d9b5ca93c0c0a73669b34018a392eb783dc62506e5263b71915830d42a582dab43c6ef153a42d68ea3cd340e641208beb2c8bc801dc8759b09eb122bea57abf7a407157c3019a3414961669941a4e1dd68426d33a056f361e98a4413c6da3e4f8f6575a1fe0fb3c569115cf8a7860fcbe4e094751728d31c1b8249979e17973378501b016e47af3ad8fcca91b5514144ff6d61d152a647a6b1e2eeb02ab425208c8337291d20b6b13f1e876230ee15a738ff46e319e1348c2b5e580c43b28349dc79ed5438d28d7c1063952792ab3dd9a9c37356bb45aca8616c81be3cdc410ee767670ed035ef46c0f265a694b809f0988bf2159d654bb6034bf4913c99c79a2985f0b6bdaf18cfd0fe954f742540b58b5b0ac41232cd890a27008b462e709fae40ea9f8c8ae1d7250791177a682b73275b93dae68a3ca91e791c63ab6ef2dd6d3a32bbda142b771632dd15df4f5ecc35eb9751abee93c39582fa21f1f463108f7deeb1e7974ca4ed0a928ae45897ac1e9a852941b4264193f122e78c861c63f1a187043437d821c678c568f45a0e98ba9155cc3fbd335f06a1135f0e95bcf69ea59add6678496c18aa056c948c5fe4d1232a6ca60d3e00515c7924ed9fe9a1a99135f6cfe84e7fe42f3648d7fc67531b577b074ddc0c9c853ff2927b592a16e51532299c5db3b70a4036b2488c42f1ac4c99123d3f3bf72412e4dc2c79623831045248427c4dd247cc97b3afddad0ff21e85630277a094c86c1c2a2e51a7fd9f92c8616dfe88903f2994dc0226d47905738b7849bdaaca7243e5a76ece3156fdb4aa09f1f0ab0c4fdd7f132d96556c8e35f09dce8daa77dd6f130204b82501475dd14af090dc4e181111ec2b6a496b9f3b7505473924f992b9da60ea74609c0daf961283ce8874ab223e58ff919106c89a199676fcc94c94a8c31e9879eef02de2a08dea9e1cbe3bdda83d97044b4e103f18a990773bda17ed59d3423b80c4b640bc473c62a1e1bb8fd32e1e6c23b07459fa3fd0876c7e68b737eb0173f34c16468275676a16d78f1903b46ea738a61444716f40cfbff7144d8b13708f23830a103750d6a15211a139e219ab7360661f94b096504ad30369d1e0e28864b7aa679f66e9e2db36c20602ea2cc2ca3463a2cb37ff1548e174dee3d5f3703335ce5d41532f7302e8edbc08de36bf9977cf96d6cf4babcf5b511fdb25b26dc622d65fe776f0c6e27b64020d5162ec40534693055b46a9936ec7c75a751706f52317840d374b60a4ba0f575c4474a938944f114101324154924f9c3b1ce825f5ba612c3abde55c0e5ac22b7830438ba6fb9faac3bab60064f2bf9aa7f58af87b816433d62f8d4d406f415c2f81e2a4846939b3f66bab912b839e2fba42ace91723f021b2c21fcba8222a53fd7e103c4ffa3aa9e921ad652a37ffc98fcdb9e365b99f6704223e77e55839c37506df3e14c7f2c9460c1052dad76af4c12dcf650fefdb499a66c051c0adcee714e4901c776ed9ab48ae78e6debca88b1758c9a98a5e7cdb2bd1d65863740fccac5ad90413b720ceba91e2753ba85178027c9d5011ba4ad73d525334275d1d2a71582153a2b60237f3b9f6879b11c8107a467a1052304a053dad10f43d01e92af6ea4798f168f228f7efd6874a56a105a6989eb7164e4e00d25e70d0bf7314e8fe47c2750d022bd867ce2f8233a3ac56da9b231d322c260d63348f81a7d8edb777b0751e2cea26cdbb064288ae9e353234b44f8e598c4aca9eae5c7c43908811210e4ea1c1616aa2063d631f1b85ba61aa64b664fca06f1b31f96a00c2ebc341b6a9926a96bc19741479639231bfc403fe55a420a43eb6d3bb80827b8eed051fbfa12cf339d8b2de1bb5dcf7cc2cb4bcbb72e5f52ff63dfb77cca69389a59a3a106ab808fca43cf50b69b3fb4b19173e0af975c5f398efc0f9466429e896997fbd352577c2b0883408f22f18d0fb54878a8ba36f52b1d7fa240d5533bf89f206360f3e563ccb418580c37f517639f0c5b4f8649fb6788c1555ac0d52b7c8988c72744465b07c0a964bb9d9a9ed8f68badb9eb207d0f7fe8e75baf2277fb98df2f3cc6566790837440f8ef0f99aa2885df8f864d65f9129d30d345;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha530c5da04cd12b5f612aafda7333e7a7fd7e23d664f07892164eeec6a15e25085afe2aa458fdfd6fb16154986612d0fae8750f5ce70107794a0da68f33ad6133004785df8439748dcac41ce1e521b44d4b2a8abf85c61ec4c9464ed507e9d8d5d84c21cbf02aa7b48e5889af1f2c2e7edc7d61fe80c84f23fa3ab63f9e09ae6688abaac34c9a67239af90f35e7e782adaaf0051db30802e77de640917c3da62b04e5b50bec645abdd69247554945e38047f92efc5c54ca23e9d05212d54aba67240b8ba49b7e922922d8f81b5a41da843cb74ba877fbd556a61d8ecc4adb61588a45cdf05546c437a86f8b2b96cb0cccfd8035b408e1ff74078cfc08c55767713bccac4d6370be3e575b0fa896a0d34d40beba4869eca80652bc5573854572d043a5ebd27cf93e41fdae91958a81a662fce130a524170fabd23dcc76329f26aad610ce619a1a6eebec70844fb822725ab79722bcec4983c1638ca6c1474a5f0088cb07ce516232fd077529f4aebfe4db13017c1dff449dbada31415860098741f3d67ff57cc31f87561e2a1109e629c145766b0da17de2749f0ecb7839e30ea0d43efe63845677760371cf0b7494581541f3e24e13677831111caa1928335e7f597cea84e89372b78a5f1de3b86209c4bf5e31186e6638e808ed55f60e73ccf76c24b3ce608b6549f820abc49b6eb5eb4e867077ee3caa3d414dfe377c3a82c550f115867532fcf558b12bf6d622024267e296a4a29b7861c21f589273dc8deea9b84aca5a857a9d5fe6448005a6d789ffd4766b2a697a09625c2b0ddc7fdf66ae368a79a47887567f740b77e71adfce39cb996f8f512b9b66a746029d6d9f4bac0245f472a28bbf51d047ba53e32ff4e5ec3c1752fcfe2c2cabcbb2967700cceabc3632b64f298f9a9455fa4e4eeba3554117e290be7e7555eed9c0ca027f336a4eaac5bd50e2c08f51ace1de5dde89ea3d6fed67ec89627d608e8323d15ab7fe08e386a737bb4fca7c477d06e87a674ab38135ad5235cefd5f4b9746cba7d9e286e4118329e2d3c590ffff4bc37ca01f2a22bc99caf882b8d803f3dfb515b45c868455d08b395550a54afa118fae4c8b51ec437b16a921fe3ff141c17bd55f75764af1abce834c4207c7ed04576a775fb797102eda466c35bb9a2db224f82285d2f6a13fcd0ccd6cce8544abbb14b670eff87636afec77cf578e5e6ef805233e84446dbb182e01ef77abc3d1c65ce212039f274efbf1cc1826d2a5d7b91e6c994289834a22351df50cc878613596d1f2f085fc4aab39da7a57a4899a716e600d725c41c7ad0e38f659dc14d6d8cf0acb0cede3b79c02edcd0f7852f0b10c12bbcd72bc9b51f3c15b2e8711bef8a72900b70dd903c356987b1f0269ce5a777da0bee538c37df527d3221966f46db5b9879ce70d09b1d1438928c898b65b035cb322ff6110b1b77aa980cdf863a7c51faf3441cefb554b5e1acd9983583b41b5ca291fa1669f94ef8061c49c3100b5574a45f12b79b2654e74247fb799274759b43c535c6118f4b52cfd709ad753bf13e271ad2e67bcf9114529c506ae0cf5997ae273a136ca0fcc9ee19ce6cbcf993e37fbdcacdc32a66daf1d631409a8cac83641eeb1ac45af108f824b1b16da7a0cc78edcaa16a4c5f7845e66dae4c79242f681b6cc3686b0357a21acebf968dc338adc38a0c032b485d9a39903a40d2df3c98ff9edd0de4fc6db0d7aa630664cd0b382a58098838727120456e6ed21b7ff01a72f1d308b4507ef8aff08a4408bb576523e8f1a9726ff2d29d5f66041e60e40622f9187d588791f715b8fb6be5ef7ab816d0e0140dc66a5c794183968137e5ebe65f6ed607e170238efc6f9c3822806df532094de0bb78600b040b9ddcf0826afe15545ab440d1dbd7edc90017c655a981df7acdd39e12d5d7643382ae7c288b748ebdc725015f899aef59985f9b76a65b2a71c00178d33dee1ceeb6d7cae6ad496b09c3933a895f19f2b42343db0e27a76b3c97810411d0c96c0e4307cf538d2abb67dfcbfcb46f4611bf2accfd327ac2c0082ecf207cfb9dd4f8b294b42f58078e2bb47c3719683e26ebb96eae30d20dcb6e542f4848fdac1057bed26bf552f9b4095fb618616a0ee5e90a1610ae6f6d1ba695e13e9efeeab52f5b95b5139f5520e2cfc9aa57d3453b294f1593397670d4a85f71b3a54ebf96a5446e98cfcfd2a4e386f5bf5f9218e211b5be2ea3557e04998e845ce4610b53aaab97e89fb4876e5e379a27e8f329e9810d43971379078cb9455e6834d9d4bb1ae8ce259c3b2a8781ed272f4892154c9c745ac88078033bcc202bdc4ef52b267b23068265f1ab2fda3c31b7f29dd3be9d5251e98e5a6583279be3dd24a612d2b40947884a24461f9e4f388cde7a7dff86a2084ebc47e768510cef631e7a665fdbfc7995f3f2611626f692e3021c06b214db2d5c26e8aa8115c9398b13b46070533259658cecd33231cc46bf7ff243b24623336a05a35e66ab0d1f917d9c9ee37bc5e8bd785c87d88b24873e208b4196d4dd0c6f55173f01714c08c8a52101a1a8b48e1c6500e7620b4e7c68ac4c89e315f5e9fabd448667cfe47ce33962c183966eedff890018656123c4c5bd82aa498e4aa1ac6707363dca04f085bb93222aedad81a9ba1a152e601a1ed96c8432f96ad6180bf96d9b9fb81728e9fc92d6e86b20ba7ead41dc6984f2f97441e80dd01444b042b2e2375edf051c890e752e63591c6c632cb3ba87f9c57c2e55f77205aaffac03350c5dc9ba36e3cd9de108f2fd4eaa071538ed25347b04112b9b9ca7101a28e072f2edac9ed968fcb9eba56a0c9f97b7285b687190d317bc68abcb5c6c947edb67855b8356468bc25a98c8d744e389cb79ffb00b50740b9d8d03177a2c9e0b05139f793c80fcf6e125f8679caa6c699503420a267a81b10466da4a73a3c6d2656f808df58486559c8fac178ebbfac4442cd21938fc9ae3848b68743804b33a7db4e37b110200ec688345a25b5c682bdda49f9258ad46f61d29f7d6f758f552fd016f9acdf647976e93ee565d5e8f046688c766d34f1e2466f0a0b4a0ab8e0a9a5250c767489c827795fb2a293786448701815cffa64c61e6f0db8f4ac015efe3b29c976d188f5e7c3030b07382879920f81f36ff76d506b942f93563a40b5b71cdb4bfd8ce89d2da8d0c18b0ed3880fae035ec7f18c90a928b0e83d469f8e0f40309d6c2e647b9dd83e87ac4a19a653cef7f5d5e0672b53f7dd2bf1a1e6070a3d0b005f2b1979cf873607a011d5d5d8ff1b497d9c5ae1f0b1fe813416035d8deae5e9c808c0432a35cfe979eb7c4df771f9e67d26ba34257bd7f6ca7c8bf73a5603e26f79412ec53c03e8d0c4197b806bfa8444a8511bfe5b09779ef923912994fcc274eb768cd9a25e210e95800a8a61a7f466b1eb3dc69ebd68f710ff43646f19869421bcee28dce68cef6c56700a38760b1e9a52e4f39963b4f931e04d45c10eddb261499ada984c403143ecddc4d00c22a149cdda5b8ccea28950b275b47da3949ca641033156078dc8406ced3e612dc913985f793853375b610464d612e383359526d0c4d720504cec1ca67923345c08a6d9a61898d3d8d8f5723767a4f48025547af224c7446f1372cd4126d6bc312baefacaa3e9a2751a02a9a725b986b24754c227fc562a7c42cad2b2242794e7550dc7e453c11d8040b1f7c7a620f3fb33c9f6f8258260d4641f605aa4a4ff234cdcf69783264d2da6c5bea7ba85caefc46418f56e1d5348a0231404dfb9eebf295c7b0681791430d42484b4c3b92fd79d869340b7136b69a1ca3ffcc2e74000230949fd83b6ed5b7b0cb5b73ed92d6f6b471726781241eb689f62ca65008d2f14f49e2594153f6fee2099f4baef0e10dde610734ad5642b6a691c75ab86e4fd20e980d75ad1363fd8419e4ec61c507029977cc8b20d09da36a36ee9c3e4222846b92ddbd0e37b6d6cf7315ffec91d870e57aac83a652409a1260db51f7bf28ebea9f68a92b37758dfc489ee754f31c6975344f4cb198e698fbd7900dd388101cad6caae5844cb55cce0c4fe607046ae915a7ebf3e443e2b7445f259e0713affb9860124159bae0f80921a5c6900a98dea6278c70cf7ade2a69a08d5227d12c6d53634f19efe02f9f58bfc55984a5cc3051bb65bbeff7d5231dbe82978c546b7a3ae64e43402bde7690dcbbd7384137671d6fcac26d69bdf1ca0fa09356a746354d7f1825edf1e3b6d7b7beb7afea2bfe0fc510d2cfa1694bd5645e1d776f97595d6d271e4aec34d0312f8d1f3645ed198465c15613809fa1b99fe1e9cc561f26a16db7f0e5532465b9154090ec4f126fb453d5dfdf9c9c84f44e873c55b56b2e94293ca3cfe7269b1ed289de0f9c462f7d5753c99dc116e1a91e8d8617e1ee7dfe8e2d0c5be030e18fa7d562609c06398979df544d7e82982e1cda93ad3bdd18a3d7778ba0fbb23727b8cce3d8034c9e22335ff25e811deb008bcabbc686db8deb046647ec5fea0edee33a56144bb7ec3dba586d9eaa74c3572c39251f660cb5752535c9e79ae6ac27d6a0e8a613b3a2cb908437da4402e15ac0d499c3a06dd71cf101f6e64343163864b619215304b1edef8418fe72512b45a93e7115b70790aea19d3f19e3da7be063bf59fb8e902a0677f7443385c161563498daaf18fe10d9150865da253d47f92042952e7fc9ef6dc19fe10ec3b4cdc57dcd0fdeec39a0b9fe2ec12b84e7ed6660712a02b5c4bdcd6d2de1c383771ee8cc992240020e15d1ec9c513084dc249709c29746ef77f0f557dd0b14e491be98030de08087d9d680e31b8685777f4ecfb2b4cae41e7da0c450c40952e8b3be59a898f66348fdf813245d94d057277bca50bbb56b569f95dbebb6c3129a8416833a1b255996556abd6c902866e7266d7a04891908642e885fa7c4f786e4b71d71ca76a6c7e945a328dd0afea9dd65993b370829e0119d8be984d148b898b3d870e3c8033b4ee65658bb22aebda8679fc9c2c8e814764eab8d999fe18a229b80ed535a650b1e47ebb657d239dd6e53d6f89e64bf51b98eee00f9663f84170ef77a0135290b8608906cbd6e90f1fa5c57441d96899f7d550f198766b36eb654a497dbc1c05c5032ef371f4e5e4126448342129d63c66d49a6bc0ef367287a366e7d7f309899711fd954ef9541aaf413a3ebefcaa3840c5c654082f061883144cd2d695d3c8a0f9c7cdda1d44e5f4fb656310bf493a79514068fcc37c76fa4df9f4e6513bbc0939739725422ae0c484dff4974d117ec3f7b5e68984474149a4dd1e4a6aba05cea76668f5cb1801dd84c27d9cd9c60bda9e806b0b93d927b2290d4ab69446e531c71bfc9d2da70eb58e613bcf0491b0084ec85ff80b46e213b63b725798beb8302128d5f7697c120255a8cdb493661b1894a2efbb4ee1a17f6fcc633a6a2f102f06f89d30233bfb47ead624f5fac0306a1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h72daeb7238b75c6ea75d5ee16912a8921dd9a663975f0f0dd24dcc29bf2ac01ca62b428cfd025d917a0bc8827a402c332272cd37c9e61abb58a0a105505ee1a8f31a56a65d8dd57eec5c5493ed719a859f48bfa5a59bb7261b67fac29c130a337e98bd98953daf9e59de48c48c6def13b1eb9e510e3bb815173fcbe81877169c222de02e4871e30ba10743527a5d86917c71292c6e2902dac2631410e1b67c107182f178bcd645c818ab523dc31ebe088b5b9c5c1d3ccb0bb5ace54a38a850d81d04d73b7af0be87a4338d287f1a8c16baaa20f30032b87371c2280fd01b33759b03fbefad132a8d78fb024c7fad4a75fb054a47a366f495089ded72ab93a7377127d0da11bf3b96c33c9caa6b11bf149521ec324301da341f6c6319eeac4fc452d545bfa9d0666b9a6b4aaeeab1acf19a5db3110bf406a090f81ce0544c7d00d705bf25cf5bc088ab63f4e7ced1b2326cd88949ecfab9682f3b3cb95122e06c674a97ee153e0a11de1cb25e7a17711470014b009afc8b9f64e3b41f53e9643f69a4e7ebf493fb4415fab5853303a798364dda271d6001ff7b0157fb5b174935f3afac01acfebb93fbdbf21300b93d1ddc7d9b5695f9df8fe0997e6ab5b388a8c8831853d888fdb7e563cfea3c5abb11b87a4ca9098a3cabcf2fc12044cc1afd30176c5372d681718981b36bd785768243bc76e81f9ad4ba2fa876ce4e811081a66ca7a8a481c1d650f9d240824e50752593df2620ca8efd0d809a5e88a7b44ebd977c110a96409373e62877caed255e1d16483b11b8a03fc8f0856a7c1873764f9dba37ca1345d17054a963cff2428f500624062ad997f552e645ed432704c9891ae595b7b9940d3455b7dea8c2b7380928abd314f39af526889d889e878eca09e9d2a79fc09d26553ecdda7f52250ef1d5d1eee337f18a1cd8c0e122e1f430628f53f1d62ca8484056c41ee57904135401f76be44cefc89a033e164c34bd309d6e8716326ef81069bb50c226173921d48d2586f6921e874ad2aac4b1f2c434b10e1a7ac584d95c6ab1b75aadd478a827264f18d7b771f680a20d8f1b9a3e90b2e49d5a998fda591847f06cfba8df6034d471857545b3b5035b320984c8504f842b5f38cd22a37fae829a124017368036b784f4788469f5a40eb87653d9c6088e0223874472738fc28b302aa2e7e0a8de9f7b0b666296c1eb9a49aa396450542e39837109ffb6dfb48f363e208d19217a324804f51b49f1bbd95cffcad92552a209dbf17aab3231aee6201d851a5d8e9005ef041576c8bac5e3221598055e5ffd607d1f4f0a59e2cba3731b51b0fb341f1f808f5825eb8c3b150428dca61eac23ac07581009fcbd75678a99b527c984413c44e9b253e03c9be66646c34f638260958b978663132c60e0fa8d4ee67fdd17d2f7caef8a19e2f3413a802db9afa7a79d6a26224406d9ddf28a0bb0cf787656f402001d6e191f1ee822f69909caa86c6ad03974b3d148cd7b49e94f17f1daf14673ffda72c98d0f400752557e40fdf5f56d44a770d37a7f7669c2a29d53592e507bf6148590ca2300bcc7cc38434f10e18d7f3e33981cdeeba2574b670d3577466c5f09ee7f748d085513a97955c0318a219580ec46dd0320b96d8bcba2b2eb8912023960b7397dd0584c98a3c8a3a43888c2a617bc029e202d989f522e6b7484b03e2e19c4e0bb0ea27b5d95ac501e8858d71d08d4b5e15ec24ded9e3aca4ff53074e15bbd5f37b86cd42e15231d8c6ed7403e5756511158470fa5ddb91e1a659e6b983895cd0cf37403aa03545e6b09778c92e936b39a920190da9333f7e7b3e422901115b4122c108b07909ec5212ad5a9e82a0f1817c407146ea71c6536e4301ac692888fca4c6c525e102030b67d0a1e4ecf17672e1aaa0d7c20160ad6404a0f3a9810d205ef9184683e338ddaa99459d58cff7533f7b08421d129e58891e917fc720167205895ce02aa3fa5800f1c58b1c6c2ba358e7defe14d0ace4f768c49478dabefaba1a6d75ca2a117658d89608eb7c81fcdd1c0569519663687378c81a41f75bbdc8a87003753d37ac6412fbc91a6f4a1f7d670328fe3bbdb1fcfd6ed3d951e316d1ebb260ad250494bd1151c2de0ef4ab6920e1b8875adbc2d9a285c4e6394e58ad370e8f5ebf56fafb35ddd6b51a6bee258efd7d8af7599e97f0df6b0c1b4f632a216fdeb3f7f8eff7f198190d77ecb66fe6dedcd539b78e4f08366afa9a104c7309a33466de58a62c421ea3a97ad2df6a4d6e354b2b0f94e500b4849a84ec6483e256cbac604b4aebb5bf3667e8fe56b06d3ba3464400dc1f8a8901c54369ac9c7137dd7a5a54988ec1be5b3d3e834f05d4c1ba8552b4223d5050f261cf344628d0786ed9acad5be2bedea165c0ede746066fafdcae9624af133fa65afa36fbb4e8a3119f871f29d4930060417bd1ba71ea1a46f99b875f305ddad868d4769532df96199ef3b1da21b2685f24e7540ce2edc4aae06465a42ea46decd926b2c4aafe53e428b5d5bbbba69e39469407672101d8129266925bbf987dd9f369b5f82d8764c7dd5fed82afdf8a2f6bdd3eb3ae4d30ffc607393e7b5bba2bd04d74a7eb69d82d0d38b61b1850e63b70ae94d5c0bd6ecf84c35365cc3d37603176dbfa9a05718361208b77b0885d1ecd9b5be3b16cf93826403c61045f463280c34509bfed1179f82e1554aa6b1dabfbe0a4be97b0cca1cd7605a1a15713c7925ab025cbd0845dd403576dca798dd2d5b8e3c306a3903597c96ebf07ed6288dd9393b59bd43b70c481e1896bc3a32fbe5bf9addcb8f10480b38b1341b84ff62c456f4bd447169fd7409d3b60167ad7393d4cf420ac6c229df28fd2bbe0e00ce100cb37fbf87d5975d0d0ead6cbff809a0f6d5777a85abfbef6b5d178cca5a7f93a4b4106fed70f7f52326b27c06368d96f4f156bff45ad14f52975ff8c27f06adfe26a4c1f8a62afee4c3a61a0e09af4c6c0e34144b889b7a59ba97cdb35d2aa9712492c604aa418278beeef7e6f22e5a2c85819a11b1532ca6dbbf97cfec6f15acda4ac9fc6520ed9ca7b5150895b39ca6a8ec7b0b3d19a2dfbb4b8e832b97b1553f1d3f3e9fbf0f24bc793afba547fab654efe6b8be9ac78110ebae0d9cea860120ab57960c10dc08f0e539e65b8f5a8f45411e82a57239817470c967221b42b745176e0587da2472eb201336eb4e4eac5f2593a7deb520acf4972c1d1670a2f8da9cbfadca06f4055c315066a6798fd070a1bdff23ee2de5656e35c65447783aff41aca97bb8461ad68807a46e02e63d26066588f5a1bdccaa0ee06b81d092fae5ebdee5fb84c27695a38ac1399495ba29b9dc7075af2e17d5a9ae158294d3b2b94ab3f9b2253a46fd4fe3f7acc766530fa49f75c72be1c88149cf8dcc6382946892e23d68ab83db5f7dc6efc35bd8e0249ca56a9ca4fab4437ed9d946a16c8dae5ff8e2f49de084e7f079fad84b4d43e7bf825b2c2292cead4d920954c955f3ff5fcf55f6e9cd24ea46d002aa5be732da515d6c217a27679e7765b671ee46a7b62c409549cdca02dd4993c0d74e0b261a92337d82f683cf7d3c87d3d0fd543271a89c15d925145e8d09b9149991734a8543ead3a4181db2ca43ad9a1c1993b0bb17f118f8c3e7f64d1d209d17fff9968bd615f9b4e1159492ca94fb832a296154692db3a77bb187add931511880837a9d73e64fff1d180be17ce22bcdab9d13be21f0bf69955bdb4bf021c6bd2b815eecd831eb9697c0b83284ec8353920a428c0da75821b2a49833f98d47d1de257c04333573f1731cf87692da7e47bd1d03994eefac060d5bc5d0e0ff78a2a72171a0c3a43c7786434cb392c09f54bc310feb611002a85eb9be9aa003fc2162ec3232ecbf167e131759b5eb5ed42609f042643af20942a839c9f6b699ef27c160476eb849194aa8d127c032e492685dfa0b3f18f9ab2cb80c928236789c230b3286a031ff75079dce52aebf804afa837ece38d2eac0535e1d993e6508fd881b851347b471d5d2d39dde48cda5d934593f42132b95b7957ddfbfd5f3e9c234e109f155f9671868ca9dd11fee62ae82f9ae6fb8c6d5790da95726987b28ac46aa4f681cfb7f68a99f17693fd5ba9c9d10477ab3d5d8f6e822f6bf5f24bb6b3a59726642be529e6468bf5e56101d06f2021d6b6efc660064acf98822eaaf87564c833dc05731933bb8609408d77a0b42a913669ae9459718fa8e8eecc32fdf9d3529e43ccac0f11113295e2355619352db425bc86caf73b24d1c334f9f69832e8937a33a88292e84036c90e972b8f2c6d79660d9b23e5ce1b74e3db44cf4f7393bf564385a2cc5bcf22160ee5fcf0924e19c5339f7270a252a6b8b6da38b44500d4acabf4190bddf98ea6da3babd05de1ed21734e1238d8e75a4b3a40f5281398d6c707c184e4c0d700cf4255e8e33826120e8884a21d93cf89782d94bb727cce62ae5c13cd590513b753bbbe16567d8f0e0339696a65cc677a08e59198b0dccd9c579e35c3338910101b69280ab9f44da950323dabda4dadcdf0b7e154ab7f49ef4855cf171eb6c929379c783129a4e0ae650e55d90fd90ce03e2e8a6c50a31120bc46c0206b5cc53fceeea5ee84eb27a2cff264c797e33ffa14d2dfc57ac76d6bff3d0b6c6a9ed658cd6daa40d0b102cd8ba6152f5db940207d7286a216676af2aa54e429903c3d5093fc588ad7a9f02e10d141ea9ac322d5be19f595b13de95ea72d0ff44826d0cf2c4de6d7cc6aa2f03a7984aa13df84866cab56a1aca645a602966a2112df31d7b991d896ca72e1c05545304fba2ee46efa7b119b17db23e3384fd1d0d4d3f47c39bd94cc7afbe9239da4ae1a503bff671c5228dcb4093b36800bd22646171f83bef37a28bdf46844e6d6e82218707fcb854e7e15f7f5a403828d15c6da803abad2bee2fdbfa10d4ce82dbd909cbf837aeee3647f5f08dc0f218c5b56a1004a2a2181f5004a4f36f05790cec45fbf74bbe96406f8be757689d42c096146a1824ab6f71f5e174e1ec9f51e5f81f258720d27720de280a34841a0bb2d723df5768407f49bca83134beb99c64f476938dd2912a3e7595c09b652ef56d22b7d5013ce46e97a7ce313961ba962496ed81ec656a38796b98f0ca70f66856fee646efcfa5878cc082bca39666cfd235c50a9ee5b7bf7d753bfc51a414b8ad2a5c70577f667a9ebd0cf48246e20561263b4afe6bb3a8dd78424da25018e43dbd92de895c7c5230ac4ad99e5bab502a8537bbc0555e52c19f8a7eea42bdba232d124c38d0ed25f4046addaee5bbb30fa268cc607e080c2abff80aee2037a75196fe5fb92f5af42688cd51047674b3dac30d091c6ff8ad7a4b6f9483e6f42b757d01f86a74e77c63659b8c093fe8daccb19c5759793791bb268f55b971ee26c67d3534632a3404779ff87d49f953b0a0b4a478cb35ac80f51618c8823e64b58f585a536c5e3a3939;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hb79019034af11625824984129d39f70532064e43553e1ec7649d28650c13083f520dd017abf7c93bef7b46fed9efe81093074bd70b6386f606486fcc8913dd94208fa36ea5c1c1f263fe25a6f2da75f988252d8ecf3c5319bf544658549bd683581d71ef7bc2aa96305cd3c78a1aea90a393a9ff0dc31725928ef9b7e738b18253e573ddd845e3b234b1a863dcced31d8bddb66ac914a3872fb8f848301af59a560109d8d21b4909123e001ef2064826d34287b1a5783da6527cc903b0e42b0f0ea7139becec94d4ac5919a8ca18a3a6825568444016a543cd7e87104e2d32b8c933ac6785d885792b301510ad2671e253c97753e02dfdbeb575b9a2e9f0fd7b919280883878d25dc1a299f4ccdaea57def558e66e23c5efb09f41db2cd68668b4a85b18aa2374bfdf99dbde0257345a497916be27e553b64e61f775ed653c1b8a56ac27b24fad9d7f17af8ef17194b8bf722c1a54c117834804b5799bf09c9ea9359f855ba21a1a803ec694e02ef5d16a1631aa470ecdebc6c89f2d58ebcb5088271486962befcfcb71821501d8eb7c09db2346f95daafbaeb751f3274350e590eea02dda7a993feb0f5057ddb623e081df942208f5e5e92d03754a32f9e8319fed79c8f1ac8cca81e35ca1f692f92523f0560101bc2a97e8086e5288868054c51114a37926e84a46642d404effae8b646792682fe5af397dd0aac8f4903a5e9c207af25075e44fd76cc18b91d39cb97d5655e06326a8acf0344c44692fe2e6a292077a35a83a6b5cd4dbb274ee8d4ee69a95d6301bed3adab606e760164ac22ebd53ba5c5b1fbf9aaad53b85eddc5193ea5b8df74b817417bf004651983aae9faa310fda054950df9c098ec9663c2b29990ad6c2707a7c17da38ef2aea9fdcd8df901a811ed81415dae52fd2683719d2dc1debec6912cb28df4430ab21b3fa0b7905f663c6254015799fed3f13af3fe3431263325c14318325f2ddc2948fae6695ba783bac1f2b1052e2fef8d3db28eb04fa89939d0d38c415815c26a0afd1454a26c8ed6ac0a3953de3fabb6d4d9b7a2c5517f8740ff809fe4764c53bcb9c81ddf0d1dda3660e1fd29dc8d9f64aebb75146f90dacbea560d04ec8363eb7c06caf01421b1ef10af186506a3ae7a394768442d26806416f103198842e59e4f67e4fb38b2a83343ae36d299f2f3067e2df477acaef3bad7791b6d4b29b42f10ee18d89d32345058d06457d256d101d47076c73d520db669953eb696da5c4b4cb21d86cc4e2baeb50b0e1147d69c881972b5078e9590e11c949ca3a3f054fc74d2db36533c578143719dccad026d119c2e48bc93c27ddd5b28aaf463f045529f3d716859002c3e2c820ca901c381fa63b28be4a9b5c9e4c182ec4d521ff2ddd9933c835a1ac80fa4d192fd351feedb96f69ac0cf8fb51e8916fbfd7bb74bb066a5ebff9400f4076fcf4accdb07d85de898930f911518a95ceabecd6761051730aa1dcda3e4a573d22c61d32910bc4845b458985f2ed62a45dacb4430c6f1c2c252ff65c38e4dc099ea3e88bcb511c096805b5aa2319226cb72f7136bdf48309af19f6143cd3d9507c6ed35d2b839a59be281688b81251910a8d9f9c78b3a17282eb5c9495df3a2b0651692f0ab12eb336ec5ca4964414b30b5896ad7d065bb9778f2f5ea4541c26b71933a2582e02b40f0738a73789956ad66f8c356e951ee1fe673135e41c958c89ed29b7e8631eb50917a7ca7267fce10c7fda760164faa2e863db70e069a5f512a943d65cb224a256270dedbd0230d13f14f7e738c28feb0020463f2d0e7f9a6037c9504767523263ffcb3d1a8c5f38680eac496170b17f1d7c1fed28369f1840be43445777487d20109e37e223492a13719f3c236f01fc10f2fd8f093372bb18475600cfce44e9bb3a209d794e15293c799535e87e83877de41bac791983937eddceddc1b7d91c5bab473ac56f1ee52f6f3014c5c4ecc0101452b1bd753fbb3c8c2cd36007e6cee8766c096b672084a6b221eadc554279afd180ed50e8b41ef9162652e25fbfb5e3cfe08751d8541cc88fb8e37476eff76bc701159989a7bd0a94e951953f5a79d3d18a34a8ec27b1b645d5bf1353095ee993bc7c392c3483a593e29e34c632b23b5320b49f63dec3fe93eb106683fc9c28d6b4073c2081b110d52f6a04b38fe485161feda8bd70fabf928e79bebf6679a46aa4c6d95ce908c3a8b9cf79c8af073c532b041f49444ce006b85a95bd91a1b5bfc446c964326903046cd23226de1c633f9b635c16f2d0bdaa306d02dcb18ae4e103d5984b7c9b2f0f8a14b645673890832e365144ba57b0ffcbc56cc20952c9e118dd9e9e23e623d107ab67869a8c307f0be7da995aa7906837256b298bf5731b3552e8b9254a1a7b31be6d8b25b788e26d41a55007367d13aeb14ce341537151c5a47319f8083899f518b30a76fcea24a99e6e7afb2413a9bbc7d9f9a5028228711637fcfa260425fd899510abd1b481a3c9489e8b10192fe664bb6179197ead6018911370fea5245b0c55f56de64b3463f8a357c7396da9fe3ad55aa90c94dfa39bdef94a68e53529fe9bf2c095b4747aaa88f5850ecf6da937b777a095d82cd5aa0a6a164cc4e6a6477108ce434d5e293fd7b734d4ed4e7df4224c938f0b688b5d8fb0032f770fb3b8f7fe06977d0ef49f1f7283ac9261158fa5e23d83c05aaf5d7df842cb28abb1c2caa4474823f2a80d5381f93dcf1dd5d68cbfd607d01ffa36b376d6bff427d9a840e35bb25a8b8f98638ac86518f4f778b9337df7efab739e3e844fab6c05ed0b8357548a8b1140857be196eaad92ba313ef7f34c97385c65390d6aa40978a082713a086b8d3ab7dd0ab166f59f1cc6c3172b0761faa77c395d5a399624ea1a2304e8327d60d86cb7ed939870c5cd8441f1b9075b4051fbf00fb625bd6686ff519d719faab2d4e5d2a58dd751fd3bf087e64cd33bd9ef8bd233f77e39fcbc487da8b3331d58ea6dd0958886e95586ff559f58c785b1875ec4ff1ae1c4147503bea88556568021d7ce0f63525c7231c101541735af137270e8dba68054cd68a7252970606c38384f4cc345930a857bedd2eb137048815b900fa880dab3d67f656df511b7a21dde77c0b8adbfa7e957713022786bba74cb057b9db135f30e5fcec1596a9ce5499cb1f3e72f90ea23c50ed4238710e49505e4a0e19ff7f5520e5061bcd819184b056c1e9f1d117542a9ee158ede3ec47c3501cfdb26d40c5ebde092fb103e93f4ebf4252c3afd4b1eb728967f389b1f42197a995ba070cf02ad77628a7c352d3de76bd9d60e58aba1012953ee301e5f31b231e4075d382fad3293f7737593bab66284d62738adde36daa24ac4ef48349c0ff1721875f4ef84bb0e6089afad50a4ad3845e214ef4e220576ceae08546c9152d292f4307110db0ba1237438f1ede44dcc67c08f843effd10af1c5fa9e64ccefb9243a6e66a141f0ba426d0aa3845ad832aa1b9f51e80f22959fd919d75af098766b5512462b171d95f569277cbbf5dfbcaf4195a7c52c64306d2794af6e6eeab4c59cd75af50f3398618ac4b04e4d6c5088e207f658231b6f5034f347a8a1102a05f47f11d29a05e775c740b59a876328aac05d7ee50dae155e6967dde30e82da77ce1d9a054cc5bb18f9599ff958ffd7708193462f3314caa71d96f9a026c8f0d5c062375158d98624a6b80c89975ac9b9b732ec468a9e715809e97e9e29cadb7b098cb98487e06283957f7b1559d1d00b8fabe5419361ffd371f2bebf9559d15da4b5765c5e0580fb70dcc6950cd2c09a2c8a78a10707230502fda5028f94eada5e7466280f0a4779f9ffdd6cf31040a0fe36bacd52ad2263745b2f137be55a7c53c83eb72b44646cea44a067ceecc216b25ef980b4a236b39e3b6ec73384be792101a3427ee5f44ff9f5a407c8de1e38c84fbb6f7f4a7e86cd58ac28524d449ffadeca1ec275326ff8833140ec6a84ee6aa7803a67c57cd783e890df8bb2c416ba38832b636f481f6c28f800b44216b53f2e1a0546d52c0ce6650578a3dd4d8f88672ffca7d86ed6881aa360388172ee5a9ca8c158c1d5c4032b392306078d592bfaeb1c03e1fa186d613cbec46fa1b23ffaad67375efbed156a9b8b9499df53c439b8e22f9f27f15031e3a0b9dbf94af069aeb1e42542db5f54ca77a6667546b33a82585014c4bb587738b37a0a15a8c505006dde277a15ef08134c53a6f2216a63f6f08173ab9bcbdff5527a875b41ee012fd3e318359b8198aa8c1c14cdaa63287b9c2be322f21647595f850ea168e3e92cae8bc6d615e420fa441e55c785257764c585b89ba32cb8fe1c06ce8b8bc31274fc8cb646668a00901b12e2fa66a1dab19c6ccd83cfaf8c9adb7a79781fbc0f88c122b64710421b5a11409d1e7f3e2a3edbfb7a315a2207673d88187fcc5d352254b459840f2a58e5aa54cabe086736cae4248c77141c3c34465beaf920100a76beb82a61934ed188b2e29244a465b6194243c51285733e5e749720fb03b101c93933a05e80dff09cd3001d3f3e0845d1ba22f013d539505f772bc40120fb4858c865c4ab69d11f5daea4e23f1073d80efbf70ad27554a71a5aad833afb0baff306b140a7ace6411d261776861054272305b426ccb2a75d0bcff5541cc8ccc18ddfff92e04ef7300b20cfd13bbd73b9801033047c78bf35437d22e197bfc07869ac51eacdc7494f26f1954342c33bf842238fe5eb496ad0f39b732d97b03bc16dd50630a3445bdbea882cc606bc0b5a6305b8e9b3e773af0078476667f660347a0aead5761542feda0992592c2b272fac1fea81bd11ab10dfbdf921cdeb15f2d2089fd71bc0a9464f5844d7b263340ad2ca29e250a617d226f5ac9acbee85a519f18893a05ffb0643094fe762e946f187bd220717703ff05bbf2ff2dc778294863ff90d77871871ce395b53b3afd4e281c8753020bdab73a1829924510957eccb2d38bf192a96be49fc8afad0c4c9dea206d0f6699147af7b378d806777c4d999a85b432f136d7c6cf6bfbe0bce0718b7ff4d2ed221ca3c1d1a4dcc7c613c58927353546596b5dad69229ac828f69c6f3d60ea7744a326ab628b2c51323fd3d5f222ef06e5b4a2d54909b1d10642b63a3561d75fdafa5cd9766656df30f10d33333302a7cbb0a186f2b6f901cc74c5d2641e33b4072fab0644322c1f873a9d4dacaeb27dcc5e2debbd74426350b5b0daf3dd4159d5cbbe1bd78cbdede57808c89ae15174b6cbdff2b20defcb38f3d485dc94383055c3706c35fe30813dafff7e76ba8ff50b600a6b3dc879bef3ba56607a63a1dc9ebbdde55f86dcbbbe61a8fe3bb2de964816388da5109b8e3293dcb0d3d414b2a90d2e5213d9f58d3bb1d5cf36a327fb007991dcac7c23f6842456d31a3f60b59555180d34e674894e6747ba7cead5c47937a4f3757a95926ba6ff0afbdc2bdd108566841bede;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h10aeb5c6c7f464a1e97fa40ebb21c7e753a12728e51dcd2c2b9a65f01631e65d9b9993cba88883130a51bb225007d20d6b5779a51d714abc46a9fdd2d86dfcb538e90e1027d1e61c5f5805b997c91c22d0c8db1ecf9cc20265c5cf2b981025637e5ccd400c8980f72a741ce05685b8ef3b4022de1d287f40a2fe5eff70a777bce3500c9413045349e1eafcf2e861abe113a7ec06b1192d9df7ae3a92613e111f9c104f09c70a6e7b3c340fb6408b73923b3881fe443003a85a216a999d7e663e3e7d366f109eb916f4dbccc1759b5267876d2a45c7a4156c14e86408a2a51dbdb2b3805acb21f3a82b29bd61e5b7f5baa87e70a3d1b85cf1f40aa851ebe3082f0febf16271f62c30d7d498ef29dcf63d0d6e6bcee92a7ae925ee664c14b0ef3e803a93d09971cff12530c6d92d7e233c73f992b9fb84996de958838a543e6cc9a0f4b800c00adb7d4b2fa0842e2339ef75a6696806cd0d6d3d9502e5bfb09f5f45534c29f086e37d962bb8d904de45ca7763a6d47fad69e2519a3d57a93676db1b4f1921600f1ea13cd6f19f4d5eb5c9e7758d4a493f06f1b64869818bc05a559dc9a5167f77140742f42168034d170476ba5fdae03fe69b58fa2ebe93b06c1afc811bf3fd8023d0b7ac2f1bf86c8fffddf7bf9ca781d888131c3c6901d97f9e6a2d67124e3224dddae093f899a0584752923eac8ba484d1e8eb6ba453e7a9e2a892ef81422300d495376bfad5f53421d7c63c896127bee13c401ac493506669382e8c21278b0a387ccf54c2df9f19f148716f7d8a972e6f3c2fe71e71c56f5c29d8cc1389e97d8167f8771b7aedd189c61d7bbc12dcede16546f1add28abb3ebf700578d88c6759910cd8b078d6131271b6e5c9076d1476fc7054f09ce7208adbe7d6e4f06744171af8f53f11b1daf9368dc4ea54707f37d12daef22657f67c4d484ada509caa87f35314d91c06811a384ee049b7aa9b8f3eecbdc82781c796f1584d18bbbc6a40c24aec8b5d95458b61ba156310f8b5730d7930e895c8b3b8abedb1b85e34f5e939708406b1bc731b76bc8dbeac4c994ad446d8899622f03cab6423bcf8d2cf305cbd95eff6d5ad0f38d1604b8b4f14f4471570d55f4400552acbddee7e4e65685cc015ca8cc027f3c217ebff184cd0f3a25778433fbbc7fb29689e66e79a2d3839e8613ce6f54aaf0cba563d0069039be1aacf7128d92c37b56f914fe665a2bd903d1f8449a7a10f1d438edb3ab3efbe6c68baec60757059c39f764ee416ecda0bbd7e52c53a9e26ecf31a23040c65db70ad39fd81b45a1d6e8db929a24598d79801b075b7a15e49b425b07897883bfe3df9c12ce89ce80290438820687e06fba4be0aa85cbdeb065bd3f38177f9b1eb99bc94b85a95b920b662c5aefe58480a23394b9559b162c47ee53d82ace43781457ecc47408c477ea760df0f8e1f27e3d455a66aab49ff20503f3ae27e1edc74bd09e78c3ff83b7745f63bfbc74612fb5eceea4944e311e739d6fcbd96e7b7129dd53d3e6dd9c272150ab827a0c4a782dd55dba9c17f29a3ff7d7678e633105d06b4e62cef19a441ddfea32a5ef521177b77048ee8fc254942b14a8bd5af60dd236b2cb1f025ee11ac63f6fc6b46457437a57004803f02a6f4f2ab3cb95c1c762905d3ab9d55987644dc0ed9cb3940adbd043d2825dff9e7a58d9b53589217a85ca7fbb2f74e36a59e29871689a0d00c1859b389da84027e6c6e56bda86ad3588efb89b999e659f9ae796c2bce91a96dc088c7a37c5bdd0fd71f14f5b09fcdf173c1d02d9b6daa4094b1f1509a9e3a2e93cdc76fb8c4d964a5f3e56a61789626ff11e16391189cb688e5a4485d8fb75aa4944ca88a6cde03c68234a09ba8702a674b3577f42962dec3015070a04a8546c43edf331dc72f3c2023b755b09e08b3cac5758eed352ac40d137a97ceebd5528f3ba8352ba4ebbac457e79dedaa56dc6863098dddbf99e6d079f022c8dbd57e19c171308eeef85ce845c74879ca6fec10f4acb709874955a49af83b73dd269afad227cd74eb9cddeb0f3ce10bd759a4a0f07dd35719f65cd2ccd708a07efb89d371ce7b59729e1a71e2a3e5176ed0da5076f851c4c727c206f7e1754bf056d9518ed2ae22cb7fd0be078c12eb07a903b77022aafc9fb1db9c07ed9410e683c66b85cb4919cc43d79efe7e98f925d547f7d83a5619b499695fb0bba167fa4cc312c47df52b8dc362092fb1f007001807d83e446ab756063bc42775350bbdde6a2be40e3e5eac0735b927fa5f1ca10eb6e243654d4ab141fa37ad96c18e909901c2aeccd65985ab6e421a7e91f310f0b52f4f9ba71867c4532824eaced0e877b055558e82db476d7a6ed2ef1100c16e18717e1d664ae35b1020a4dff8ba24dea36daeed493890d0157762bd8790348761d547541718985fe953bad84ff5113b8d0bf0b01591553cae33849bd16be36d9d34ce13b28ca114f6d90d6d80652a05a912d92fbecce8df08a006d556bfe31decca94715616f293ec8b2c2e15f070f188bb3f76544908456611e8685f73167867c50237737e9be06fa878d009f09eedd79386b1f07797fb56009e851bdb628c2f14f287f506522bb0e53f9078cff36288245ac58e94ff83e301a4392bc8707a77ba59e5729b164750a4c4a5fb9391008ab6da5ee7d02ff205f62d28e043b2efc9ed525f7b40ff2f2d7f7ed031a6a1893054a1012314788fe7aeb1e519dea6b6455527a3d444d5ffe4524069e5aa0849f6130760d0bffd8e776a1e16e4a05caa8449bc734428467b92f5792649cc20bb68f89a68612f1e8389954003a3d634c0691c3bdb5b5400c388819cf9389c0284f47b993d43a012b867f848270ff0561d0528d55865769ad13ef1cc3dc9d057fa905c6d76cbc2811e0ae530c892176fda6a6eb4f05bd73ebf2ae65cab09b8aeeecfc2bfcbbae6b5a3261f073d2750fcca5fe939fb7ddcb8f125e713709d8028482a6e707541ffd75065b3966771d38982de0dc27bf4c34b8ada5a8d070167908fbe990ebcf4a26e83180dd77c07bdd55f8b9057568ec7b2f24f1fab8ea21341dadc23d9af00750ea62763eef02c6c6fee03b0f1f041552c63101078b452257dedf78a025f7b3d1ccc140e7b3e44afbf4bf77f8ced5487384f85a9da9d0675c4d18bd277dca7408aa460ac09291f99f885220b9efb5ca897c735ea5975c0d2d97efbb6eace6a90e50db4f0e3ad6fad28c857e629086cebd69b5f126cc8c09fe656b5a36afdbeb9a8695a68ef78366830f2e2b5322d6c0bf64238db4c2120f265cef4ac47c5a59f24dfbc577885578331010327a6e85bd23f06e2ba3502ab70a1d8d4675f223c7dfad7cb7ee4073966ba7426840db75eea3b9ec8f74031933ae2f3aeaed1b591e91b3e5518f936f56d16d22b86a5c9b339409ba0fd81b131ad5712362ef246d7a08e9c04e766d399f6de655698ff20a4e52a2ccdd08ff34ab49b2493b5ae8f1a65132e2b28973415ba590849cc938482b1ec10f0021f489367ec867b1fc1e783e52a1a2a85038e910a0c8f3046545addb22929138e896831f399d933d8051faef4d0ed0c7af26e8e2a641033164b7e41b95f55d0f66f5233ed693d2f549ee33ab976860f607e78385159955bf55e85ae0971b5a22100c20e21573fccbfc49d5d267a2c38d0ee1392e8059d5a369b16727aa60cdefbc62dba50d582d0dd0236afc20e895c2a85e6892026932eac2c0bcdd573556a97aaed1b46a725898ba5c90cbc71d0e606367c1c2b1e2c118708006a56785d070556196ab034dd52879893f58c31923e4c62c12a492225785cb5e9b061089cd0cce3c63799f17bc767c570085f10c51e0beaf09edddb509a9921e1aec32921a86ce19e23a23cce6bca71bacfdad648ca09d3167c6caa7103aa8721576f23b4c66364b6629f3a416e0aeb734a445cc9e76ce96609275b45b55b5757e6b5978620fc712b2f8ff15f747f462c025c00010298a65bffb866aa19ff7683384ea22ef2f959a80bfd7ba4c667984ab5edfa47d130d9b95dc230e37de93a2dc849128398e9b91f87cc7e003a1dd52d95061cfac8308c012f51b5f6b844176046d46230619be0e14cd44c6ab8536e103f70c5e462de496bda0325fbe0c2c0d4b623968b5812ab2a702e10274c75f9abc8dd3e0e0ddafb1c4983a9dee74e6368bedf59c4c311379e7e897022a38dbc421bb168474b309ac8af1b17b9e857935a52d719285196ce1daa22a5bce8ec71ba31379ec17f3e69b2623c350a6ca7545e5d34b120245fe7879b1487e7f36532973f235b4ea17da4531906a716bc06c0fb3606c23ef65875b4501bfaf2a45d082b3f795b0cd56eeff115f5625e7866d85a14e59723faf40cd2c219450aa171ccc9d10b7ab46e208d8e53badb6511951f12f0851830a69e69afdb55642fc631b46c950dea66619630a853a65c550de8bf1e753af0c4bdff0bdde7902fee8c1b4b942ed6c26d4a3800502024942648990b8220bbd83dd716eb1d492551a1db147aa87828cc6d852c58bc5949b6f058873ec7a14c4f7419d93cbe3bf51a1a913ae39039ad9f3743716940750a6b4cbe4e8f0f76b018439aae73624cd8c10761b5950de2c7354e70b5527f2a40ca6b55acb74ae0e38da02a62be6e757e9bce8a3efac5b43a2859f367db8f67f3160bfbbdaa2213701a259be533d4905a84856680678bad233de7460bcaf076453d3e3e189895b5cf1cb10a6c8747d454d57e993d309c75095f057320f078b71fa1de3f273a33f188e208a33a24e4ef2f6fc377cd9fba50f13030f3c1c4257d3041c6ddc2910f66f0bc0d5dd56b46bde2478007f58bb7b233acd0d39122820d715300998914263f6334e5949065ae461317588f71c75979cc8fdae300841a9f29931e97299b634f6db27f1c1cffd2c2d7ca541dd91414ca000bf0c234d09a0a3cda74b784ff9680fbad8f2563cddc51ad937ed091320992a1c9908b837cbcc068ca94552ef2328cfaee413534eff93ba96b5e9b5fde241feabff739adc6e31afdd2d3b0eea6853c2992cbb369ce6be023ce22c31e11a5578696d7e893714fc0730f063a9ec01e6654ce2f5fcfdc5f99c2f0853a04e3dae6509d02d85b39d5c585071e9d20bda7bfce1cfc8955f0d199430e6fe93989475df51c650c95ff5f809dff7c703465d4e72db08334220bfb9bb7293c59063e4148ae80785778d2de1fbd327e291f318489c3b5a6f5aceacbc91c8540744ff133590296266b045853448dc9e1dbc0d02a499aeeafc40b9091003461f867079c817104abd50817e12dd77b77096c3133d004eab19f8feb7ceb702df7c5e7194678019ab4f824dec3184a4dd18ff8f5bf3c796943d1863c9834f3bfd235dea40a9e5c6e2d650e242219fa630660ed3360ea96fd11642175d8e976b998d4a6d6f16450c5133fcdf54b4bc5113e6c2a6803273386b2db91e7baed118ae37267249b99cdc5d39e23;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd99252ccc83eaf00ebdee81eb4021bef0223d6ccb8c061e3ea6e85926c25a5d7e91a0d339bf8848b6eea5d6d769bd3e888400cb6f9f1706262e7c8f06be96c86d159e010f156f6fd35e757a1d59f9dfcf82f65eec5bdda0c1de1d79a00b2e24d9f143c72a0de5bb4d11dfa9f725e3416bb3aa7e425d3dc8bc7517ebd364485da545e32f883055a5217d7cf17a04b3c33cc44af90d1d13157efb38dbce403ad1a6195565625478f0bd25b9b1042522e454b151ab4c80a0d86cd5fd8ad17a1caf6bf607396b5b07255b20d3b9c080ce19e2a4f2ccfc0adfe411192a3a552f0d7d9715a4f0668c4178a555ef924b08e04313e1643705fc2393072e59a3f571b9921954e6aac1dc5f6ba401b3ce8d396a1fc56e9f7c799a4df63119beafdc448f1ac81a23feb22a142a35793620fe28a5eef6d171fc964490ab0eb1c3241fff9c3f6db4cdc6d7791e0032cb00c815d7e916b54abee701c40807cf9358341cf4b42b336831636c95e60c3db7241c083c03f04d12ed13ed75eda1da1f5a0215d3c4c3f6e32bb0ad9f76daf4cedc6a097c3eb741f1aef45b8c054e5e54cfe761a6478ac3546d7c272307c65e8c0c664649b94199443d89295f2c279b2e5575e027d25625e909a248480adee9a08de9c75aedd1bd34bc1d919761e843384eeb9eb8cbc4d831e8a3a41484288bc2d7a49c4d3093c350b1282fa786991d7d83fe5c08e6dc6f9912f0af40c52536cbb15280637ee6fb1372ac30b56180b9cbf62033caedf2ce3c3daf933906d1fc68defd227e6956ff7520bb2c38752b9158d4e85f3a1a64fb6024bf1e7b3e1bfcc36594ed5673c31cb2e7cf2e124f30de69e777e615843600667bbb7b8262a9dbc300875f31d579d15675028052946301bd7515fb08475f99bba2ba444e44b1836b4dcacd0176099e085276a18455cd8e0344c3c343fa70090f1e679778845adca6d1d88f7665bed16b7604c4aa20e8e3ffab36074cdb315be10d6219568947027ffb8ae1b31aae25a5fb769ddb44dc27fcf865a4e0bf1c037ef76acd219ca2b9967eeaaf853bd3dbf35bf04a25d24768c2542bffb8d688b3d645040bf11e5a1b07d10b0bf09a5d0aa5634ca6a1bcac97accf98aaefe29e1c8800b496feeb29404a53b6170479b939c1e71e60ccc3f40495ced7e4ab44dfc945689280a50f163012b551989985f2bb152edf14c87f31bf621252b1617c6161eb63429c2f134771619c295dc4f4005317fc037b71e45f73213f603bb76cc3c5a3c9698739c659e19fb400dd7fc39d159bcea025d88228f7f3d8b04d758786f648d802a0b67347c8f46dd1d5cbc20937a524500913d8304c3926c9e6c6d676a591c43567bb39680ffdb294952cf4823081ec37da69740aa4335bcd1ed6e4bfc17dff9665164c01d4afc3ea3a9aa07e35857507e3344ab77a43bc5a29e23fcefd106f8e45363695876955e7a97c832bdb8157bd7aaf61335c1b0d0c990571eb83b752bc8b451b163bbb81c8269972e8ef7c47f2048f1f0058ad458b0c5d1bcb6202b503142bc39d08aa618122f990f09dd2856420fb5e76551c66de87c60eeb6ba8836197c41dea13bf4c92dea574e9a7e6379a83efc174aebc3231a31966e181f5f9511fec0819843468313b36ccabfca10f20e797ae4c2aa64d71a583397c86e9ece2e828314744d7f31e054b5280f39b575c80e01882a8fc5c88355f8858b87c1d56bf8bc1d29e38c1160a7d9d0f540fdf9e5d6ead56b3ac3d659f508280f45ff624b8b4b713bf5a28f2402e3592c312af1954d12da444d0d6bf48c5f5360a8afc41fb341ab9533b679312b136b84984aeddfcc36106022320436e2f398ffb6ea0349368be210910aee86379843fd5af290962905a1a1d704c84feded9710af370d400df60ff6fe1cb49611e8c512efe44a33c3cd09aa670205069dd6c80b1c5ca5cf015f574084a73e89ec917bca855517cbef06c23435959b15fc2bd6982599235c2aab0cf12fc6adfb540ceb7d875867788a26d4e44130ae343e2865f2b6b24737f1e94d852a8a5f7a84d0fce9d7dbc20e67c0707cb95723f319798ef07af725a2fcdb6207bf30a6a53cc9cc5a8b25e1e296f9750d37c44a962df5cb6469b9643a41a945534f35fde16aa1a1090d750428e3ff9aa0d0e23e7522bc6a88707d4edd29d884d7a5deb4f4ada7f29c6aba1d44894ae6e5dbd710e3afdddf906f5b8a0241c3ed8afba9c6000cbb298c69a0d3ad69fe81d9254ef2ea3be658e8871c1f4f4331c3abf919b018fa67bfbf71909eb5a315069e10fad76fe814f5cedc1452be99c7bd0cdb2ff29671fa7a3ea819020bbeeed06f0d33ea2f280f4a7870db79ac88b1f2ff215492134a8f3cdb7c06a5fde3d31f652d6c39927f1fe099f2bea677255698d804374d667b509d603f8751941060d6f9e472d017c831537b86ee784dff75388a8dfa1b3921203311a0c0e3c10caeb6368080e5fa44c4c4ec7e03fe1d5cfd09361f1d1f4bb81dc953bb71c6469b0f83791b4dd4cd30fd46af0598bd0d67ed9317fce2891a96296ff78137d0a8dd8cbdf5a49e2c432d74b489a9f0670e6311692b051b85b2e3510ec7da1cf4ab505acdfd2c1e30d8d1345d21e1252e0a705a04f1f5de9e583dc8895655d427f32107d3a0c126268f0f1f1899e1803e7bbd952dd3d87c2152a360b4c16fc9ab55d69acbd8ae15b66e106e7d8fbf1a1f3a4480c2647cd398d0c07c524b59388cb3d3495813a8e9640583256ef9463cc0334a84cf0d10a2f3b0873201e30856f14147b11996c7f317f0d7c01b2316aa198a9a4a0746b9c38690cb9f683da4a1779debf196b4fc65aaf86494bdfb3fcf72508a57f00d130e9748e4fb9a39aac3a14d3de5efa0bca8d8f9eb18ef3e83b66a5c0542a8023f9e590f3cb4ffadf2b26fdf0b084eed8ae0d15b1ea154081a2dbbb29a16df6ba43f1ab342d43b50544dbeca79be9861b2e78b80cf5042e509bbd5155ffb10589f447a3094393fc4176c3d3bb5edf998ccc72ef03c0075d305a1e555f59b8889ab608ee54591f2877fba68cb702380ea517f5a964774899a492a0aa21d6999261d71ec399878876b40dcec20434a7fc13b8e4dc965cd69619e23454b60982f2c52a3494bd65135529a7f298b03bb52a0ddfc3cc574599825edd5c01d4240376b0737c25b1dd8b4e7627e03c767330319b064cceb99809069e696c59b7ddf138ab6b26cc93c298372a66df6e64437a8d91147f8c393057d03b1ab44c54f438416c9537121b10f28580d58985a4ab9880d4a75fb5f55ddf49b63224b0d195adeb1015a52f62252061d095b91af842a4c23cfd5e591582ede86242a79184ef443c7c20ce2900a0a096aaa964a35fb6f89247c1efdddcf24da06ce3fce06a920c4cdd7bc615ce296708f75171a128ed6da1ec2f862d3670de0df4f84947d0dd5d651b381d04a570005468c7bec4ad149912fc8473fc9016ead04efc47aa74dd42025d679772c212d950275b5e8063f8429da000ddfba5dbe44e28ac1e1e660d9d63e1b1f620e373b43344e76073a254fb20b44948301ef2710485f42e60118743eb773b46b96f6c8cb1c9b549b4a602809402bc68877467fd2b2b5658b6f1542317f0665688424577e825d25a93f7f5cb49bfee239517aa12b46086a814be03bf3e1c9b470a539ae637059a47e5c182f69ca4414753e53abb6381a949927623d94da9ad34fbc991f421fd22a46675236e3c315a658964e383ebf8d3ac2cab239efe37faf25d19ae87d4e7ab8ead09e07a38b255ca00e3c229f4a0f73adad4083e40eaf951fedf8ae00dcc99fce44f88282c0dcdc0fdcda57c0b985579ed18cc42b2ec3a6ab195338c15f334d765ee0d380fa51c9e82bc14c1b7650edd42bc0328d7a3cca44069f58d9a4eb7503c851af6b74df38115e0729069b6956d309659120673205ad7e0647d063ad0e3f224320c7c8ae96e8a06c5166fcb800bf7a5ccda14afcf2db868fe16cd62ee0d81b6ebec4f714e849736b25ffde314399c6301e0bad538b7af682e508bd971bbfa86f07ffe01b8b90284ae630a7d752ed78db364ab36b4ac73cb4651f0b8542ab9d0d8b225fa28e53527912dcc6f223b20e56796964708eccc04d80d933ba70461e475e978ebffb9a26d84f2451ecedc1b25ffe3562dcf85f41cc4d956bf612ab959ffae5f2e259008a35bd4a49adb9c0f522f162d2e8f51ecd0180dd5668765177fdee6f6ae12fa495da4ff8b30d96aa9995853e3652f74e1b54af5d5507cf43eb4d0a296529743971b9a5e2d23251a392dfd4421c042313e9037fb54f2fc519eded9d265b418b9eedd4888582e32076b9c449d760ab3b5e42c2f30c7da45f53b6bfc99b21c2062327dc423f8fcbd13725bbc9063f0b1c5368fd3760731407f5e3b6c11427417f43e952b18653cdc1a07422fa9153e6fe562a927ab9d526f10607c9316ada815b870e97d0f4a8ed4f92c6747426e59a99143d2975fe2f7ce593f75cd9d2561f843f90320cfe85f01e20f1b4387a8849db749b83d52e0db7e360c384f79707cdb2e452feec9695a6e2476a1df4ca33ed09c644df804716eeb212dbf57edd07110ed58d9ed147e499d2de469e522be81c352dbb49943274bb88a8cccf406e391256297e710d307890b9d01aaad0b1f50b25b5c8dc78cab3b6478409709af548894d9d6c741e30dc6a02688cbf82c66f2d83694edfd30417603d5b52b0a28bfd47db3c491cb41d9e3d0265701cd0eb66a69a08a5cbfaa49c9ad755035c121cd29009ad979a92bb63a85ba1afa93bd205e99a62f24bfbcf9fd74edf6c14da8cecc91b695d24342e2a191fe655f1ded1398c25bb5d80b0bd5d504d7e8247afe243876dc5671f3910a40c06ff473ee3cf850367a566b113b88d8dfd8e44902bd35e23e94e3d24e5233a731bd5920d68a68d33ea6daca46f4e772d501cf3965eb247dac1ef2486b66e5cdd4f00a9e8827e1cc342f2308362f51cdf12b43ee690cab668d8524ff4336e6b9af85b794e3075a049ed3727416eca5f49b8144f3bece8d859f51dabd94f310392f7623a743943691a504d9b3e9835193dccf5b77a93c927123c6144c9dbfd8fa118f4de459ad6f5c0b3ef15fb2cf2c968639d02046fd86bac5330ac4d43f6cff5e85f5e02f2b5f464ce31bc13da6bb161ddd52e886cc3c1e435257c6e5aecdc5515a2dec2d02b44b1dce052ae9aae8e39b0e64f42ae7a109f7dad7643051d6388e2f7753b00f792911b2f43ac67848ae569bb1093619fc78ce13159955f5778a07dca94cf9fa729fb47aaf98823122bd83d7ddfa7c4cc74111f20e2008d3c335758b1f3722662172d142510e3b114d3ea641344fb34f9ad1e723f4e2cc2e6db9e9b446bf17d87cadaebff6a147df9bf5b5b5c54504951f8f94c982858872498e68645864df893e58666f8adc3b89ffa223161c3cbd3ca91b733eafaa9ced7b24b9c0b2009b25d1663c5180982c8a68b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h171bcbe8c66eff950b102bb3cf9d8b494021a7490834a808abb1aed8addd4fc7476684efa847ae5eb521633f81e8e5d1499f836cea80bb2d129645c29bec02c40f87d73a07f6e3294d5df7d8f0331c3aef2ab673069e7cfb1eac5ccbe0a89363240bb6802f6cb91076f2e48ed39bc5d46ac1070e290d6a9174c5a5c471777b2104d7ad83bdf66e45442e51e7f6986b1704b1b101eafaef6d1df4bf294eacd5fc4bcc01ed16acdb215b08d15eae5bd4daf5f30378620f266f8610901f5352ae523d44ea82339bd506bc904e4591cc81436aca89f06eb7c246cb09d799fc55de188cbb9debe512f4e017315e3b5d7b8424e28e59932b527d35a1169b95d197df39cc27ec1efb7612d4de48d639b3143991580212859741593bccc6af81169f086dd120b4bb69e53a90c95f94f893fbbbb849b37588c7d472453e0a58db2792a941ec896b0e8e8ac6d23776c6144804fdd74d2d59565c1c27ac53b8c84cbdfc8621a5810e4af497960cfe0ef848db408e5b10a628a6322169ed57f4ef9701e4124964a2438ce4eb57eb04232cb129cd09d2e2c61e33647f67e53a6c99214d299460f31776e725cdefe5ce3935160f1ee37ec54d7209686dc22ec61a279a2118ff437882b9972b8ab384108d19fef301b60ca7fc5cf7c3d89926ed0548e785e29a6dd556b856aac2a714f3aa9182094007faaeec0771686b47e73f5ccd211c325ace406334a6f2b7266cf2f1d8c0ba718b5e316d61c1c604e8c5c42f0739a90d64b97180f256f5c06fd5e369028a1bd64a96f5cfcd741108083c55d9e592ed9ca2f2e61623ddf77cdb4112f29a90ce1cd924974070fb98dcc07f470f976888485429d0e6248e17ec42a91f5fa5a1613aca5728565ba5e07c50bfdd71a6cb3a5016c2edd7b8a47261b79aabcf7115afbb9e1ab665f4563c7e410b2185b2e61d01747a62733696af19bd13441a5d83734ddf0b016e3fccc45d85a3afebf37fcb317f439f39cbb2dfddf93daafa840b8393500d20bfc11e8e7eafefb8edf5af4ff0fff2042e6f1442cfd4b3690071884f556956f9013007b8d6991de407c18e8ee5268b3488a5a1be06ec8b44b79b08cc43d87ae41e8fdac0e493cab262aa1f05debf93df1929a94b37d50dcd254ac0aaa780d4c4f8775e092ba6ad812a26d9ef23a14dfd194c9b3afa7f19ff2d8c77a3960333a6072d352a98cb6907d2f7346debe468c5779ea9cf56d199f50c23f6867ffe2b6525f48f6a2581819925597ff066b5c646796d20e7fac8f2286afc019b9907571682dee24f27fb7a8bd15894f6d7293bae8db9846bfeb71801bc8923d9f70cfc64b678835ae597ff030a14a38b6da7e0b8694271ed21054f6f46974c3096b252500208ab2806d1ee91ee68cadda65b5402efa2d21005c47f475d26fedd7ce5ed289f2aaca0df28c4db6312da99f396f534d2f97594bbc8a5ea4c223504f860d142409784fe3e8fcf00041899dfb48548b41286ba200ad89d32d3f281ab80beb55f960e645f34c9a38b914e3369b680abf5520025c2bb19707fad192b030262fdf6d8448f51181341ba0a9dac404c5e260eaae990bdc8acf0a23ed8c386cb317b8d788c88100fdc98da5733a3fa3db5f85b28271fd306899654aab612daa07e0969d840441d8c514a7d7cdf25e922304df450d40bd5c7f505df5b75c3d9dabae931c64259a77c9ace6a7ec2992067a5d4c36fd0d8dd624e0ca505a3ede2a31f7ec8a53a0ccdcd13a5fdab85f14135e5b3d37a1a262fbfc88d7964509adc8eb60dc76cd0787d7a0161ccf71d2608fbcbdd2ab5a25871912c5d60fc0a593fe1aba9952eb1aca885959993da9be648a8afd6a42ac595dbc7d2b5698e5d77c5bac0c047350c45e3d614da40b38e6477dc248bddc4706a69a521caf508f072e814f72d3f96fc507e54712af5c834710db7fc40f747a9489279d167a5556e3e6deca6fe8fdb41deda2bf5d08dd3543fc6a58e290fb5d2eae70d2e265258289d8a8dce6028e6800602c0b48e191fa7eb9f50fbcbd6da2cad30cb2491aeee41dc6fa87d015207e3daeece31e08d72caf65f18d8cdf35e53bd48d57b86c0d18775c72d05bf93d2b40a22a3cd8eabf578b3e092052e377fef8d6d2a6fd258df5ce6d7db6dd9e73ea61ada3097bbb13ae1dd50491257034a9405bb631d869f1fbf0853fcbe8ab98e9e9ca5c6f1ec4ca5889157dc3a5fb86fab970021dd145c1132482928138db741b55bf4f828619a2b393747411d11c5d706edfd1b590df7ee0d297eff75292f9c64a85356a664754cf9424f8f306aed36bc9d25abf566478e02c296fb24d3e575a64712256a1f64da7d480dcec7023d7880b24a388572c1abb33b9d27f5d6e75ef5f2299623bb785f36dd40f70f194df219a67b95907eefecfe1bdab791da243a6ffe0a5c3bd8062bc5c509ac4543f23ffb0948fd9c375236f2fe8d5afeec246586c1ba2588fd5fc43e5e25e65a97a21608c6f391e6ff97dd6ddd8ddca8c4f8bd694fe524858be569331c280c301f8a2610a2f93f1be6faa20b53c611fa2c050e5f08e2444966045c0646a66165b5a4925501f6ed491e2c9a5ea10722e3c2b450544be19516764612b9531588f2d9451f431332f3c87f0fec83a4954ff940960230f5ae0d6b0de2245791cdcee01e382bc9f8fdc9b48287070b3b92afb3fee353d9219b67ec9be2e7c7a3c0fe86d6c0311c920cd363621f40eccdf3f564f3a702edcc34d18eaae607c8bf0ccfd2afa8a35b09d4de801495beb5b29e25d0092b293940abadfddcf828222aeb4bc9cb7f4a56cf8a4a3b6d813936ee7dd8277390be5ec0e32cb46dc34be1b97120013b3e8363d82df148d67014c9110def5abe9dd12a1fda29cb527c48183b7945e144ed5d3006c0e7d92dc4dc7affc8fa6ef5d72876c474efbee41d8a5a77dd49aef683726ac9c8563a338496f23286921a7ef413996b061f67fb94e427664495b624e96f972bb1577db49ea6a6f41700b4a5285fa52a9cbf14e0ecbca61812c646eeb654c0274f0d6cbe2059311da0aa3bb2dc5928ceb4fe124a59c734e0f6239a33d259d2435d69112f36dab5f78b88de0af82428e5eba52a932fa3cb8d2d8946c9967da3182e68a335cb3e0deca1ecc778202d39de5b5e03c5b9867d80c509b7bbf7f45a00f7071e85361d256a613e592dd9142214bf35cc7870e7d80614861b07798b784f78241b92efc67259557fb8a72892c4bb7928832ad117dfdcb898dcb8946cd7921025bc5f47418117da5d43ed68e50f6b09f8c4576993858e1afc660d258d57b273900efbc099804303c5fa08ebea31b71b228735150fc12729d4254ae0b041081338c38e0ea654bfce9c10e8014b6c2568ea8c8091999d63c16270574ac54bae2887cd3db39abda492ff15811eaf67339b3fb542c4700b4554038068e2ff3824c56363b56722734decfca750bdd6be7b7b3fc800cd4473750efb7c6996233398ac213b69a504040d0006e687a0a6fe1db58db057f09e5b229cbfe390b7c04fe94fc833e8ef9774f8c0133c9a5100468508db61833d4c4f3913d5681a1007ae421dea4b8ade8b5e363fe017984bb52b21eeadc6f98637d2c9195e7b8edef453d1d5822b21cbeb8be7898e02787dd0730da9fa655154182ed559dafc979cf7433cb5fb9ffc81e5ba9883c3c91fa7ce7047f7418e3fcaeb749c43c753c27992d92f8e5d6a4e2da03e3ad346b9c14b7807857002861742cc02f68d43e647fb085846f17afdba52ec4b1f5cad9cafa3d1555cf670af05eb2e635433608a96093b1a7df03692c14286269da49b60495dca21d0446a85294f46f0531289503bdbe6801d8a214c5018416209d5c5227e6257c76fe3e62676a17ad896d959ab3af8110ae0584898050f9b83baacf3d5ae97909d1fcfa129f21052c02b1dfc7726b505d2518ebbd1c1f60ef3039b651b0a012217bca038fd144ed2cea6e77e2caaef0c537a336e22f6b4712d148f305c98ed0ad46529bd96fc813e95e75dcc38e981f83f6ade4e17e9f07b81bf97c387a9796d15fa04494635e97268f08984cd9879a9d8878d3ae55fc57c1aafcd937f985f7bd295332811364fe6ca1794d0b9be72dff00a599b139a0419ee767b10c8095fbe6021552316a4f4279bf120d2c60aab4d8fe765c09d35a5aa0666bbb0f83492d697a61bc4b25cdbe2d71782a1a0b7250b5e5addd3ba03bac6aaf2608d743604e7e24c687523ba1c9fee275fa61d00641aa1e95860f49ccbd650a8c92c33d3cc336833515c38750e3e5334303a27a7a942f83eef1bbbd30b4663d166310c87c09ce68ee1cbd95db9aea3c3cdb924a4d728b98b5cecab2ff688466b810451037d1c0df280b977c9d9f3c63aef6632e9de80e63c6ff9bf6f551aa0d36dbac584379b0608ce893fb1cd432be31136f70506024f7ad48dc8d54ce364b333326011c7c85d50e6b2ed9a9b819b1f8df966f797ea63463e9a661282097948b87c1a3203492e0bfacb892eaaf16a1504d7e660c994137c43eb4be13050be76925d49e7aa909d657cb4c89cc3b006200f3bcc39506ab8af7ae72d97ec711cf5cb3af730db6c8753b688004453bc983aea62d621578dc32f701a43e324392e4e642f33f952668cd8b055473e6014ee0d11616e68fb3b4cae44e05235587ef87bb6b467bcb86f6aca91712eeb200c036e84319ec26dc51c8fd0ffb43d388f90c2b7c8d94677d6357f6cdb7a9368a22fca5317fcd97ebf5d766be3ad16b13b752bc8fe24198c02b1d4ff4df2fe2d5a308c11501b6b84a8df367045fbc9dabe9b6f13eaa237816d9bf6fa1b011f715617c684550b5ccba2400a0af99700a37e3de136f9b0152600deb793b1272928b10376ec3123fc5874327844411ab77e1c354ad08f692ef3929dde953c09de1523a85412b856d643e53b7dc7cf20a4b2b9bc6c4a323f5b897493878f9398de7291581e4452e199eb2709552ec06652d0d8270648a1542bca4c3242860f41f5163839ff4e83f2cfdd0003f8b3391f5849c1f39a82700e3ebf3bf2a91239a54c7109660fb3b73597f19a2b049f51511892f110108edaa122912f6a2774301f961e86f37198253a7665eb6da893ddcccca602e640dce8d5bc81ab4d7f1847fcd4f75d8728a29ee81afaf51b8eee48595cde40ac7923211de48713422ece09fbbbc09cf310ffe2b8e024b539085e60b6cbfa9e80b587ec393bc9058c90b8d15e7bb0e6e51994cce5ff37e348abacc7baf78568568b9a98c8d3f280a57b22bc0270601df06cf123451a1e20676e6a064bed2ada155ac586a5d0a03933da2a1230d926972b733da23ed33639723797495a7828f0f254c803c81900f9aad2c81945eaa804172defd0a4cc67f6c04dd6b29321bf97a0fa74e9dad86f565ef07fb60e679a1214a691cbb293a7a3e79e95791a47f534bc63d9609d6de71bd970d390b5d4d75759df1a67f648cb43458e42d24cb16a19cdad9e95b448;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf95a74f80f04ca527f836408b66b879e96ed68d51c45728ff768fdeebb0c57bca072fb291f2a5b727b2fd084e7c4687e2dbbc9c6cb2877bd53a60c08e071cd8ce630a74a28d25b1a4ec845bbdf1452eb0a4957ce651d153ae586d0f640839c53967908a4c3cef1f3e8ce82b35d8245baf00507d3980be1e24d33ee726af1ab267474b438c37fed3e300ba69d8e50334a0c05bf3e6902872b66f391d8a47dac7b53f22b30cec33de3a3b0fec4cb20573b6fc85212c3bcebba00f5c02d80fd985b9b003cdfb68a3277ac6531f452b16f098562ec87380528db7ab3c04dc7dbdabb17bcb92665e4ef9d9263c9ed697e7163cf81194c8a8b44046d28bbbc3d1c198cf837c45ec46f937b3fbd31225d4082d1130ae8c891f1032fe869555a4505f7303508f6bdc49d2569df9253e824b767014d333c6dce2d86eb9db62b85c90e4bf6a9dcf5e1757f344fe5cf38359dfc3fcc1ea06ea7aeeaeda7242b04a5c1d1da2ed7a1eca7543891cfd55a8773c3c431485a65e00e87b9210aef1fa8f9b87630b033bdfe1aacdce3a010825be6b5c6e472ae0bc997015d63b42869deab12431f4fe899c3098abfb693e7a11049953bb5d62863afb9bde32b1ac2ba4d5e1f1d8978d9f32f636186d3d3a7abaea83bb0c3a2ca6aa8893b86041c907cd03c26554ef60627d02c0c7b13eb91dd5ad9a685be24ae20ccf2426595006495eebfe607113a1d1eaa526fdf0c88a77861f9a5dc8e844e521ce20fc5c41086cb144a515b2a44d0140c5db91f39814397f3be6b3689d30aac522ba1ee242a18cbb017e9f332d056b60bc4f90d067aa885bea35636c95dc58344706b5efb2373e55cb1ca94a8d6b5b30cfee8f7f96cdabded0379d391865baaa5fb6c9bd0c78ed5d94e389ac73cdfbfa4c21dbca859ed4efa402fa0e539154c3c23f806e4b1c2c6a92477759249223630f2b240f0600a3b8d2efec87590107f3c7a8fefbf0611311258b4349cc6d8fc580603dbf62b5a2c7fcd8a66cf4f72fcbf22023ffa5f0ff0093b7c0dde13aef8e44945ff82514480fcb5290e522b80987d2adf6ceafeb6947fb80f9bbf8c50ed5a2ff0fded7b2b4f80ef9fb169691678e20613361c05079aa523ac57533e7dfccfe7439071511aaf8d6ec8c36de91e1295832ad62c8fca0886b87a15c83566109319396da0947f4b3b141cc1a049e8cc947b781db096277ad5461ff0178a458c457e0de3f2f269397e1656c2ca936203cf7f3499b025ba5fbfce05e40fc22926338e692f285e0d82d4246cf0a542e20b5fa70b897f3e3f738e7b3eee3b4ef50360ecb0341e3b33401a5613a971ba681642ebdb513c29b562dca1aff26622f4012c3a39743a4d306d99060cae471a97ac41eac03760702b556daf26703e2a0a2fc3f2765dd312a6ae8085684b92d15ee943a063027987cc00777c7aa7a5c7a4db3e801d84be06037a714d9bca5b12d1ad67e03037ce8f8c9669dd924968d3deb15ae5ed8b5620e8fe6cc0b5b72547b083b0355b0ef7d6642709098c8f02e52477b5da3f521794e7d49a8f298dde723cfa3ea1e64bfb64745b53016752c75834c2317505a3a45c677ae8dffa29ef02f6a350284bd1cdec6996b25f77975a9aeecf0bb84db966f2583b3766b6f149960a6cfafd8c4c7514c665471d74a624a129c040bb250afc653e41009e2a18549e986748f4ce8f149f46bf2cd3e8e0c971b013bc16a0ab68541e32e3816149cd6220aa2756fea43c050d4ed24ff65619e2cdd4483013adacddb38efff5a3c0236886e1677e83ae171fc95d7d8b0252a6d000245d8a5b9f7734ea968bb7f149768cd114a46c9ba2a4d6e403fb28e653de7bbf56ba35072eb74c154bb21d3de75ff8242b1972b1e8eb98b4df86af107d278f5126c5d32108aa4f022bb412195c9f26ba764c6dedabc686f5c495664a2d283169ca663976ce4e7b584e16304aef9ca634ae46eb7ca534b3be02e4d99c3760879c4915db8de562241687081ca97ff15e081e811f9942e7279c891d393a7b532ecc4b552c92ce67d59a2f1c8582e168c87bfd0e46619210d26c6787258db73b6bc0d2da50062c9909a4af1304206f948e4c8e66ba8413e7e5fbd6b4a977aa682842d1908ff8e08da0dcc6154f34e91223c1c4d62be2d9fcbd4a41f2a8c2c06fe3ec76961409fa5a1e0083d3698c81aca6bbdc7cfa523aadfccffcfe7ada267ee8b913ec38820bd7039925250bc1554eb36dca5dcc02944643f18e90f9836aa37f96903338b244e637e08912cf5876d112e46cc7f5773dd6a502a220a7156538e6b8ed672402a342d413643331fd5a41b59b6f18156afdae068ce9b68a5164a3fc9cf7e5b56451bf247fcf23475a8740bd00af8549fcb8f9feba28e12f5ca8a608c90fe7775c52180912014a0880ba077675b77fc3c7af1e2dad2ea074cbc8e994ad868439db48f6fdc8e139a8d510faf4dc22fc15ec5a5cb5f80c326cf9411b6255c4b78a88ad401821c7490c61c22af76991e94c14b3c368568e59d4df8e2e3d71c2e603c61103e2baecd84287480bfee14b671f143bd8d37cf989ae0d30518bdf2dcd687f03e7076fbb98cc526e4cceabd5e1883c81153541a776f5bbbdda0d711658b5d89181f32b3472ce075add0850fb396b8bcf193629432caad2825b09ff07346d3a6d3f399840bd02feb34f62bbc3c5c6690920fb355c5dddff3aac6bfd2ee7cc8935a21dd6fa60881893b7c5bf2d2deff8d9a2c57e0deaf32857e116e456429bcc1aa1f1ae0c1d899e778d94421569339690f29a0a5b8d82ae18a30c4038a76d5b22d1977efbc8153013105a34943f6dbe5d7043b52ce29ecb85e600f02c989b317dc7aa92d5c5849d05391671632ec6d6ac3c054c8e0c1f3aadeb8afc5f35ed06292cd4cc19c965e735b6543f39626719519730eba054970370dc5d986e65314d97b8290f4777546545a686198817c9acceb1a0d7e62abc29d8db8b2a05548546d2a9bf3a7e9268239e21758a97d4e407d5838cf2d0f3b294134d9b902111f3bbaa8d1288abea87fd469f8aa3479ef4a0f308ad157fc3518263240468b825d8b76b0871e3e9417483f001965a79f74204d0100a2699a31fdc7d0731c42be1d132a1a29452adc7f774ac31bf0dd7162b45112aeb5fe1ea155564c4b8338f7dc4fcbdc5cf7c60ca3065aae3e15ac0aaf155a7b36e4f41dffca78f8aef4365708b98408441e28bd7b6f531125fe2da1c9b1240b6d9789b3469f72570260203229b1be3f67fbcf30e31bc9e7495f57089d62a38799a255ea6149deb6b7810805b0f7240f4d9b2a182ff8f94df209df59b47a48f6e2186a0685e77e88179b2391be7a7784b4f59c94a1e46badd0436f008a5df23d232aa2008fa0755d4b5d275d7989401101d5acbff9c525ea4b5add12cf5f14628399f94695c79a139088068dfe63a62c0328230c60a3c576e23368272d83175fb0bfdbf5b892509126556962f7566c84d71903223a88b05333af195654278578355e3e1e068d3866e521a79e9f2e2e76743b5253a1c444f9a36fb193fb1139be263b860886b0e13ae4ee13e62e32feb309e806f1276229564c82f6d09d359b75d1da6d4e1afc4eff7548b16e39b1a1d197c4bd2465cb01c03d3d0d6cdaf87671e6f0155f0fcdecd05c00c0533b48efcb0a3d0e5d866dffeed1568448b2f6ee64a8a127c6e1f6ba9f2e10aef746f487338353e39fa508ba7b815dd05f5053f708402a17ef77ab2bca16347c3777c0584d61b68b882c8c41ba0d82f4735674ee89009704c302fc711a759b9da386365745178bc4595e7b5e2d8de09402cef4277d5a55e0e6b1b98295e1a97cf733be93fd407029384a8539a9c407610995fdbde95b15ce85b7ccf55f6a6aab3ff32812b58cdf30c185bb8e8642dbd0a6cf3ee45ec5f3d3726323587252e0e16d5c38d8df6915ee7828bdcefe76ad9bd6d9832db640876319efcfb2889070cf267e4dc98d873265cd25bfbf4dc0df4551f24c9b5605fff3566c7d0f6a18067311ec2a12d72e97811005c06ecf31df5ac6424d90ad98b222b6c75fef08778acce20ceca4971e349e3cc3d59eae70f0ee16c3f501b81f840d2ba07c3d3c929733d54c66025070e53b8626f96f998dc2cd358c4715ab9bf4b8ec5ad05016b9c92c334b56b7e4502faf74e9dadc420b1dbfe6912ec787c5a7d95b2f64f2f77a8288d6e5a4253e96ecaf13017834f91b2883d1cafe11716cb4a765a10dbe6ca5097b28d31f0d21d06a3e3fba930f7082302a31897dc87230eba075d2b9a718d5eec5ecee96d00c68988537dc2c083403f067a1fe7bd785110271a6fc0240897e92c5230d5aeee6c7da9980fff0c50d0b077b09572436b277a7859e70cbd1e59513a3bac8bc34e2c9daaf95c393714f4d3e6457fd302563db0a4f0ce1b1da615be1b9c2403865830d54c7f66a4ce9323145b818c6b80498f291bb7cd41cfa9c4cb08ac1f2533fabf61fa0228e3d75b82d7516fe199b45a4561999e51b92e8008df05bca209795f728e93f685dd59d26ba2ec0b171d36dfc4d22d4c7d3135821cda53a2cc3bcff6a92488d7610401e29fb89019514f508436682510b1eba87f711cd345dd8ee4412b5a4a2330c8c61d45e079cc1e19dbbdb95fc1fd1dab2cb9242f2877f4b9fbe7f5ff972a0d15cfc32321abf35a38d0644db2774ae400a63f69c68ca83a0fc755350ce3b97cc209a20d0e77f86f2aefa20ead02e029ae27b65ed903a6a7addb696a6336d97b1ebacf137001a2fe8837c4939cc37382d9c9b51da81257e53614496a33462caa578400a845c474a7f09cd0b5f4b40d112c49f5031dcb2d0b5d1b540c7272a7902220983bac9fb151e5591bd30917d3545d89143a1f0adef1bcb96dabebcd93de604ae7ce7b4ae0f41a7a686bab9245dd585e8b47ccb66d366f2b8d3e4c43040ac1e32d8c3466dec9248f94e0ae7374fbff9980dadd9b56f0407823a449208f89828f7eb95db5483459d8706e902834351a8789ef628338f926f0ea1d2ad89302d9a70b78ef0b2adca708c1778e90e64271ac75732fb7471253cf8e03ac4e52e41ce872e9f328b8a4636d1bf2035ab650d7ff0b0af5123ce2497a53c4ca0eec4dc0129d34e51abc2cf9523b7e46c73553f5e674b72b9137c6b5904e2f187d72da779d9e0d28f88cbd79435a00d41abd76270e23f131113d455738873c1bb7307676f2fc318cd778ffaeee0dc2eccc06567dfc9cafb52b93dd9abc1df07d3387699ec313bf90211bd4fb994f40099f6647ff3edc4119bce5e38d1819e208057908720a1adc32d78944f51f6943a697ca33f4b740bd83c4e4d9b5fa56355fe6e479647a96beb82cd2cf7f8bd7894f7e4a45f4abd5289cb40f33b1e406a3d2447523c5c7e4c8d8339c437ea03f916d2d035e30ab0f8e73436f0750ba71733053e26742fa18266dae20c966f2fd0920aeb049628abadc9f143be8d783332e99c19f2ac3678cbe3c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha64d33af30e826c4f2e665e10302ab806662e59c9a04027f0e78db773b29c2b12c2c6496a6eacd99a5136d3c3ac1813a37107510a76a3d000abdfc62eb98476e361f2b1fe36db9e181ee6c50e457dfe387d90dbb6c03d388cbb610f1b1de5134faebdf1b39326c2d81d3e134afb81e57131fb0d2b96071bc105d0c8e5d5a9b537c71a653321b9994f5c0df1f5a0e3b2fb8a0cf65784bba44b86b0e86287e9c5415334940e397f57e00617d816e855f10caa47da1bd1cb7179017ac22a0fb2f8765d20a94d9344aba493e7d3be98948c0e1dffe1cdb00caabf1da8942e4069582924babbf94186c03003da1362f2a3045784c2ba2c73d9939e752958d4cc82f495875f6b7b836e6110d5b95f4aabab4f5904d1bad40254c074514cab72ca0562fee4b986cda49a0daceb45dd3750fb04d1a8d5a0b5564b9cb6bbd6265f3aaa735e9f42b8fccc55265958c80b0bd4d5d37656435a0710d6f901a73b8b16a7e2e7018dfbfd3bf0f2aea76ffed1aa49e1b1f60d4f1440ab54154fe576cb1f522fc155bd25af8b89a0170d9f2a34f8f6e47914b6ef98e11c2697e345039fddd1703e32bbc78b8c6a5db95d1c80888deae0700aa341555381c8077b2b5e56612311234d9aebf2a229dc6af18f80be0ed63bddc54f1042549a0c43cbaa9519c464003e82a0355859bd478041d0596a1d22071477d48daf296cf6e89469a59a02d7792c16121634ebb5a805e31cf5b6ed84698f7187ac031dc7eb3c1de0cd657323cc6690af94adb3103663fc181002ea0dab42186c47ca0c1b4a0c4d774cf72ef8b15e2d79cc1db86b623894d2aaafa0403f21c1094ca6c00ad1a2936aa540743fe30d00c3c3568e0c3dc2ab7a5f71bebe1eac2882d383d3638513726d420d14d530e173732bb53fee3408bc6fcbe114be562a6f6599ff1019aee59014b6c8bb2d1ba3deef9ff1ca39d9554ac1efb5a46276846e61c1d4bb79c492bda688acaef08301fc159447f4439374296a7d9b8f146fd6c5a199b23104f2bff40619f77abe16c96f8a23874d89855cbd5cc510b6fd82ced2705088309a926afa18b7914f0f7376dc22683cae452898e4c6e13035a1c15e432d134d655edc8ab48e27000df2b041355fd970d3598676deb45c8fab7ca4ad672d37611481db7e03eb06ac1da192b53a99449ebf8fafc24bd72609c92abf4af46bd4d8772a06a4eda217497566e30b62f80f727acb47c4be777c19f156fc68731fdca46fc848d27e02300b319111888968cc82fb91c9f3a9f4bca3eb0aafb1dacb97738a6bd559f3cce0f6a527e3fa7c93d24fc74cde53d5fda3d2971ecca50b1b7d2813da95be8cb6cca34b24226ca3991f76d44e9b92466c67e5cd76503ec6c743abffae80475da90ee6b4b220bf8852c183a83839f5acca98b770ccb317b5c5774deab635510855546e3912e7059d61af2fe29a198d160f415e641b4a46318d8009fa673d1bfeecd2a642e8cc16612a17d7fd9a579f60cc289c8ccf74904c1931f545f9b3a948dbafdce90acd09a20c231a3daf57274d0c4b591da53d751186f1667e66d51c27eeea53bb25849f0bf9ebdc4002b15c842d1f044c0089ff48be13a2430f9c00800f14481f47793b9e744efd759f7d446a7b8bab8f6531edadf8be2667334aa99ae7465f6db14e71f63dcc42de5d47269148ca4ab658c8a64863691517310f741432dd6f52aeabf96e1aebf5b8764c9bb936e96c45ec821b17e67f6df42f222e6ca38a794c3139f57b939189ca5a0b5dc1ece177e4ac00d71daabac5c8595bd403026784ef508c081d9ad9fced175e2d020f9739eed897f9c284b3e08b5da5a5fe87098a7ae339612b61908a8cf4be10c6d97cba4b59bde46c6bebb882f4271279e4d4c4b3784872795976cf4765b0c4dc41c45568a53c7969265fbc80a7509ceed8ce7c9e3bd09d80ff1196c6c80b7f3f2155318651057e676abcb53842961d272aa59dadfe749e0957af2373bd071c2a86763b9f862b96a0cfda9d6d7b2283af534c642e6e81e4c518044d9440b05f52880577e0fb9bfa193cd19ea50ce8a3a0f2ce48e239486213352c1b610948e2d7e495e9a37c2a512aef915353aef4c6139df241a8fedaa7317ae706ada9807b483b18727d10f9c21b5e89650655a0e86fbfb6084fce977825aefc7291afd4301746072f9489be95901d0e24f503f650229886b2233c5323baf7a1c7ace34748dbe23d6ac10063c6395376e163cf22f51560a0485caafa5632aae3ae0707d02f864f3834124240663e9a038c763e0da4ee646724cd471e72f5da3c7dba3507458ae2060cea42680c77d9dec5dff34e0fc0b99037458c28d7b517f2531ba4041d46f02cff3d83baa697b450a73e0f5cf33b97d7f0eb354856ef182830794a665951dbc86f127b139e237afa772c794159941620928980afa388b82a42f0ce49d343713493c0e7dff3f992d0b3bae197555ce0a0177422836034a850d78a3dbd648d56ed6381380abe0df9d0c0e636cd99a9d256df21a181f08f15adc015759741b44d1ab8412c11b455e12f9f75b5bc4c8f33f6a89c9159350f4f522efe0518c5b76107be25bb46ab48dbf3838a02de692df6021e9e1c40151bb10d123d3b972e5ce76408785488db23153180587611da15e7fb10a09a28398846e5bc8f6f5692d9c54310b23aad23ddefa8921a9ed6e632e5de28a46b77ed2ddadca60340fbbd88a925646db57d14231d1bb75d3bf1fad2e9d8888ff31e27534c5b69a4f08dc85df1811e77bebb246add798fdf8f1c37986c5b8039368efe3e6866dd3c876d018ab15ef593752ba3581fcfea843db4e6340e5885f6e18a2a3076154194216881e0f1d80ba7efa8df75e3b125df0973716e1c32292c4e2a62d107c3267ae2c2ea53df669b2b9c2261156167806ac687e6a167abacc77bf79814f914ef5fdcfe0f18656dfb158b25f7928250b29afb4a286fb4402a9576c653560d21fad1c064bfe6df611f6f8c1dd92981ea0c422fee7380b175aefe3873982693110e23ce76220dac6a1427205bfa13e27e5b370e21a5923a2bb0f7b1d50fdc748c1219ddbc56ef0984bf6f5b41b93781116f78d5370574288a0af5ae1c5810d66d366c0474294deba31bc30946a3cf3b879bb2640cb99e045e59895ebbc857be21b95238c7acbdc3035d7528c6c429c4cf753de1a774fcfb5e879b504cf6c9bf30e081e6f69d3eca98cbee9ea175e1089e872ee5c58f61242c42a2a9d6c4113a9d4d460ba0159187d8dbac5e69a591973dc5629e3871610af3c9f92f4f4b9bba92698ce71caa08264d6f82385762aac70f625b8d5f656e41a46a33b6cd29c779930408be6c6e0bda1f461805213791984deab4032dccb67126ec8fb6e0e5fde6d49695c77b1d876c4eb03d1e2db9b940d394ad3216cf4766f269d00d22b0c680a0ceeb8cbce33196614d1ffcb07f9d4d3cc9044bc0e558d01cf6dd2f9bd7088a686d3e3530c45aa2ac83f9c6b96569699e354a2090931bf292a184f0502566b6d7c18a3de0a273775c2efd631a375f58e907853d836b980c34d78e4a3f8c51c247916ca3ae9fb9619495f797d12d131b6e7590b899f5748dba46e7a6816c0dde88d59a22825c3a4818fc0484e81e9c5a3ab1b426d895676a58d953c0d40d386c488642bae9ce8a1e3647544263195804eeab94ba9062b9ca49d07b21ef7054dee6c9fb88d31a895cbc516cc74ec8c49f6cbeda2dd162378ee145de57ce435cb40bf950c3ac9599f08e1f3824a0d723ef86c2bd8cf456e2500ff618e0405d8841cf390372eaa10a48d9b67e0449418e344acc0a1c19b9c2d8f0317263813b98e3ed9bc8895102841d0dc10c700f5f9b5862081778bc0b43019fb5c104d635a962286b83a5bde693d2afcb83997b2adae54992e928fef7fc914a3480032187f5dcacadb76d36dc34a24f4e9a30818582c019dd608bfcbff29f8997fc02b6dfb421712209035029e60d1acc842a17c7cfe5b5787d6ed0a1be046525569dbf73c5a6411b5a2571286e04d2c7fd6feaedb881daebf748d3ff0be0b23f9a853aa6216be7bb67bc8a3544a1e8d765670f38b60b6a8ec9ec1585f2aa721e6d0ddc5d9e2c86305b58c287955f33308aaac3905d234b95c9b9d86c7ab01e580471c0a411b8b9ec228256d0091d0baa9c351391aeba763e01fd3c13e51b9edb786b421e371e3046826459360ca6d6b77d6e37bcaffbdd4c8ca470f63badad5dd8514cabe008ae961ee9386a0607cdacdd789af50462b5a44485e38c3e386cc82911c8581d88afaeeca29ad04ccce97975861e033d656c503b6958cf8adbcfdfebb412e7f629329e95512ea8301de20861726cbcaa8e0f63ef77db433472c9d10eff38677bd42a1b1a54ef2858e217f893ed620283325bd1e9ecf479520044fc432167745c12f02da3371d29a1a44bf2e1b16758c42f8db1abfa542483fbb9aa7843c7b9c176d008a170eb6b043916a67c0075688a3e28277f2894acc44b7926d3a483b95d9237f1c52784a516a51efd5e16176676ad45c9976e1d97e0e9a31f67ad8b081fcc94d9c8bbafeeef93a5a5c84439c02a4814a6501e04e9de73d640995e938a099075631cbf6adc2de80a1c4b4203428668b8cdffc0f9999737ad8c2fab522d4e23d2b2a2982165cf993f15ee7194ff8a2e5257b5e7ee2cd0ed8186df32e4b0569c5ae2476b3cf995073217d988af2e1baf447c3655141168d5be54b63c2fcffc21f818adc23a59cd7e0a7a44d4d9fbce7cb2f43d3f6f41131f93c8657906b84f5b1eae2750690a542ebe3d910581e0367455f068d5959fbe1d6f8c96b9b46a0180919b0f13ed551f2f0c59be9ff7d66c2d3877e4838ecd56858a896e06afa49b478fd93320e2b2aea82d872ccdf2193d950ae6c3241cf2e8501768e283f6f43f395fcbc102d3d005fda92ccf973f4a64a5f54111a294dd1f9efec8896936ce8d898c556c78906c32d51a7845a93b084c9d75e7612cf291223ba52b4215f4981b553467a5329a1a3bfdbe361661f581469bd8bfdb16c74900679a9560a276cec205d26aa77eb12118e9ef3e1270382f39230c73d92f9981a9e3170ba87964b31c4b0808f4dd8e4627ae36411b1df7ae5f192e1ebf928aeedfd2a270ec63c0dd3701c98643e40c2cffdac7cc187a0cbae905c500fb61c0446dfee928649b051e09e49e878dbd204b350ccd25f8b00f336a90a89e831c75872b7681206f64f05a492f7bb6d3f382cfec016455777860f3922f689d495ba357ba2ca38726b3fc3aac33457d1020085d8d5542c0a1f6566c04f9c18ca2fd69f58e6a3be0f94f9e00969c3dc8cde0126546402e0f52ef366fa7cf82001c6d6c85bb4c8b1394388258c499a55e240b2fdbc83b337adf101a0e37e8d19052465a96b9752cf7c9d4635b17846e534e083aa82faead117f34d5db98c09245fbf52cb0393ef0a3c9fe59b825227f51dffdade8f6a1a7da5c5d3cacb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h985ea5f9f41d68c2d30598ea0ba091411cc377d0d9ff4b3200a64257bed1a012a75f7d7c8cffd13fa84a8c5f10e9a9df680265492e73805acd7031eb06e973983a2519b1c469cd4c06774b452476f590cf080e36607ba41eb2cce82979bf2979dca590f6f33ebe69b5393f150acbc5c76e1a0d09f4e8edfacfb433c5da884390e7d607f28c29221ee58e5511be0ff767fea46cc463aac6efb788f1c618bcf953acae5d447450de5b01980bdf6afe093f6c127d39cea53199fa6faa13df830bf2f0e52fdf7a8bf0af5d670a84c1d695115fb6a89b26391a104204d71e5203dc08ab45a4825e641bb6527c224b1142e7b8e4a92600c8d2db082eb68f8cfff4b3e698feae6833e70528bc991264cb3295a9d9184addbdf5ced02801e6ec06a032983e09bd684830b50343f531e51b4f5c0c87cc2de00f47e2360fcf75138b7f3335a0842e6498e240ce8a2f222403fc29030c44989ff0f5ed8640e2c0d441d1b21728efaef70970a61b0e1da49760307f1eb0f72c27c60ecf51625c01c9545846340d88e776a6cd4ada84525a31648bdfe5a5f09ca0de4e0b5ccd489e7b6b6b3799d867280122cc161163ae9c8cfbe7e1d21444e60d2aed08729f91f727ef0d372735ece08e01852a97a9d002743f19266f53d8968182f2e3ef14ce1c3593f5d31e793ef33944e681f720cd36b3a0d7714b102168fdc1439215cd087a29a735e16d411fb319141d1f1a80eb06f2124da27e5c3d7c56e4926ef6a266a4492d959f72b88e181e94f8345b4b88271370452df1aceeb7709b4487f7b7100fafe6634df31dd11f293c34dae53c6f0614869df9f6361f329e1e0ff9e657ff8bddacd8969a15ea71e960a8a691b40132267416f85b5674443240103cedc6ed42a90ae33e7dfee4059f11418e0487e4c8b43d05ad869674c9aaebf1f6fd011432dba2d0a6f0351e8413796e5c7bf034708608f9dfebc2dc90807409063539d3a7e35fb0a69694b8fdddbbcde8fb6a8f345708eebc9a1af8fafd97b2588a65c9cee70153e9ce7317f47d84b8892727b7f4f095c3ee22c238ff566deb1d9414c2d0f64d921420f3a124356e518daefd95f9c94be8a8ac9f8a3347c4f9a037280db62c9914d85fede63072ab5a948949f59cbf96caa62feda9e7846bb7104c5e87d67f0c7903e39d2c44ed49a97b4d33bdcdbcea95242f978f48e4f91608e8bd9325237026deee8a2f023867da8e6251515e14254c4db391571fe26857e8a0a6d8aed3aa6428274bde2e0754edd56bfff38e97bc04df67e9b8e258cc3f6c3c09a7f2c7591c012d01f5b8e72650c569b9c09d74d051c89fd8f40ca0e6438c5a5c3e609e1a46f0635fdc2abb7bb59d7b33fe89112b2c613bbee4cbbae773285efbd7d3881ac8cb6726fdb9f8dbca90b93f8fbad5456d4e41853344524a7d29584aca93dcb42bdc1c42c95aa0ffea0f15726f3b370a287a777924568dd2e2046a9341f7329d737d69e547c384c7aa020838e1dbdc20e8cf0cbca42f7278c44e598cc8b7a2a1c2cfb16e2b728c5f71532fee291eb98239a504cd53ee71c0925655be750d68e6aead8344b117a17d0aafc5ce784d7e4b8e2950d446ba9ca9632d18d7b15c1d5768bee5a3eb90c8b9113c27e714b086aa949b65ae4b71d16b2f38ef7bc8d8efeae3b8c5c209abb8cfccf4bf74eb7ee41c04a2f6ce240c7bb61a36507cb968a55394e9b9fa8f33da7e3a339289e4425fd4eeda560657b04b4d5a48d0bf46e956527fc0bdc1fd604a0ca5d0bba5f81c84d76511e35d556db05b729ede1b89a3d6ace18df57f88e2eb2c746e45546f353635abfa936f494f2d1eb781424aa13917ef2526e99ef1b26aef325b3930da9c47d0e33211ab66a3869a791e6d028e65875d520bf7549679a152b89b83f9b7eafda6db9d02f4c7e0160a9301d17bc434c69aed0984a3d4fe95d40f124376d6ee6e493cc52ec3ad6b3aa9735646307d4489850af93ab5e52915f82b999e2030a878e20673b91a4697e33b512adf4fdf461fe49f6f4bfd3f123f716e0162e92c513aaf226fdf6ebfecd997db25b0db128fa653da714c0cf9a1044150549b5cad53994734834cd807da2fc061504f7d9d3a8ebf1b7f88bd9ae29e28f93e8782a34db7c922d9e2f4db7a029610d0e3e73897dccbbd27560e39368560723a32d378fc27f830ffc60713760465f9bb53f1aeea124131d1066d6b234a0f79d7da56ddb70ccf1104f3f430bf4e76cb6f81d0a7d87bb8c69dcd0913f8a3fb07c1e41e7cc26cebbea75eb6fa9f2d9f3a4f2f8b2e1e4975f89cd5f9ea7f1844cc7f69ef961bf70429ac7aa4f2af89ae7f3d00e3d36f86b9c62ac5d74497425f39b7aded95eb43234035cccf02f1a1ec20033ba6bb2dfa021b19dd57b65f3a7905d8b8f73a99147d14e4ea244ae2a2f060d1cd43fd1ed5e47e1df011872b6a2f86e7bb78086aa156243590c134a8e0144726d472138a1c21464aff017bbceed2e5c548ddc7d2a410e26ac673d46df66ec0f6d5cb03298dd3debdb7a71303a04b265c03dd04774027fd7aa9958b1acc985586d85db55e754a81b244666a1704ff64e4c25382729bd96fea1bf7b93c2d280e2ea03ee004871b7b8ee24fa2c9117c95785a95c63e7c26c25fd4e3b1cb16f80eb60d192a77957aeb44397e1a53204a6541913e1a48ae3a1caf908a574b9da33fb10b4a3a2496b1d0c81da744d0c6913816e8fd4c09f9d1ce163cc6db1278cd1070f35a08129db57703ee90add0b0e99fd8d2703a1a11681a370c93631e9506b6bec8f60a7b89dc00fef16d8c8243d5674264958d313e9dd637d9eef10a80b05420aa93a459688fd89cbe9a1b33801955229af8295d9634c03a8d188f3892f7d5a87fa922d3ac8f73dbe3095e884bfc7d2b17f0f1eac23b3464e32f0a2d52eabe295d5356c130800fac028b35a962bdd2f2487ff22c3eea0aed05d243ccf56d15637cd342e083ea80df8c50a266987589246a30051c89c81695f77aa2bb43ba571ecc7b8c5022b9d0d547bcb456ba867123fa3299d25d75cda662bc28741b12b16488aa445c097dc420ccd18ae808cca882ba977e8ccae042e5d75e7b78380870372f8ec63ec3843189c32c1640fca71434c91eb021c6b5e715a0c153b1b2fc655a53c9e12224062ae2b39cfe06ed94aa4082de6213702bf99ca98e6bedda08e6f8b950826bba28aa7b0472e39c0e8a77a5d34e24c33068bcc12c6d6a960a70883361e20c517c6a802ec3016e2a27765cd51fe5961cabe1084482229f7fda18bad95885ee90f58368c59c78a3e0de8e61d1b77b02127db222bfc4f2cb5387b7834ffb776367225065d800ce356d0fa636f2ea2a9f3649b75b5470a2bea29b73cd2a6ef5bf6baa3751f5f446d3eacb82e76889cf95bf92ab5482c4020962a73e06489d522e7c9afdd3f84cd1917308d5ece347305497a5b3b0511070ce41cbc49e2d71ee67e8b1529bd6286936c385d533917a29b3bc62d565f7c57907645dbc0a3f74252eb31dbac84123bb8d46050efe9e1d68bc5f2165845c753b34b570667b0798d254efd1cc2d434b0f6ce8f20c27441488ffe6566d5733a21525e25d800b83c135e049f3ff7a0e4ea6dac89dd1a1bbcf4cf5a3ced331758ec49aeaa8765beaa6ae966c7787c6f2e98933553c3643a5bbc88825141f2cb2ea12f6800afd5e1dd9276755f69cf6504889ed02c81c7b7d4ddb9e22ebee0512a348ae8b0a8f945d7a09d6cf456e21a03a9d0ed278e278debd60ce65005b0a8e29482ef6e6371435a1bd84bc2353f15024d56b1898e27104d7d4c32b12fd1e337a34d6b413e283ad0283cf24a2b014c4d6d5b0f33ba1b9b8d4ca7bbf2d3467f433cedbf83833ae017cb1d87e47f9265ee6ccbd6599bc8d10fce398829791365892cebdb6928eaad46b1e2f2fc5b925fae1beb567d63ba0b1f56d3f72f4f31f15d88e0c03acb0b661d556ad5da1c45ea8d52a84efe27f66008b9c78617a592e2192815fa94b34907159732c496b3647fefcd84d2957a8e8661efd319900372c70f7d4926913a9c1b3ee5cc07a2ee18a76b8446eec3745f1206958dad7d5f6879459ead3f10700ed4302235540b1e988bb81097a3736287c80240eda9f3a0b87c61e114e1148c6ef07f59175e4b57dee6c785031aaaeab768db6e553c77b31e47d7b9dcabe959fa419e4e11e08b63f118b784a491f2d7462022c5318df9739080dca87a5c4bb645adcfbcd7a32f6e8518859d829cbd47ce6593ecb9555ef8757892d698f2eb5169d4ff49f15bb889a76e8489a69793d88507afb34ad9eaeeed9b9548ac15f9b8c532dce633020ffd4309b269444949d52309e3c823963fed9ae3b44f26121305f543a71ce25a1ef4d0994b11449fd8d01c315f284b79c2791d4be596af7a86af862a460a0a89bc0d7952abcd0d15f9dcfdda6a5413c43b24572b227f7c1445350b1439968575bf80ea99c6c1f4886847e86dad107a902f747aa7dfdb8453db1d0fe2bda9d97a4e5790ad6c6263398a906497fab6ca4dffd80df50f4607303865a024d8c14d71ea4a0646b080e0b856874142b12707504dcd7a1cbb130f7bdc7a652e35fd609f94680262a8bb06c5fad1181e25eee76260b7578fc235691789977d5594a8e4c56927b323c168f4d809f973f13f2884e696ee2b82abf151ae412afd193eff2d88e0a3dceb30d654570c486977608ba0f2ca74a8d07e2bb57a36e078f440e53f46899d652600e275cb4ea3cd7e07fe7a1cc201d5672a88659c1b5da638e47e7f9e4123c5032587940783e98a9c475751d15bbb0f76c0b69d1f33dc29135dd692b0a7bf24e2f272599a91a34fc62e30e575cfdba0809d31f746abb3bafa6a5325ccffbfaf7a3fe8e34ab557ba4e5a81765f994db6bcbdaa5d6b3bcbd26c1316f8e148b227519af490a2c567ea1d7de163bb61803f292011b6353f9e5999677f52069a2e515536d2915ee1430145fb25d360c895aa74ad56b475b43005eb138642fe8cd0ed69499af4c130c7da9a8fa6feec313a0571141ac3a928d9444a8d91df378c53d63351f525dd79bd7c6ee68d3c54f6644aa3c7165476fac65bd4c89c87b6df7f3350d3fc94d1cbe7182c326087c362368eb244d41c4315b6dd7fa15f031e59d8e44fcba34377479a7324e3c13706d17c328bd5defcb63657813ead490cd7ccc7f39dc2668b6cdfe227e5cd0e2bc7be792174b39ca42825c9ff6b97a02b0689649cd4ce4ac5428e837b8561036e9e6637682e17a852cf469df0cbc934b005e7244a68472e1992a601cd8768a88a746ff4acda3912f4fa8107556949cb466ea28debabc322410e6f8ae93788b5675cb0a62c5d050e355b07847cc4f95f31400d01d30b5c01e963511c53203a86a80c74a79eaa8377e8e8c606a449308539eaff0e46d9fbd502a7f51cfc67f50c2fd8ce3d933e75efbd419e1acdf88c5dfe54a74fb16c7827bab5a4bdc127527291bed7a127c69fb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h707fd64dfcafba46951e876a2533895939d87bb3f1714d36e68218d6d314c1245478ce46d70274a5bab13619ae68207ddd1ab2992a512df3a337875479b5929e75886f74e603ec63ee794e2afc2bd6fe85da557a2feedc856146343be1a90ca8cdae470afb19152336d3ea564c089c53b93af7d5f636bb485aec68dfe8f3aaaf7d8fc751876577e8f414f4dbecadde10b3a739c780ac035884d3344b4708dd5a038ca959268ca99074221793b66d0b34eaea69664d7e143b8796f5a5bd3d604326fea95a13a00cde5a52287484f086b4387b5acb0e237ba73b06c396a3856dec24be4cad9d28465c83051f0662114fcd23838dbeaec9ceefa0c5fe499464834d132fc985495fe87feca5669e2f736810f16f0c577f25f09cec1e4340f509ced5cb6d476c0b8cf6b7137140cdc4e4f1154a11d9cccd60ff5f355110bdfe9940258e3a6be2ff1a4ba2e929781f3471452515e671b2eb5f10d202157e6110c172c30f350be7e63c6017653d71170b0ff04b0ef11b8691e28eae21084e647899c612f804ddfb4baced75f812ed71f81dc6a9b1b781338b4b7bd6d901cba8d74cb28d5b6eaa576f0ac2355c3f85b5ecfdceb19235c290487bb95a43ceafd7402204a34155e0f6d81137b45630c17ab831a2d6b67014883160d22ea829f180b6205e88fd4fbb854bde297f6268dc131b2f9f1dc58ad78a93d2858de40124df66f84875e7e72a974225f23bf99ddc422f4cc830e559f182f6654cf3b99a32f6e60099b533e1fb7de192a847c1e018318f61246fbce5e581df833f0bc7e7fc426d6c7aa05926842933da8bd7d76604284ac51c2ea94860f03c29c778dd9a67c003faf2e15c3b4277aaacc9f462fa1086cbfc44f3fdfff30f82c5ef4c24261a2679b816392358c79e6f7bc51457a1cecd8d0b5954fe56aa31c4e58b96eb24141f2a417b41d8acb5383b7acb0471149c8d4364ea43da1ae56f39b7a4d0834f6b295c5125da4a21b73f6296d3df456de99ea199846d98a9a789eea2bc60a77447541c0039813963137198b7c8b9c94cb2196189a31c75737469fdbe6446e93b57cd8d8d07e41c9705fe55099e33af1d309346733ce8e4d60d1f170dc297a897fcc1b08073fff99f62e2fae418e73301dd8baacbbfa6541b3e28ad4e7ec98a88f14b271d8fc637b09aaddc8b360dc932158baa67647d0c410bad79b627efd9acad0d6b41129c5f61fcb6f04ebb4874f269fae6289a236f8c24de812d2aef4844877aa942089d9327a4fbd19579826bd21f35e6ac5efc87505a118bc6ca78eba2906414c4ca71b35e33354d4b90f0a1d8119cc7c62add2f6696f5f768c680102b3709c77f7575c7b0cc365529970d87312c42dde95101a898b2ce1e4bfc93088bdf65fd8e711114d35ee8e853fb714c7010952967eeaafa16f5eb24d6a1acb139e8878b48c21235e693ec588679b69615892444e1e6092f1579dd47056801705a2b784e7a379e55a51e2cac2efea57a40d375397b6e678483f08c6b1201ab040e34d1352368aff7398fc592865ff02702b1ecf85d18b756929d20e45ecf1e3b088e5c2dc8565f0986ae4a6feed3ccd453964224c87145fe3d53e2a8137afd182df5cab6617761b45f5d079c6c1ab0dadccf012deb31c773f37191613d035a6c56c10165590efd715c1b6ef04086eb00d9cd250f6c098c96be8978b7071495b4a8f79e1686e0ba7ccea1e0bfe08bfbcab95eee275ed87a2b01961df659da559a7f936c57b1b4949245701f6fd53b6ae9708d1223588b44dfcd21a8f5855bfde50ea5c0f04f93271e01d2d7db4bd43225bbccfc27bc0e88301eae7323c3a3abe4492e530c3bb811f8231f7d12d35a663a8500d9b5e8296576fdb24bafe36833b0ccf079c502e194916b6ae0abfceae04e9071e65694b0ec7d5f2303a6ed9247929a07b3acde823c0c1b4a1c9903689acad00769f104b46a444df950db7c182b917040bcd367d6c64f72726bf0c746d2630dd8b484326ae20e394ef2873bbfda59d4e2afc9f19b7178d19f61d08ecce41de43d3ee79240329933af29105605b03433171fbc7965e034dd3a70cb11a1ff01034afc3478c86d6d7befdc1059c0f6d7db6978b972630f1d6777ffe4260168d239986b3582797b08ea1211dea53fa2bb44050b1c7c097da762f0f35e6ebfdf3626a27a921d3524d9abd2c68ab4bf3cebfeea46e66629131fbb1c0aff008233d5cf2ce1037b4391f3542897be39486d89bb4a1fae48ad79cc1b41eb8342b2a3f5366e2fe555ddde13a11fa277ea38696acea4635ce3a590a4001beeb8f4c1dff8d90ea192ebcfe70450dea861959039df6905a09c7f276512470a2b68e81fbbd54093fe488a24f17f600005d6ab3fc096db0046c90d37d8714d269ed599590f15a825d68ed6da3d8e17db52a5fa692da4cb6f075c80e028a6bc2de23378b28ecb6604199305e0953a916759e1e2089f1984a21912ae3b807f02af1edec6edc2edd0012eb335e7c9899042e3d98d62c159dd4f0ffd7ffb323d9527ac53b28fcbfd945494178886c6be2717d5df4fc2d559d386a7fd7e28f3c4b9343ed5987587dfc9be57c018127d1a26e32c5f865a89bbc75b9aef43827eb0afc858386a83277f1c5e6307338f6d55fd9f7caf5454e87f84d2c533714905c9341b7010f4f48c4580e7623f65e9bd8326e0d6aa0a66aa747ebb0a258bd1a3a47116e1e06eceb783e08c2a801aa41c85ccb6132c930237400881f9e351cce30b433f4f19848d501cf7da70187c021dd88dabfd2d7c2495a1eefbb7c72043702eca46920c78792f7daf0c84e268defce98577991096110ff681f75c6c322364e02682f5721db049d241505157bf9ae60254c62f032b676f343d6a5a422e6f2e4dae63c73e36dbe6811125880be8f2bf6ec9dd1ea566179b80bb1bbecc04d504896929ea588d390eacba07df638d62ca46225a54f09effc2e214d27b813e6557143d2e77f1f54e193aeb5a7351868e34fa6ecf260d80834d565017608ff21cd9311e7482194c04faf4c01c729b7d29808480bc707fe82b24a2c3857fcd3c3a76f152b1e97f4ca01d2ded71c6e7a34e4c0450f6cbfb52899b686715797d109a5833ab8f833765707e3645178ae7b66b792eefdb562f34c7d6d0b434b773deb75e6d40dccad43ede8a0d5cc4629c3e13a1d091460118459c1ecc6ca707dadfa1c9f60ddc624f60e5687099c624ba375a9851b43fab819fa4ba0e6e737bef4c009ff23e5eda4a83406c660a93455ba3c06c464764152ff2058458194dc3569895b35ced46bd7e04e1b68a2b8332af65c6a724a2137e51147859c28560b0a4b8504312798212e2586a6bc48e9aa6d6908a3b2142dc26cfb0171469c9a08abe65385ac4a40e73d84fda45e05c0c065a37abbb591513eb27ac7259b391f02e55ef632d9a4284e9c5a5711ee4609bfe21560e7a301c4fca5dfb754f30c85c946fdc884bfdd25aaf24bd50b468ec22d761dc495e0a45aa6cfb6742c6c5c7099c6843c11aac877ef0fba00ba03269233ae23e2f964d8125e23644fbabac033816037df037a2f63abdb90d829d09e69330734b6fb946e8fe5207f1e3d23b85f51ba9fd88b653ac05fd44e13d52724125e5eb86349c366db65ef0816d3ea3588dc13181bfc50656a89044c074c69f7e28efb9bde44bb3e04c589df11408644d306493dd9a63baafacead44d4fae6ec80d8acdd47ba88420436476ccae02381cf5fdff3dafc950f0ec02c460e2f017bdb987ef28ec3d8065a146e6c5f693835bee175e24b991c13783297e228449fcc6631dce8dbbc19af8ed24a98440a122e07c1db80824e886e0c0cf5706f13c9011e5143ce4f0e561f5fb6675f199da42812e77ca98cd53038defe8d8c17ae65f37bcfcadda4738939f9cbefe56617f3dd4f27dd79149b62f11dad132af54329a63e8bbd93fdafa9dcb7148c91dab12fb7539c94a496091a56ca23a5dd7ced88f67124db279b4f8e729ac4e264a4e6470efa6c019d7a9845583aa744d83ad7aba0f1a8660177c98a2c5b52194a1aea46de5e1a7173eb6e6287e5b4a21ccd22f9b53928bad2ba5db98d7444534cb71c7dd81072c66bf7b89e55856509b79753cf752ae5c99d602667bfc4c100d2925ae07dc85255fc85626bab8b566e3378f4b71fd0860e8c3818f61483d18f80144a05368c06037e90e1385a9cdfc3895235e8cd9eb5a2b1c70297a0f551faf03be2a5640ed7a16ba34aef343a9cd254f23223f2fbb2bd9acac584ad749cb159f1e48e47c1c69c621feaf6f406bdde310839d0af099f4a4dc08a88c2397c263e825fa906cb1958fdd7d438da0e72ed9db4d5464ac2c09aaa0544a384acc2878ca8cbc5f6b333df3401c95f8eda852148bd5d6bc81259f6ba2ef5e3daf93558b88dc27db49d99afa51e8c3f8654bc6f7d9630c4df20e31919c67a953b4fe6876999aecb6495d073804b5aa6e4120a05aa1737f2331469b5955dd42db59d676b360f5d995552d1e5a43cf7a7798ee957fbe945022871585d1ddba720c734b507c3895cb47f41f50ed35a7a52c4522525507747ed391266d9b015ccc4dd3c8c00d94d1e05447b8439fa524ea079b80be44d56a5a671088cc62b129dd5039f6bdcae14e2335017395a78c896bf488ea23144c5c30463675dc2fc6f2ae2cd198895f18f5b461f05b6c36ba3a050b46017543437d0222fb4586c9f8cfd3058228cbe4b34994b7105be8df317e8a37c51a49f5797e046e4bbf303ad7a815b92be002b7e479e009e0a80027bb7e506c9ecb51557ed443abcb45fa1c53555437b0accd1a2e58421b3989175c34753fe87c75118bca497734137118e46cf29efc06a8d2e41e1c68589c16ba53b80999a14f1bc86c28cd6c06258cb6c0e058493be39201723fd6f1e26d387b2d05c8315ab46e59c0d7ede5d86051d42343671c9ebc0a745df9f12614468fb4d86608078777a3b2b26bd5fe61e81f6f75a4d9a57d564ceb28e0ca14f6a706b25524c8c74656f175eb603695a6db3f5c8c80169a7acd1a3e3b2af28d078786635bcd343a4dbe573d4c4f4b9e3d66ec732d9ae12c24838258131e0ce6883eb9d73c006bc57fbc0b740f37f9aa11ec183fab3ac55e8ccab2988caba5ec1ad36acd904896ab3fa97a65d721cba132cbc4fb7e140246c62831c0121f57f5270f46643a7187afbf800d3c222f8474725df44480bfb8b174df727ce3dbb9d7864ef32491e6ef75d4b1474361db292d963639ad8a8b9dd396c9193fbefa7898e44a607526f0ef1e4451218acd21a4e966ce9c8831a450ad68b80e7f5c389894232ac9cb58f7205a441be3ea262eb5b07b348d4296d36077a5b24b894d7a2413f09d7eae086de74bbbb3899261461c05cc7c3b94ebdeeb4de434833dfaf979b2ac8f0673898ac6cb604225777e17269e6f40a87a68d805f05f5c3aed23618213c7625e4b17b2f4f23416df3d230809d1639cc1e3867a6f12;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'habc886e43beecb6f1544a5ef3800b63928e1eefdf6f6a2777640873d187c3f95334ee1f422e705680c4fbbe9b7d5ba034076c2a3b7c6e53d513fbcf0ec9436ef5a6f3ede9aef1fef7b4c012946a00d35c2839a08880951a2cfca28978e3353dd7de294ada766a6afab9f4e1a294f40fa66e210faebd54228d8d4f60f5be1856c2c1c7c1fefc5f95adb066e58eec057c2b045ff29e30b760cb566934bb68ec35f23633031fb4b8f018d2b742fcc60ca982ab9187103f307ccd8c943791986489c42c4d4871ddedb2e6bb078bbdbd6a6d8b3735d1d44c5fd58379d767f456f8a19d973378caeedf8272d2059619acae254a6b7512b4383a06fd15ab08c38df7abf06855ea1ec09e0cd699e43105abd7c13c19e0c428278a75699bd1ee6c912728981cad6b2f721b4aad896721bce70c394d873675c58a3bbbdcc44394c4b34eb2767031197ff22b9d9ad2fbcbdff94289dfc1b6abdf1da91a82b7bee91170d6bbc55d39e79007780393b84237423e3932baf15a617d9d51ad621e361c5b5923daeb5576b4fffce228ce1143cbf1d8be12a1abf779b571e510356224d6a132e29d20f2908fe145762b892725bfc9ad1e42ac9b13adb1ba0176a0e2ea0072ecc3d22bf49ee60a94e74c66a8da42602ced4455ba2eedfe053d65900311aaa1634266cd493bfc32d1ba20178c7e9eb43458ecd9c29e6135271bcb74a26c0491dad99b43d313f2fe95555e625fb298e30360196ba8c3456777775c510a1da29444764a33c096610a898bc93f87099a1e421ae72e7bc30008c0f55ad02a7c02295735638888eac8b1d25d0d2f6c6d62f3c437a411a02cdf22e791c4f522023ae134d6d8e6a3bf358df99fc2c73e3382432621fae4a181a4a2b10d84f9dc98327b983bdd8d1b28e1623f7f6335e7415b9dbcadefd81ab3ae48ee8a7152bd616c16b5eb97e1d2739f20e6688e1434312e0222ee195e7935aed70cf0f3cc3c764eea868ec23dea6c9c1d740b968d91dd84462adae151281aec948df0dbd01052db57bb1a6f58fcf4200b5b0bbe512fe60f0e7fbec6a97678c640222d2da19f4aff9f81afa54a27b3f1c767d562c68e35f2b54c1641bb8d41a07bde61b737c3e2579a20b9c9c64fe822e5d342f069a477b54cdce2a2dbce58c465dadc61871d8a004286b272c6f58553b5a1a49656d1228c1ca5d940478e370916bd1433f20a5675fe0486e0acfee604d8cbaca324d79e188b9c8f7f00a2cc53e97b9630d4cf12a84230fec98a4b5292f7b099dac6e0216f67b85e7278f12a4ec0bf17e7dc38a4e563b68c5d7cea9f6aaf50687658d17082327a48c82283c17a9eaf36e0127ce6c8c7cb8cbba0ae5fb3bfc6543a3a3d74b6f2f9746dbabe3b89298ce7871ef3ecf7cf77d557fefee31014ebe7b924f512a7ff076a9aaa00e24a15c7060a2d19481c27a9e59d9ce2605f293b4ccc66f4474f0a91b84e1e95bd21669343df63a3249780213034ccb1d47dc4f0e47df7a2ce8d0e57020574c32adb26262a8250e20faef32e497c36da2bfeb999c2539ee2fd4e96441bc04c0ad33ce8f59b7bda43e6c1441a3e88ba4c5dc90c0b188f2c780428066781f292e5cc2e537ce3101ccffceaea1ae557ce15d567c4e69c96aebbc90e708969a2e955878b17be8e3e2b9c1da38fadaf9e1d1c22ed964f87823e392988f2ccbed9a236face1e2cd270f2f5f21d130cbf2fcd6d219d5a1395e1c8a6617f58ca65c24e028df04668f511d10cc10906835a98d6a11e4cf924b8a5f3148d8b51d0802d8aaba1007cbc2450a9b157f3c9f98e07e8f6a3e663b9e9c230a5d7995088e80ae90ad7dd0aa15e01178d8781dc1b05226190963865a9a513510218eebdc0365e9eda52ec4847fe1957af6d06d79c6675f0232f8509dd6cd62a9a55b454ddf033358ff1d4344a13854893c4e5deb98961cfbdd6fbf0f8b65184345934a1f22581c7984a4cd67281c506aa721eeeddbf280534db30490bdd0625609dd5a7ebf8dba89294687994883899f1582e015190063bb2e6404def53f4fe1adfb9d1f121d00ba67b8227c17259ceb48104a54bffec302038955ce0b63868dea477b57a3f0ebaad38775aa4ead69f64634691158e5ace54c5a4f684de0a10038c501babc5236ce4b528e08e6364c2b90bbfad4023a98365a58be31103d19f916ba291af21d6635279c02f3edec350a138b82980eb0faaa3f713de7a032696d03f1749967c56158c92271c54fefe120af1caf12b4a30190fdb77556f920b86bda982a23663d8004633df8061dfe66bcd2c23a77efc8d9ab8baf0bd42e764d34fbcff02121251f8b846d5884f91a3f47694393c41cf84ffd653dd25f91f5c9afa9bea2e66404ecbdeae3a4d66e6990382fdd4810866adc7657c8bb1176b0f3d7ae42a24da2517e0353fef2f790431c8d74a75cfd42ea80a23a2b9e7eb44c9266b171ddba618f0283c7c6a7cbb56ada2fd8d7d9cbc06a5db0ac9944173f4dc36faf834c94d960628d9264a93aa4966e29364303bb6c2f28a15e4ab1a20c88653f74bf8d3fbc37542979ef9e3a4eb2c5dd4f84604d369512586240285528357fed16ca155fb754a47004b3175970c254f864d707eea4fc6095ff593531603aa5077ec2203d458a151269d4a7aaf2eb60cae787fa3a9557a76dc23e273372b35228e2d3695de07503e2a9ddbb19f1cf066adb3ef0c570409e0d532c2c6d14cb8e4fd927428cc4464d0fc0b1aeb298be41a0ed60aedff31709687abcdc49f1b62e3eae981d142456345341c5d05d6b8804bdd47f57055d27dbe057fef2a5e420b8cbad661724d164e9d77e46652f64b90044d0547d9517a5e45445d56bbe56e69a66b70a7d8e0db727e47c87cb701a5751b4afa3817d10704a45f55f15358fc3254c8fd2c207c74ef0cdaaadc2006b5ee1854373894e24327d7da7ec0dd91ef3a16241e55c0a03c1180e75eff76d72652e4bdcac81c68e4527f46ff675c2913b3a375667bb775117128951869a05a9e884be6100e0c5d822aad2f18183666ad6903c096bf7d1cfcd262a01d5e9ba646dbefa4173f42bb0abe8d25e787becece1acffc3ad40b0a4533ad4a484d63e40ded00d681a4fdf33a0c4bc679d578ae66ccb9722e6a137d8dd61013ac9d3b1d671215136337fcc43e302feec6ecd712f8447cd56f91c912e56a28d69d35cd92e79ad8e78d004b440a0254d42dc399566e2bf4f1e0796fb07c167364416c58a15c7bfc25a7a679073029e69b70553439a419475129ed5311acf13b725188a415d4fe9fbfe20cb140d5b27d355d78d26a0b98e95272c37bdd22817bf836ab973ca36e32dc9950974610d2a30daeb298d66af0c3b58416c1595aee8ee3288d97bbd3e9b09134706c8e7176c9928967d3067555a03ee999c1a29977b3467326ec3f95351e06a23e036064da49b181b4870afec914b617c7eb6d482b6815f2d4ad6cbf08aff2322a54d2549957e42e3fcfdafb457ba2c4abf736e3bf2357be20db359d4d05d2642885d8e6c4285437f3b4fb11013553af2c6c8cdc63188173e03aad701355b9adbbfadb8b37747c3a18c2e9f1029bbdbc2e476963bf1408f5bac82710917b1a2a0c808fd505b43d01f1a07ef5919d243cecc6746f6535f07dce79c33fa2e4f3d1928a8891774e6768d2613fb826be72aae4432a0a8d02547550ef8879c10d2effc503876e57006923ff359f5a9ab4496c4291aed575bca7b77275948abdc2e217a54e4e3fb6e8bcdb63a17fb124e2f42691eb32b1e80fc014b66754e60f86ded4345c38fb33547af161272bbc8d6e4d7a1d86a0449d616bb9d2dc14bf4dea50ab8153690e06af72ce296be76a92bfed8be580fe6195a1de91ab32a8bffe55b6448cadc0a5107f11c7b04e947998f34adc04247fb959b59a1cd2ba98a094a3c840f7e69a93128aae42809a0037e17d2418a0d3cacb924f554adae02b710214ff308714360a46cd55d0ffb29ee9ff875992242ed102fa08616972e9d9553f39de7ca4995612bf76e77670691027b1f7c44d2d76904c4d5d367ae75cd173cb73e15738759658c77bfc226f81849f04f02c280e482007cfd3b0e4cc36713b5b46075ad681a88ec994194f465dc71a249c044620cddf5aedd1cacec84a26ea02c0fbdd68612d83649d04d95d24a6627f9c3c5a139524b971beff9c4f481ebe3d1829d1a53655263219d170801a8ef8ebb186f97adec8d22eeeac7be5a16392287ea697687827f1673c3b65c11b10aee07b8cea6dd8e2ecc2b1a40103e093fdca9f90671da9ce371870b476bde31db163ecab5abe88e120791c5f3348aa6d703abe80196d996f4d96a7c82b1151d83dcbb85a2f1bb527faa9c09c2a2ea9fdf2cdf0e8d09077dc5fe6e46d79698e3c630223b6e01981c205921bbe4612d48ab303a54898999dea1d4692b44d4db232d479e48e93aba532a9cb610372337246817702f6681e3bff0f4e9d51293215fe84f6cf38e3ec4ed7cf0872a52a80d6e6723b8afa0c3a3b5b6691c9d3b1ffee752f89147be160eb3d17af095cc9127e6c735c6a3668ef6bf6f75806c39996ebef3b8b2e1fd6ec5af469b3b6903e2f285469f823fcfd45580cc06dd5ae7f1e2644633a07fa13338453aefd0b413cf4c96d9e087a5c97c5d093b33407147790a94f5b95474fffc813503a80d0b4a2607fed64bbdfc32760346225f75881b606c073c642a32c1225aff6253d0f5cf443beef96c591f05a1bfc028ff4f2eb5070f8cad051a5f169dcf6187d6ed8acd882b4d1218eb4a2c311c81490bb26f8a7c3f94a9676ac144d43ae3cac91c08966647b977f1cd7c10b23f64f5dc2e93e55f0fb252db5b7393569c7818224a7dfa3d90d21e1102a2e18efc10263f85ffff6570bc792913b6aa474308a1fc7910a86300f8f372d428cf18d166bcc92c51272611bde19fda80eb325958988c67f6544e98d3689683bcb00239f6b17b3060cf3e4b62384290be7cb2696936d934cc01c8f28512271b6f6149a536f300e33f207ee3273e5ac559c42d23aa3a4b7892e7f11ea20c08dc367273023ea9c797e5f438343c1c8ff08a8f3b9823654ed062fc211c90624f23a79b4c8035972d7ccd903570b296ef4a4c639a2222565f7ebcef331c4952267b0c358860665a714304ded106690980a47bf9595aef4e50f5add64f8d97778f9207d86f4160b4785c9f8dce0d69093ff1b63046b1b9dd350bf4b4259a1f47bff2fa7fb7df6be07437a2dd158fcdc908f79ae91443b03074bbda49cc1177d1832776bd4245f0014b2f0a0322dbe0aab438a08c435e1c6e7ad30aad0594edad57b7fbaebc3a7272f2c2bddad28168590c92db66fa7b160c8876d92d7eec26808093ec30b9d827b2d35912ac7125d779a9318477f2b84cb0c041ae8c9348ecea4e821864e0454ca9b6c1f809f83315cbd174633105703ef7ca2fd8c408085e72d3e6fae3646f6e78cfd08ba473b590f3ab6de2c3d0686102698e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h198da127555509ef04f62d156cead0a427b00d43204ca3239396e72ce25de4ae5665b2a8d3828d019ba354c041654c0bc33f764602ad460efb183b0642fc6ee95770eae6eb4b1ffe95aad65725e893fde2dbe47283081039407d3a7e2cdd47e14f7de25635c4c05f0a991c489c1ff8ba0dd6d62ddf9c46ee532f464ba0d9dc7a3a776b8c58dcb4bd22d066f179eb47a828196e8af26e809290b56c55d30398b8aa47c7ba59ecae9fc2de84ea72fdf2d7e85b8de4a268f588eda0297fd45b5b898ceab1b94be2165b549f7017644d02ab969ba745d71fd26c1f7364b246edab44d6800edd47654b828d5012f1c0027fbb072ad8f8b37a8786923a6b7db84c190ee959148927c18bf04e8bd34bbb6e80bed40175906a75d993b197cf5dacbb450702d9e5f775415030717da1432567dfd0a536695c099b3e9125ae25ae8b90068848633657a1e084da135b3fe4da37a7ca3fae0efec1dc557e947d75ef927b5a810523f63316405caa12f945f50d56c7bfd28f55cf3d37b9969ad656ff2f8030495c889df4cc27d20ea1f4758c49459af79317cd973fec16a88475524b3d9de33545bad3a1da112039aabd118e3b384856ded4ce433c96f8a64d974ec7d871a76653afbc747f9cf8e26e9d09a4c33b5469b70b7a7fae6884f5f304af1909bc67de84fff245e4a8c0449198c6401179f6340dd540e9832e5e904e4e6b5af2a92f2864f309758532ceabf2f5cf33e3f33f2d0deb980dbdef60a6360879ee10247ae6d4826adf5d9b12df4fd5d34198203c2b07a358509f14eeb4bd55b6e18c0436824869bcbfe9ced9e0b57f90ff80e10cec6d90b323f4cbdb7e1a4e97c90f5c551b5cea88645b961ecd022b48016c76369819daa8016c578b1b64d51ab176a7b4262bea8da89fc36b11157673cf2cef772d2858b8eaf5bb5a71470a06979e7b5ae92173c8c474577ef711045d09c25d4f0359bcb8a60e31ccc4fdb3f55c2f8ba98eba00ee47b4ca0ebc105129f9781338bf904006844dd10d2b8734eeb165dc780b195c2d6a785c49c19feb631258e2032a571aeabcf77e9fbfabf70353471884999f072dbdc18512429662ef9ba2ee268b0884b9128d795f7bdef63284b6255aad25ea525ca98621add544369bfc4e391d3b69a6177efb6e6d95a46a2353939f022718dcf6141d801910037d890e4c91c85220149f85cb220ea9cf356caddf177508e6a2039f9fdb2c6c67cd30cdb3d0d8a1ad24338155ae9854372f4933bc7b96d3d70b748c61067730a419e2deb6044a3ed4e89ea27d42d4718133e018b0d391dea6c094e0f8b3dde25af68fd163501f6b7fc5193689cf02f536069f9902e119447350a756dfccd0a58397cca49d97155cce27cda6372ac473c31ef051d00ce3aae8ebffec448a3b975c5d2664c43c7d2c5406298cad848a35f6f2ab1f3b3a35b139662de26d5a97f3db822382ee02049af2afe8c672577a1464218b975376665e3e547fa2b0ad48630b1962db2f3d9462a3251cbfbb8027a14db5fc9c41bffa3da276edcbc93c581ceefe6cb5f46f9fb0a10d9abfb992b2a877cb8f5094713bfe8238b859107585079fa4f96f785979a546858dedbb5c8f7b2bec1ded4f26741edbe487cbf5480952e59a9db1fdc0d0671bd9816dac62c011307439d11edeb69d946b7c4a309edc78e88f106da3c8dbf1c50d68703c66f2222edb9f694124d5a5202257eaadb5c97e00cfc9e37b01eb38fd03edc079f1074fe60d435fb64bafcb2620a4975dc0d3942c6532c0d26b0d41194f756ea42440a522dd75b32e76bbc68960265336d5cd3dd1f58d2835dc4ac9c139e6a62b390df3b70d41de0231d35461cf3c89b60128423f95f02b80520132bb91c39a429ccbea5b35a0bb10e97860a54c4ba8bfc954153d91dafb56c8482028d630558792e03849ccd5b4834a66dd31b555cf5d6d4023a822f9402db8c46d76266c0a120fe36d7922c640607b06eeb072a423c1326a699b55f0ea49021b5de34a77fc1aebf2b23561d3984fcaf06f86ce82a6ef84002e7004bf2d5ec4561fdf7f2bb9ea11de93ad84c9968121b6b6bd821162f5f6f8add458c472a500934edde084f9648d41040b02e684e54acac81355625d9e7c1b89835b6bf460b20ab9f8d994a9a8dcae240ef1ca9e123cd8c7ac7d8068cb847bb359e2016d2107f6b3176391a2b17f26ef5ff7cd0c247cb84972cb7ebc18f398a96bbd1d568a934571dddc547bef743cf108e9d7257b544790ae263f3ae13d66345c8a2b4e766ff3751053f6e509cb2decc3455a66a1dae76ac37e1e97bd0933b84e4a8db6b18fdfc500ae2f757c1dac553bdcfdfeea0748cc89397e6e96da87884e8b4543d0e85e496bd00f3daccffb8bf2d083fbeebfc77f10a10effb38e75c2d6f444e326912bb89aee5d41fa993696c0a69c212f63d994c4716c3d97deaaf0f2d919606b0e1ebc56338843fda332c557e7f219d7bea01f66c72aaa4ce915d6d68727884c3801a4ab917602cc363dccf199a1d94b2da2f93900924eec0278962d995c002efbf1a465145cde4fc8c36696e87f8f761e5b114319d94a04cc8f2458bcca21d87e8d94f75741c00cdedfd72aea85224eedaa7e1da18ffb48879504ef8523985448bd125e5c322f75208c0ea58782b6c3f9fa8bdaa3a072cb516cfb1a0b0d9eaf24ef3b7ec20216ea5bafddac1d858a00dc702150ae10925d5e89ebc364eac0f5defc7e40a947d45a05cf51116ec1a7035df5fbcc9b1c0504e0501295a44f9d35d1e1bbda05c3ff25ad03de6db0230005d7180753f842c7648adf85c39d353ad01c1c2a8d25ffe3dc88e3376bf44509e1cd5264b688d70813d6064769639ca93d4007dd920d985d1cae2d91cb1982e42e0e65d2a5909633bac71ece5fceceaf73ebd45e78d26f1dcf9810de5b6e412d61141378aa957f3c4a35e18502726baede6b59be7a31d11d20a6d7f925db525b7337d74f80bb09ed4997391a3f0b55533966c8d6b566b8a16da84f15dfd2a649dccfe310a01612d0803d74473775235b2395051801983491cfd31b04442cb2c80fd669a5b1bbdff7d7c57527957feb3d03bf90abf0f404e7f4b8e511bb4ff00986af0fa1bb161b15a4669f42eace5f6cf9ccbebd09b223fcc2d241ef755f5ae3829193c0fe58b574ceda089f78445c619300a0bbfa66f38aedbd6f177a2d9b69c1482750a98c726f5600e471982ba1b199eee50cd476733c68fe476e5ac5816f2200cf45740718a1f2426f681a76d2684f2ec431ff46b9976d5c26807ff2ba62c001a963c165087de6983d639a26ad16e0e56f12501f541c864cdd51a95b44d210408e76d25475969ef5ae6979d7e21cf20eb62b1d3ac59607ab64a61e3124683c4887546eff2255750613ebb14b249f69ef82d883f04887380ce4d4bd13136b7954e0a045721f8c14a440c53f16cf550ea46d1af5b24d37d0b3f616478fc8b14a388ffa712368be4c67bdadda0da70bf9dc671fb512fae35a333e5d608b6ebcf1257a400495b1af8044a79aadf4974da4c0df83bb7266e5c283a515a9623981f8b7003f5c60992ace803103d24f75d3cc8440821157ab61fee12208b179d8e071d19e31bb96d9dafcc5c59a22771484817a0708ef5b47261a97822df4c033e600b2981094f593df978efa918bec26878eb0b6ed24279dbae8c7a28a6fcdbabb380b92c522bc756e962962629dc134c51906296c599d65af0328f806cee191ea02e5fadb3c0ffd219aaf4eb4d289ba461c57b796737f33fb0a3e396ec49f328ced62f93d62d47a6e11c3dd25ecb4bdab50ffbc5799e70126ef40f69e971a74869e08137e46920df892d22dc17b2207b9e8544314291fcb6f78f2d020efc3c897eeb20862d13c297eca4ca4e45ef62469cfaf30a3e2c644f6d1e877d64148178735ddbbd347563081b0adbd87bd50c6c37d3ee4824ea7433eb56be393720e04eb7a7a2abdec7e8879fb412806dc045eb51127780737ec9754358e64b4d873fba53250dbcd9dd5e788dc7df2e74a0bfd546e7b2398705030a2bf003baf449ae3fa59f5262b9aadd78fb8cb02eacb42a6796822cab9c95b9c4ba342ddb95f361eebdc47b835e2a9cbe7b14118cc6f69545af220281970430c7c5e58373fe50c34c743ec464cd6daca8563885c5c813be014097c666a2351f69e79760097d97b201d14c1aefe776c2371b1036f17f4030af318efc22e3dd53a35dc5ad1a2608031db54a755ca38dc4db95379328a52bc8afd6c4073faddb14a914dc4fda8336206a600916f548b6d7adf5bd977c40ca7935f1e061ad1f8b2e0a503d43042c6eed542776e22b536ac8cf589fb8005470c22b70c7939f0ff14ea1a24b35787af5ef76bbf11e5bd1c71d02bedbde4204e8998d62bf45d088438f8a8e558a385d4b7c5508bcbfa573823a440e24a899fea2cf188d6123da63bec75f9bbe2f8ea01de6125687e2583424541c5685d44adbc9dffa4587da5bc67ed20d39b2dbbb23d55bdfa056e52079ce31e3d4051c63fc78cc1e52da17cfa73d9ecc833554c728596765d954ff95265bceb91135461ae77b3dfb91e4ac5fed357cc45ff4867ceb3a12c677a4d619e48f66d540e132589d311ea19dd9afb4e1dfdd89fffeebf5847203ad15e72cc8b0ce53f6088ec35d0ec7feddba408c53014cd19ef4464c8ca34ac8a8d00f63bc4a2623d8fedf773fdc92d99477ac149bbc5a26e3228cf2a99f0c84f95de1a34f1fea6d0f712bc99c4580ac52f948cb50439f02c1114504b0fda5d386dce0b1741460a847379d269187a58777d7ee097191a2bc203d20a7a1170251f1bffc773fa56b5b8404c109931ff72eeac8c25dd61004910ba8a591af64a7a91daf8fb19cbe690ef0bc23398a0dcc58431d8168c1d4598eeeffd1d50d34b55792da86d7b3392848bc5bfff353d71d18a98326a06d47a5755a44fea83e9409c92244881458cd1d182c80b261a3df085890e071843974649d029f0e1e835b1b3dc1dc856d91e96681425a426aea5a430356756861d20fd1c1345ba75bd9019254bca584dcc2f5dd9a9b3511ec0f624d160941e03247cdf8768be5bb724b8553b37a6bdc09d576f7d330aa529d30b274c74d783b0841b235bf5c780e02f6d1fa1bb094b9eb27a48828be571bbc16975082c8a1af78dff3320b1b7a63a645107bdf5c1b53911914b9b6cf9206e22fd8399a2ea3e082ae38eefd866641ce63b02b3ff11ce6fc08d000b3ce10641fb0d9a5dbd5ae697267b8678b44171b693e66ee0c35d1b9487843f84fdd823892bfca12b0fe89195961ce6649e862201730d5c212adf75a5f4a9638e3aaf5dde0649c570c367e7ac88e21697615e28e93ec693324915c3dd2b704b405add738ed2392b7795b8085cbf0b4e9562fc404598c91c23a961dd402824e92dd679c7aa6180414521fefcad761a7303bc567d547331b6acee305e17238af2241ea228b70521715e7e2bde741a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h49ec0bb3907d724034aeb2ded3b94173aabb55aca0db9bf7f3c2bd0cebbe7a16747c9664f68e508d74639e9803a2c2d22e1dc3b8bc02d943735668923cda01a2c7bfb5435889e8bca79659b191364d3ede02caf9db7f26f19abe6ee08e3caecb18c63d5bc90fc40ef9caaf4cf8cce5104b254d33faf91850b7962cd3b7cc9f2f7115f49285e428a1575f220c0936c5b52faeb13d68c3f5bcd0819dcb0d8ea312edf6430cee2c1d5bb47a38d98e2d1142f415e24f463d869b0c8ec285fccff9d721aa93d2149c0f1cf578c53551314475d35f3b1500706df410b2d1d1ae94cc832a39de611f150f5ea1db8fa48bf3fedb5f4b9f4303922f02764a053ffbc94a69fb5c022b6968cef21ffdb268839ac2ad8e30c43ab05e242a1e0ef0158cf19f1fa54e76fb65fa8d75afef79e509285fc239eab57c3e29bfb9758c8e9853cee2e4d2ce4880552606c3f2e0d05bc4de7dd4fb749f0e62b4c28d7540d6bce8b9d4de8b184ab5223898f9441cb4a4804f238052d162c3e97a7fb9d6e035e42537eac18185fd1a5d029e62922ee863e459b6e712a1697e7b0453176b43a54e8aea41f3fbbc687f3d0eb10b2a97a7a7943572d4f207195d936e16d876f8b593dac4009d6d9f1cba773f8c1b5c43bb461602321c41c133534b3fc92b8a4cd613f3c1658150ab840fc59c6b7e0fe15cfed230395f2c11af7114f8b5617380607d43fc80b0474bd85bbb98811d0a5edfaee7d835379b4aba1e1ab5cef39eda1eec24f1f68628f4ca23d7453ad66f4b241d9fdf055c60c4891a5c49d96450edb932436324c0bdd87a12b7a2d7800105235fdb7ac54198861740f3950eb431b3f76381f4a2c6796b209b8df0d61bd515000172d0d4b862892ca3dcd7b9fb2a54d3e2fee66121185a874209366793fd0f1014fa88adaeaad97c7862ac007b5090ba76daa8a3da40d3c5189c17b35c73501a8c3db7f608a9f2b30b01f97a95e37eaf8cc9db7ccff556d03340e71bc02a385606ce2d2b3f06942cc6c3fe56bf33768364837718f85dd0237e8ceda0f4f5ee790c1f922605fd2a5b1134f33cac79990bd93fd8eb3417b97942a0102c60e000d7fa5c1f549d025599dd83ed2d4863b82ef3a151c8e669ed36cbcd47664efb8be6e46bc9e423990a9fca3c81893be3c1fe4a044ecbcd00febda27a568067f3189e6454ff8223b6f43d778e3798cbcf080e1019376e1767a0ca0efe55f5a0cae1b96f5fc5029610c3acd6dd6e903bfc766bf5825b11011cf5bae857a2f17dad5842d3d356428ec3f572cc18cf21e99524b5daf7f99de7a865adbd9e76fc02aba9bd9e7a75c44f6e922ef84447b3eca0df7adf2f2559320b285497575e722adb1897c03c18d176403ec07a992580d0f85d555b37f49111c582a2e6a803b6549044d440f5bc99c65f1d4e19c6e66e8e1a788c11c21bbccbc89ef535c26ec8254e340fc9cdee5cae9c24a233d0427528a8567c2d1e749c364c07e08ef2ecbba1b51e39bbc2a61f4f5b27aae4d5d70769b65084880d9d9e35823700f956b78f94ec889df5958b2fa6cf356497de78808bf4d6457932b020294440f7a0faf4b0020c51b25c375eee35fa15132dbdd41877a0fcc19453c58e8a61cf52f9ea622c3401fa31fe8b6ae7fe760e0d07eef2863927ec09a508b8fc8eeb3b64630a5dc819a350004a329a65d4ab7479427317ca927868182fd4477c95e5f0732b4d59afa8fb896c5566794264d719b49d2955ddad36851c4e27ea751eae2edc54b70c2ed28f27bd3b863be599d763d48d7f5dde9ebe8669b2721389bebc186f341b3f1488d164d42e6b758ee07f100a1ce0b692ef517d6883eca2d0f9e00f1cd617e4c741bc110db89be76550e74c4f5804422e943a095d8aba66de58a42d0c1ceaf7f4e8dafd342a9d27fa2a9bef12d665f6c902f4cc54fe97e505695f6dec5d7e512427d9f37f7618e975709962abd9de7cf628d51d1f57719c951758334f02c24302c048f75e29422a0f6c63456becc34b71aca783cb5515d22f1e6d28fc9ababcc64b774e8c0f6c112c761f75201d0701a4fcebb98da3d348e697ae524eddf6c71faad63d50cfc0f3d1ad762df78f388b1b19353be1a986859717a1d9936fc60944f1f06e3bf74a9c9be413c9512d90fe5025cc6f04056e25fd1fea9b5c6c42c45c0223a4c64973b203e6ba688a117b60f19f6cc0526e59688798b7f4b52e699c771407acce531c7a48da9c7f71292e98fbf572671b8e5e8708e4ba7b96236c1fa6d9917faaa93af01332719ec85885f440b4695ca2c16c2dc718eac028f09913c22c7b0d15f4edf8f7f6be7eec57f7481658702c7a3e29a0c2cdd1d11e6a8b743637c1ad31ce0b3f7fb8ad5cea4d8fbb930e79dd890422defd5f42917c57f9b858c8c6eaf8b8fe93cf75ed0ae52dbee1bc59436c3dfa5bfc5ee77dcc1683c42be62629f3961dc16f0285f4c3767566e61a44eead1ebb88a2470d37df22b100fd3798f5951b7f887b9ed5008cc4243d5cb75b6ceeecbea9a4ac9ae5a8ce5c1ee412808493c35204ef6a465871ab77bbc1e0764e439216b51348c3315e365309fd722313764d6c6d9052c15e97995795f9a741a29b2e447a758cbdd6936900a015cda525b68dc3fbf4b62bef74075e7eb37e9dc3d2f2012453140357840af73f3fcc694c366bdac30db17db04b0625a044603a62354d5e0e734a7fe567cbe2f3a37de48788ac2a73560cfeb72636378b6a11e180c1a492af088dcc7569bc08e5fd25178ea83f53f19458eab0c0882f64baf349838a7b36cf499cc850dc9bb369643d7c3874d020018aa6f43a7a5409e4d8f1572994f4d486c5c35dd66b77ede3f532c536eb067949703d7207938d4927e11857f50caef0a9f49a7d52cd3f9df1d1c6283b6b2450989a9d442c0beeed17c82471b9c2e6dfadc88d9633561d217bf112dda70d6fb5afdf49bf0db17862976ef5f3d5ecbf569c1ffba8e6fb5a578cf5693d33d621c32d97b99ddc7e3d2311beae972e69e0eb1ac09196f65b4b3e005c153a8418b845228f0d79c32c003f42dbd1da137b84e3b66864e120c5c4964b7443d4c7ee07c89724dd6f022683d0b34427b2d2b688832a3992cd8051e75ff27758c9da257b34dd6075dacf6b94989477cac4aa98ff0d5ba877c0bea8e36c1661fbf2ef43ec10c3542720dda8d53dc132c113a03bc6cc560da08bb466d0290c2bffa77c8e674fb191d2cf75912eccabf8c5c7247d6d1d3957e4f46cc6b0e7baf2860e26dff75305c2466a3e6ee8cd88466592682a1c74421e521e49d4441eb585700cb70ed6503969589e165057d9d46107c0ac7eb67fe65eb9fea420a69faa77aecd25f3d5e627bdad31617876c640447f7a541bf02afc9ead1a8815719c140a8428ff1ca6663ae60357d70e376720a6e42023cd0c3dc161398e3b3444b87ed0fe624c1b8455c06785f87f485e418216a82a2da8bf6d11b3cd922cd0fb066c961967491a33bf802ed7b615d8873113556c142a306f4190658bad9c4a65ce0e4d984c0301c05defa87dcfc598b82d82fa77f9bda789f22769e09ba3cd89852403d168384e9ea4fed6a92e677b43e2b3f9d29980e3ed1ca60244389173711844eff5a110ffd8d3ff0cede978e7b1e813165461e0e330014d236fce81640fed1e911237b36427810508f63f0304582abd6a3759952e8368d3e138fc7c2087dfb28ca2653ac1ed3009afda82b85e95116d2e37a94b8972f8e7d1e6c9df8b7b9965476e7561dc1d4fd1ebcb5918966b77284bc5bec62c42edf1a80581682122d9dbfdb19108c9c0cb0f6c8655068a2c01457986485bd0d0a9458195698be6db9f674fe8f20b36e154ce12fc50ebd298adf4c4a0b21c0b75a618b64e8e3832cd47e81c3823040d54a89a1206a8c9796c6d1f8e65d3e62c4a63d075e03bd1592bffd3ce96725eebfad38739464b8a64d5c3b8f99227155c8f04c6d637a693ff50dccfd4de4251aea6f2e25c526b966966770615e97fd01ed6823f3337047894dee0bee80c6eb661450a038e6ceba8b71394efd7e7d042386cf9f2e2ec3491d88410eebdbe69bce560639e66cb84d0b4652bcbcf892d46c18049b32ebf383b57dcd2b90ecadd521b2f376b1b297d7d6542e31766b1a8932d172b94c8495d5bee471aa28279733daf015b019a348129714b8baa5a6462a51d9123db8c78afc7a506583aff025c200b6797fa59868f5e67143be64eed886a6a1a3f5849514d410a085cc0bdcba1ad838788ccf09f63ad10fed9b5c3340cadbff6319c44c2da3fd21dfb67475f371d8bce2f6006f4dda27ea6f2e1f4574ab607b422c3b3280634b526672fe8c6b0636d3d389481790f8c857930e9da3d1c2004b2bc99c9cbf7554feca2a398f0db4749fd77868b978ce40e8a998192a8ff2a7e717dc27c35b1026d53318928d17931c3ea55e68cdca8cb33b14b3e9928e440a30e2ac40fec52cb1f5d19c23b579822878645c2fd0edbfce08a061bc939fbfc301781e39652263cb572a1a73c924d4c3612dbcef4c24e6448f19357ddf04669210dfebf943f73a70349dd8743e4391b28596246c8d1dc1dfdd9f100edb08218ba4cf39c351c291dd3f709c12c947fd94df6002e72725d8ec8a1320f69fabfa2a1a8dbf68e0772e9cb5c922f46ff1f0c4b5473538d6742a8f63df89c31f533c5b0a712c7a5ec6f214af32f661380bb44d97daf4156900a4bd53af5fecdb94af5b7827fba0e59d9fb537322d38408570465265c937ae975ecdec91a47f4c3de97e680a9623d1ddfebb87393e5c5f4770f64d6f10a4d9c6d0fdf81d999bacfe3a8c432f36a6f0799d0ed1473256ae84d2bd982178ce71540fd511ae613ed226becb34607d833809bcd1aff3ba12278b46b40225b6a2a81dc014a1b5f430cc8851c3f747918e579db4390fc317d2f153e9d8adc8574e7e7d18a9c922df792ca7002b602a7a5ae5d0ac2e1b6b961e1de14704a5a6e629f0d5dc0399a5b3456c9b50cbf5f0ae2c4752362b8dfa418148320bdd996807d0e8a2d5d3ff4fef416fb64290c679d6b3df58a97d50e287fd67018ad8b320960d7c1d82a11824035c1fa8b88902e297d7f16635e3b6238f4d31f7bde5406377a9b8df6412a00123cd85b596d5a6826ad30430ef6d67ba1f501fd55409a00b121a9042b73bdb58c7af0fdc3855982fab19b57bff11ebc54311f4faa21a476c449d33c14de0485eea85960eeade3338e2871d0c3769ed1b12c8130bea1df42e042dda6df32da7d052703a157ee43d35fcab357275ae010f3e0a21d95838a8237e6694347707aed43d0be009a0e57cc062c09ea2a22da5318e231fea4bd24ecee069901116a36c89f32efd6b860673cc1149f799afdc36d9790195fcc54e93b3ec55c3f157450fa83fda707adc5599dc61467e1ce4e7f2a09e9b11779468857e0db15958fc66dc397e42c10d8893d08a49b208592f8e9d61f24569560c7c734726fe99628;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3da22a4606290ed3e367c22d25847a8c2552c4caa8e1593218f1d4d369d66c16036a05c6fb9a7d33c836b2a1311d09616b3aed71eef8926bdcf4d16dc4d30f67e252ca79f526041776e5412001ed5bee2a49df9df311b674e688d164e3b87fbdbd18e89f97c4f363afe1807fa7d9f2ccd8306ad105024384c4bef2486b2c5d0537e1a21446d6e34c07bcbc5ad1956e0888aeb1738d65bc63c96d97442d17d92ae27b53969b040b6b153ab3ba4363eb0f4a12e8bbb05c0b7f4d8caf6a8cebd7ae07bd95f4eab91cdca496b0aeed11aa69c58d3c68abe29bd2aa1a010cfd831e06a61e9f87a827c9afaca903e04cd55615678b2940772907ef7ed5115cc2ca190678112d2f4aef27baab03448129856698e0e2ebc59ae85040c64ccbe58d28830b452c7d795a375971fb34ead0d6a9a059d91a3e0c6b9b9be252f49861ca4f5ba9db2eeede75ef45c0c435aae9afd612a26e40802685be36c85d9e289f28246664d07abe020316a91a219a427f3660f0d51f594cb2513b0d87e554a5a0c20f15ac8f44a711ab1c4e23316e3a8f8753df4d518967a070c75fae7a4d6a3be11607898f18f89122585797a88680ef6813fb803b95edfa3ea0c92d04149ee67bc43fdf54f26352aec306493fcf61049440d1491e87a5c0356ae16a7336d75a5141600ed8a17c41413fde909b3998a46bf7cff76de56eceaa44917a8a28f2560d661d78a63bd3d380e6f887ce4b6c6cfc2d121d584fa5237c0c0842553aec927e735a59e022217ef3bbc6c777c3476e15b372a8a67dd20c38f2a3a5a11f2a4cee94ae154d04aabfe752995c162e0ba18eb1229e857e3aafc366d87b9377ed1e6cbbe0f1aec8d9e6324e4d93390ca2b6b599577719e4c0ecbf34c555eed72ac7457ab8dab53504941a58cc7916db4d6b85eb3e001f48737d71f4d4c88d8430a3ba0fb843277fae0de75afdfb0131af5963db3629c127e884ccdba0b811016b2cdd4d2eb99145f369f20e1de997c9482701fcb8cee78504032edd494fd8be21292fb029078ab38e3bdb826cd994418c584b6e9f72df0e629e829621c2e73d755f1b9ffae31f0e0087ac79be377297e5614da365e2db65311094c73e6acad81fd6741851bd24cbef5ac95dd694c41fee74bc9837a858c0fc7f5bce8bb27a6ecdb6db1605da570d1a5fb08a0266e51947e5ccc112fd9caf1636a2c00072a87a655188c9780d7cac2955a1d5b7e71a384f5bd774bdfc5aa87dc228781338190415d8f5457a3bd0e0dc16e20a2e98f454109ea73e58a85f045228c12910000cf48bd6220db084a285555032c5eb49cdc43f4d70194046403688f451e621078f018720c4710d08afdb53ec44188af2dcc8549dc3afda5e6d0c78001fec138daafe6e509665d68e07cc0339d0616d449e7e1ea1678c45185831568698580db8ed09831052232a264ba682804f2387827a502b5b38c4db771cfeb0244e3a94272b886337f58ec8bf950572f4ae0851abcc17c5ce03598fe157a393f487f64ee97303ebb0584c43711a7b1bc7c3284b519e5562ee1278ba38386fd4fbd97563fc77d8325e8ad570186ba6a40ac89c46e13b7c62eb1b665b3bc05a90b6b1018c104b92079b02b0f6ae8291ba194af58bf0b229b06083e4ce92ec8bd943cf0993d283e136216de4e4b3c2d7a3e9d399c2368e1bf77e90d515440af795e6cce6e93705ebb06f35fa84787b20581ba29b183490ae1c4a611e2545f1ccb0a7c900a54dad3631496d4fe918889f7fed677179558f7ce79305eda3ea32edb2312d7682b57552f5b341755cd5dad7745dd4ea3955ab6b456f944201dd985c786a38d1e25fafa6ee0504cdccf06d7180999f4a24ed297d1e267365177963556812f6c537a45eec9ed55c6b19eff06e51c52b46143a0957988de3019950f182b0a5f17b2ee9a2dc9f44bd1749dba8e13b0d5f6df59d1bb2eeb784b4c8d4779d215d4a03735c0740a2fdabd5e38a0be044eda0bd3dc1522d368e997c859bda6474daf81d92934b5a7510edcab2a3fd969b8ee65bbc4bd9f9a06aef61a53b6bcc3426257c0dde2f07161cc8a74cea14dfb26ba9625c8356b3d84383f2684a4ddd67bdec4ee927d4d67605327174b8deb6e39b98ff01f33873c4e46d7b5dd2b5d93e37b8f4a9bf3bdd7c8efbcf7f15160c1694d74f221720ef98883b2b2a783627db1d5413e9cdc12bb52edc1b9f3ec3865a420f10bd9ae65532a2fc5cea0b9cbe6298bbfc98b1099cfbae3e0d79d74f64749d4fdaa8ca1419c82714507c0056a441ea90d05bc597ff0057dd75bcb153384937450d021ecf3831ca786d92304c70ffcf783cb9d4b0357bba51502f27d24a224ee156baa0ccbb06bb4a624955bbaa58588a56ceddabd509bc07c53b524f59ea2e9929fc1f80a4a9d1b75998b1279a58813975eb361f5ed887836879f75fbe3c27ff88d5ba8335572a2f8203dbe1b284f445255fb8d193aff86b47aa2a265b8cef3ac751d94dbce059c9cdec33ad0e9a2fef86ea810d346750c43d83e42a09d7d07600f036d1d91f5e706c05e7392e432f1d554876301805f4f7b28671b10eaff777b5da7f117b1a8909f63e4e0a5c3394bac709fb8c0a4795db9506ed493b713ec4574f87c0a8fda3d842b1100df5f1395aeed31a0a77e3cc258fdebf6ea4f529c3cfc791aae830cfc6c4ba17c19389bcfe1d88ff171e1458625f5b2b716d860b6e5defd725d7d0ba1bf7749ff94d2ea032aaf97344774a9008430f657a69f6bfeac33a106ead94c0e246b52d600bcc7ff6e7ff3f319b307e1695c8f4cb8ff62b81d7be1992f099e2c85faf22469b121996465185f7cee05ebf9ff80abaefe1a636d9b5aa06cb024b9b7d23fce068f21fac035a72a3c936d7023a0ba0943b01eca5b0d5cd1007303becaca1b1ac209fffd46e86ee2f39e51baa54358a5d4b55b8a76e45edfa5b533bd3eac17b716c5c5e504f96fcb471274301710b647f5c83a48f389a00fa03968c24ef968b6b7cd4c7825edb7e5960720765400a626b6cdd28b1caf8fc50354193b1c6ce7f22626423222b51d961c8039aa2c8ceb24abd92c7c1dbc65ff17b5a63f452f4cc61c1332246cb0fe75a54722fb66336182e302649fdd821e381ca235a81059c5eec3ed5e0b143ec7b2f5ea601eebf60af99f26903840e5cf0d5c8bd43112ac04178676881ba4d95e9034728b69e8e24e0705d4e843eaf4ea7fa6349fa4ee6e493f5005f710b6888f325936b7245d11b0f2034940db5c6e7e81d8cfdea2c59f739f2c4954ef65c13a8036d8a48b0af76c387fb29c7bdc520d1f6eaa2af01354fd1de8e74ed502f15e5e1129267a10890da30486f0aa4ef50b3b77d46322d01974625af7f8328f844e30b0481ca78a69af134c5afcb7f01cafaa80dd4d1efa6d280382d2ae440f40294d92255f5c4d518e34338b02925afb1382889c1dc2847105569f7ca5f733a371feeded4367e24e590b20d4be002faca56b4a920ce0f75bf571a2ae37ccd239b21be994f704b571054d9ad7099976449376f248cd693a1b54897e5209d216992e6159a2a59d3aaded36555878c4a97ab019b5ba7db72fec3faba89c6bd63fc43b747c93119daa65e194cc83e08d62bac47eacb1d55743049bd41a57a1c174a9f742b641f032c3b1f4a22b33c1d26ffa06c3f2bc209d6c402570bc58e2aca0556c876087801c4d30d73fd1656812b706665a3e1949b32d322afbdf8d6f2dcddbbda82d3aaef03af73147b8a989d577e250c45f14821cef2d794a7beec8df85f233310930cfa08666ee25edb7c13f72aec8d0a777e16c3414e0e20405e825fe382f22d0fa0751574530bdc0fd01c7ce8f79cfa0045bfa9630718237d916e3255835cdb5a65f84c088a10709dd2662e81468364a8cd6a53faff90fefe35e0434bc88db7399eaffd8325f514a4f4f50ad5ee804fa2b824539d5e7f81a1fc4758f52420efbb214bbfc776df58cd556c93e254abc6d5c700afa281125d9e6abda4ad05da8211d14780751b9518859a1937ee980a552e941f5a40f14865bf6dbf3473b6a9bbc621c5f856941cd26c58288956cfb908ede6c2fa7dc39d0823e83d56f8e9909791201cc4de80cae82ca7873e3915b98f801834acc71a647c84f18454f91faf11558138bffd7a8217581c3c0fbbd8fc2ac14476ce5ca2fbc454298d5f461573cac4e829750bcae39f4241885dd4790a85d86e38dafee43c3ac46cdff3cae7858bf27a35c7f5f8dc833e0fa75393983027492fe0faea2a78d84bfb4631d11665ddd5c1561df47ac56de74a005da430d6bf6301f97d062673c17d2747e739637d2890619a8b9188f5c1aeb9fc638bbadeb02bc91d2b6e1d73e5d4d05df21c088a7085befdd44f84a372491a034c42b6feb62336ca2e81f6c7e768a2569ac1facf932f863757f6e4aa2274cb6bb55236ee16df2b0a30c6c50ce5976fc84f01d0798d236b274e283c16b860d4be2d04e2f768d9a61af0bd789c79553d40aeb3d30c8773c3cb2bb41da693ac67381d320304d138f4eee69b5f3b20e9d4aa59fcc5c9cabe18f0a377b2b6fccfb8e77acb738742f9be821d86f1bcbe9558c049036f8aae99a984b8a7fd282549d564082dc2817b3af6c906dd72f1b89fc8e0fc47607b26082317fc4d719f88ebe9726cf8770ea0701eb384d446631abe012fdb7cb535734e6da2f5c811bdda8aa888f7fd6cc946f2d78c8e64a146252a0a2ff11fdc1ae1f080fcccedd9c67ddcb80a53bd1404bab9ce5785a991ed2fb7f384af041f8ce81ea0831ecc55040d06cf3cb37e410e9eacc78141199c2fa421947519fd029ea23ed6bd1cf4463861e9ce0de8c37dcfe4d41b9b98f7065e8507e4cf0758a4a09a5fdcadf1aebbcd52ba774f092744d4d5e0c2312b1a1beb3744692e41df7e6d5bcec5a526aa10e0e1221ad24c914da86d20e180db2961340c059a7c2fee81df8b1d0d05c04d7f84ca15027690a7b605f55a085299b25ba3059e567f4dc1538982b4e6c3b95b13c51b9469df2defc9f236cca3fe42a04f325538f96467d4d3cdb755c52ca215405d34b1be776a3ff04204d24c224b8fe2ea3b7983a6794781390edb928c96c792b0e2b8653bbc0f349cdf6b9047e95884d8897399b9338c664ca8d4f5d79aa885e48590c0910424c4b6b543f53f3f62ecb66d1c472171a082b653edd335a5c2bdca720f202969c946ced27668c14c9bc8e0ad4b3d3a319f25439d7b0c59cffa012bcb022646474a7dd1203063b678b8a0f193867f1dda144203d2112a2e85879ee90ec74a472882c88c1300eca050542f01aa31da1e3758facb48ac7641dc0b11620bbef59523700b9d7b490e2ff341ad39c7cd18aff621727a0a7297d815c290c40c2a6bb9873bdbeb181138e8b4c15a2c7ad39d730f9a90cf7a13d38d4ace730a42e033dfa7a1ab3ee3e83b07b7e8d3e5061ca1cf22eafd5770a4c750a2021cad38ee9ec602d6b6d04a816e7e728b53b2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hae5972b9accb6dd5a0b3f71c1c8ad84e53cdaeb0494c37350ed1a188484c574d61701e590ac8ccd672ed9f0abc7bbc6bb78c615c4f9faf08e2ec4ff33bfbd2e979c89a3a1a17f4c82bec4e5536959ede321fb7ac94c84f03c2170a6bdb99e9683f06ff9512c320897a8d8cebe62be0a3443b10ae3f452e2baf79a0bcd21836e4e46aba0c3b7a8c1701953802ff16478edcd8de4fe36fbba4ba89ad2dac3bb27e003fc0328a1ddc33fe13e3d94ca8e8f8be40ca200d64a8a8894ced301a3c1c7f02b4e16a0f5803dd9ab7e48f386c0916967678435288d06ec8af6c0696e739409df4f1fb05caf195da1d84d15ccc1d1b8b287f6bd5283b35934eb1d5731ae249d5930630d2460aa0aeb7f950f8bc466c468b3863a0bc0f25f2baa4861be6fd97f4b42264750626f62565692461d07e3a636713a2d47a51c39b23126bfcf496361018199467e40fedb9cae91de9b50b820e65cfbef83a60a429112b9b3ebe6ffb63dec91335dc02c299e3e9fd488e4a10276b0f31910a4af44d6ac230c44ec16f1f4e4c289959479ed4ef140773c53e50c34412adc4b764102567bcd942e4899e641b4989536efdae71bd6dcf4d59c83a76586b9bc7c54e6d9a2d65007993dfe13bed46010b8d40ef22b43e0d34db02e2f48bb1b1c65b37b7e00aac1559cc8e7d9b6e3da72d774222c69e27f6b905b985d571f1786ce8f718686004546ea0711c03c3d4ea6a00ad7e5043e0267e3aa2f9e84216446bfdabef9b4a8dc70f351fc6e9f37c23d4e1d41a480022fc92ecb540da99160c3d3d457af40127d389c7042b32d9150a8dff7024da1baf4d35bcac71a3ea32ed7664ffebd78e0e4514efd6a9e0d8a462d450d06aba9b9ac213b382847f875e614ffaaec1755355a1c4be03fa5a14c8d5abe4648361ca0397a24e823683d801f1d85a80ddcc7774f6fcec05bae458c9365453c59c2347547e697b8c8e2eeeece865350f86478b5c27f7e6300096ce501082adc7e7d5b9982fed79b97e3b01929b2df9c7bac7076bbdf4da76fd3a85af651b41263851163f1d2d0cc1dfcef457be85839766a129af5db19743dfc8dd58319f35bb1cd11e991639a663f5363e7dc497c072ca2292635b9a3a74f768b939ef579a1845b17d3af64bc7fcf7e33d82efafc35792545779effe5d1fa2cdea3a95cb33e3b13d7c02e4998c544dae05cd69683567b7613c00dac85616488b8a45c44a76e9a47870e5672b84173491bad1608123ec21739843bf62e849e241726d677b4e0cfcd5403e9fe41cfcae8987bcd9bb44d600eef92d97631213670af438d03e2d399a5afeebab82fa6b9c784cc8d3c7519d46d8630f4fc882ae274caaacaa407b219ace045af40ec31d4fb2a7fe48dcd037008fab26cbb4424fd76a4f65a1ee26a254d89fc127ce0dab8123392fc493f2a4ada84d5240ab3836ad838a6ea7fffb6ed4615a504372473fb3ee0c1dfc7ecb60898a3437dd066f539dcb4f9e2f5bc250c26583d3ddfcb750ce55122537cc498da467037929ec05f7cd07cd3060fcdcd61ceb6ee765eacd67550350e6c3c15c7196adb8a774a661766edc8acdb85850b47ee9f08cf854d275c785f21a38c9ed5a9eff2f394616f7bbd175984ba99fdce58c4aafff11f215f084571d722c66abcc891a085f8f29c88e9c12406fa64e0fa262ed68014b7346d3709654166f9e865d496446f83395cef40ec23344090875b240a974e8c05a45fa01de1f60c19207ef3f67cae183e1ea595c465c63fa71d8a0b4fb780c3cf5abc2051fcd9925fd52654a0156b259f807b188bd0363ae0db44218dda9245d5688f74183014ec88114768674b8a3e1bea21badca88b2502b3e1c24981e0f185cfc65964977dc77e0ce60279ee92b11840b2338501a69b8f35f1df46a8e0169cb5a82c771c1dbed2900e742b20cdfe0c429e28ee870e4604643edd1f4e3eaa93c4c6b5bc5bc13e791f808586402869e5ba41756cc796fb96ee36f9efe0380076e2cce1282bfc1c71f1d2c45b4d58d511e3d02ad9e5737b9cc7aff4e9de283d62076c7b2b2b2ff6edced54e09253ec4dcae6e4a3e0220ffc12c3f5b8721a626514e14da5bb51e2602b3206f40ee80509a51dc68b28a375ab71d888459bf4fc92bdd357f7167fd9ecf869a029faea0df0caaa6e6c420a9eba5947875d7356f85ef047822e4dbe3783d5887f5eca59c191e8bbee0449aaa73cf2dca68d015588759494dd22c539f40665efad0e633f0d89567fc92dc1d16a79bb8cef6abc122b088e22bf53ed3577c785b71a84d2cef167e6f161f1a07795099f59f550bd736c4fa11e84d14c62e951c719748ca4e51e90f580b195b503926a2e04bee141e204e919d5b987ef82ba6594b24670c992031435a08c71b7a0cfe8609b09f36bc9278e128581de3d76ba80013a03be01dc9f04cea7d283312f56d506f2828b4b50362edc829b28cfadb639b988ff9a3b98e03e8d1a7ad7effd10cac2d5bc5f4dffeb5d0fe0ad1b9df2ad852960f0ff77ef0bdca2037314bad74f1d9a05f3a0eb2a1d6c653de6e0671075e88a8bf802c2c0aebd2a44cb41d793df991998201f726b6975f7e3c890db7edb8cc58cd4084ce252e851c9d6529b357da924ace73feae21c131f3f67bbfedde0365542b62c7054a5cab4b26c120278a46ef6a559c750f7c512fefd1cb5b6a02619f5421fed7fac9fa6d5c2a8daf1bee05b3f53700ba117cb2f7da8c5bc66b525c77f599b69525fc341d18feddb6a5a375507d9026cd5033777abc635eb5d39297380c26f32642ecf99a87f6b15ffb153d1c14e7fc7e89b3341622fc96384d5f3d9ba72a5d6eeef02a3549f4ce1e04efd8faec1f7af330fb1c380310e5f871ed9f3cfecc9d37d101f64c03e86d68dafdc787917c7d10e1d04673a71e3b8bffa2e2cc5c3d825050d21c4a60c28e01e8e25de492693ff7c08eaaa1ad2d486b3af74801c947a26dee84a86d020b689fa1ffd40278923820d93898c5d45da675562df293dd1e09377091ecf287b9b060776bb0a89bf96794f1176c65cdc506c4310914fd59328635c347e5a77b2ba71cc9d0e739db52382d75c7d91f8271b4586dff5a9fb173a8a2bbbd02e6d1b0778a6e5c24c6c9ab0fc1a295dd6fb0123d5479e3a6e564ffbb9a0b93052ef65f9f6c856131634ba07fb14c6c7958806976a40c443c3ec93e6a05a241b8239b8e5c33a76bcbc0589e3f7fe9ed7c2b21f0bff0503e6bd9091fc463416f5434a4c01e52d18a4fdd112f0cd30a6fe7a91da6de298183296e0fa51bfaf93d231ed01ffd66e3e33fc3a723c3fcb454359124aa8a1b5bd2a2c85a2b3d93605c384e16359fb51cd0908c8744fbb6b2550b58e6ebe63e0022182865fd433f87f9fdacf56ba829c3da917f9700f43ffbb9feb5210ff04864214be414c245b4964aff1b35e3d9e9d013e5df996769001caecc14744593aec8e3e59d9adcf4c01933d46557d86fc657d56dd91fe22fcda439cef6d351d2862b22abdbebbf751822d46716ecda0bfb917457a980a08c021675b529ecfa4f2d2aa81bc3d86ed2818ac5fac82c2197f9dbfd5b508699cce67b40cbaa05131e5e0b4d5722ad12c3fdd993fa278227b75b35cc50e0b22117d6d676d6c7500250a016fca4eb091d94245c5a97eccd3d20a2a81dcd58fc5fd51311457a2e080402773839b0c3719f15681e12485218c1b994fcbe81ffae4e88025ae48dcef26d5a55f5128c1e1b8e98629bce47494dcc319be99f128470abf1481c9ad852fb62194815176116b481e426148bf5ca557f0969a29f2333d556b12c83bb7a165d556b701322e6159192dc89534eba4441eef7f0db3b72aba23a8eee0f563649603ab1abf874d13eb5b0e3f2caa9c409fa908c17cb8761b5dd5a15be206301d922dd554efa09b9058860cb30a3418e1df0e1d008228f9104206342aa7654f01f3118ac89f393cece3e7cb844e95359a022e831d59f4c6d9fe1e77a47ce1160414ebde38d79d4c7ace0b9039542961752ea73e2d864683c5f31e6f63f6f831523fcb7fb7513e087e7c63a426dd313ada31f146cd7a03a213b1fbdb93964614df8ff3951d22528b19fc0d92d5a7c97182f5bc5ba2546fe3374521913394b7c92214505efbab0b6f95927f2adc54a56a367126e50d785d04b4ee3b2e4b9549ef3c1e7549a0032c0a626057f92bd294b09b78d7b3cfffc3f88cf76eba3590006e3531219cff78241d10a99ff7a059666c2c77ab7e7ea7df75c8cee93c53cdeff9cf44cc315e6b7960a64e237f11940f7549d8fcb64dbd61c90ad708300d133c948b7d7c212c098ab8e0e08cd7864cd1f85534a00eeb7e7028d0783225f9d2b631e41355b4630e1b49e56c5955bdb10d252b92b1be02fdf2c4e7c2f1d401607233caf80c468fe2a5beb448b5d8dfd4cbc38e9c080c5d29864d4d7a08e4308a3c33cb8f3f6014096c1c61ca93d887e2837c6300add0f7d227bc9b603f13bb739b894be4c22ff2029e5b2bd94766c91568673139a5a418baf4d8a3d615b054b88d32d8ba50d72acfdb6345711494a2f60ef4b291206c6db987ba232678c7bac4677a731ddb241b65fb40b4ca4fc66e32e332fd5ab22ed6fa9d371c6b366c453a705fc5384fbe36d9ab669f907cfa4ba642769a1313f3b8e40050ef35e19d584f7163256ecdc4b47957c8be2c54fe9c4cd051aa09372a8334a68ff6da982e331f2fcc27bdd7a806341aab993549deacd5d9760926e2b821fb781d5e682cc1b3dc73b1eb01aea44cddba4efff23750fc405964f9ad8fbecac35a4f51cf197a991fb810a6da7983dca4f2a4645d454463bdda9bee3beb1171d642a286432adbb55972f1390e1eca4747af0c078f094ec5bafdf366543f5a6635f9507474410083d8fc3bedb0123328f725b4c0351567499ea0cbeab72cadbb8fb60ca76694e84d1d8cfc7c1a97d3e5b4bb1776c893d6aec50025c04fc329d61a0fff10f20d0fd790a25e52c106efdc583e4b7eefc0dc6452080561b1d6ca2b53ff0cf240192078c4c3b2538d815b81f66f930c2f72aca72c00c8c4a82b11fc64474e8c568b2bd8e96e0926b42b0329084ab03a77855f794548452c82ffc02da525a4e60c87516af866ac3e8111227edb34883278b9399d45e9eae3a99a55a34ec1bd631be507b503e038660b1a47d66cd6cc9abdd3a58310e2a43525157b4d367f548bec59c4a04d560c7cd917af329fddfea985ddf5728b2a8461a7a80a1e21f5b7368960022dd296910dc16485f651b97caf9c9b3ffb74f2357484d11aca1168b749782220c2ce9044c70200b997cde4b76c03310e0a54cab23ec18d22b5e45df8c1db6460a88e2393ddc516e7a8db721da360c0a39b06fe060d57322e90ec2623cddf6708325b7a92f52a47f088a4352b30f64b287ded7243f232e9cc915671c2ac8261e68533300f6a17710eafd7cd4ba63148dd3fcc79464e8f18b2dd7a6bf2f147327d2a05af33774629ebe4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha99ac0cd8b3b7824915c7b069bcd00d7a2265c7c2a1cebda33d71df71c9d178bfb99436b8b07f4635eb875c7cdbf316a76b63e85d7122eab49fa991e4fea1613f500fceffcc90dcfee33777b5ec3283365a668ef475febe986c8e212e859c46b0f15b232f9f09d573f4998d8509a01df9f8f482b6ffab149964baaba069e5b84440f447e0ec4defe53a32d5938a92d11900488ca6e4db3c866acdd5dbf014cbf37d7183babc704f95887a9d7a793e3f8c51ccb58e906c285dda4a6c2a8fce1a512bae4c6b36635bd1d329f8667ba21d794382026c321ec001dd4c07e842c6c15ede1b2ce0c5396939f157e4062efe9df58706aafb319fff477f7dd42e86eef6576d2229fd8b44d80210c0eef2f77fbb993f557f1e4f3711351b069d823e8d6e849ee685908c92000b54842f27f5a4a3444fc99d090bda18c421367a83c175fb65eedf6991b2bf8797228147c55e2d49d20d91cb3d2ef3b5b9004f1d18303bf3624edb81550f1135f0ded4ba102a56daa0d94579bd092ef4b35b8c5fceb1362dfd636729c50203bdbda462a60193eaaa7478922b753723c92ff6f1a19cd30fab251169687bdd7dbe9f461055dde05d7b066ae96c9706354a8463d083a613255888c6ca31de37a08118e4133e3f839af2ab0e57e03a7491232181bdb20e62ad47a10acc8ec03cd04d296f4ec4664c98a92f5fb6672b464cc6e7c00fb640dcba594634ecb7c7ed6c49d5b768ab516352a09922ad4293eef00cb4dc225dafd0d38401923a8959f94296cad08e8bfc005e7ee6390d700bdf61c9d221e3a37774228a0225f077e8d927330857ca9accbf5dac0328bdd2c6ea7c730fe07d80e90ccddfa705ef20a934a87895a0e926674ed84196379696ba66107f8f8c850c1da01e4aab5046a1d9cac11800cf58a8d466f633858c5427392e714387b034005deb64a24181d2727f33cc32182e9db4d9cff99dd8c2d8ca192fe93b395fa94f5543b50ec86d02a6b624d8914981dcc82cea6c29ed7436b6801ef7aef30b7e8d6cc95093fa82a1325505ea05166d1a6cd1fcc86f329d33bbb10eed648358cc115333c78c0b7d5f11d63c1824dd56a16932e37491f1fa269fb7a333f1c16ca351a322e425b4c4f835180b2b48153566c339946ecb87ad756ca1d0c7c6bf7ac00757edff630575e34c31c3edf836ce1c0b61bbb31ffaabf488fc5068cbaafa014bdf5e4d047623a840a45f68f23d0758f71a50c967ed5f538d2eeefa6bc9fb138bca8ceb5cd22ea775592968733d47fceb3c437e53308f46190f91042e495cee94def3ab8684097d58b18c5e8af0e673f0d07437b53a75f9cef856ffa028521c1ab53ea9335d62590a7a1a5c05508091fefe5e19e9c972b0ec5949122f09e476acfde935926f5d425296d44de83ca8b38f2f9e40419749b65e71361f10d78feb59c4c32019c990ec894b3f20eff8e1f97fedb51dafe3d70b21252e37d519dd7c6f3056a8f94e96c4ed1c5f34ff4c929c536f99a4d7a447250a5d5c3648ab005341036dbaf8bade547c5b8e0c9844725e2333897bc4e548ad164ed7a7ccf5316dc04b3fd86e903aac437f975c78fca7359224379e1e5dcb2051bbd6ebaf6edb38e72acabc4da90a8676f748c42df0295a44ec930b6e4732a256116547c2ca5affa2b874fa2965d24ee066791415f14b5b960ae0b4e89b5b6daf085803f792d69175fa04f8ce52db2035f20e52683f0e197e1b33f28c2608d5cb5a18c43b033b169b41865766ea3b1bb2ae88ea09fc0ff281019f50686de35e80303ff488baa828020855905fd50e8cf293ccd62bc0ae473afd36c1967ed0210f7bba5e629ef2a1e7684277dd6b402086435fefa6a708a0e65f4663aece887ca975f83c37d1c202f010b2c572d093b72e918a8c9fbb5d6d168b3f30f1c77d7b4ee9928fae089ffeb13ccaeb4f0f6de13bbf4b8babe62011c54b7dff61d97d5e3c30bbb052ddf53e06d4bd689b4d18bd23148acd555c3a426aaeeceda19f29823b5965a07f5ecf782804724ba8d5413c285f682e58a368e3cc6267ef4c16e2ac5a5e85f7aeb76e9fafab57a8f67ec97c8285a9f6e9e0d3f36355fba001bd7f2331e41fd30012a03a6c5a98eb8089f91e4d3a58f190e714e9c210f50f376cb99ae27a78c799f74ec2f9e1e3699a1ddb8961f09494acf70ab1691bdd212789f94c783207435ce470a66c40f17990230184b505265f503a3be6cdc10d98ffe95432bfdbb5441b751b3715e08824e8ca8c19cb49eb264dd50ed10788181e9a5a7f45a5018b186690f9d050d0d40fd3bc45acb96d0bf2391b1e49b0528f06a4f5ab6d850139471526c1f11e93eb1da126661d6b9b869da5ea92636832e68021eb93400c9d1429c1247f653104129034f6911bd84bd818dd90f0330ad9a4b7dec9d1dbf2bcdecdf10abbbf42d3a4dbce1747fafeaa3de3d503a043f61f20c306d15025e37ee11f84da86d559f46dec886318c81186f0e6c43d5394a224a45d57ad589000e8c589c620b1914d993947ef6592756c056f7d0d8e1ea8b6c975e483a1a6b8cdc1edb4a26007009df5bb0510eb669c2f75f808feb26688be71c96cc06ce23b5b4d9d1dd11635f8ef8330606dec4ce49013f684d91b7d4c11af59faeb39779755c8c0ccf0485f60d989c8ec5d05f802cbdb15084d6b23af6d7040c643bebe6724ce84b774f93cad337dc63decacac0dccaf658cbbf4e48881e9124cddde866a7891cc4c952151a0dc0f0a18498c61b9d54f491301b36a911134435ae17d0f002ce4eb482d03857c3caaa129ea3f6fad506a94352e8ac4525279632ae16f31808041d9ebb494ca15faaab6dae2ecbeebd2a03714c5515867dbe8e4ad750f4981c7d986c63aad2aa3a4465d59580928262977a3fa1b5d01ceb7776a352cee9639d73f843c9e3b8aeeb02d7f11022c266559b6e7586cbd29e824b53695c103930161aa385bbb72d2c09515e4bc4defb6b7a98885abdaaba0b6b0d33f3d2c2e134ebf84f6a2e0d875722424de02c295bba25b5f217c9e1657ed3c2b611d035a10e64c1e03cf4ae0b11e90a810156fb9a08ab66ba3f2491994fc9aa43e6db1bf0661911ce4d460900ec233b4044595439f5f73f4d5b07ca473b583a3979a3f813869e801515fa7538d0da075c2b9992ea887de26f3ee60a6c1ab539972bd90eb04a0b23588deda17423b387ff2f17e1934ab9cff1a0d574939bfd2eb6607d818f00b3c7fed8957805ab803c5119f114659772cfbf521fa39d0d7980fa4470e6d431cd487c27b5a1d25d9bda3e7536e036257f82910136642a3a0df4e7facf2a7e089249f1fc2961b80e1689fa88593f7206592011d3e8b39391ee9e5a090a8178172dee98dc2c0ed710f7ac95b38da23828e343236a61ee4bc45f74fb2814a405f06d483b6664668462bf7f5148e26ef18e8a9644bee74993ca5191ac5046be177d927bfeacd22bcf2347fa15edfcb0d365f828b76dca1a7e5d708cf4cd1e5b550db181214b8ea1a758228b40ee7c1175cbcf6e5ecf424298de8b10cf9f0ec0d7b00f8baa1d4dbfa92b29a870ae1837b37912788c8f6143def87361c51f1b08519ba965f725c0623a963e2c4978154920d6c9d192961162b503f2e9c7d96ced4f75b598f0b92158b50d6c194b311663ce3e0d48dbaea8d46b545ff334f5cc9ec30bbb902f89fab437dee8d1c74f90fca12f0adb902bbfa944c6ced94c9bb53f3130877c5e9119d935d7a6f2d21b48b0f6ded35418a1d2b1fbf11367558c87a69adf76c6b7d9314ac06543caa8980da1dedfaf721d4b62e41d251eb965b17d107c86be8afe4d78b3517d9a0c43dce8ed42408c62cbbf82bf9bf2d489bb65cbdebf469f2cf021c10fec06c92b68376e8af099d9b81af30a04bd372a16d92e7cca64cf1bf306b8c0b02014173a161292d66482fa6df16ce62902539349ac39892f915baf76bcbe0e828824dd4fba1f4fd907add4a169a87da1e7b82a879c0e1ce7794c678df7eba8b0036156eb68d1289e8f05fb1bf56a96065ed99b31cccd618a821f3b6cffa48fc028f5b2b58658ddcc7a10764cb2f456cc466953324c26469c6bba2a3b87e1d7d7ede9b5890bc0d80c210d4904335a6ef40547a9a00f1536cd2512eaeb2888a5f91f825e4119eac024d8fcb684035bc0647190e4f4e303f2027e76dcc4afb34f12ad27d901173e829561146c789b30e12ebf1b5de7393024c5647d544466d12693893f6284c9b0d7e7df1704b3e904ae4485bad78e3979b902e569f9b810423a8207200f85c88ff5b7163f06426d2f9cc8fa7674c3a3dbc95f83b8aba6dcdeab255a437f97ca6179b3cfc62c9d2c48309a6f538837b37da9873181fa2f4e075ec4de4d9cf6e7963f9b652b9fec433ac36ea4061e1cf927f8fa10c0e80163df5d38cb8592c323ccacd2364e8a1a2312e011a7f960a70b619ed2d3bfebd30367a567adc981157b02c003b25d0d90ce4868ab606e1ca82f9aacf93b628549c7af2e9e2d9bcab6244af435a35dc602e1782d5f1bcfb04934527ca1242b19a39856628cf602265f971fac6c22c9a55688857d3c290e948ccc210aead7085de7810f01b59a63d5808c63e1c0c013e176af7854db93abbc072bd781caa6b6161ea7b0ff5cc31591ac8ce2ee53322d371a8f0a604ad3175503ff7e21577f2bd5f1c4ffbbdf7fd22f292f69c9bc17b7791b7a62ed16cf2cb360af84afd0b334cd4ca36b8b63fde949de08205fd6229d6c421fa5744bfc194f42fd3d4ba5b23c7e80c8aa5453d0d7e6f6dc9d72b158da95968196178f1147c62a49729143853f4fd5caff4847b39d17c3353d7a466ebe686a19b9d80d20b61a667645c0dfc11afe0237488391e0bbad7d9ef9d359b4708573dc253e5c2108fcd25eb01f47292d194a93473769634e49f7d733cc17e224a2d58f1824dc54c9aff90a84d0940f7b7c93e606081420e902027b82d3e78edf4f10bbc8c0c6fdaf5e3359e8e707ca9c60435025f4fabde29b0497b322cc26bf8048eade7734132d3acc07bb70537a512e91bc60c74a7e87cc36f96eb104ae1894e8702253a072d58867f90c8c25cd69e35b2fd74be4f73bd1dde2d9a01a0257b806e494eeba1e13a92eaa0ef69522c7358525183d0e860ec0832077d04829dacbcb4147cd72c5bcb3ec1c22cee21fbe0518b045c12e9a0a64d0ab2b48c01e9eeffc812d866e435d2ce678b9659fa9bf26ca6b4c47b2f835057ee5ac7f627d096e5c671d3fdba33ddee8c86886940e603a88b75135ac8c19bcd24e015f7da2bcdd41933a64c16f397c25dc89d448d4fb2e1ecf55e868b36fe8fe90cc74d19584b76fc0add2204918b7bf9dee109f5f25955fd58277a1fba2bf3f7cf5ccb9c023f9728389098dcc7f56125085a16e5b9b68dd10c204bbde26faa97b108611b7f51cbc523c00b1cadca0fb5b86c6901506b52f77de2d174c4b5f27d37f3ae646514ea91f2e22ec1c43697b894f6788;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha515fd1c5ed70de943a47e2c49e91d48fa5cbaea994b360c9706f8ffbe4060b82d6d2ee7147b4f7eaf10c6fe63d283442774036fb83d0e6a4bc5bf43fd7932b2634a4eae34ad17e1e104c43cae2e3722f602e817736fca9d0748333fc9481353de43027b5081ddf109db9c6753638798059ac87ecfedbbfee0883e49c3985cf428fad56560fd8f5bedab363e46dc32046ebc6451d43eb713af61d8d299a52662faa1ce254e1cc004f0b74e93b8d572bbef74593014cf0f3f654c5e7d18376fd57f01cabc572254f3bc71437bc3c853ce6ad11e2746b4949e0d27f2be20611e89eb47d5352daae385400cc0c4091865a4756e1d0c62a4c3640ffd6f569cd210cbe3dfa43adce433874b6a9ea63c3b6c1b12103b1b56d1e6f1bbb1c50d042979457555215d5196e96d0d354577dcdb50d72dc0fb97f889b5deb81befc5f0295cd47aee8728ae61f0f3a5cf0bed167aca5755069516398fb33ebbe2c4d9556648eda1ae24d8c3fa5e907f3cfdfafe7c6644ae4b0d9ab12edb487f3a7ee3e0feb6d504627c29e482c67a19bf3b0a9372fa73c1c446501e18b9da982e5c4cb4cf21479b49e07eecca429fb4a3de9aa88d2fcaad182c95aa125f0a69a2e3cbed3dc4ba2471fc0a34a4fe32900545be30f1cd5adc349058510bee6ce17de071e775d3f0175f42b4f360e6e8a0ccb68f7498d6874d5383dd7c98e473a016fdb18cc088316866ec80cb77b2e3a1f5db2fa8c88ad1d84d2523070d4b1f901670cf2a4b5c1eadd620a57e5ee5f947f56f5171efa473b889f1829114e6f768fa0a52a3651cc533f801def987f37ade1082065f24faae71216afc339c5762d0bd9fb31255f7d8212b08fa8b521d7a482c250f277a4d9283547fda5eac9e158925daf5aaa17d85d037d4d2c45a8db27ebce3ed5ac863bf5c145b1fbc7a2d403516574c09b5142b559d9999d04fe94ce19ddd96e1099a99f58c3725dc730ca986ac341b04e72eaad0175e5e771309c39fe4151784abb3cfa2ced6ff0d33d05720a7a3368b0f3be263f4e40433446890cf919573d7019c42e228ea0dc5a925c9824cab3b150270d7ebc3e497323a8a47fedc8d60a61a74fd0f2d01c1dad093e07e7a6f82ab29ac314783435471b23b739e9e34be3c4540f714a2ac74ef36c9a2376ec373cdd83ac4f4739a327f38989dc671121e54eba278764b45a966e4531f6d4bcb47c65d9315cf9c2f22d25e8dc765ecf9063b82abca29757f99d84874132b8930b0916e3ec0b37c72c4549213e8529685434dfb30e323423da805723d6baa3756bf420f93db79eda38a63ec484989cc606f4b92aab2ff8ad2bb8461459d4d7936f8f190d54fee4aad041c7a5a2943c924c43b4b226a052dc05738e6d58468bfb2304f07ea160c9b83bc30d92e0d0278e69a3def87a2f366fc45b3db5f83f686cd9ae42489b00ce8a8c217ed901ee48664037d4a3c944201bd098fccc03a94130a97d45180df1bb400c64ac6bdd71a28142e4a283b4eff2251f85c6cb935e7b34c91686f6ef065783554d01f6fc3a74067032f55b4e18e701f44fa06881d5a486961dcc976de24a9e43b9b7d4597110cbef768ad2eacf34db9ab7f98127d98d107f8c46e8adb80790f3273939355376bd4d860b65637356dcffd76e117b1d76a1ab527fdf5143fa2a7e3f2cd5075e167dd3c4f57aaf9aad640395d93f37eb5ba91fa24267bf0dc85e36923d975f1615cfdd455efa99dfa2c8f892a31efde505fc9b4bbb9b4d9bb88b465258a13302a7076ce5c9eb65b92bc22d673099c20e55bd337648492cfe0936997666dbba32467a0ca33fb1e9879aea37a85f6c740bcbcc40f49b2a273742bf2c4fb23411715335567f5b15090508cb6598ddef9fb2912f21b79eb3931e04a26aa6794b0960c6cea0f9e4553de5263a526c50b56d485e1494912ed02bdf72556c6329720c7f2f0322827291bb970666c8f98a4cd8d1d7a26980796a0e323ad37f5fa2b06c1ab8d99afbe865c310047eedfffdca14a49b9b45455306b01ee8fa937c7390f4fc6a7a18760f28c9abffbdffeb10b208692c332852c6444d9e99d0e70c4ebca9cf035a8c28806ab88096b37ee7a174434a429d4b3d9650cf5f334206e83674cf5595223b1498ab128a02eac02135f055f38bc9742d01d189a4bf435e3e4be59689cac8ac347797ba31e339880bfa8360c615cd9cf9f3159a97b465296d3ba07b94c69b16bd4a8ed2d497439baf284e907d472b9444386152f0a3913dc989b7ed8211d1ff218ab6806ae8e66b3ba4a534b3b3d5bb5ecf1edd32c8d5e7ed4bb0c36e931f591cb966f68bc8d67900a8807bce95f5e72e3ad80eb637c513671d32acc25613ee91651bdc8569a81f2f3eed3326f08061dd1277007bd7d3b698265cbe2db0be31fb601a79bfb2ab70109e649cbf2edd20e3c222a9dfe227c5cef8c5e02a1835fae2b61568436b848785c8225530f91f8d1e04033e5c7b4c6f6fafd8e61b9554a702b6403322f9a65ebf5eb044dc60cbbf4852d4ada3fa0e2a34b4f0f1b7c33b27450a16cf219bc72e574162e171f65ea989a216fda970a8541b80c2a05121a8de69f445f6c64f0d3f7db73aa99e76b72de2df28066098170212ae025c418037d8ad9150fd1d3684d296f695692b7dbd393cf4bdb430f8dd7ddd8dfb71c0ff45e36d01aaf1a595d0a26b275f3d08d2059c9118563ece6115be172f2df4625f502a8b2d5fa86f81f761ae45a34847c2938d7386103c81e7bcddb155e1c8ecef5873f49a70c2aa0449ede682af0912d77b914babf9169b782a5961c45b5ff948e6f7b41f0ae4062d157a20705f792c14839f7c0a6d0b75d98f1bd8e0ecb04738c471e810a0679fabe809d5267c97d2cd2343f41c6c232a764276654f6d537b0fac9df1f5ad853ecd3e99538a8c05ddb16550381b9a8a2699ab0cfe76179c139a71a69c061416028b4bee823fcbb98ea534c0ba170415085ca22242a229504a6060caa26aa449a2c89b9fdefd6053de17e769f4082a18adefad93223eadebd7d79ec88b9ee3e92cf88d1c840247dd60e52030a4fadffec7515f5139883fd41a6ae48eeb2dbb19b07eee58939bfa3301c10a90f6d41cd2227bc4650a6a51d3a211ea2aabdedb448e9c68bdefde0dbb8b5e4207c78021d682e8596e419d2ed2266035c3d7a85fdd1aecb22044eb111796bcb46efc9d2a56f5b9303c1382d0344d38c4f258ad5cc76869f645aac1dec35023ee241aba1fb40088588e42b5ffe81c34e8b7a9808c505126e2ac609140cda7340eaad86b55b70346c1223c39646e958f8b70959e7520e0116902857ca52b1c19a09b00114ea2bb2a236a6cac39d5c490980857ccd98ab8cf4edbabd89f52bcdfc9aa2fbffee0dddabfc54b9ea4e4c04de29cbfb18f40d30b0b40d64e20b935e3b89f12dde023b304fb9a2f7d2947016cc135e4ca1003d59defec6623c42318393e1e68808e117659087b117fc8a93761ab942ad3c6bfc538f145abf9505ac2b20b1f5a5a906e2504e6ada72ee4b5fd18cd2e293d5e8ac4a00014c272af9c1654c33babff5fe29be1bd8f4fada75dbc1615e740975dcee18be7bda1a8fe6a9aaa9e08ce5d56fee96e42306f1a0b36955e2ad07f999457423571effb7d7bdcb74e51233de7f7ffbacb593255a25ac41af24163ff33b8d9f83017da83a72c012f01c6e671599e55cf714211fed27ff73246d52c99e0b0269fed384da78e1adf3937349109c9f5c34736c37ae0c5449a7157e253896700b1165ef3464b4fcfe6a12b3a2a98223df0b8fb5d838b48680450e6d121687ea5004c6afa07d357b13a18bd8b82e505741529568edf56571fb65832fe50555a37146f80fb6c156f1cb0dda6cf172b6f6b800f20ba833b024b2f0504f957544cbe7daec0fa40d57c8db2ed320478f7c4135d98cc58c39273d6d0e0d43443b36d313881a4c097a4ba1ab60cd63e0e2b711f53d6136251ed142105a980468d54e7e47de62748da847d4618191e9e6245f6c64d7c989125f146ff0a64071cde97db9a6a2c4f8afccfd884b5b4a3d866fa984274ef52111cda728a4696881192d95a793152e343a282b1299759ac5269d7b667beb694ffe7cfa6335f779fe3481c87d88bd1b82e20d40db02047b36528e1212bca4681ebecc4633d74c0f74e1e17d418e77128d87e1bffd8f672ea3fb5bfc5fe6a5459885b840b8e21e36773ad22b64624672f15fab3ec1af4e97b1bf6567bef9eef8b370df3ae8be64cb6a66e979523d2fcfaea86844a00ebeb4df0273010f4caf03b31d23f127d30b24b1ec5634cb4d736050b74d9eaa59acade45accd3827720da67ec462ae9675da804d1bd7a27fd2b80e1efe6ef466723d1171115993d9b3ac7bc06334d2995416d490091d41723326ec5e6f1671e30a35d4cc04b4d8fa4a6df59bb1466fa116441cd68d85213e8e86c077da1c636b9b0dc4fec7db5559eb46bb82c0c5e67c7a56c50451200abf4a821763e939ec3943f542124d6f6bec6c0e9a81b44aada07d85000e3ac9e8c5564c63b7f029d0ce3df12c232dafa526feef103f4b72bdf4464557bad1009b8d4e15df0e769dc4b5db36094be69988e515573dc20cd8599e2495a2437c1bc10e38c73691c9fa24a9ece73a1fbb7dedbade8f9b2d0d7b36eb60c5e44e5247dd94fe415703eb8f58ec1636dce9f0a8957a630bb36c955a4d11844f985369cdeaf39a5feae1ec2aa25c38d5770d88172aa1c770d4174eab0b6b7aa1943e27804838f99604c6f1506b6d418c60d3dc4ca0e3e808f6e8557a7719cb54fd2355f44acc37ff2e5b5501bb1a597216624a8ecfc9ab4dea5fa5b7c4019304366c76ec5163ec36184f568019bacc1420077d144c94db7fe00b6084489fa4c811abfef9ed71ebc40400c16eeb05945823813244700a44d4272260819b6bdff56b3a91c2673d63f39943c4534482b111e387ac4ecc08ba60b5a22b4ddb8260ec2bbc08bbc2db638c8f58ab716e0232c5184df721b3a5e9fc3c82a2111fb4f81d5d468fd7fce2d0cf1e42848707b80b967c33485d21322e8329af70299abd7ebe368276a0cbbf9a2baee4d3514895b4b271aac654ffecc39df6a94bc85a2bf4949f28de5b78c3895950f6099f47d3c123b4b70020debcba90ac4a891ccb58fd4b3dfcc5ce8b6c4f95f20959b4430bde019acdfae095543b3c021038fbf7081d86968d52f53abf0f913db82ef9deb1ad8dd164ae1e5a4108a7af9590ee03c260bfb01f80d3b50a705a73f8760847ad6d623c7d9a18f243e066239907e40d359bc48fbb37b1eaaca45ecbf3954c927335aa14cb597612c7864c95cf44251a895f3026f914149cb44260ba7d36c88f5ae5ba2ed8c4c2f649ba28c9fcf4641ea71bfafb1f00df4880e15c7d994f69bebeafb5e5543eb6440499395f846e7a45bbf1562d97901b67122c5a492ffc3de55e4fb751145d711f9c7e6e7fef1c1df89062fdfd3ef8e99563dbb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h6fb2a1740e5072f4b75b99d43a79757e51ceac5ce5a1d73e14fc9d62d1177c4d290432673e91d9db86304526b48ba3387050335133f5ac004c92a9ce01d9902a602512a7fa600c6599586f1a185a87a60b8924cfe31166c56380eb266cbf89ba26b324344829bfff0f05f5e5d5069c9ff4f77f53a74e480442d1e333a685c0e9266d5c02cbbe87faaf5549b9d43370d8408aa1ee972688d11390374c8ac67e54f4858758647c3dfe76ca6612496aff0b7205ed9b7f90edc716000bdb480d672fe46336415247ae1bedddeb901d1a73ef20a33bd34cf94b8ab533c0d3c5c68957dc31d8b23b165046409b87cad04a453f2a3264044b9125c77c68a73237209becaf0d00551a04c831bccd4a9b5d63804b57ae609153c0be01187e74e109a2afdebf398648bf3329cecaac5f08dc27591feef065dffb61019cc36545d723d2447d1cd677a7c27e6f8216b4767c682963ed12da61c8a0ca187e912b59c1fd428f6135ae7e11d58d01273b92aebca449137cc3e2530d7b35e03a3b2ce7d527e731227165733b0de4c065fc3ea2028579f45b3589715592ec94b4e2af8f29cdac54a7a0e3daf0a7f81e9f488a04d8a6c0bd69d12d07816c27155a23cb2743aa5a3d016f80a1ba80bdf2c51b3161824392348a579336782dd5d36dffe252b513f998595aa32775acd3a22ad066122ae54d0eff24b1c8b7576d5953ac732d80b935e57532b8e0655b74dc61952848d1d47538ec3529c78ec2d37f04c90b9f4201b087e9fdd0e5848902e576b25bd5de2c316f7e9045735139bea33be4cbde3cd907d1e7fceb6a130763d6e08384d47a7c73174b568fe53fc3fea9f75cbbc9eb2ba0d998643fb935f3caa9df09e697c5899350dd3f53086c4c74e726ca7c293457003152d9a9b97a53556a631f33ddca428d120e59dc5c296bbc4e6f384f727a846b740af337b0f45368288939fd0e44fdbfeb50a9bfe42066957770ade4d813624e4fb20a9892064ae28cb37e75ad7c230caf0ec80f264d5f050984d77790c3f1ceeb7e1e2794c12e62e986cfae99d2c2b5707129fadf1dabe4f90322fcd87fd4eaec94b2c7462a2f8f285b99d0e707238fe301db7c20ad5ca0caf746545f22ccd0efd68097b660d3be01bdde07577a51868c25ac1780d2ff51920cd05194a80cb27d78b7b2376fc631799f026aa75254a7b40c61742f83f5add680c347f3c2a660334991561058758b4f97c1dabc0e11b7fbcd58808f16c8fbaedbcce95375b022a4f92fced2e605a48b6c6a2828d5a86e5fd2580d6ad6b350b5b1d1c9feb6907809e3a66d9c2ce982a467699a87e5f721e2e68d4f9a3003510e9c543182bd5b8ac8ddedafc7304fd0c3eff6935caf013a24d2273241ecaaa21991baeb6de14958a767d0417c4acbab2ac7f50ba9190bd3f5075323c805ac55cd31ac83624a42c764e6bbf056a72ad6b28039e8aa017942d8456c33725be0e7c5b0e6fa7099089c9bf6e1ce8396a29b0c6a87ef4575a42f77bad9e2f4441d541ef27390754c1d8ddb3808f91dd02999ddbb98efb33a98b96f6a34b39bdc07e82a71f5cb9b35738bc0df0803c0148eedf794431a5d9d8e2adf3d95f53dbe9530bfa2307ddd4ee587648f8fe2bb0cb81664af4d354b926a281554e591a05b0902e083b7c48c59fa3b3ac5c1738583ad76fdbb60e1c1d27c0724ead89cfd242e268a67e59a0dfe8b03b472a9217ee8334b1b6908161ae45e1ead8b9998dacf8d8571cf248762d70bc10bcb5f415883d417ba3b4c107fa793fab73e8cee4ee2b8dbb52d8952137c198c164c62cd73553f6560990f0045f644870e9997e332b10f4b657824978e254ff072b35cdb1cf3d2c76647854b0cda45f2d3a0301a95db7947aab585c23e6c52751f6f46a8c7e52542c87c5a794512dff102588a23e187bc931b217a23f2b758cd3c6ac20788a67be48efff1fa5c8661da4d95526e19b971425800bd5138327c314dcfc2f0f1e04c0bcf1ad09eea2e403b56de666bb0c8eb9827ea3e31b8423586cebf0a1e395507d7081e4c31280a4432ffd636e937eb5dc608c59afdabcfe082b21773b1812cb5fb0a7a6dc8eaa17e992f63e73dd0fbbb8ed929747c23e3350b9d3a4685fd1b52b8c2a14628536fa25fdff5d36654e8ef1506e0049a87e69db6c4555458d692ef75e3c29bcc4a53968b8c1008223f9e2f13f74c883bb5b483135d4170250b272c1db76368302b8075342f04d8c4d0efc9a0ba08ac26804ca557da570c67bd2a855a66d0a73973f4f78deda73fe3580e65d5641471caf4d59a1a86004d5122ec1010faef216588c02412f59f29788dd64a092e93056fc78c331cac230fb4b0613cecbbd9f174469c4e5e6a6c2e725a0d10bd0678b7243b33e4313d2c6fd16d3ec94b0743b200115aaa7770d8a8526f2d0db5c0841ca57db51a9b87b097b58fb9be84db4fbf6fbbc9a6a0e58560befb1a2e55e26240c07406f9381ad9074edd9d5143d4ca3327ee76eb405976d81fb7560cb054c58bdb308f0f4e889fdbe3b88cbe49e8b31cb9f1b93cf5aa230c5d3b8dc07d7b3b3f8ae63a11bb06c658d01e5e3fb1dc1917dbe3653f51a2a75588356800d769bf84edd7f278758fb316611426ae4e4327277baaf0d4f8b38bd4a5090bfb8ce55f8920ed58c9483d97872b43687d6d7f06cb47f00f3bafb200814da863481bb997b5ea05362a5cf8260de61741d2bbd9aa5f607670c8e89b9dd1d7e0951cfbf37d9ec2a288fa2add1d8bd86afd9084eca6c62f3b99a314f515ab69384b6cc76abc565995f681f0380f41b997ed3cf0755eca9ebe74a14ae341a06393c7563fa2928a86ee7d2665d5fb9f5f6143b49413cd47c40feb3c820f2cde7d441ba01e9d8cba2af616fdfded0561648aed27fbc7f1bee3a5a1cb856002cdcf543ccc16dcac7272c5c00d08fb84abb7f9549d241c00320c69f129ece320ca9864a4e2ac47e98e0aa80452a5fca82ef03343a67ea0e9b32c41f883faf374de4e93eb4b68c195f228511940c41361bc3cacd1fb5c5b0d463d58e03698b0b7d18d247dba44aa87d1c0734068a20130714d1af688bd732d9fcc499f86a8b3c194d820655051280d815d03f646e5670bbdc0d880c1170f6d20a971a7d751d3d3c82698179451c91d66e03307530007757eaa04208726ff7edb5fa460efbc9ba6f311c34bd84a55eeab3f9477cf7c594ef246ef50c66fa094ff39641dd4bcbf2e736190dfd1159c3b294cb387ec40b706829b2e6b1a297924dcba9c0a4873b7f8be68c835a2571d198005858d35ede716b60613b902b777d802327562da06e01748c93e3544725d9637ba5811e12887f98071a80ccc2fb0a6b10fc2a5aca65604558c4a92bf5e0b057834ef04737149f869e7203fb13cc0e284902e670d4e6bd3e3e70cbc2a11a489761ea1bea9c2f290dd20c79806c861f32bdab4ccbffd77e400499bd32dfc2816ed3eb98b6df2049c56c63f469e563d6203f361b7b1fdb2b365418ff9afa0112e35bf2aeee59a1556af7e0134ee07e15c4fb63237768c87951f48d191f5f66b484581b1f71b84a3e2e5239ce26ef02cf97eea07ec6c9b83d26345600f2ad3cdc437673c77605876f30cafcc82134401bae71ab4829c587abc3f7af8e95eb9abf95c72d080871f7e112468d36a56b035ac968c37d81488d0506960a1c118bb4059d4eb7f4fe1f4f4f7ddaaaefd03b15e2643b3199850d0dd0e775849ad5b0258894ebc88f8c9ca5070d572c274329e4ba975da0e163103f4d16bdceb7e2b8658fe63de12be339b7acf64d23b41cf17ad9c23ad47b6cb804c7f5fb582ad2d9cc886db41252add5dfb567692d1a505401954650321b8abef4da526a66614553811d8fcf1d94badc548734307d74da7f2afb84ba4441e242d397a9b9b5128ca2962baebfe8ac6f016924d266c718a874a535b81641f45eed09805eae00d70ccacc741c167931b4adf1d0adbbdc187fc9c8658cf9c86c5ff8226eb0bbc67d1b63e9af63f544763ab60323e2f5aa16d7a70ab9b74c32aaf49054ce6e1d2e0c4a86e1fb4487686c790ba1f9ac18b494956aea2f63dbb49f66b5d3bb5c6018c95e802e37a30ced8bbf1124c6c490a9429cdf56dc0e2c56e3bb2cc6442eee4f092080ca5ab003b70aa8ef9c642a9ec68b11c9a6ab036f34c9fbcdb1eafbe4a546ddbf7076b10ed2785d63fa4e0d89465cfad4d6f075d069cd58bba3fcce82ff1a3b4067b9b8a75da6d294ea67634b74363443580308dc08f1d2b5002e0adaca1af1ae4477c2ff5717a6a193b40099678b812e452526e1ca8119bae0c97cb89a058a1c8c1f43eadb1526e6b5bd078946a3d32c4db92ac030e458968039258c04f545a08cd16c181024abcc8d982f596ac4e40ec3b1a415c62b680ef693b27a25d170913352cba3def7977c5912731beaa2f8b3ae5d2424cca2f23743c6bfd7c1282e0793185b19e7d5f132308a985c59dea2025c3bf9dffc0194dcfc3fa04e742740d4582894024913f9d7a469667389027db5529d5a6d6dde0d3f4f6ffae500d6ebf5ee93d52f54886749c91006de521c7bea0486ae42fbe9c007ae89163d2aa993d56e511a693847a42c53562d4f11b7d972ce0909c98a605406f05ac0113c76e660c4ccff5ddc70759d58ef488814ae524175da0f12b21faedf82ffc1f9080fccb0bab754f6ee6c5732f1b97e79a2eb9b8b409d24e590ab06c14f497f6c510e828d404a61806ffce43a6943e0d2904028c158527bed6ce149a251befb6b0198ec67b15c367a7e436fa3b2e0a015d7e69041408727f4db6706bc41f8aa678e3930297e0d42b19f69b42cf8228a4bddcb42f336ade6c7a2bd0ce982b3cd7819b9eaffc37e6a6f1218d202774477db41d8da82a0f77f459628f7c20f143ebdc82c1a8890d3db273cbd0e3ce83034951abef05edd77d6aa99ed451715336fa5bc22fddec763527c4598e1c3d5c7651b69cc773cde79005cc2ea8e3c48ee322ee822da01ae8558ff547fa6fe70501434ca5698fd68a72dc9eb8174f0c0fcf80685f41e78ed4f6fd7a16cf6058abffb675940b356b32f0eb37a9fd66be1e8b79845fde92713e43a41d0e49c04fac23823c27ca9e79063e29bae9b9767ad2ffc30119e69e46432d83b89f92e00d3faceea162f0ba21326463e3377df88e84d1f11424b1c3e607a9d5652d38006a3993296a8881430496039110ce8d1ea7203f59ba96de5cf386e0c108a553dd1a7001c6e9153c67e324a44da7a75708f6e75dd263e6783aae3af335f8ddd66166dd4f1fd67a276e09fb6954862fd2743cb18d623799702f5782135936294af1c0a5f89f986041405c4fc8dfbbb54e8705fa24d5be2e49f77d650e02f0f3b9da844cb74a18684580b5a2ae01d733b3e28e27e1a5f11d210057a8c2e6c5ca3bcd4edd5f12505a533de17c0a6b66777342d1d988503878146a4bb3e11ad66fa1bd1469886a69c08ba33a5850f0cb57ddd2aa6550;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8e6bf2cea079be26dff39e450b8c1915313d035af69e59788bf94b2fd07fc230bbe65250593fb53b333103586d9bc36d2226f132e48b0daf6b86eb898e0c435fb4955d8a6ebdff9729ffc6a1e0003a27c7e14579975985d691facbef6d7a21ba677d580420294c24075548b91fca38c098e62a95c75dfeee59cc8be6f37f987d63bd7875fa833a7eb91e78a98680f3984e6dee099866d11b219eb160d6fa58e74a26b9f332f0e41edb2f4da059927be4bfbd0a4b988354f3b537b7b150c852fed365dd3dfbb62e9ec14ec9f0aa33d01fc69e3f9caa40de9f8e2c729bfea934f0f30b93f69426b6467e4de00bd2dde0f7e2540c1a455bd26d5a6d6152e54f7434cd803eae4cd96b3bd810aaec76ca04deefed5b33f439a05f5108e3a822bd414fc85a6b1667180a87b961392d65b3a3831475e0c2194a49628f642d76d8bb95f4f031900d3ba126f7bf3db51f6ca1fa72bd128842123dc98176dbef210368174c8fb6994a3af16582f32f933b5afd88070b9ea3db788142ea1f81cbab2dd7e17ec981ad5fbd773e99152a08d9caf77c926f254814dfe0d07a686d80a56044c4ead1788086527be417350eee865df3a91253edf6d2739a21dae26578d334ea0b51a97d7e0b609087b77be4d8e4235c869ac5abef7cea9df692e27340bda96f3ecfb36074ce2b00395947bede12e40cf1351d0e7fb1c6a98acecc6f7d8de606be7b09a1a7c8d5498e7caabae4076e6d0a84f845d0c58a9a6a7f1b2685a9af0f951bd23f7e6084879b5b78f2c8e7d419ed553c2044cbe5c87caf6a2f6d8cdd90a6f10206f835713c50c500d23026f4e8ec4bb223a708575d4db234fefadfc74e724b6558f3ab186ba2df2aaba78500585a833deb47c552a76efe2b32dc852405744372c3ec88a1899aed9aa80f32b80767a5b643ebe4174203c7017c8e30f700460e92c095130eb3e68f90301795188c2f65b83cd8e34ce0c65a9c5b92d7686802e57080a9958e9d4388d1eb6f321065601c7a015ae46447db059eb476b517bdc06f044441d10d46019cd2cfaf4bfb8a6b0510da828edbe734daa2048c402e7f142f129f73754bbad3cdd320c0da21fa8079a9ac1898d83aabc1fe07602ae5df71f1a0696841d8b20700d8fbd8a8a5283ac0c94188d588a709717ed34f3d553fec291650da2649759e7361db518ec47bc4b0883d47967e7405a7526695611f033f085ebc5d3ca5c46743c9f7af1df9a1e16c8c764abc9c5c025e9e39bee9372e861cfee2ff430021b92042041fd9cf3e62ec0325bce6f6641d580d8489308938e097efa08bfa5f73ebe28e730c91f671666dcbede8d9019576a1705aeef778cc006a367ccae1298d23cf4cd7e8aa1a7960378196c1092d2cb52aeb4266f445a2dee81964f2d2ce5bed6723c87e24ea3601f24b85c4924fd8ed4e7a30bfb7a29b85d5d108d7e5961fddc636278338f878df36b39fd292ede0b9eade091d21747e3b971e38412b79ccc0f3de13b5947d8dd14a17856b7c5545b2f135cc2a1858d7a6bfe9502bca424d6e9a81d5691fe72765786ba92a223f1ff9b33aa3252c498c02aaa0c2ea6664bf371cd2b182c970a7b5ec875a54ff80f9e8c44506c2eed43e607d1314a936ee2fbd5e19bf8490041ee4565c8feb222b7e2a21a5666238b57034f50b20149653fe9a6ba7775ddb28b2c1eda19a56cf9712ff1a2cdcf9af8532b3e85450f54cf99c83053d411da930030e62c7c5ae8e255e5e2a6f2fe51fbe503a2f7c619d7897f5ada8c9d3175987efea032408bdc128ebbcc7f8e8cbe4c725950e989d235ef71da15a745b6372c01c91c932b590057b5d0f43f9c38275b96697de6938babb2068289311ac10011914579f617614938705b20864e868235f252ac00a7b9c2de8dad617112a8d4637485c048ba485fa7b065e548b593b6489d231855eb5d667cb050cec5e3485a4b5beca4ad9e5d987a7fb7e73ce4e865e2dae317f75d19cc74ab05103082dd5b08c5bffcad5bac7e9c844d0dd461c93b0ccda7fd952d51eb14dec8780471aec9913efdcc6d02ab16e059ab8c748938b422b2fea09224641d318558c17fca13ffd5b3b2392e2172a5a6fd12dcd543d4bafcd3734baef127044b29d8f1d7c24fc93819c291ca8e36529f5cc478b46bed5aaa7260e592874fa15816288dfcb89e4855ed6e4170ba2bd60e83f597be8e6b9baf4bc04f6d9c6623354e568385b4cd80481c092a4eef7da6313910e27e8b486b5cf099a9842ae13c55e6d716c5b183dff9903f66050946e1a99e6322f4bc61b9055cdcb1e71bcf27b99125cde069d61c45bdd785d7ef8d6148ccc7b2c7f86c3821f6e83cf091b8e840714b1697a9c5f24219e78b2be80d5d602d857f0afbc639994961c5943d0ec1c8eac1ac1a92d43c39bf61be994b027d10c927abf2bedf4e2bcb42210ba0baee07089a18b4ba31c04bfff205ac6715bacd30c6aa79139f4057211c28f73ddc33a3975297eca612ff0e0deb11316784f3373acc76f748e637a1ed378f86e02db94cb986e723d6bcb1560293a0c0b53e845394e3034fef991834ac9b003491a7388cb50d567cbea42b9028631191fd976ea401d434d0c409df1aa7e8e670d68676972943259b2fa9299a4208f9511d92ed922d220685cb8a4e85605edcf757ce8ad33d68b08bff40e365bd6a0706d266aa605c52ca2d170939c20851016f338540b4c77c51d1f69203738e1d89026deebf889797f4100f8960bf16b8745c298bb3f0010842f3b52a4f6e29eebeddcf263ca3d8c70930680a7998b1dc1c22ace693c677c45f1028240dc6cd71d41cccb7a7779d2ee305d8c6dd088103a44a85b7ca21e54101e96d8d66ac449ddb16b5a20d520eb47412c047e0635a0af9f28250ddda93754b14946dd57170f6a948a905d176bb190e5886ed46e0083cb33d7fe78aadf8f91ff6f876e302d29e26f4e8f79e49ef175e9aeb21d2059862d3ed258272028818a8f081a806a1c0705bf4c7406ca5077c0fb8ef8aafbca86185a32ef0e24c8c39126d0b722c8b17371618c2f595574d2df8851ed24a54ebae876587b30be009fe25455fd82e99257367e57c5f2d4a1451fa02033a4e0a8564bb6c3f9c8cecadcce53852ca849899702bafe1aee723641adcf54beb941523abc7fc6ad9e8c00e3cfc8fc8173b6c271e61001e0f97cff93e98ec8ba297c1e9f9ae245ef1231586dc25e56dea5eca28e99b5665e623f1cadac83c664281090b6f113d9dd2fd9e106da8321e4acf822a821b99ee12c61af2a724e65239998fb787fe659474598ea9fd70c3b82caeada4a0e8cbbdf3c4905b48bbc37236801f84f75ae610bce23b931767e3422d3ebae28541427110d964702558005730682fe322e47ee63d474aca407ba54c0b27ef6f0d7082dc9da85c6fd031c0b8a6a502b0e1cd8e5ef6f38a350407d8d68ca797cdb53de9352c74993d8f10a4ee0bc691ee947597ab21fd6e4ee570c5b7d2a633749a7d280989e7fa124b73c2fd4ec25cedea3cb0d1ac4e97a9417c71524661419f436f68c52a09d9a7805530d1b93831c5611a51a71c5a27d78bdfe550bc985d6a3186cbb4dba357bf00c67d365c1de6079550155b52cd61958d828cbe56e6d5b27e14a80b0823a067203dd98c5efc7e7a66ca1a332b6e46498c59d979af3e752050c3fee90f819d4254d334da5b7ddd12ee6bd0bc7dca715f5d585a75aa0f3c8defd1033a82fb7bbf581e0747b0a0d07177b708c2194762b4ff845db22c81ef78f3d3ea0ad44236e11a3ef42cbceed90319fa60c671afdda347aa27ab32f82c932fda8effc8ecc2bd057330d2ca1a7892b3dbb2328c594c80e3ec7877c4501e4288371ed514dd77a4e87b81db900df1ad3cc8aacb52b3577fb77d2d9d41b6f6e6d6b4a1a5af89b1c828f5d7eb2866051417053436c230bda3d86d9da4c55fcfec3495596fa707ddf0d195932a0aefd4d24cf1d4cad1deb390fbc19fe168a18b67971655fe2e3a5b16e1b5e0fd85d80421c29b800dca5de4fe3cbf16e48afdf914b3736f30ddf372e6a7836ecc3f86f00296f7ab3cd5e2b06cfd92f5347da040ab98c1a8c913d58401eb4fbe5a6da58bf488444360a559efd7ad7469c06297da762d48b797d52415fd5a42386a0bf75707c959a2e08fa82c38db5f3eec16f4eb635d5c2e7ca598d56a491b1e72f0db1de4bfaf435aa35b7f9cb7e9261d9fb12a2524fd95942307fec91fbc48d6121489f88ad9b067abb4d8d189a0de1ef362b2d76973837a5b240b60e19b576a8992558548223b1872bcf77eab90e73234cb165afcee80696039bb851551e5b6374d9fb734d8d7b82734a348caaf4e29815963dafe4854fe93623bc6bbebd77103c52ac0c0d1c2dd66fce8a09dead57d9b857572060963929c1f4896d76d49da9d0a1b464b02d90d0bdbb8c225e5145b645b1b417fb5f617f0ee6110d889f8686b101ef75ada16640696a399b45c11b6bf7669c7c2a73a232ef06913fb0233f65c946d8458f282bb54ddeb0a7cb87b23296c5af4596c3ae75108ee6998fb181106b91b1ff79b82eff7ef03cd5eb7a62098b0bdbd3f83e252d7589925f86df55e7790c0cd48e3b3463c9a101c11659fa4d4f7157ea09e476267c466015f71598ca6e2eafd41a6b8ae4141bf31b9bdc9d7def799424916a6ec014d710769d4ec2b436aa253a59f21123d2f51a11d22e2897437d853bc46a332297b454dd03814a579a47f517892bca1543299f15299fd514cd6d3ad24aefa2e258118395d882dd823050968cfa4a8ecfde532dddb11af102bbeec235f4a213620dc6ce3969d8d6cbca8697e4ef3f2cf4506aef8d637ef577a7fc954c02e785df140b5515347fbbb477020bfdc1ab1f9de17328d96fb0ff497e0c31341c099795c25121a5e6db3df07bf906cdec3d462636279d2d73526da07a05d2a28b3381ee969290831245b44cc1bda128c9547fcc216ea954449b010f146aa0f2c8e899d9dcf273acaa6955b4c52a66703ad041c8150c1c0b1c43772add6bdf8ed741b79d0eb95bc021fb62d90b5ad7f393ba097424c5406148c5f77073d820f9b2bc4ae993bbbbb3bee150094328ccb21f472ade12d7f37cb7f06f116040b4ff5802f814e9cb9c95ae02ace16f5149273701dbfac521255eea3aa8074fdb07c91e44760d8e47127b27e53c71ccff90f921c8320596a69e0ddb3652e927201f2e7ea68499dbf6fcaf0b566a0cf392d4dd12fbe7863a193fb718523b82d8bdcbf3d9f4f73474091e8e7e2759904ad8645a1dbfc6ec3d3ff3e7e2dbb137f88032be0918391a94ef47817428d55082776ec2a6943ddc40868aaca000e8ff6168e98a28e633397f0763499b8248247203edf6723acebe4b46b2d8964ec5d6190ea133dbb3547a86c2dd584097f241a73cdf6d7f3702f08b77eb34e680911352de9e5401b8ddab88468708aabef1d0b233091a3bfef9d5d76cb2253d989b8d73bb6dc6ae70;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4388c08a5f115fa8b230770cce65e3db65ec4cd22caeb50cb7524a1265c499e5d514e15103fbdd470035f4356214c999dccebaf695da9b3f4a4a47a9d1714148964cb7da1208f3f462819d729b04ed60fc356fd97b2e3efc6e0f67796d779fec5434752b95fd7775ac04c612b53b5482be4df4f4db3a2e305db335210965d3a3ac1cf5e4c47716f1099add0982e42e2efe05b4a42c7a67ed70ff49a5dfc616215b5aaa0a31a3008f6d6aafe6d17c667fc6da39d1eb01b539c1269835467f843be307474027c359a9be711c58541a3e4a301ac99d37753b02fb3af53c95517f1e049fe94412125521121c20ff74dd36a1d39158d0dd786a85e6667c5bb9eceba0f2ad69acedfed9fbdd41bf307401af9f41a29bc0068dba381e02ce35bce7c51d5c2ad80417070f2e4857252a0f3d81f2df5299f5ff0d7386fab03c48844af7aa474eba38fe3d659d5e2ce553980d26d709bc44e4fb26f878c960f3357299b26f23ac6cb6f68ebdac2ad530b37df26b31c94c7dcad818df442ee40574681f918cdddcab7bcdd9491800c9a07d131ea7b7e8a2842bd9f81010243f5609c321406a231d195f1e1fee394ce5142bb5bb16b737dc9e64e5704806cb9ad698e04f7fd9ef653b0fd72861b5456cb2fbfd728df3f24f0eeb94b656dc5bb4cb69a96f623ac01bc7afc6824a9d917a6cfbd9e09dd10e626563ea93634a03f47e0542d41b6a960001cbd7c6aa89e79e6f4890d383fbf877716d011439e3941e4a0e2a3193b82de022467346e64cd047eb360114f880aa37cef9348b3ecc07248eb4cf9e999de8531bcf92e4dfbecbdf883f54c23f4f6f298387211693c45e290f2ba3e5cb36a82d536449d1aa7f24d4fa50b60c8a6b78e4fd1628c86909ffcd815b77a95f6cd083ecfb053c5139994927e6ee0b9e957f5bab01720b6b5ecb95af27e6b445720a2424ef803d4d62a1872fb63f40395688164b8775b843911700d9e86c643d9c46249db40a7ce0e0f5b786390fdca38fc25535eafb9c69e4730117bd06673f5c017be8f9d978574bded6fd14c2c46f34fd5168f0c4aa851c24b09388aedcd43106118dbcf215cac16412fa0d538acb6fb95866a8807e11231fe62b452474582c824eee834f6f939895f56eadcf1fc15dc2d4cf3969f4ea3f8d8169b8b4e1cee54f2eb7d44e76359ad5be2f8e2b81e21b2f02977fcc2e6248416da8e2dfe6839a6d2c581d671a9d26e288dd7664c7f87bdb007aa534e77d57c3f8909cc8c0ab151d3eb1dacf7a9507f42f74ee55b172f2f4d638f235ecffd9acbea3b1b5fb89b3150fa974528b7924bd0e9212eb18595971c3b7877e2e8f84ad1d6f83c7a631258ab83ec9907f94a058ac2638c46a2e656f3ef108a8c55e39795af3a89eb62267a7537a83cf11c0a2d037667601e6ee36c565735d663ab0b3d4c8e82857476acf38b0f853f5ba9945895f60781e485882d26cafc058694ed5f4c8c62d5de3f3a9af80bd29d563b6fbf5e725d4867ce4f2f296d80ae58d357ba0f16b4bcec8368f995c37ba39d43e4436be1a23534c112f5c739b8f8e70f6a3820f920ad4d17610d6cb8ed78177b36729cd5f122e75689d8191d3228d230a913b6702b2762c94f75a828c87c42800311385dc72809b6ff436dced16a07f75b69d8806afeaa86f0eec410c4af0af5979f1e04230a6ca7a8349c980a713b56a395bc613dae389fe59b9a212c4696e84ff500965ff02392b1816c9fa608e49b6b530d1caf8dd7f7d44c7b3066b98789203f0defea0c74061b15e4419c89c01c15fdbc0c2a11fc75621bb177fbccd6c00628a95225ad6725ce94544fce5d868dd7742bd185f1db38bdc32ce6f390c8585c95f65e7a816618aea18f7577afad27808043afec28d72c1e08f9176a575fb34709eb5f672328ce6dedf63045524ec7c5ebee81789de84a0ca86f7c9c5c6fa0d790e83abd7a75edeb89a850829b8023501984e0b67304435821c5dea43977d0da70a51ea5aa029bfdec26206a6376c7dab577519a90ddf1d4c70cedfc3ea49f50174ac422acb905d7ae05320e1e859b558e1530dc1fc4d6ab878849c51ae4f75dc4a6de1d1032886de698317e6d735202bd004cc2a7fc8f654d0ee18f555f95c34e1358543f4da8f720f7c3e7527f898460bd8670533635fba7816c98b9debe9e88eaace3476190af2135a2b581f560744b44799b74c08f679a5c3a146c0d0cd944a72634228555d7bb1be226fce41912143bd38103e85e43b072ab792a6fd52cd46736ec1f5d63faab7164648dac79449b6ca7a9d9b995bea4a01ac04a1326979343cebda9035a0dfeaca2c33a80b2a5a51ab392b75bec25fc3b995346683a9c5c154549b5046aa7e5a8956dec9bda7119e2e8a44a2921f2010ff20a5dd7cfaa338ed1210b7de3044c31d2da5b9707784ddc96ef36ba6c8b7248fbcb035e767a1af6e4fb90744f8e459249efa66618cd14d3843dc06586bb576c895eda7af504464ec9ead92f59689e02f8086cd5223dec25e24bf6c5ef36c4a56d0b89ab7bf549c8ec18fc70a9754b1a9ec3a80361765be5a7bb8b1ee374db9f2ef5d7748cf0fdd0d1d772e17ff43f9ae5cbf7b86e34d21c18081d4d89fd29f7db61b07b899d1bea749b60c2e8889e82ff86c3b66c87514f5f4e1a54d68f36507bd03c844069095773eb6b564903baf7485246a7218bae637e2ea697e1af9a72579a7226a35380019eed6139063bcbd93662d788abb6301b56b32d5e45aa6a1f4778aab345a413266440a901be00917a419905d138ce8f423bb05b7cbfc377ca2808e00607f2828b0f63000ce71bd3604d9a5e63674b3e4d3785650fc1bff5ff382e6ac94b30a9995659b9a5270c72fc37b0a4ad077aa1760ab14e2f46d022a03a36a8ff7d0bcdac37f5637709a28e52d32ebd29e81b9fda09eea08f3191fbb78a582222d4b149279fd33cc348357247849daf0383dbc4e031225e9731ab4f6f1a98e97ec109451d074723351636f9fa26624955ede0e1f153de531a960b6af6d77d0dde2de640b74fde5a695021436574baa06d2b8b52e3406637a7737ac466f84560dd21660cd239d347dd24a8bb9b84277b8eb37e19f7b4c1bf5101076a1868679802ac4ed1266617d46c2207672f1d52eb80f59086b576f0e93d1f9010b2e04a7adb8cefe9ad2727dd334ae523acebbcdb536cd6141b3aff21adee8dcfa3ab48f5dfb9e7a3b486677db143f106cc4510742b7573898c6141c7f910005545ef307cf5176430fc328361b227300aac472b236d007b0db9b869d76a0cb3e91ba86c9973c1faf42e58238de6916a04c66104fb0fe966a207cfc87e128000b55ed4a12776099da91278ffe0f23871ea6898a778d32bf4f2833895158e0283618a4e2f4e559e0197e855d90fc57ee6da7d233a7906a630b4ec5ff60019d3647d39f5f8e0cfd2748ef480a1610e714094d97b8eb6d45b9cfef45c2ed2f6619146a328db84a2d7a5970a570cafb9673a6c5b39a0c56024ac5e4e8c3fdf4b2c352fd048f96a69b59e2b21d26ad9d5fa51e40a5479be6e26d382f9752fd431417c0f74a9b4e1e771f6145ec8159f0becc2e3ffb61a271e83461557c1cd00d5b2b3ac8f8385c4b1048e221469f6e77abce44a76dcc082082ec8a816c24dc6fda8db630c945bc1b91c7ab8391bbc9325adef641f1cc7efa1550c898e5501243cc03069a660f6568e3b5f938216d99a50f65b830cbc2c71d06712003be8b94020ba1f385a0da6a68bfcb67377f9fe3bdc90cd5755852ec8f8eb9eb60df34e6b78d438ba8cc3a35c0e9864d1d5c16cecbba67830290c2c387213bca90b291fbba57db532f424e0515fa3f3c3fdc398cc4e4d0bacd5a273c78d3ed54c1ca4263fe5b38ae7c23d951c4f5d3afeb414e7460aacfa077ba26fef51a649baf476b092a0b89fcac6442ff081ada5109e11e5497d86e4392a2acfb1f1e1cd54b84fe78e733c0b71f3aefdca6609d66fdb1abddcc75d92e6709c92f90a3dddba4f4ab00dfa06711fc9371091fc60550eede409c7aceeba09e568ff0bb93c61f61557ebde1e52b0ac7d6a7d33fa7d8be4c37c40d5a9040c212386f46043b58d29ffc164a1bf3d128b13d24bd0060294420d7119e225522d83f8fbfc6d197de0427c6d7491f6df90c50174a73db22b9516b7997e69b61fffeb15f12c477c87f676a0cabbc027fa0818f7ddaa6a2174c5f0fd557cece44e54132b7df5872f1522efcab6808f44a223f086b1217084e142c0ce36f4e329e6531d6d79398b2c1f784f85860ee24e424790317ac1504172b45c13c99fc150b3dfcced6a99a408580459cb6a54d765d19884bcc9d633e08184c95ddd15e338be7a6b04b898c8c9988e313939b75d9d66830227841cf8203dfa8b4c05194eaa393321d595fbdf9c587975f8832c1e0bf8cf05ef410cce9ae99a0a0083a603ffa0427704c6ad432f8aefb3b4895d07f699658a80d664b500c5f5d8862e7eae66b252be887c8eec7c125c5272262f908a3fd6d1f70852b00fc9be6ad3c7573e0cd58c66199c8e9832afcdb5ba7b648e23811e53f5070fc6427f5fb53ee31f2508f950b573ade16a1615f48631d66d6584ca13ced116f342fa814040cddc6a00a59e5f0d9f3dc23a755abd49f8fc445d2b3b06bce61a85b44463d80e653f4a29f25cdff3395b5d5febc7f2e392259258d29d00d62d1f5dc8e10f7461a38fccea29d5d9fe766f073e620ca3664436ce94566f20f5dc286aa6468ca347d159781439742d9a5c18ef60ac709153a24f81a6b0ddad6f4b99aae753d8ac72601bdf396b4694fad292c5fec6e4c1cd36550aae0479b61de0c7b278f9cdb1d3b9db23ba0b4b98ae8387219edc1f9865013e9b139a94021222b56a8d62fe37423c9f6b4dae2e065822ca90c13a34d97e0e1c669e5cb54185a10b6ba09b11844fc2d1e48923403c958cd3795277970aef114b6ca0d93822a1682def64f66d49763f7d870757574d4fe2209f81e2b032d5f2d0dce05d305ebdfd5d2c09d39a04ce959bf041ed00760ee51a669b533f5d192a614797a615e4d7d5546fe7c121860a193584b557aa36ae82178511114f388d5218def1f55efb9b1592b573223f4651bd4367ee9d46d158f8390867c0bcbd73d66777ed4227dae785313b00539b0c67d039361ac8a3db4a13c97b67b78887a9e9cd5276dff157fe5c8e05ed6ca30468292158cb9d9f38d11fb13b2aac369aa4f0b67b86f934d58fdd1e925ebbf8f26e51aa82aff7870d1c0558acc9fb5cbdf7c56b540f9ed57046a3ddccb9d9d2158cb85e1ece9f97f3c69090cf46e627b017d162b8f696bf245535be9855cac05e2f9a5e89b27ab0ae635bf1596e5d972d9366ceca1fe04d319df45b036cddf47024276af5d5ffcdf092ff85adfedbf3445f702c3b8f1e61a57872f692bc7534221521fbfd3512d4d878d89bdaa943297f098e313a49a7bcc45c02fcf7bf3a8623d7c90b4b33e848473;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc612728dd975fecb10067481d8cea420d6a93574ac31041331aa08ef9b187da33fc5a79f59ec20407816eac12b924d06e67f3d5e933f86bafa4534a49e23a51664476333d22c9f70c82e915a38594adc17ce9e5a4ee90d5cf599c8845194a5c18bdb4bf1979e6f18d89e3c1a1f5d06f4c05b372b213f165cbf4731810cd1c822fe02e1912af45a7245f656e6807b461bcc942fc455b82b0136833d08949966fdbb6168afc5c18e0c83ddb27a398e1077e9cb7d94689c8d5ca5bbc790c078236b67a3239af1de9b5a67217b7d6edb16038e993a842e692cc735e62fd9658c232247fed1fc2bbbce4242bb925feb314feb0662097bc54012db54e5684be397bcc35ad6c034ce2f490ba8ef059213f03b2717dbcdc14428aff87c480d4f85a2675c304ebc6746fed5efad997abbd746c5206e40d9dc6bfabe2cfd7538740612d0abb12a1b3a08243a14ec569d07826bb941bede81a4dcb1171396e79ee43caa9c882c00129e0fcdb660cffd7fe9c2adf00448daea14ccdb9ea3bc310cb5021b7713efb4d2189efbadf241b91d03297ee71c5bdd6594e0897a85a3a73497d422eb13dc48f6ccbc93084cbb013b86961f3488e415120544a06430cbe69637195344953c0911d7010575983d17b7eeb25bf82dd23c50acd41b345503704e9436654cabbcf9f839e36b3ccad51a94da949cade3d2b36923e6861f6f48726bc0310b2963efeed2c4868e619e14159685cec096c0ab8f02c259f4591bc7d1a93cb09a78d24239f5d8e377412adf786737e3c9af38288932331cfbcf832b19ed9dda4fb6fcad9d9158ae1c6619226c7bb82d146d5fef44148b8b9ac9fa3015d4a4d9d204585630f08de5be2fcd4295bfd1a8c0b3240a34a2105a741591325f0602d3acc68a38cccb40d71f115a65c62456bec1cca7ec7ceb61e95daccb3e029308a9b21a696723317ddc0e077d19019a4e4c02f3737114c29e322908a5b06d1701f1c9080341e893113360afa1f15ba9de033a93d59e2096c1dfcc72f453d054ddd78a498a1990315fe0a9d12e38e42557a658d703cc687b998535d1908e003ad350bcfdabdb7d8ee6d2e8f2b012a5ef059482c0d1137de7e5687aaeea3ac56e5d0f1a5bc13c61cd83ee39a2dec895defb77e9cf1854b47f82ac81417289e1b2572ff9a3c960cea45e7b85f71f60cee1a985be27d29465220fa0cee1892a39083a255692ff040f06c8450c4af155254217e6036383dc206381994bb5896b67049cc79adc443612ffa1947f35533772cabd8d1277a4f4843844328733ebbda8998c2ba28df22a44030a2bc3b7b56ec4655169eb30a22b65eb8fedba9140eafa48f852fb2d8be0b31bcf1f50f105fa15a13ff55bb6cbc4df4ab5c67149e6a3e01a0fc46727d9e980eb652ca1d0395c6f4db4d3a0746fa1f4b72482eadeb58624c28f3c11d7dcd451c70c904a1ded29c1c35035a2fcbce849ea9ed6eca8fab8a9cf637bed51c6dc1f60ebb6908537768e1d65d34b0a00c62e0e516f07b26b46687ae2af1c9aea6249b5b5bc2761e87e85f89bb7e28535ddfa2adf0af3f8b39f84f18111468310a6cf6a96e73b8126a5f5066cc35458a561a0914556c3cabc11c6b2781063d16465eb6b6c2e3cfdc5fb4561afa31fde440617afe6615e348db78c4acb92aa8705a8aa12ee2f9c5bb9622a3a5ad7be315926042f9fea2fd2acd218ca9cbc7160e6bd2380276d5bed99500ef4cd6bf5c08df07427d585f0e2b5dcd17947bb19ee76ca94106059b6694c91388af95b736cab9a2b988a7853304eec91df2026df86a7baf1f8f2d8a712497319f4c6a29c51910c4c79a8321a5fdcc62959affea762cf41f128c78a4547466932dd94db868df2fef6181cd1b22e323fd5ba084d3bc745d992c4d1461a7250cebde170bddd052a2035412dea1e2a1d59ec6d959c71636076b31d1c7ecead6585702388b652e46021dc03cd11777d94b1a98dfefafcbb27d2444c64520bac19a1c281530b6554a05ca6062d3470b7ece7e972a7cda4126af85a46cea729982b641a60b866ed5b00f1cfb84c7b9a9d1c054b65d19a19fbba7d5f7fba8b6a873919753e83992bc23af4e2ff2126b2d5815b18da504446319137b1d147095a8014c1c489410c85680dd98a5c686c7c7013d3b907f7c82222b8eda0ad1ad0bddeeffeea8e4d4067fc81e56d053ee0c407777b442c4044c2efc6d1578c1e5bd26b20429f668214aee6c4317bd6fb739b5753ccf64c60baf2e9298a0a05e8dddf6b11de95c13b62ab6ad4f1f3f17a5c968e49a640d127dfebfeb2d036b1d9a0959c8a934f53c964b27949bdb3c660e816809332466c5f834b467879fe528ec158109e877a41ff5bc607a3479f3e348d1bd61823ae21405d5b58703ef727289cbc2ebcb624e3ce6a08d89fa44adaa3be48ab48975647d588857b6aa484adaf1e00b7a5fae0f5587f5a0c666b2dd377565ca4b6b7522a3c66724cd936d35433f9517a18a15790e7e41f8863e80432d8db3f9b1ad336f0bf9fd06568788b43107947a319a5b349af5694b0fb9eb4bf012495d6bfcdfaab129f8e71727520afb7c23696d3bed2d9054ada4562eb377465e9d740444b2f52c63f936ca78c6855fa99bc9d5c3d0e58302e7c247d195ea290ec8e9f149b961c043e1f4a9cb9c4c99d2c8c384c3392944ee172efe95c3f782936e2282e2c216c12976031b5fc46e3c0532bbcd1c5563a94ff29a1b3d087cdb604b65159cb3884dbbdb635b4fe23b0f60fac17b7a742905821e213edabd9111cab6324c2f8254310e590fb307e059934fce52e365acf3106d36c9c94f981d3a35c9d49c897cc8526b211ddff36e478dcc1838b154b15ffb1a5f34e1d59fbd5f237553b3f731cb3d30140bac090b55249e70a58942b47109deaf827c65ab7853903964b5717bf0d649257e942a584bf77afcf1646968830ec2de9f6093aabe2e9cbff8dd5497038709ee81e9e8aef4f9d13c42bebb02328a4d0ccd9bc1ac6d89510d1b907a1ce835459af0fa1f67033d6ba9f23172173f7feb8925a4ff1024c1e0f7eb7c897810dbacc56042fec783aa6d98ef2d15c000df138e3e3458cc71b6f5936034437fdfd146100353a90358ae581901b0f0b34bb7a5a93be60135ead6d4bfdc97ad929718fe7f32a3373496aa89c0477c91a540afb3a1e2f6ec4024ebb280ee6c56574f981618ec094e94c906cdb45a724a9cf83f977a5e4daf434d3dfacaf9f5d858c86a15cd99918deb20d464f5dc27771f8f199687e2f2a04d694469b93381ad3c9145873ee4f9cc18fefd99c56034278cf9dac667c975be616a5eae4f65721c625c91f7526df2bc5a89853965d38706368e3dd88dc21fa9e6d7aa150dd64cad1fe389d42035064eb1afdbaea53cf91b4777151dbddf8157764527d4e16eb8ff9e764aa4c550c30168afad3f17aadbf08a8f86c138684e457a0fda3e3d325d145acd74aebfec8d7ac9b7088aee9a70c396fba572a7fc58acaebbb3706be9f30a3bf85f5aed86d647735f5aaa9587fc2e49f62deb303e3486bced77ae344e84247eb3862e3a8ec951c6c23d270e5287f7253b44e9b3cad27881bb3ab990f3f0af07826563760b6b5f62b647844c66ff5ee3d0d67487c82de6215e4c2153148b95d594a405796c6e59dd32e3801dfda9273a41a31e401e7ca23803864f8a05a76cb85679e39b410e7e9e9f9fcd13b5b7bdb5a135db709316931acdc6d7c4ef77683555c7de4b4e967c38d93af8c16f6ca6153f99f39f2cb7804214e2274c7c60f01f64071325d1268a265d500acfba04a7b6ff8f0ef9e87321764b5299e10388691b65ecdc6e7925f33f296fe94df84de7b46d11f1a89a61dd0da8e8df8ef10caa7a9c75ad9071756a310819073e0e91e73ddbd02c7ce7ec350532af9ea3a3d8887936bbe96878ea4ca2cdf85d403bc75a3d13d31e0c2f2ce2a7e24645fc875ac38d80cf4b47c940c78e76b80dce6a78f472d161a8978dc184014ef7095fbd50707d0eadee50a9711881e26a06187f76b598274b7c87cee7b73aab0dde7e46f4bf6c1131b0174014931dd9e9991774820781e1559a4e797a17cccf38a6568c389cff2437abf20935283a10b69709979843214d47281a755fe100a41ca9d06d2629ad31c88d790d475f47f5e7f691498b59e8ba8897a248537466512cda8b02a820acf046c01272dbc4f24a69dd1ec3643e34a3af30aaa42973e1e08f17e615e97a5d533f0df8668ff4e7b6bffeb5d7ba59dbb52b56a042a443c91b94b2d5cf08426dd7a304f51350e51492743b8a0789c9d1e6b478f8940b869ce79412bfa378e122227783241189c1ecc78ae2a303d832665d481994ee3666a4725ec605cce50bac6431b7414cb4c28005bd1f66cae78194fdbc85a76bcd45244277e2fc279c8978e30cf5fb82f38180fac6148d4f776dd19164a39a3b86bf70550fde18da2db5b5eba16edb294cbd205bab6eebfaf5830047bcf86925938b341c8495b4ca02bd390b929bf375ce7c36b7437109efdef047f1d5476810fb1b477ffbb18ed6db629c86e96435ee46bb878268f53b9cf9f71409874f9becb3dc4af617321e903de270d3b89452ecb0fa103a2734c2adc6fcf43f1641c3547b4f628875b28bb40c3ec39578eee90b8a819e1d1a96e9acb2f15fae5a9e352bf1cd1d452dead4b02550277f7a1bf764a740862001d484ddb7681ef90c212ec731dd940cc39647f0f7da3c91550793c3b022129260e096c9f5e99188836d7c3eb4845fe863f4efddc242320909836d65843d2c7c5f0bfa7060ced2e49c1a6447e792ecb21d88960bb28135ecc003241181d95a2c82025a2514bef68bff1e78acfdb34581d9984ea21c3d59cab6af4edc72a33a9d95418ca78a9c2b72ad4c12854782d6da6f6d2d4af046ff16da9dbf08b1d3cdbd45824a24e5a5e1d22ae67393fa6323693b063d2174f2ff4575db8b374fd8e30a84f4bef70d27507b0d060d83e0ead50b42a19ef7dd0065cbe6f30c50e5169a8a68bda659032f3b593e914a017a667bedc50aff82c109a08f0206de51a3b06880674d86677a068f7711ebb4a4ef4d8d221f3df5d1f6fd916532fa80c228bc157c50fb239076be022b5d3db6c68a1a681137018f41090764db372324cb8cea3db5a5920fee926dd39c35ec017247e7d89a2fa0d5aaf6cb2b1206e28e6d1445397f5df81568233f41199a2489216d1a145a353b7a98f6b1f51a0ea94de40766f8421b612c1a5d86cc42a1ed31351d34870e909c34ef4d4a9452566b3a148a7385588f8c43bc7dce178350406424af7ee2086cd260cfa6ec23b7acd5131b2b8952d44a587a7527aa50f63f94e0cfd0114ce2f44bd2cc356c893aa864dacab07dd58259f9ee1a590ff8e775c26c7687ee0c2c0f9a44752fa774f4c98d905c8f952f8c5e5ba8ecb913634fa9c9be556d6ba157acf434a3cf788bc68d0919fd4e08347fb4b0dc9cc3666daf7da9ff8dfc5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4333478e1b7c8252288fa86e88603ea9244631b9072049b1536664806a6092feb514ecc45d56188ab74dfc2e1439185c0d4b1c4e181a2dc66e587bce8c8d4d3e58d403324f66d84a7fa2694b51e479e3c69811f6fe5b1bd0f78abc57961b795cb666173461b4b8032497e70c77c3c355644e155e17e9aa022a48a247cd7e2f139ae5dfc34c77c77eca5ec773c95ed194fe5df34814280c02712b249ccda67f53ff93b0d21ba0b448390318f2ebc752c0060cdd92fd2e15a50449ee7e981d400a8615d5a875c9e35beaa13f6fb1f0797b92e195c42d7c5cbc17bd662a79e042ac34d904ce7160a051dc958360e7d333c3ba17c9e7f943c5c5dd0e8dfcee3436382ec06cf81c0107b6c382a2260b5a2f5b3db7f213dafa97139a1c04984a6a62185c7f7ab9cacd7a0c800a0674813a8a452df019413c46b4347945c9d41926c4be4bcd51a4df7cb22164bd5b02bc49a85da4e4bb4027ffc0d7ec40d0bb5865000ae3210dca5aa3d16488e65bbe1882bf452930872663ee95e77f30ae8aadee035fbaf2683cb1043f36a3f8149c9c2b3b7b98f8473622d4bbc3f6f11555303c6c223a0440979ac65ee45ff62182d5c81924800d7a762bbc71d497f16f983789fff4349a031e8fabd7e62ad2dadb875deab597332226565c35aca5cfb6b9fe8be0412fd8fdf651dbc4a09d48a9392788562cd63162f83b9546f58340e978fa0205019949769403088a09087aab5a757ce337372113e3c6e05f5ab76304331b40425daf71ed20057cf05b07f1630f176f475732776e03fbff070edc2fee429f086a14cfe85ccff4ef16d51da06af5d22e34f7b2b34bd977c741f57c55267143983f77f9d5478f51263698927fe38d698a60d1cb3216fa7be513740369b98d02ecb67d9bc04b372e364bb277090378f00f7f9e2b340d6e4549b3833cac56c9b415f3e75c5a68a3dfc8dae1cbe29b15bba4931de4115194d892e6d2e96c06518b78e632c76f803da9c38ca3c9b0a1185cf148fdf2ee5aaea42817587f5a2bcdad165bf50ae31fe9ef7f7ab5578ee3aaefc727abb9701d621580a7fdc524a1de32ee8fe9a2189744930a73a5105e1f32ddaab8b23e122fb554ebc4b98dd13cb2044122dbc1edfbf54619a7a7d3b9da0614fd83ca610de39415c71e45fd9014b38bd9b4e7c98e549843a2ca399b53c63bde4358875b2ba5c7ea1c9ee501b0ce9245790b02556e3b3dc1609eab2207d5e3eb7b09fb2c1422bf682256f1a5e8af1b3a4f521115150d91cca13519273bb496ffb92bc001aac6e22ab3ba94e1b073670ead7ef3203016185b06c294470bec985abeeec3d6000b22b8127dfd350e902128bb48d48116b171ba59488c19437a4fa73ac798bc3645b6add7a7fc8064567e88bde232ca065cf919bef49df0f9e1f9b0bf4713df189ba70b3e8bde6f8fe2dceefa3a6f7884d7f7ec408cbcebc8f2eeb0ea08112ecf4fcb994af673d055c3ebfd9e9b97685f7e22312392574ce156d27a9fae7e3c26095fe4eb39aa543083bd146409bafe455649b708685dd9d7c2f1343da83afb183c8092f39e233121ddf39c169347911ef1fdf2cafb6c781500549866151593d4468c37bb142646497cb63a74c3f0ca5c9f89c5360e08b5a6ef8b40e049139e470efd06795779d7f07dcdd717262685925290eb2bc685fa19d68b2ebfedebd65188c8d5e9b375226eaa071f7328a9fe183c246831f2cf7e0d9499af825732049b8ae593a6e67a47f6f6d52c51ce2c8206e398e5f94a2fade8416af6d051451ad00f382f39f3109a5095e2d4fec38b1f040c01d0c228e29ca590b54fed843caef00a691b4f0e00f53e5225cc93a9e17c209328468b725310528f718f7ffbbb02fec6ebbac198e1ab9b1a1f78cf99d47620926797aad2dae99bb3819150b127f4585b6d6732e82e9c7a94d7f34941b83686db7263be89b050f3dca4bc1518b61bccab72d461d88ad685744eb1783cdaf8fa068058cbeaf060138bdd590fc565700c3c28efac381660512f7a6d51b928ea24636538f1e06e59b5140b0dcbf953bfe049a0f2e698922984ee43c0bd9128897df9661aaf3a910e6ccfaf4a85035099dd86150dc041fe3983d65352b8ac50997087b9b9cce2cba959f7f20861163ae854e53969604019567a3d07b9d7355a62bdba9d8bde8ddd81177d5f32e5e612280ffb5aafbf1972b38fc40b476afae18873869c2d4626eeb91c144becdcd321d74232fd9e14e7ab0af9a5f3e9299431c7deb47dc59b03751943426349f83e2acd0e5e1487582c1d8921c981540b346097ece41c7064928447cfb55011035b665ae813597425f1ca162a3af98bfd6351ff99483ea448bb8b37bc278722a4d4f78da6f0e084adaec438678fe6cc3a1725238ecfe281371532ff28d3e7e072d83e77a0f7e5399d61656b9ae07677362cb2a39d46ba037e66cba7cb27c66a1bb78bda1ba03260ee0756ddae4afc54095044d605a898e3a8b2a529e24d4b1a9d1b66792d849d8ee1ab200f8a38c469ff74e334c3ae8eced286a8ab50dd9dd8dc44b2f6376840f71a3fd43bbf665b30b8bff421e22a71aef1ece57f65ee3ec8009bc91eb3df18a77f9ce3b4321499f46694d0c7f01853464a4d49fd83fc891bf543e5e459812e8c78830eeaab55e541d228758b2cb1abb2b6a81a328b6294890eb73c721dae191063d547390874ba6905d159c5c091922f138083ed104d5f036b11c8f8f7f94e0f940132f024139616339a3d230a2e7d1ce91c31505833d02591ff8bb8d1744dba6fa1432d68ae3b0a57977c3c92c15bf7dfcdefe7a06f7c0bf796b1ea09b32cb99d09772e4afccea40c288af3a83e453f42cc73e678b116fd6a09e86f05bec2459297f0df10f1a89608148f29533541efec63b047a761aed8fd0c535346a6d79032bde3d8a74d3dc8c58ea4e4a1a75b2e6a042a470c2c84bbafb6a51500f5459c865d8c6dd202125fbd873ec833d1b8353f51d0892f78306c7d72d3f1bcee3aa034a7bd20256cb017ddf577e93cbe63a20ab8c5285e6e6dacd95be46bde5671941270b2872df8bcc83d7aabb8ec576442b9b6fe42d3c9037c8dba96c68326ccea555a1ffb54a44c7380d628459cc99b104f60879ed617377fab3605bb445c63e13af2aacff6e41942705c648df9131a933894db00a3f9b25ec8903db3e6b6a39a2b99243af8701a858ff1ce0f9a89ecfd6af7ce127c88ddf9325d188644fc4895cf6eb86e2723e89ff17eeee61733161bf5f7b7f831fdf286cc55a8b1dfb10ee39382a48b22e1c302e2ee02595849bb624a3275dd52ef7ae8d07a987b17ecf73fc027b60ba75c4a34fb0c210633fa2d9d8daed2142fbc94b56f11e906dccc805af7bf8ffd0ebd023532f4720bd7ca77a0ad1bd47f3d0595dfa51a9df13d4f5abca7ce488bc06c4f7502221ffee85fa9450f4a84bcb4a7fe5b53a065cbe5df6b3289987291eb78ca590161f75976107758ae0ec1578b00ceaa5e4b5ac4eaa4f90ab33bbadf9f92d3f118d29e7b9b78ff7af8cb5402ba15da96925e44b65f0b5e100e27896baec89363a802306210837e1918615de7886a1094b67ce1c069b57302b32dba349e2b23856d067846dd7b661e72ba5a159c4b1c73b71577c853ff7b297d4c430d5998edbe95fe15be92bcbafc9daa447705ab675f2094f070b0fa7050d8d345798e8551af8b40c194ff9e88a89c202cc38ea118e378430133b10c04825e4716c9cef15299f232a2b08cd4dc80614d4f266c17885d9304818c23f477e2611e7e13ee4b7b76fbc41cc9ee42b6e6cd1f03e81ce8ed33135f2a10aeba0b2c15d833842aa5000ae9e4417d2dd32a56b5473628d25793eedf873b50a4b2be517be5aa52b359838b01de9467b290586863335af38b2c08790eb96ae60d4431d93bda6fdc690d04a274becb848fa9e5629cc2c7c79d50da727e2e0f3fb81ef31b295955e39ac2bdf3dd216f7e16baff84cef95c116b440646191d17862284ea672dd2be915b3cc29f70e73a2d14b4578823f9bae881de94a005662f137ab275bbd1e55d9d9fa0961c4a058fca8af5e6647d226e2c7315b8b53b93550e8e2f0fec5fd6b54aa18cb9fa06037644c5ecb2ecd6727aea8b4bef26c32015650d206a9f246ef38873c76c1c0bfa940dc2b78d117c4e450647b855169470249bcd23232b7606f72d6adeac09aed19fc62f7bb79119f92693deb9b5ad31373e58473e5ea57c298b390f0672447a954c867994df655175a7aabed9b0e9b0f2506eb27fb0bdad99982170ee8afb6b7df249c607da87c0175315bde233cdfece5e272904db4e0049f44fcbf2367b0940591e69980347d1bf4005857aff768da934443ce85fd04b07aa2e235ee2035003e5ee4db969a4b9c088eeeeb56e1422e23a17bc0282ee418d79e28b371a5fe412b3be512fd9da6dae47eb56fead38222c2b78a0c30bd9cb645a5ace567cfc7c50cb16dc88d8a84eba95f366302ab3fbca2828c0d8491891e005a4a97394edded100883c5614221b0e791b9966f6031c7d297fcab28b6f0feccf85751afa76e509c5cca6b3ba91489bc71e76e84e103a712ead10235ce77154d3a5db41834df32f57d8e4b6f6514a94d5a3fbf4a347ad604d306bc08c1b606aaaba32305388f5be767e8dece8bba0a4ae073a1804c1dc6e34364c0e41560acd852ca59ae2a7ce2f0c7cb666e7a74d54d7583dd01c6f585fd2863bcb6bee43e0e1274b3b1f05b326b025d9a32f06c650c48530b24a0177cf83dd8249fd8688bed92a26758d4662343a0b873e8b9ece70b57b267dfd5102ace46d84ed913a9544806c0b397ce06e6d3382ae5869e3faca32d322ad293b57cb0362f6be1148f2cb5d63b389ca2c9f8b7f8be0dfaf5c0a478e7aff858d04617d7f58d9237637c538519d20b30d73040adcfe0ad7db2f3c8a7e64d999ad2b755e3c3e5e2ff0b7a3d20b76495b9426cf78ba3f27d6e5c937ecdbeb2bfe30cb92afe4850c356c9b9d8e8c5438427146248d2e3aa3e4e544a8d4dcf201cce35cda685b1e79f1406a919de5b41a2a683f4164f8f7d71416923270b7e99514a41b0129ccff301cbfad6d7478a541f9d77e62b21a9632b93642cf60399099ae679f4f92a9977831e505e080a6473a2289b51571a14390aaf01b535a5cf6c7a1dc1d7a36bf0bb103c459e0987a67e587a23c55626170eb2d3c3898e8f4bc4a90c49b871769300efcf458f20aa83392ec7926b4b7f0639f9c597438be5a6590c2337fc949675e09c26ebc522a4b8e7d231bc1b67f69a61f663a06d2dc791f7a8d4028d6a0e4a09c493609636907ce5b8d0228a7a7c3486bdc75f6f78110edcf185d744d5229e7de513b261b87e8c4cec52f8fed2365ad4cca5462109a86e456a61563e6c6b22642d7681aac8ce18a7027e75dd06735e9e28a2dbfc88a6058f392921d3edbf0a79b5525962b69a275e0b4ba02680b87a6e232b4655cafe24985bc5734cdf794;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h31b5988f11763937d8e5ce2198ef66df58e0a4581cfe8e2d7ab9622461a1212af919c8492447d054cddfb758bd6d39bc10b1a270ae9302775a8014e8eb51d837cb12d27ea23305d46ad54a014a4dc36254a3396a0595e81778d37c9c22f06d95089b4c6cbe38e0b1b6cd3236c10ff0580dcc54cc4566d688846d86801992155df1ec5464c7b5cb267911f5f94af32a2609bea07693db7fe1ca94e35ffdf5355c3a6b64ed0a1ed985b99cb601406edde15fafe9ff629132ac33bb1a186993f7b789992668320f111a04182c4051abc07d3ce969510e03972a8fe87cce8cea9383120ae4dfdc71652a09b2f783e9fe1981ce9b858fbd235b53b4d06acf5f6bbeca407e5309e5af1ec1a35734b9016c8d5d2cbf369628a4480979e4880a76b0791c801ebeb0474dc00a90303323732b622cf46557d4b48c42ee6379cd23c98a353a4497e5ee1615b711757ed403790f2cd67c2fa27db8f353971fe3a85f4f28188ac37e7c9b0fc44a473035dabcc798faeff9f9d1972d6a794343dc06a8ec619f443339dbc20c9dbf6485ea5cbad4e0db93fc9f9b9d91168d08d6607cb1192343f9ba286ecdaf6f085d15f17757209fad5caea451f9c34245e9cb9d56471f881eb5dfe09558f27a0e8bfc004ae74b272a42c6f08a63de961b00e6c2f9ef15b48bbb45bc5b0f31dce185c16e0678660afb14e47c6218b36638205bc2dcfce3531be17d2bac65c4b61ff5c00d2981a7b746685b813c590c252f8a6bba7468e1ff8cad35bf6e8c3dd5a63369669c9a8b4fae6fd1f5c1a5dc165089411f82b6f1cda5ca530b8287af787bbea7ce7659b0e94d655f27559d8d6f305d8e6e3ff02a3b2b7aeaecefdd23fd47b859a04ab3ac5d3baec7bce90f9640b197e33fa300c5a6446d2a88ca11006ba8267f89aca66ba8dcffd8a745975960a091c974a2c329ec8be13157ea025c9267ec0962fc986fc1c86736f6c830c2bb41db8e18f126e2e4611efbd21a8cd0441ffb3afcec2b01078ad217aff0f895ef92e76b9090da2e1ba44389ac3ffa5e41655bb4a64cd6bd29da65980b9050dc0a482b917d3555eb9d183620736d44338e516d27afd2f2c3e48b8b4b064515c77e18f28e24ea4aeaddab1e748095088cf7bd054a00dbb4875f89b80518c9c1bb143f48fb930e0bf728f10841c5a8a986ad45f47da2822ef8e917d1e250ba272b8d2e4af2bcfd328758981f848930714d1c0f34d9e427cd94c7e95d16b90319dcc4c69efafa5d307e9856764f2767aa4f8593a2fdd999e5c56b830f782184d10b3c2556a45d4e52dde40c8d6b3b62b69bca0bfaa488e09542f128d4bb4c77bf4586de78405c75ea79b9f2d0926ecf9831c892b030199d6208f0a9553d13c147d641bdc595254df62e2864956b820fdc450317151423d8373729b651244096b0889942bf22c3101f93dc7fa38984961a0ccc887a3502775d7b41a314b697d2cc6faeb3663af7408738975e16859192f1a91f689d49044464748bc286ad91e68f6f79863e45899bce900eb1fdafa51ef51aa114daffd9dbb83ca4946c1f1d2f255eb3b0184d5c3029a6364084cbf7c084bf85d190bddf8c884063875b1f230f991f902e5e26eeab3ec6784e0c16bbc86affe0919e240cac2c007a42b336ad1d656dcb76c08a77a5db40c60eda9ae9208ba94981b1b5db3a03a97df8cb0ceaff466b88f5051f6374e59c19452af17bc8f909df452646cc49b15294cc6f1501b6d1ef18c3a0281dcff8e67944c6e1ac8135e27baaf57e6d1938a08d8d29d018b086e8724952affa0525925d8d8087c7d673d2d7794dec4cc0d6423323c4ca779e70e775b774d199fbb61bd1171e4f75e6bd85ea417fd431e3849bc84d708768e0e1dc5c9efaa441378c3cde9a4ac564eef3cbf7d812f8b18cefde2a47ca13004a6d974f886931a6b4bf340c2969dfe8b0f060482620a6dfc5f594535a12c8082909dbe53cd3890d801be9ab46f116cee22b598146e722c13cfd16af936ff9d87b155f753b518ff5e6c2c8613c9449f64ec40f474cd7cedeaab6a7ec7dfdc1156f839365da5ded5325c62cff0ea8fbf6d93e91c76d229176266cbc4c44f986e2b8109e3bc6ed228c53d66392713a6b35309dcfd1e9acc3c3c9f750f54d7f574c315bbd4e236848071f9c5fd279fd2167dfef6424f303c5f3cd9ba66e42a94b283f689d9734878352e361d38386a7efabed0784d9997a16252e1a39df6d53453ace4dc20a3800081be07f18f296d4bfa53ee2eecb8ca55fd7e637c575a185519d8e6194b7c8d444f3ddfd7fc8a7920a6a52967f13786e36745a5e01ac14221012539b19baf59900527a17a058017b4ae43fedd4b6c543a9ac9d38b217a7f58dc50919c939fb18e168be25cca8bc53004379da1fee9052e4930dee9a9442b363a2c23ddaf05f5bc138dd3fcdf2b79178d2d188da09c429a0e094a896a66d771c2623f7eaea7310e092d3fd1716ccb6e567d168f48bac3a0d853e73374885932fb9fc9ea9e8fa3bf385b69096a5979d873ceb84fbf426993372b31a28e4aa116380724bc9e03d03a89d1e5181dd641a0da59967232b6a831c92772f695e49fda4ce11a5227dad33b01725ddf880670fda870f56c2447ebe0d0bc4fcec30699594b6d0e74bde57aba0d8c94039fe577c8b9b942aab9d33a6d5d542ba05e687be520985cc82279a0015b21e4a99acd7377a5c3e8580ea548a55422830e791eebf38e03aeb6fb61508d56cb11de904ecb5fee219f690f356464053ed45ce59bc659c89e04850208f300b22b7a71be26acad79695cf9c9b66e7b1ae7e5d4023442d00e1fa82591455ad3e2f348b9a505db7ffdd03adf03cc1add5097b1b53655bb31d011958e8fdb98daee88b6dc792410e9f84f68872f52a405f7d2c43036da58d343e01bebe0daeb5441da34ee3b3775ce48f673618f9a87e41ece40c86c79c4d411c4c304c0db00e9a5e5236ee1a924cd0161e06ede9eb38aa78854145eae6a6609355b4f5811be50d4abc41dc8c0eb195de3293c4bbb13d220c75f18c8b76f04be291325db599cfb25f9c60484ad4602a9a90e8eecd630c7ad973ccd66c041436e9df3a52bb6e450d1979110857ced4137d634ee4cc37e161de440613c596c2cfec12cd1adbd67becbd8c8625ba22cf938933bb3610a525ec58df6b5a28076a59df5d4b67677a455f2a7a25db7830176abff74cdf646d69f222f066c85dfd409aae2400065d5e63827ca53c66a10ed08d73ad9c65a47e2eb65654a4f8534027da9f852abb81ade5026ca07e69a12aff620f414c2321d2fc0b32224c0105ab91cbf63e1682153b3082a903c3d72e21f4b2d393726329f2286dbdaf34ec058c9e5117c45bc15dce45d0af82e6aa29b295eba68b14db2a180e1fdee0819249532190d7e15b9b2dfdf9f63e14975c6c84b21a56523e34fd7ada731434a703544c99ebea2f79334e12b42deafb10ccb241cbcc6a595f5568ebf0ea40b4b87be9b9c13a760c74586b6567a65f5f47cc5a4df9f44941f592679a9b7bd070b6e2aed81153b59c39b8a40fac19e39692381771cb5dcbbe2036b0a941ca4cce26b7425a14b4fb781fa12cf8cdad32cfc3a846eeb75d1869e3635eab870b08594d148a5a19eef2eab2d158842dd33235f36591a347a77e9360e690df1d972e47b0934d3516c84d1c5455349e68d5a7a4b3a1d1d8c22152a1912089dd5196cb0b60d8ca9bf4c10000575c0711417441c68aa43711ab72613b59e96bd0c4252fb675732c211f207c263730d7e62e2aef631312f1f12a29de9b00d1f2b08b4ce077789fb85bab04a9fc1ea77baa547c687b171c0f902c79d12aa97091758edfafce1d97498d25c2387ba2b0dde68c3604aeff0dd63b82bc97427fc20609bc33d13b67f8c02a15a14e31f0507effbe1766a35336f755e81eea7df08b1d1b57fd4a7fe4d068445911b158b88bf6cc3785d6c5406be2c3fae0a8bba1abe2728c9bf8c1b81354cd9a373bf5248feff3f14a0c6ac4c389a8ff1e58cce93c753fe3b11456f21af512d379910ed31e84936e998280524886f9ba5e7dff519034484dc20c89f4da1e6fb5411e019c09df1bbde8f9a54cefd74eedd5e3c902c3ee26e5904f30dde00d4fd807af474cefe88f7723b4acd6f3721a0f162b2768271360ff3e8fd61955ca780b0b537e8ad9fd23a5a7a67c40951f4e984de6e419e2aec938b8a706275421a1a239566a0598ee7bbfb96c78ab584555d4d3c5bb15273d0a4197ebca8ecfd3a90c136fbdbc262da9987ab4160b3fb562b509f56ffc28e439b753671a04abab01f5241fc2187ca30a6c1cdcdbb5c49282e8bd29745b48e44539364330d71944dbc453615767e5f906186e73d97a71c047aa653be6421fdc46b6d6474c4b8cc24470e339edbf3571cc44a2de3b62919a11f6f69dac1a0bb882301bf0ad3d3022956864b6f9e4db68b57e30c8b2335887efc716fb11a98500ec56bc3dc5c0a82b0252d5a5ec8643e78b84b560ff818a6beb5b709f97ff9be9b2b2aebef58a1a186f60526f4b3aced41b0f8a1ab399deab9f0917257cf3c4d27eb6dfaf01328c2da6f4790043baaae788f0dec2fd268ca1d778ae1745db80a2cfb6150795c917c19d2bb8f8ecf03cced966f98cf4b65f03f53d5162f40302f471898a33d1a336ceff67d55938b54b65d6d09c55f6239c12a61b1c31c4dc5e7e3554b012f97308cc55b3fb8d3f529309e7db31615eeef1267f7e0db956e9e47ea8670e1c16bdbf78264a6b67ee02d3954aa322e3f615b7ea2d7f9127191827b8d1ac1edccb6309fd0f17bbd5465a22b40a342995850944f8949a811291f9c50072f713bcd78fc8ed922fe6de5d7861429d7567144f442564837ee8d0e4a5c230c36eb5694177b4df03378fbb24cf04b97bc10c4d81a043a02f0dd728e36ec1d92e88ee6c207319f02305c954b843081f22ab8958de3e591af0871b9480c2494003212438f80a1ada4c0d89a81f7e469b4ab4f0bf046a88a638640579ba3ed881359bf10bc1464dbc6ace2143dad7dc0e2b4b8b5965c73b47163170ad053a0bedefb76e40f988175ae3d5b134920324d96c0f491a0ce66ed3f2920b024880601ff20f0ed59f8e0dccc984b36cedef1b6f562b1400879dc08e730790e851877daaced977587f8c31d1ab1a2d3a4f008e8910bdc6697ca202165d0ca7cf565ae7724a3f0d549dadbee636d513296f8304bbbcd0c2b2bbd8231b96237a484a1076cb80af93f3d1dcfb89a96596eb783f9ff327b6acf4016913375554c8055350a196daf5957c77a5d14120a72b06bbd295adca31bfc14e2ac8285482d8c21352d1e11c24f96d5476a67cc14666ca90d146b9912b5e9497125a316839d129663f7d10d24f1631165ba86c06bdccdffe5ff71be83db73ccf4eb564985f074472e5423369b3972d56863ef0ff74332c5579f4e79b74468a23386e11312de724597a1827d3e41dbfd3253994e502;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he58fc237726184dae05d3b7c4bd89d049e53f77fbc2e754ed91e402a56fbbda739134d32908571b25136d4fbddd532379356227cd43b3ed742d7ac3762fbdc390a5780eec24a494944e59dfe57fdfe43fecc02911424bbc770c2bfddd669656e334f14bce5509b6bcffa4d7b114bad2e1881ccfd161817abb8a9f50c791047baa01a67e66e2017da9942025ac6823cbf91f147723535ae28e15bb63bd900d7f3579f416220d6657e3015488495db5a1133fe49085ea5a9ce163164ae2b826be00a430a3e3332beb36fea8042d0e7a9f70ae408844866106fc2606239c30c674b0cb1c9518257938c0beaa7c4ce394b59bd3dbd58f24a781e9ca8ce97e9390d5f9db97ba9e5c3c70861fd7708a23303f2ad44a0e92155f1111adec598df8ad68bbb97d059eb0de81c9938bc277e0ff3edea736087139aa1939623b72ebf1322a14b5004f8ec1a5406622cf4bf561e2d4518e15e2c508ea45f8f2b482f9b3d3a6650c2e943674c0e1997f5ea599ceb5a36043fdfa7c6667bac9a12187643ba0d63c5ebb034f3ceac983b6245f35f3e843dcb6454d57068fbb6e91e626b9241803c98affc9398ea18e8bed350b5d0a9487354de8b2a02abf4e2c615db8255c95625974634930fe20dc772e9b69b1d27394f85a3e4452629436550fbbe90f7d03086441958c02ba983a5cd78fd7b7dbb0b2123830cd9e713cb5dcd892c30e11cfffe1d4d2367b434725acb3e76eb00094473de927ffc2125bc98d79769304dfe753f9346ddea46d53eb99d7e7618861763271b72f48ad22fbd6ed20e9029ff672a2cad3690e925ca92c92bfba57a79b82f0a148b3b67a75b2f697ec2e3e81b86bf005214804695019092d018674caee24e1ceaf145f185dbe868d66235ea046396553c830c1b7703939cabdfedf928c9ac2f900e03422fc9f81e3dd44ad790ab89dd43d5a96bd56598cf0a0e08db204f25e6bacb243f329339b1277e833b91174aab38bf98f369fb06ed93a0012777f916e47aa9ac6a5aabd819163680ba8496aa0c971feb09b595df33c6cc46be6bd39e2cab3f9edf6a8129627be2c96a6656d5ecc219b63fb761ae74bdd9d1f16e75e9111b834ad690dc380d84bd4f13fe8b87343438cef85a896632f6a967e0cfa996c6cdcccff5cc6cc27dfef05fdc8abbeddb747fad0c53c87ae90e81f74a7c7967f8a12a2603e2c9b0f5f042b14627ce014db9e6a2dc6fa018fd0695cd5810f16c35a8623b5fac1518bf6dfb9bacd6ad31ca9a730e4d9b2cf9c26049b523469a7040f1f413e674feaa5b3721d231ff18b8a8d06870ddd3620743841f0bca39e338e1d931439b5d700fedced241aa0f11b243fb3884f8c7e8a374f46db8bba1ca700edc72d5896bd558b7497619c8cf9a88b5ff349daf85a14989c3e664d9dfd6e1238d90c1eaba658cdc5cf516cf25ff92d4392be43b18eca7335e097bb22e4d2293e10f18a4cea348873511cf70c9e12b365f21a3123be421162e2f4b7c8d797d21c5c08a04efe9dcce48b352a80e68c3603251a11caa8cc4e2dc3731cb3222e7eacf6a48135fd5bf5489487bb6a0ef8727d134912998617c056d3535ac29651c5ca5234eb986a7500f3cd975df8d390aaa243ee88dfa1a196b680c76f3679fde07364941f8c6609b4d16bcb47d3a4a955c33e1454939bee780d349166d8cd0f7a41769d1817c2708d6dcfd1daf1fe9e139e48d897bef481a2d8ac962846af0e71682285e471a40cebd6f376c4bfa7909ae95cd1af78624709d044e157c2fa6630ce728ff83a3ce15585a0dd32945c10fc27c80ae07e3b46cd21e07a82ed010727f157609a78b368d344677f6d87f8024be50128db109a2a218b4f16323a22218f15fcb325e6f2c30417ace14d706731d071cc8e222d57ea15a8d947871c6dbf43e3107c23bf03b3490d05fc8254d7b8a7797a97800ce084851baab2cadc0699a33ff7bd237ef717c814d0309cc21046fcf0f1a87dcf3b5767bba700454673b95d7278637f3a96941a67df2b21e656a501db063864b04b6ca7a4e7cc8e422c79feef2b180277aa43fbfa03dd000a4b610f217c04c94f6d6ead03724c606efb848dba24cede659e4068e5a4e445bc704a91a72b909e8c39aa9da242821f115512807c59c39e2e7fd16882051d8a14744265f07ed1d922f045c7f2a328f49a6725af8aed3f9d2a7a92fe12101882635231d4551ae1cc54b1274d5a7a90050a9bc6b0329f52d4bb5981954452a67ca9c06267ecd7b12bc5144695834c351a8f19fb9c6cabdf41f91f716d83afb3e114d1cea671370ebb7d5666192fcdf64caa025ae74d71e44baa107ad731706fc05bc5e90cb1c73693a937a8cbb7050898444c56d0606490706e3343e66dd8a5b3bfaeb2953fb47e7a4b57713618a5ca75ba273fd58b9953ce2fcf33fa3e37dd984732b68e2cbb88d4a619750732d21ae2b217e79fbd08b09fed059b6ef35f794cc8047cb91c354704b9947ba48a064ee407f7570e81a62f68422da51b88952671c482276fc89ed283fa8d60856c3d09da3095ffa1bbb1fda6344a6a5e89990d8bfd133685f58ff1551d8ba288f7535eaddc0a066eaa67ad80615085f3cf6a5d239e99774a9d9857614baa56b2f41ced529e1e5f24485396944d9b13b6c598b57fda73cbf08894ab8988808f5539fffa452847e97051de0cdd2d588e6260a05a1290c0547bad8b1a7cecb70920c698114c0709bebd9a41e374cdfd05e8d0b970a119c4e02758eee4634353935b7f9e3d79d2bf9445ff39887f6483d5ed91864ffb91f41e697505af8ba0487075fac78597a1eaf17dc05c712f75dd8a04f73fadd62f4a633bc05fc985619adb29c10c931ad43c8ed4513ad7a72251eda7cbc1a2a2a6765e0ab27a6cc322a3a084d8f053df451170c7588c1743bc4875b2b893a84d9f80542afc163f1e6bf39398a72110e964eb45eefa6d9b29b9b59a268589fc3fc914b030da5f1a3aa97865986d6e612c08a55a1f1c6b0d868c8f2bccd5e6e15f2383e7df36396a6a2a849bb18ea4269df929702ecaa59ea081583fe8792a67d8a7ff52a653a946880ec1a368c5233476ff48380865a0c675876ea9a85df69f0ffaa7b0cf08717e70032883337c0aa2ff610cd13f2de4cc248e84d8c8a18f00d458fcb048a26823a2a1aa7295bb958381fe1cd15e50e8f0ff355df26c9dfde1565523c3d8c200d8b9b1b849c45984b09fb0bb6143089ce805b66224398f4bb0cded2c0463bc41c081a363c0cedb59bb18caae18c314199da29d41a6c7b14da87e498b4d255e119ee6f0609c93e2b00f7f12a286b179f281b27fcfe49c0d622f96dc86c664cd70f07ca118b8f58b4f0fad751691d23b5d4acf3a0d9defbeb55d56e3be9fbcd5e1c4967887ef1d1b3dd9605d92073679bc89693b2387d8ce3574f479260dbf71045b9735c99c25d0c197b7f31efc7b7de143cd7776d4d2148caa370b5bb344a311d16aaef068410f9d5f17fbab8522b667b10abe0eac2f06c01bf16e1ff8c2394d1a3b34d45bb5ee384a9d2015327435f01eac23362060f2b44d763e87508f44628d10eb3f4adc2e334775302983fd441d66a91fa37aa95eb0d58826d061e74e97b0cd6aeeeb6b9424709f88ac4964ef9bb1e0664ff3e0c01d391cd7ba3caa3e419795733844c418280009c31d61e91291513c4bf97c284bcb14cba7c0ef2c324f8a05032dcabd58d796c23695b97f5f3b2d2b4afccd1db046c3abe286aaffbef76d6897e6399cb824e0e6a81181b701e0f80427c55a1d97ce910bd9c7099b071123f275b74a0fe003b2848a906f139c39f9ff6c69621fff46816ffa78de913490b53959354d5e975dbd037f69e0b7fddeebd7c7d172acf00c4d7f6ab1785a0816e6542a4e8b34510c06048fc079ed542b4386e840d7c9fb10bf3f0f8a74278353c3963879cc29fe17e7c9550f1b58f8579da2fd1adbbee7ec5a42da78bbeef0da160e433e3edf1196ae9e8292ccd2cdb14a003048e35f2ac2f329abb7524ce660c3a85f747a0f73a6497c35184f578f1b86b7a9cf74b9ada59face86dd97cddd856762b0144c82ab7d73b28eb9b02c7df4735c59797eeccff7e7a256d6403e52639a6f3e0cdfa7aaa336c0459b9c76758827d5ebefbfd6c3b78060fdcb2fd8facf3e34a63ee5c35aa8dbe383f958ff8c73fc2532cd5e53fbe76935e570a7bf00341067d344ef1a99cf0acc9ce0d05fbfe2b3c869bfb9f6c78eea3abab4e7c91e51b4213c2d00aae884c9348cbeb917ce75ffae06c6a6ac9f2665b01529719a4d0a344877f9e5417afc0bf095378372aa5ba38efa35d900a6d314e4a3ef18eb46f7d51ce22acf4b8b39b4b4ed906e54736803299e970d60d1550e6b297e9843d97e1cfb38da3f7dcd1d38554da5caf08907b8adf64d5a08235614ff6faf235d3e8647c7c7dc42c6c7cdf438c81bdc8a3bc5f0605a5458d64c01939bce37326515b8c116dc01e3defa9b8162377f22258d0b4b9ba99625a3cdb51ea14f2ac52ed1a6a83527894727c3a1b78cee808c6cea3a61324379b20d706a549d2ba252a0bf04b8b752b880c827ab6bdd694e4dddaf4870117e9310461fe4143d3042003d334dc78b67c6388fbd79c2ff6323ce58a4322b92a29088a7d7ab975131ffd80f5e7103b06b363770f48505c80e24b2c3ba65731524aca1dc3944735fd8dffc778f3175788fc96ee578170ca06d2a69effbb9f75c300f269a3588819f7e9f31a36dc4356df53566a6354adfcd1a6a9df64251d374f6b0c0dd6aaa01e7e7e279e00cf8c54b927def67237646b4c44bd61b9a4106884c0fb881cbf52b0bcea46e8ffa33fa8506b3a9e85dc5a572494bfc60b3152c75bf1221d44807da9fa7fc01e6922e9184f426b569402a4bd877e55c763d800f585234a5171018bccbc9f9628e5287d02c78bcb8fbacf888f0277644880449ce44ba2a4cccebba90ed22acf3a3849da6871a877509e2180377d031462555354800aeecef0577e794a429e17fa61e529e7c657d102dd7b52a40af64afb62a93b4a7beb3e37258a8e30c3a68f444fd1b44c5b3030e1144268dce18d27c96d3d5dfec63fae3e1eef4f79f1108d4d8d158f546b1e67ef8e2a907c2c2400d90fe2e6f7ed8ebe678d9b4c9ced1f6f71b2a67b076c88f3ef4c726c32614285da0782e68c25c81c8046a341929d141c5a7b84e8b9ea9175f6b4edf5133467406ae0cd388065e5f8a7e6587132cbdaac02696e33cfef9ce1adcb283ea00ff0b15ab91ca28b47b3ddbd1452d108cf83e0d8f000ada242357dfc5988505a9c83105a8a03e171e863620f175e35fcfbff9cfd15ca30dd55568a549c5bdebd876dad086e061da78727f35261fd6c6e187eb743f193b4514c9f0437f25e837660dc916df9a23e7b1452c334bf690780eb984bf656ea1fb044e0dd3fdd2359381642b16d0bd538070200bec0bd1d320db1e2f50d29a5a944e775435e9785048861b1f180;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8003b8e378e87096d8ae98a5ba9900afba763f5af18459a5984ce066688df2c87629d632612710da2b82acda2ce26f72428637d09f156ac0b389e62f2b26da73b975808d97f362a364678a9be3cb2084ed1e4dc3d21aaf8d9cadd268ca5dd0c91e7d03c649cd6f6378b151708dca46920cbffcfe3880f8b8da28f35c001275473c205f5b790f696c721dd431cf1f75e8cb7f54dd45b82cf2cf231a73fdfc2737345b8daacc7b8fe7e73aceccf833d29079b9e6cdfb88bd65cef677323b534cef9958506f96e914c7b3005bbb1128dd74dbd2256bb20f6a1b478e881f556f954a98670cc52dc203278936c113b3050cf35eb4f6e8b2666386929f066e3184abfc2481f2576e4edde3be8ff8d82819514c50b10df689fdf498c5575fbb1979f76e5d2c51b6ce313170eb0181dce014bde2995a5a9aa09959c94141dfc6a24faff232bdc0926a82b940987b20c0b4d55c14c7151e0afbdd43807d6db81f290a743e354317ac331e19727963b6e42fdd685dbe7cd5891b8ddcd3c7ce095ebead80bb972bdec1b9e04af296571280cad1c182ad823099695b2f5be1250d5d7a2b5417a850dc0dd069dfc3698b50812326fc4e3536306b8307e6c4fb53080ab2d8c68cfa67d9ea991b383a6fd5eacfe0f2f4c43d5c1864d75c4d3a9f3f3d82042c3df7eeb990165c84c973df3bedb824362e498fd55af7158b5d42a67b90b12c1d97776a3636e1b5da8eb81bb98d83ccbd39ac39d4f11cd84fde3c05c0889b245efdce507976f8048038a4dc1d58419262594f848dec4e7b0abff2f9de326643a1c748f07708f633fdad47393c2cccba59f2e8517f0a0571ef9405ccf2580b22ecfb5a26edf9645ea22363ffdd345710a025e8d9c9de2888600c648c2b222a99081d20fbd06d29bbca3c534be2f56e603a9139f793959bce0bcd3e98824f3ec3a09e8a9750ff6fa682a7a0f27d43aed845ed6863b58fdf0a883d30805bc98ffd48c6e05957622c03d88eeb38d3c6fba5b6c313450aa1eec9e467716fcfe66d01eb63d0c9e09ddbf97331fee9abe0ad4f2819435ab70a44e2d18ba0ecc17188e377d46147893b7078653b75b575403e0b0e476924afa658a5fc48ec53bb9dd0e5cc98ced014c7ecd2e72e52333d82b5444eb6b0f413499e77f7313161df66b97635f39b4eb8e4236722eb723d62d3497c0c26a196d3264de75660422d61c4e45de55ab7f2ecbce7f0dd76511098bc1fed3b2bfaedee1dc73c889eb9d5c6a8415bc799f06e95249660500370af4aaa955a83c542335e1583018bc1e8f8e0a474dc076e1ca68192149dcb59ade23d340380bfcfd28f0aa8bd9fe3f693de2b327d3391c769ab614efdc422ab155551a9a7bf84d23e5b15e2f0d243a935d77ef3ef2f1f4e63dc896911d3666d2bdde99a0316d9dae35c5a5890bc35bf68ff94dcf73fb7048ed63d8a03a54fd86195183243032900d6bc7e2ac502a07f94c6966ce76fa251c509e5bfef0d6e583213287bfc8e71f29550b9389588a95b1ed974dc80b0f1d397ad4579c834a1285c374a7b4f7b7092680a44660967c8b59eb4340dd3ef690c06bfa77938bc0cc417d1363228960668e7269dea030f40a035a3e97205e4e2718d0813462add5b8e3c051986d2ca47023d079ad41a0a279a3835ca5d99498afce9e4fb8b900b280708b197b5c33e31b638610f6a8d83f01f889636a79d57dad32c32586ace6e344979a754d69d8d4233492c7a908843f3940ea6f5c1d511e4641d4c93762d288e24deb951370a5dca6b20bfdd0dfb2847a95ae417a4826bfa55efbc6d169b7f2ee1e2013e4bf6682230c4ebdb4c17f1f991d84349b4eaf227a5851ebc2faf0055ef5fc82c94f5d94f8964f3223e29518da0de726383a6b2373ea17f7068da3490d19e32dac8b4d22214b859cde894a539167d8d996d11b1f861a0520b8c18bf79f0b59352c0183d5982fd200cc77482566e8b9a0c824433824738cf2aeeb313e3de3f2c177d03fe5ea2954372143ae8c6b0fab72dd53f858272cb7f9f0a081355ef3dc82f575d0b2a4f332a0ae68e7d4f817a0cbbe7ca78b92d87849e5c7adc1b7bbe480c12c403b3240e2a66f3894d1848fcff6850a04aed7610a98bf2c667505d2eae4ea6cf82fd02d6504bb36a4d96f773b0e05407a0bb1b89a28e07f4e568898b0179589b6d51190f3a78d05c24c448b970fa424b9ac5375cb62a72bef660785f1691b95601283990daaeacfcb0fdc7e239455eca7a96aad8fc6fae8d1b6d44abef02495106c70f00e6caf856b438c6a962203eab72d3282ef8e4ee6171e296e8ca1845786af304bc59dce9f833101b6e7b98ae0db310901135c43f434b836e06d83789b0386b94cf7dcc20afdd4fae04e65350725a0a8109919f14787c6b0dfdc6053b7919841a645bb52f16e6b424e9ef46696471c109a00f7d71531d273c2a50e8956840ea1a13ff797ab8094a6a6c6c8565073171b4a40878b8a95d4ebbdfc6d73841a0aceebe47fa910879d788c07a46fb5b2e790a03cbbeb815f0f76182adcd46a21acc123db7778f4af25ea2bdb5126f405eed49fa1fddee559e4a944e921a212054ac1122be54d3d824ea7c423fc9c133c9d40e9a4f8c9544d3da28077ae3a50a346b83ecaf08bd2be8c899fca50110ab5e4f4e1df76b7d567a52a8a0c120f5e35c313391c54b1ecadbc858f49a7da60edf7487e31b49403ce5892cf13a5fa4cf80e8d4b3fef179576142d572c5d072c66afec0d27f57da1ce46d03822b163428fb82eb16bb8fa6cbd784a097eee20a356d3912df9892d3d5c2f591758c9b95785cc6ab7a5d66f31471506524370a8c93ebcfbedb9b6314e186a213fac6446ef167c2e42ba6a52caa160b768dec2281a8fef78b079e47b07520c346cd81862718d6f3868f5e75340852479c82b9daf98e670a856089f146b5eed86711f3f772e2c8517ba6fba446a51c6c9b32b3fe8e2f31b6fad141f1c9161423e1a86322d7e994766e4c889a81776eccc1f39b47cac9085a29ab01b1175a45cb666d4c9c994bb1079ac2d02f75b8695ec36235d01b0e165fd133ec8c240f0c12f91088f5a79e0ad16759790d62fd7fde80c2daa354152d7834b60161cbd999f687fe237897a9e0eed0c608df8be7b4a3d3c6eb882ee0d3cca206c8920e08431af8693dc1ee240ca723811450df6cbc0c03e826228cae05d917b5df15476bd45164ea4ef16d4eb877d3e2bc69519a1fe5074b8cfa8c35f7111782d1ebd9d9f004b19e93885050e528179d2bcfdd6e58941e702859ffbec372304e544d1ead20b4102c16c2d729d41cc099a2f072fdfdbc1737d280f8c306d0a250937bf8d82f891c8db564ee9b54c11c200d8a01e7837310be3111acda57250c722d3e1fa1ea07b37f264c4a677c8e489d5ac4fab0af356fe6b13e3869872c281df87a5f7ccf7afeac77cd993947bd976c000479689033952da2585726d5ddd3c9247e7637f7799d4d3320daf6fbae7dfa2a1e8a6c34e2074c63a75bb87990096663f36c9e9bd99b6c5f17bece820b0825b5a88299dbc68eb6f697166b833fca56b317c39c1b815a51ecc9a25b23472929e89848e736e11f8a9f4636c27ddb517b241466c2a569f586d99aab78bf950ab6363fbf7e32c40741c6496fcf8b459c48f5bba9d0d1813312ababd50e1dd03f825c8df618abaaa3a309d1e76a863b298293e5d3001d11e250449ecefd01b790a116426c16da4f62247865c977ee33caf502c7623551d6598b050accc0103f610c1bd5bec958b7cdc8c244fbdd785a819e842988527cb4591012491752238083e7613b924ead38261f23a774805ca862df345da9708b62982fb32490d216cda6d2bf9deb968e0b37c42661a3995cb4b888a753e5dfa44a7c073c36394f41932fc69ce426abb775b0179a1906389d7473dceba98b9dda4c35d16735063020940d1a3f44133e46bd496b7f7d251fec5cc0cdb8654f67bd5d038e588ded30238fdfa6df827d9d0eec4adaa2c0c4f4318f082caa3e7cfd2b7d0da3619a2e2ffefbd6b0051615b719726847fc9fdff4e4d1d93bd41f99437638787a202aac9730db785d3606be9b75aff356241e51534260a8c4435c99b4c3c0f5dea1c1a51122385c9a84aaa33f3af7baf4a48b2e413c1d42008653fba2751108d770ee71362133b70444fa41c3e5db913abe0accf1c4d18d800127e09127c349a1dd1050d08e809c14dccbe480a1bb642c2fc0ce8e9bbf2e3365397f9f200bca5d2e647f64939bbf621b953de441985760e0ca733f78abb88685ba616d930b2d9d413191ab88ba7cb58756131cee5693c7c98d7fad1354adc7e6dd4375b8f4654f910342c90373e7acef31236b714b695aa5aced111184701e25111da302560e6b571edd394e29ddf198f5ecf9c3d041059210c0caf5a77f76c61429505b3740703230831b898fc3c69bd88e7471cb7f52f33289eccc4114530d399b7255eeb7318de4b52f781ff00be65c068c1c8139f2c30785066b1c27d644fcf74cb2ba027e67e55843e742602e40b2291e8887a52e0c1518bef4857d6794f36c6678ff6d64dee442ef5cd40c5e28392a42dd4962fda6100e86a4c0e9ad5ca5f15ae851e2fd51c204e8ae91c1c69b7d6ed4eb2d54f820739f175d49208ab88478013bea7114cfc0a8cf2a2de10cef10c744719fdd2e6c39e69560d143fd4378c4f4910c840e60f174a6b1a5db6bf03dda4f4d8986113f99de81a6ef8ebb8fb8455c1901b0cab0d1bcc84a6d9eca1cecd0f9c25ad91aa4d25f8745e91c929cfd27586a47aed90571c011b04550281c771cdfa19388572e07ea65f7a37b13212d9feed4ce36db7ac064c8d3c9cbd2776119d22f17585bc9ed0a1611f7825a30b78657061de56f124fbcfba50f4935342e7dcb6e8f98b898f1ada35ce92b75387088c8c43a2fe349bb0ef5542552f8d194f16021cfe471e8d8a0d2649d6d3e8b6277f8bd37380367fc34a39060cb65c8f85546c5ebc6dff50c14c36d49c881b6e429a98169b4daaab008b7d08d37642714325cf0923b0ed444d7fba79645d316e45d592a4b1f5b1c207dc2a037596d8e34adb51bc7c8fa93d12e9fba521193f952126990e7c7fe8b2f0f47a19e9c5bfdead678bff566ea0a673693e59e2dcf1d342aa02f7a1751400f8eabcc89988d3772eebe926c7403912c9670efdeb65d92225594799b7dea2ade5c7fa39231138e29f537e3e92608642e71fdaeb4f8bf730abd9b3b084cd2d7482f4239efc5ac56729186b50c833f9eddfb2624c047b67f788b42c426394d5e58ebc6a12d6d1bf521a6865e4ba8a78eaa67ddbff07ea7ac953d8a0d3e41c588d243d6e86d421a88712ec0111357a066d38dd0f69ea64efa3e69bbca1e92262c3fece4fdc9075a39bf0e4dd9e1abc88991bc153913680b82218c1f3701b512cb776a7030ae9ff1f680bb9aa7081fd0c7c91c38320c27490d28480e955597a98291a6f7c9782aae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7b529589ccf10587fec791be8b58970e7eadee01632232253913870693f028c11148c1301fd6a8fd364f858fc230ada263faa1dc48e650d061b6884ac2f8626974f1ef6cecd74d3b28000eebd4ca8eafcaa50aebe2ab35f0f0b4c1db29cce4e284cbf38216f2c348ab739b542a271671875eed5f95193ad1d9d462f0cead8ad72115c5c1215ec4500da71081cebfbe134143f0187d54520c7d72065e17b09a0acd4ef2d94741776dd352be71a36b768cbfec504c54a7c961846f5839ca6a792687e591437e85995bda48ccb28c2b36e76fa8f2c9604c0ee34c29eebdf674afdc3b2e16bbb2015908e9111fa3036d6b395cc27ad9838e3e21dcad170a67c86588922898b2f251b0785571828ae57e5539570f0308b73aeeff9b69d170f376e7967f41830824c0144ebf1a8cab601789e5aa7c91c914660898ed485da638d1efad1c3fe47ca43fde410962a8f857085781e5581fac35454efbbdeb6f14e8ec57aa9a62d9720e92bdf0412fc5b21c66facd396922c1d34b7451b7d5cf0b3e7432dea0b456ffd856f3dfe9d39a98da1c7d7e1e45a13cecd23ac837894c4f669e35dec780f90d674d829f1d9514b8b16729a3b0378654d91465f424aeeeb4a1a09ec6d87d26b91cf7f314190282cde5a10478c868d4dfaa01c3b61cda6adf5bd6900177fcdb8cf5322fdc493eb4d1110d72db762fd7edda89d3580048cb1e8ee8858b45127976320accb8b5d97e39d035ce918274643243ddd5cecd9c33ec26ef0a31757d22cf650fb596503d73ad37fbe73b217e9ce2099355665d6028440137fa7442ad9c24d383ad430fd058fecf6e7df4c779edb2f0002d9e9f29903696c82b68023db10548bed388c26d7395d7e282a9437cd992a3bf4be342646af0c79cde899604a8596a80c0fba09370c0747f25bcf083cc0c90bbad989306f395cb7907b4199baa9c4b50f288aab62c47ca6090bd3b500e2b9ebc5891afc40958e746a2a666b8a797e03854e2042eec28d415eb74a9416e2d0f906b5f62ed32ca24a9a50da45a24d33329f909d58937f5877c39d4cb136015dcdccad0cebb67fa377a357ba7560837f117796619069dd1b4821665fad59635e90d335208142dbcc8b9f2dbe63ddbb22ed7bdc2f3bbdde98c5e8013b92a6d8021e8d05c4b93f4445f71be7235c64199b39a82f5e254e73e23d04854532328aa48366c01db41e4f8a35ce08f80851c79cc18466454e6872d0ee63cc6fd6be84a79bbee09f2650658e3063940c707cba6b6f2073b13985fd0db75c4eba493f345584e93bdbb705506e8612c5d44d566dddc6b5cd13e7f51fd0a5ab1284209a4a7c65affcb1a0898ba0dc88acd54fbf7e1cbf816a8c5132b43a509ddb5279ad2c96f58c11a3d7dbdd392b989ba6e576a289a0c114ed6127b47181dd0ab63c664c505e64ade6d1de122bff51e068018b647bbfc6711f37561ef38df3709a8ea93bde050b2ff4a1f43de8a8c79ec3199785a224a9d13b259dfa61401d341af3f4f39e983e02a1562ceffcef6b73394a03b1bf4f479a11767b9ee1a78390e395b762a62828a251bbc75c9e8b530ee6d09c5c2d50682d80ecbe870c5ed15e742ed2ac34276d1388ac848a3c5b81ad1c836aef8b7ca19e61f1260e477f281e99b42836f22bc72ad7c44572f472b8a3ba15303a7724243348efae49ca582cfd7959b604930c69dfed4132dd3bc5e0ed8c6d810487869b79f7c8d55a9575ca64e9339a165f384648147f295a6b4f3f0224801a2746925be9acabfe4b810242760543d3d038d36d40ecbb1183a0ff65a19bef2e6f4ffa2fc7a9c231be6af2ea402d350270f0c95cf22dfb304eafff659e5f96a3428931a6ed6b2df486788d763a44b33a38d76d90890cb08666ff999e57392eae897b96d6fe1206e41a7e42ad70893d359ba8d52c67236f6574574c2df4a2ad090365e1fd1c681afc676ac2021c4a2bf032c25d09bef5f6c91471706fd6ffd91b4f2efdbb3650235d9faac765dfcd90ea3cece9ed8987a34c8fdb8001f42180a9aa3d170d8549063e598163c879d9e467b795d2266fe134566f6ac4b6287ec0fe85a873cf8990f8137f32587b7922a523a3475acc65be320d698d634adf8c6bc874b898eeee4dab3d354b327c93b91d6f30738191501d7bd9ca4258c9a85f941cda7c84285dac8dbb37a99e75e97c79b5e5950e7dcfe4db8cd2e5de27c670fe6216ae10a1ecb09be6f190aa98bddf502b14b293de7b423b50ae059990e0e54874059b016e35916793358c4bc1c15b00c284573d604f4fe0264b722249b95b2be70ba82c7ce44ced57efc0612b4b097998a8c3707831eb2e7d01e56ba3cfd10bc5d255cdfa514a2769c955b58409b34c425a46046cc40037e613eee3f868220914c0561bda16217430e292be669d365cf1d0523dbd80647446b898ed307468efd60df510057dbb12e463082823d3eb5eb7d1407005ab385bd8e8675a50090d4cf35c44517b767eafae0db85def1b15b75379f3f34368108e40ca4c2e3c77935e5d473a659a8a5eca001000c1f6bd451715a8faab9300989a5f720415da28fd2ade16d8c5e8ce94f950854601f6339771c5a72216193f17ec7f8f2ac761f4826024821102efb283b2c509d11ea930c699bda4cc25f724bc96f2f5147201ec75a2c1f4b15e387374a27816a6474cef091766c84f24bbfa801459c3c7e112a50f137f4e121a3068ee8c57b64c3d6cde64bf9b4cd96c489f66ebe0f3b262dbb5e5da956eda7731a614c58c52b1e4331d37e35913b39290663e58dbfdbec420db383fee207339a01d7bd34f908625e797a0e8ae4c9ee1671f488e66c291a4a1e0b28dcfba4c54223c15ef91a5948d4f42fab5ebf8ea63d2b2a51b336ce86a3b132ed353cea2960746b7bc1085f16947fa8968d4009e79542baf096b4330bd770b47a2ed618977cb62069460176dda6f0ac3502b0795a0c28eec56fd4d4968140ed6c4d0f7d57e6e0ad5ffc6967b0221dd1285abd14346a8db446675132091ca8888205f828c5c2320a9fbde287e5fdc6e82ae94a576705a542275582684d97b664e16d3251591cde3d25a6ccf561272e5e876eceef4660a5e502d17b01389adeb4f6aece9b9de4d0c496b1d6ef54379966f062bf5b3a5ec18e7dc1c5a39beb08a86781038777c0fd79c058e14a379eccd47c03611f16bb6fbcb5d48923804d9762936a76a8e65c3c9a25e4fede88d3445b21c6af6ec2903979856479d67fa560452a53743578309968c9ce01c20e15fed4f88d01f40a7857830b0ae2889a0ded74451dc384e32e6767e4e25dbac027f3353c4614f5ea2b41bbadbd6ebf370e7044b0e2cc1a337658db887fbde57dec65632b1e422a0e30f894287099aa2bfb6576aa60c04eb002743c5cc475cc3e649e9afbc3b88700e59b20dcf458caae183ed6f047b83e6b767a361d5d93af86081bae0193e830dc23d08c8104236162737a773313d8275000271e3b59a7f5848338b2179cf02084af6d854124993d381774c035586d70e2152dd467f0e46a80d4e779b66a169060eab7baa78056df6e5c2e2fc8d5ce7c0f192dd6918553dfc4d8490c160977ee2a39936cc27112ae88760c5355c88d2353c0682c10be870d0d88185c8a1eb8c8b25860f3fa684f2d3f137cefba599b1627d5562a2e8ddf9987a1280e6ef6b98331dadda0d8dbb42bc8bf615bcf4c58d3893d93493795d5ae4f3de640626a8bd199505f41a5b422c106e3063d3d85a3656f3cd1115d874d021e7e2b7fee9144d3bfbb8d00a6b1cd3bb3311898f6db423b7f938c3c0373e5d8435b371613dbe497ba509049c12ba35f08ee9362a98c458350a99e2f1d7f142b9105997fd614e1f8035a993dceaa5f9f0b48eb88b673cfa8a61841bc92eb5798010320b5c2464087d4de0c382977b81deb9f46ab957644ff402db4dd0b8ba30d12d92884e671f971e797560743bcb65bc62f194cd2fcb0f4894a6440432d0578d4d0416eaf0075eeaf92b80c1885f3ac275bb3d028e01d1ad2eba8dd9b5ee9c0bb635c35dfbd6f793735440649623883ecdb4281c26e6e2b63c1c9b41ba08c97c000e379e6c9c73cce4d7e7b054eb901bfa34591b2e7923173526a22a2fb3a820d97ca6f47b5b6d57263f1d218ebea1e09cb5fbb776c8f06abf9a1bb63715c1ff2092d6e7a8249c8c4f7ce6d3d1ea7141e84c64d7fb8fe492d68e2d127a3e9e09189ea606aefcdf17ff883c0a39c946bc9b93fdbe379c3a3ef485821b9cdfc3968f7fbf4ee557337987ffc98c857bc019ae5dfbd8d7f7aa48ddd7ccda8c8bae50194f1268ee3f08f91d3a2611627b3ddf6382176b5a69ffdd9e70c0dbd3394b2e70228f242e447df55077ba4b432ba5bf2cb8fd0201474af0ec359b1180343275ac9eb76289433c01fcbbf3594e8db7eaff1f31121a4e0b2b78ccdb65d29b98c8601a4e677bc89375802cfa9b4c28508a42b0882bbb546d16a103eb5747016ded31016ea3ae37ba699a6ef90e1db5214398babe5e1564301dc709ccaf28e17bdc30f7f018726e2952ae660a25387bcbc5ad6754455fc89ac67554945021f61dfe7304c49ba790ec549984e9ba2367bc46db6dfb26d6711a77604c30315a810a3190c24d8337ca6bf8047bdf8314ef1d97982ecdcc681d423937234b38239ca36cc3da66ceede2c287f9dee1053d8a1ce7b7dada171ec7a130ef1d28dafd45ff5604523b52fefee1e2b96e870c7d0ac0f669d5a9b3979e58c533e79ed75d1ff227d476ce0f01087de73fcfa0887571c94ec31aee56485e29af925cf78464aa4edcbd7b994a42d824978fef5e5271b81bc8492ea88f4637c7631e7cc6e76f2cdc7d1482720845ea57d51552e705be6b3381b8ac4314dffa38715a18ccd5031be77d9c6dda3fe52f21ec469708fa08a264db59452d622d0e61dc7ccb093be60fb9bd249244103daeef3a47ca08b755e560b2649eea4c3f3b6c73a747ee54a1f80c0bfdc6b535e088ac8bce80a73a61822f0b62a52f5e82cbf6540ea1c1b7f94c717d96a4371060fe1f4a6f73691feadb22e94c6000cd15f00386a22d796530c77c3ef65f8811b39b1701ab995d3e86b77c093c4cfc59e77c18fbae87ce6adb61d116158cc007e66f28e7e4615d5e1c65251ddca61109ec03e4da1d4eb0ad34e9f54d7716020838554c3e856af84bac9fd1edbcddc1e0edabc9f52a44e2464d627458d560191bac3047325eab2ee10250ab43c368c4394f01b32988f926b1005d0651f2e3903428f58b02c6525596d793aa1f099a37208a3f0d51da321d22364ea62fd2acf43875f12456a7777c568e95acae7f67f503049944db8a24f1dc470c2f73d0940510a77ac612225ba7e86e2b39cbf23ba7b09d4204116087882d16f40dfdc679a3fe634e60f43e55830b4a993ab6b15796b18df3b6e2973841383ece453eee3144786051f299d90e90f9443743871ef8c205f2bec65ed0b24c2275a6e5063ae1bb5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hed18579f8ccc1f003d9f5f735298aca3a48ab751d065f15dde59649d65aaeb4edee3c78c329c5a1c5d801741a7a554d4ff2ddb0df0238bec735319d12af76f74e2552b28fbe5844b2799154ec48b35323337a3c44d1ad9d8104ee576b39f8c843bb24c66829044496f2af7cca1f7ce29063f3be677b06bca657e0b41a542a38d302c887170ed6ecc1e67d6fd0c5cfa338004cc14548ba6593593cb3ab38dd0c35e214020c0daabbd5bcd6f1491e721b6cc0efd8f23862a3b72bd285de6d1344be561d0d0f52244477f0182f4ea8c4b2b43c60eed7f93aa09b9d197825dc79e680cdfc57b12113377ed534411dee47004f618786cade0ce80262d881931b360480cb6e620f0dc73a343d997a66d25efca6e38263340f78fe00738de2a1359dd825b8fac58f8b96c06b3e19c7f8343167c69db33fc10895297fc0c48b900b4b2fb3ef29dc825b984c6ce46487c9aaea3922a433610747dac565f475b84879ab671e495b5f5c0554d6de5f6b475b3ee33e96fc0945006affa80e5b4f849b7116f4d76d95a853fb64a9bb8f7a74b78487e9852d24148b8a06c35d7df03ad4c132cf8487dc0ef79df8d5befde2e04f1026a16b81a1d79b415d05409c4b39ddf5558c9cbb950cc57f4bff7e7e6f7438e8170dc373f17ccfbc30e8b2fdb8c30223e7b55045065f3dae1589d1e49661e4394b82668d79f7d026df78c27812b135a294688bf2276d9421549420b3ce618bc28bbc71c6dabaca7e9fce22228461cb14608861fe15c489967908991b064b5ce7f12aa0c921f54fa8dd403deaee6c359c7279deef877894833407ba2e5dba3fe5fd9f259fb6db0571992373a511914d881f7855be29f2f957cb1a3e3ab07130c63e07f24bed3cf997a5c19526e3567b5bdc3f6d3e123de6f77ca67efeb176885ebed6f9d530f318fa0712983fec92f849d6196e11e66c4d46c25e7b71b0aba399361d611e67af3c4ec152470b918bf2e811afd03e7692c225644523364f358bea5a875e55747875db4d1d6cca52c46f7f0e32f1fa3d335bc2c04562860dc73905569fc3e3b3c9ff8b4432283cfa4b835fa850743cc38c25d6decda5f909be4b9eb1b1ee2f61072eb29d573efe4e95a98860d033a1bc0c6ec24756089bf24e00608fc922e0edf8fceef7df2a1011e7ffc62c14230a216f88c09078494bc18389905a2809eef287f0910e5489f70c1c193a64bc7cb846f6c84370848a9c584e6c784709365c286926f9dd6608cb1b7d55f427fc5c3091a6676939a04c1aca2fa9b4e4260c9d98b90c7e37c18b677692f0a5aac785ec9c1c9add9afadd67c258d025cf89f6107ac2c830b96606579d905a27a21f0ef8bad13c6bb9841feec0df8beae9e6a5fc7b27d71f11ef55294cadfaa2ddea1d15b6378d0fe360a90b93919ebd3daf3c749b039e055813abe9cc42cf586c591d31aabc8c2a13bbbfa89d748602b56284e1a8040fd0ed89e5d697559c4e2e1189f0da51013852532e9aade57cd27cd2fad1d4d5d426f1363024ee3b5c5673f56c7c89b184499644d9e943e5dcb755250437d1d7bfad9941cd482504b6fa8d506117785688cdcef75a5c682dd6fe1154734ca10f75d384229537b5fc28547e737789da95f85ae26e2969269c60ac3bee7ce2caa3539e20c8fac3e2c1c32fa5277c54bc3685a60733ab27de245f6b01bf25fad7eae4f64d8635a8ff894fba63920199da75f20d23e3a31df5371722db2e0af81216966eebaa660c328b729eace24e929cebfc3e85e7035e56073e8e95a38072b599437330c8030e3510d99a227fd106add3ece8451127e529e75f3a42a21072353055007c29bf06af85593f1572c49300fa4425879be095633f339a713b392668eedf6329a3f357f06b9e9ac0a5ec02141a926c67b11e00167934371c30ff52caf8801384cf2c1f382e78f18d43f5562fe11df6c177bdd756d73d3456536fe2e2e7a077f2f6cdd5072d70a850c6325b1ee011726a8c679df4330c167244aa0d37156b6d9d92f518af14da01f66587459cbda9f2bd775394b28c7b0321592237156f0d44e06281b85f594d0355837551004b5f506bc3ddf499d6b131c0bc70b6f76197d4bc63bc4460b7e4a15262bae7840ef2d21dca1f937e1a6812603308cf649241d12524680522947c04fc0c3818fcfd74b5cc4d0079e2608a5486c40363899b2e376d02c87d0e29a7a263bbde965ac81fdefe0997e2feec269f8a12b9d0772930bfe40eda1b37fd3481caeed2de7bc4c7fd3af368b4469c943c9eb95e02ba9b20d727d58920544b9aca50acf9c07df4eef62545d954893b425e61241dd6261caa7cb41e34792824f43c682fb38c788f5190866ab48e643af7b566463dc40b3158269032e63e6c17758e6b7fc22bafc65c4f9aaa219871fff36e4818917933507efdd39ae225a6899cf6734e63469a2dae326ff5815d0b6ec6b39f0f6eb849768642cc3f5cc902e5834f0c0a2619948253c23e7a386a17a697e0b9d740367b1ccc29a14077015f17b1a0711fa53aa68ba3b54ef36fb0d483d5f1948e12d1f94990313793f1dd2e9640ab948beaa19db207f08acdb13407504ea62f0845cad8bc8bbec7317071425d14802b7fdc5e27fe253f82a56a9269b3c82762c586b450e84417ec364f39b27bc55b45647019d998dcd54e12d7e3a46572bce4a20d7966cde0e46313403c4a236442c06b66c80e79ae74c5fe06409166277ef7592474bc1463d8b59975ccac1c0588f068f3591efedd609875dc47142a1d5f3353e50c92618c8e0dfb3b7e6f8ffb6b5747b996c11cfe520d28dc65d1e2a3ef392beb3f8f5d54ff87f6ef0f687f5b964751095fe16b8948a6f8452d068a16413962bdba318122118f6fb5dbcb4deb3b46ec65a6bba681215480878ef6993515c5025446ddaa26277c168b41dc51a760a4a707ffa7585302f31f905d3a85ee63c6ef413ad511e9b1ea39d1416785e9e4bcad9a863cb6a77f26617f48079ef08d169670a3f65368b39833adccee7c1f0eecdddc90f4383411509e70e56b96b0bdd18be6577cb8ce95cfb38aa474cd648eabb5a0fd6703872e4904fb0e612b54317100baa2bcfa1c165eb762f094a9ad03310a5ba7cf758be5329be4a2904653b888c005659e9018ef55f12fa13c32cfb1c3e7d8d06aba8a17036d2c8b7773226f8a52b9356edcd204c1d6200b64100c812f080085a660a86dd331b02a096643863c382ef831317a1a52811ff7f32162752dc8aa5dbacf693d73bf8f3a0e085b10340d5371ad74e41cc517e407514701c161f03c98ee00d32b2d56014a0ebaa5d79e5cca5d55fae541b741ece9b187c050ecc6b8b85bfb974abff562497380c1c99ee44fbc3a5f10252ee501e590309d03400878f65e7e4d0b451895a8d0087cce12ec6803a9267ea8f784b5f61016bebd4a17fb8e511320014b647c319e2667ac39d91ef1d5a9445ae44d2a4111b2c794f565b5fa9e4e2be0ebeb21b7c10421ff16d112211ddf60a7dd818ca67467645050807270830fa86aceac2f969f4b5e75c416cc861ccf49f1558e4e838aff010622c606df26fc30fe16d7f969f3dead320248b55b0c64626fbba6a7a2c3b9f989b1adef50e39befaf3c06c3e31d1586da60e2f4dd79815015196f4fc9e769c2b7f46c50362abc7e936399eb25c6ca86eff870ce779c30f3cc5d738d583231da9a485caba0f5d60df3a633df8b9ab60f978f7b54bd7bab64232b5046765d371c723a854c2dcb986eefa54802efbaf6c121186824a9d32c7e0c4a2820e4ca89d341efd9f78b3bfe8508ae19fc12d191f047a336c01f0b1cc97d91d0c53a2608265fffb99e1845e0d66a46f6c98ea1ef98944ce5a57ba306f273afd6ae4703b113e0384a6ee0cdec456465eccf3b028df9353f1ae0a29d9d627745c4295128058491c299e349492ff0af64d4682578aa3eeabc7be8636a4057f1b4fbd07046972cbb3b240d4e59afa07e6238b0816b06afb8a764df6176dee1f077a6c5fe49851719f17c30bca6abe04283a10ca3f76d2a05185ff61d3b479df240075133c890c3c83b4446da00f1e854f1519ba16451c833e4416fda4f18333afa31ca0670dbec608e644e8a9738987e905fb71fe171f2e952422082deb6a5619db1ec1465ace0bd67304d3ab6fea48bf142395e0e6a598d26452cbb6d59ac7be7e301141c42a91e92de898ba0907dbb613121f0afe51abfbb7ea780127668047c7e9258fb17b5e6bec8dcbab71b3658473fdaac148e6902e6ac8cd60e4f0a7189f0636ff2828dfd8d9aa3eb645c776697bcc91f5c0fd2d97c26306cb26104510a16cddddd05c941a10e922fb174674eebaddca9ee321072f9c993d5035476c9a11e75a666084fc40a35f0fa19f22fb3bf3aa3713e9acce25347ba79a12132378ff3bc855d2f9fca5c85276d8143b771a1592e84bbcf72589a15202a472884c544df0271992b77e0c653c128ca4ff7d57dc9a46fce8249b52a107caee5d7dcd33886bbafd3826df1fa0a3d4c6175d70bd1e253b3521058fe0ad115e029ae993074c87092700b17da882b3f9d1ed782bca6f943f3e92589755fc621619b991d15e3c81e1a7e0b74a11d7185bd90aed5e709b66f4610eccf3c8477427d32e039e436d7cd3d98a9d3c5998e527b31d6aa582f24db53f8cf0b2013967f3e1f6eadad61cfa96851f3666bc73ed2762f3d5c1d996253a50677cd221ea3ca14eee5f2af0a5d03ee40d671372223932f16c1cdc0a727d401b401efe573726c67a62a2511787627a544843236183cd84066b7c0f11bf9104bb3768f5f32811e4346092aea28ced8f98c4001580de2f52f41ccdb47a4ce23489ad9b270aba63ba48857059b5988bc5f0b959e8ab3ec32230aaebdfaeee089062093ddcc1587c13fcb22abac63434a82e617f42f246469b69f95457d8d8533f7e4a5f922a393534c9f40b550ed5a15ecc0b013f0d020d94b0f231511892ea8674a32e09356e18bc3a7527c62a2b2128cb5489b32d3868b20472f2ad21e9b678e228f863cfcc78a5c94ab947f900aa6516e82123f9ec3dc90049d3bee0ad6888603681e7fafda5a793f2bf8ee83520421d0c75c382365569d3670457682e794e8143bcdd51011a1b07e46aa6ef548aaa88e0ac415a9f51a4c381505dea4c47eae6d8acd855e28d60eb22b02f657c08fc12d0500bbceaffe7dfe9cb3d9618e43d8c38e8ae972938af85d5622f549b7e131e80cbcb174d92c308a0ac8c0c4ff46a2efeb9c4864fece6b8a68601bb90b69f5c7a97852627a3b562ed7c7c20c550633fb6d7874a9abdc43ad50c12dde4b08a30c53f76b544790ca0f70b2e307410c6e96d899c04abc9b3c9885bdd443109daad24c6d28c63253a991ed8e09e2bb40a5bb072979bbafbd75231e19df106bf5aabb56c7840f76b35eaa1196a7f0e485926aaa6a559294a74b4ec6d69188a3bdb372635d00349348bfb8243eee2dd95c52ea3173f94cea8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc9f7a75387204b2e964bbd90383527bc571163fd354c244193a67689477d8579bc109a39df80c737293aef692e4aa09bf63e66e502e20b6e71fdc2dd124e7e5dc54b08bc6df5c5f9c985d410144cc5d96957c4668246031a30975f40d2edea6acabe6c474c1fd72ccd89017ae45708924cbe241d60e20b894019666d63954e97ede9339722331bbc60c27e0dd79f677bca51daa6189f9e1e5402e5a94c24ad7b74bb542be477011245247cae72d6ed72c7b567f2608e3fc46025129cc69baa4082ac8f133df32931e5573ce8db852a6d55e31601675c3ef29594a49916d96859984da9a891071a562e54a571c2920400644d4ddba2b05c751fe0843d0e491d2547c1de86f2d2a8d5a032960930a6962ccb61d7e911edab067efc1aa95e88b0dbbb3caefd30c63a11173c89c33e19216ad57d270fa53ac21d1fcc8f7acccb8cd7d7b288bcf62a33715336816da03a6e53345c8ed1fe3d457bc32d9b6abb137715844a55408b2b3b9db571fc92bd09923b2929b6207d482576ee5c1e51129111fc3f57b10834de9ddebcda35bd4c9717ae6d45d5ece49497ce43f65071cd9ea8065ba479b7446fabe8bdf655a7a0e5d7754a32871ec852fe4ecfad19d5fc8396e4224663f0eb161db48101a5e97afadad8f3024c53e478b7391e169237150eadd07e8f82bf4b7b5e7fcaf39302288af0040ff29393da4766d689d2b7b8e4e06d0f458f1e9c50abfd98fcd93d43ee930214a812086d7faa3d68de962243cf7b03e9b04f18370b9e6fe7a9fb73430aa3cd69e7ba9a848b4e047e2bb933a5b70be363a5df5fd360e6457db8207d34ff6352fbc80ca9912bd8925a895e1664eb21184e0ba363ee5edb3df338130d8c42a0896a1c8da693b997587bc9184e241b4376b967f5025f4bdeeff2334e6e15098e2b19540082b5c098842d0d396a16a175b3923aa20744828dd0803f8528680e9fa6a03a0e7743d280413b086ed463718d863469345164de96f7ae3f30478fbe8e0942edc4a863d9e47604c9ee0d2ae209c4f1d985b950a19578ec2580ab3638e4216a03dac22c0045670ffbad2164d6e0b3f952a1f09d39c342cc826e1e115d1d52546890895198b5d7472f0fcfed4b0977686689c810970395e1fcc9e7bde48e606b04415199d41de218d34df679a4abd443360437fd9655871763d5824f030852f6d562d511c28eb9abbe0187ff5312e03589ffa867fee330fb506f0831b878d72e100728a7ec0ebbedccae97bf73792bce2b5fbb7ecbf441b06a3bfce1687e0ee89f4375028aedf00f1e04a00ef9d7422e9c54aab6711a04e6c2466fe0023ac3a0fcdac15eef55a65f52a7406bdcf245765f34d6bf5c3d50eaf2f3b8a7d5002f00552819e0595adbb0e06c2e815c32fce480073d98d52ced05f6a51a0f1626cfba2099a77d238861f57629cfe83e54d8209d4d181d023c28cc4c73b74cbdfcd2741b09ecb484752c15b5d9efd3ab520cb126be302577e0aa3ee629391eab352c2d1ac289f05207620359ba26bca1e56000f13ba28c8025eae9665af02549a210699ed5c52013ab82d5ffef77bcb99858477f49b59d960a68fae6d48bedc1b3bf2989ff9f35b172446d3ba8fad480f70474d754dc2b8d574453e240e449d90c9434eabf6f2310fe875f70bedad690715879eb9536a6767952b25b2206d882489f41c5f317682f409fae655b0dd05fee428a9ffae85bceafef864167c8e8d65a1d38db33fa65af4cc950c02dd8e9df226553d6f04839c4ce1a8d1fc4a7860051ecae1670e09007f2fe1360d3022da87d23fcce40137cddc413e993dbe70c38ded4a0b97da026ddf919e79ab1d66b1420378c83b3a1150f939b722a12c0dc4c51a290494f7f6a145b5448dd30bf32098f0c00c895b62d3ea681895dd16a805e348a22367c8909d1a3c59f17ffbb7d8fbb8f6d5a22f53d029f52f9220b68ba1b89bc5ca255b117afa9cc4f8522b5bdabd18c893e7f1b991aa7cf2cc21cc67139ec742bb5163916a8ba518cb0a950ac20b2c97d4c6be8e8535c00fec1b98cfe0baceb37e1a5ed61e2a0afa9fb97f8c1768e8159318f16ffc1f636440c42311c4e88ef268ac19bab750be209063a0eb811981575d668c440e1f7b97b875f11849d910e5c6a20b662f576a951d4422ac5d736542340f866b9dfef9103be0c7678c6d2161695f6048c9e88ec74ab374183b862c1a1ea99a718af1c79aa0fe8471f7c508ed15c84416f6cb30dbc45284133b2fcc9b0c340a4d6ff4f0ea2e05a54956ca3f2fc7f03faa3228d729191f0a80e34b44cdc05bb6dfa766ab84da55157968a5bff04c0a423d3d726148ddc2d294dd4d5bb4ec3733fdc46795e1356acd22b87860257f1f8f40ff50deb395d9ae51a9ac1bf53f25f29bf2f0dd861944c5296be30e7faf3e527a4e55ec5e890debc43beab5668edd67a780800b0b15f2a4fee84615ca1f2f627fc99c95e953df2237693b3363e82fe3613e9095a7d0de2e6206763cedf999e47ebfa95d989839d6c9355266e39b0c46ac7ac77d5734f4b6c301d785e579e6127a3bef0bff9b44337ef12cb4810822316f5bbd7c9caa217f42dd10e5962f331245c9eb54d0f7e55ac47607c9a89d0e08827b9ee85e7367159c0817cd737348f555a0e9d45d9feee13dc8942be6425f12ab9b62981336bd8061a93deaff903a92df4a145b9b231abafa18a1911b760cc333b09abc062c6c9d968588c9f1cad8c3a9c18f6a2abb358cbf70a979ec236c4e68e930fd273429d9205172a1ad7a855eb2988e9ae116f61fa323b244980125bde9c4c6dfc44a6bbcf93dfb9361babe0d24e6a108996c7bf7c0e45d791d8a8ce45d708855a5c22ba70a4fcbdb66cd2e765cfce4cfe59436f69058a2f71b79f66c0ec8487c51982e762f68073f8d6a1f295fcc5c9c3217ed3cce25ad70ef3fcd3c0f9429d61c513a6f85d699a23ef0f5b2a2d1a12ce44ca2e3f6023f0f18a357657b0f447fef8e6265c8e6823632c03a3e37480f0f629a83d7202377d410bbf6c5999b762229034b981bfced7fb62c29938645a154fd710efa358e97c61de15d7c28bcc2d60c912747cc070ddd79207054df8cae773b55c0905b46ad239d7345d4bdce176545fd433897c61c1cd49ac53968a36903cc70e1a25de61e405cfc8bf59ec67edf57f250ed59a1c55ac0e52f3cefa02012bf55942cead07a6f269ef3700924465d805570ad0feed4f2d6f448f8ac6dd678af081bce4ee92b945a8224f8d90b08640722e79ffee044a353b4b3c66c7b427ce28ffe39fa2cf76084ed4de8306feaf7a65822da69333ec692979c482c46fa54a7bcea200f70ded8baad0aab2a9a8fa0c69a130854da42393138223250cd31b8ffc379962b43358927745c4cc1767ad8d4a64a8b12ccd1300f83cf704a22e837e0953548c56c61bdb05706ec5cbd1b955d1a11da02ab11c11b9891a6ab3f30ec2063388782b47160a0148d979fa3d5bd29fce919336c03a2bfa9bf74d42d871bcfa3b9196b36838232e2f01283a5aa95254609e5dc9fc792ac9f2d544560578545fa6f5ed13254515644b2e34b53562d5836171acca75a86f2a7bbd2ba78443d01fd29f988ce0e8d566c552dc1b0bbb25d3d015c824d67005ab38f46098075edf1395d44788024c11367b6cb8ba0adc3f28a04d8ed9cc27f1075143553c9502b1106218bdd1fe1d36cae5e0eae70a290672b8e6d45824362531f6162e718e4e46ccae2db447353f909623c1ad6e5171a08530091fa9fba660a4508bc76822c1795a9a721336b6122ce50ae2309a20ab8d2ef1f9bdfb4169c1f91ac615764dce69e9d2cdb8dd5c058f6f5b3dc9f4983e99379bdc5ed0f394dce7305f95d8a12ec15f521dfa5b5c7e4c9c1f17ed9e9b2cbd01fcdf1ddc806142b0f5782231b95480215b5af2174a1c0c455d3a07a7e1ea7a1fa30d5585dee2187b1401ddffd1655e029d2cb962f0cbedced8c68307a1e5062c60857e5f0a2179321c0ef8e14f598869398d5f2fd58c8fa0644d3aa52ae2f7fab98100213e016d9230ab92a94c3e4b32d9c339b527688bcf4ee5dd0bdad72f82bad2ed3fab236b3bcc787f3a8272e93a1bc41d027d461b77cb5b57c3329db8bce56b862d9c5c02678bcce0d6408a210d7a46e5e28b7866d091d06328b06e9ea7896a379266c0d20293d26d5158ec12f04ed5a9e387cdafa4277c638a839954c3d411d83052706ab88a13081575d50f75ebfe5defc29b93ebd838cf5e36d3ce093562b5b5397df0ae7ac3dcd1b20a649d10433edf28cf4942c1ec2b783118cbac625f09cfd8fbba8ca866e37bc6a83dcf613bc895d7186295b8e53d065c16df799bb510d4310e7b52f6f5fe4222e7d352c6cb268a23ddc119413d36904f78df446c5384bb3d9eb64955420d625d465b7608acc38e517a6c5ee215716d730a3df14632a5e4ee5fa01d73a27e82bfaae8806f96ec2359ceecb3dfeb92a1d0c0cf830355902986d830ba296dd061a7bb6e7d768b208b0c245c6144f550fe6c6dedea57b8305a81c485a4b9e17db98c1b948b0e3137ee1299e17280473665c8a8459c9085b4998dca9b30af42e16d46aab32f0eefa2aba67ec60b91ff64640b4040a2fdf5ba228aa0a5055414fc137aabda20cae3def54cd583aee316752e16ed1e49c84aeb79323a959961d126d140d308901cfb8425c30efec8fff50ffa302272204a29b7e5155dfb6156e58a7020e6bb2b057c0b0d86a20096cc50a58a6087ec2dca087b19501469a99b8db252b5ac621e35d10d02a72f580a9548b13f3bbcc83a13857363a5b3061eb5d2ce7408a63349b4c47cc4f9977d61a5b17a9e0b003a660f05792ac2c150defa3d0f37e25effb97fc7224f85aa575e078bc5c9345d685ca27ae7516b7cc271b5563100fc29e8cdd7f1db75bd6511f6182fbcabf782f3f806262af8e2ec097c43f16c504c0a595783d0b5abfa37a36fabfb8214e758fadbaee156ff577f0b6f27c5769f1948ff78dd8e5e7f46792c22cb5025a150bc55420d83c7f5295113464881c3b11890d3ac0e991fafaa74c4e041e826d60e34d74e779901b43468f16a7492f6005f6d6ebcf98e893501c44e69b3901e792ee1050e1013f2b32220c577de6d291248ab53b40746cfddbb3e7c2621ae5cf5899f96e1381e4d452f6d39dde915890c740a0aa6a86f7ab9f0c3fe3673b282c3dcd635078ee17fc85a01ca44b7fba359d5f370a2ea554b6a5e477b12205b25e6627aa5d6ca2cf0cd96a6bf40b88546a380b54579eb9aef600629392e09823c1976b42df40bb0ccdfcca14732d70db7f27232d4bb04cb3bdc3e30738c3032fccfdfcca30c0a3f33cdad356bf8d27ab63ace0b4b8947849f1a1ea06e28efb879fecefb7e49d5dfc24e6b5f935b21d3075d31d03f80095d1da2e466f43fceacf9670f74afdf29bad24b7ac2e29cbfd27136de0e42bf156b8eb651949564a9ef820d664db3306e805c5fb10e3ed9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hdb45ba6eb2ab10eb6110111f79f7ea4ccd5c49d078ad0cd510c1e1bc68c5c0ee8f59e07525fc9db077abc01bf99980530559c5393a49be9db6fa75a80c2a0fd2693b8879c7f8d05bc405e28f6f8321130516e8d0bac9d522492d3cc71c9ccc6ead096c6530f55ad3f0ffd80bdd15e80f700785e597c05041454ea56e7a1ae2296e0138fb11e36c023d6b3136edee0cef5c217c4a8137a1039246d717221401eea0324db1576b2650c7628a1aeafcd95d9f651e620eb4a92aeff1340da27dad98f511c8c64340ce0cdb5a50308cbb8ba881cf5d1a4e26bc1a10c5689bf808993d5a5f9abc456179cbe1dcb997b9972bf64cf3269d2393ed6fcccddcaec6b0ac4c434e126f56066d409abd4c2aa13f211e01669d5bdc1894bcfb88f5d09574839a9caafd6c1926778705cd6c3abd2a6760a91e093601e9b2390e6e8e31300b005d5702e63ab9323acbe030bf15d485e6033f26bffbe746494c25512acefc2b3ad723f471074e75f37707a62184c5d5d5584dfea87e5963e70b19b00e6c4e3d8094794e776dc441a624988d542a0500bd61c5b8b965098f6bb8e34f75eefcdc530e112a27760500df1916c07f32109c7165904803f63828ae5b8432641db365b4f4f49047336b284926d6b3e60ad2fd7f518bad50f9a79c8ca5fa21a5d7f988d641713e77e6ed0ece770c33f03ba0a6955aece701e52790b2d24834c7a69b319655ea226fcb04880c05e4ef8e4f74c545d6dbeefc209e78e370feb8fde9a1be779e93af6dae6fc1a111e778380ca1674b9cc88bec199eda620b53876570461d204c802483a43f23227dbc420ec9cbd9103bf5fc1b097dc172af6002c150db812598d36cf13783b8f70ee536fb00bd28714ba483f71ee32c3e67d04fef0d36356fc24e247ed6e4c1ccfd2de059097f26bf1af15237cb495af5e4079f1dda3e4fd8df5dff7ac7a073eb5b12b92be54574a2b98609ce506c24f0069d757cebc71c72d834c18ae9098036d372b0385b8e914fe7bf9f650b688929acef0c75ab1d1ca164046806fcb8ef89cee6ed59b79bf6c6fe5346a23aae5e221acf408b76a531cb220f350e9cdc7912b91224536d1a8784f6b42a71143b174bb18c85a39038f44c55b3d1e06059bdf845f92e0b9391680a1cb10cb509bf8eaa327c4e36e3808a686722e02cfb4392492c127df82f7b59fb19625e95de0ffc59cd04d5ce8d4c89d14521845f02e6835efa67e99eea88e5c44a17712394c142c833557076768af21326957bf80da0f58150bd5094184d297ce2171d26b70906c446e3246c99ed49c38307807c59a0c142c05673accf512d1c1b6e6b680042e6a3be07a47df2dc27f6caac7c248b4cedf4f5faa46cb5b681c2b8a6ad6cbccb12807d9d7ce1a9d3997d22a7ed3007a03d4595d112ae40477b9753c6a81e604028e867775bca31253407f491a04e07612b8bfd45ca3a2b38afbc237a73968669887675a7b7cae66c91890a313d2ffd3a2b3d0fdf4e3efc0818f19b3dceb29ffcce7e14e6e2e525560a9c1d758243e7faa7d7432c2cd074ce966d2cb34a6e354452fefa3677ebd8ba106dc5b4f61b304c2e38ad9070432e8861d9c43eef8504fa95d951ac037bad5617ab39f3a1f998793bbc3504bdd3e834367dba6c2d7c7f9c9442dd6f3c24fc1df4a53518078afc0f1cbc62b5f140bfc4e10d0082f8f1b838e37e7680ddd2a179f728ac8026711dcc45da14e77331fcb0e9c0bf97cd4b6caa84113c2f74bfcb1d29d3d10fb190c8a261cf1371085793d3f5737aca76f88d039473298a22c1f3bc036b36a8be0175de4d8e13117d7059661278815febd0d3024de30c8ac9723d3aabb247b3773568448479acfbafeb12a61af1e6cab80f487d22a4f4ed0360463b7e6c611bc4e9f7f1e2257b484e271c1f7fdc833b6a80986ef19b756feb76c592891881396ce58b3372e8c78aea60ca279da44ab932a03ea7581fdf575abf21b734d3eb92ea0b9efe56cac586c07990d0c42a4e5413675ae63f555d0102d9ac9687d1f0bd7dd1fe1136e192bf221c29c46ef9846bf1e298250bbebee7dbb717c9976a4dbdb3f8dcbc93b40a1ac577632aa12ac3169113e7788b81934d2359608bf7f8c07e7b059b6b697cd193ab3e2563853699e47e6a2fa811e040372991ee6348aa32ab6f837d244b557b4fb3d85998cfc5bc0be79e849d1a6ac085c91877b426d0018690f66e29c9f6755bf24bd43c8efc2abd3e4cb0416e2bcba892b4d25b9076d2c84f1d7be24d8a5bd783cdf7f5506b8d593b1a1feb23a9c7cfc497813a391a98d51a2d25bd41ceef2d413605c57c627a73f888cac08649de3c0bc45791922f1e17e2898a6472ba1434b607582ad61e198f4798c78fda6899222bc633258b94f3eb6a3c3c3ce544f3238d8596e17b07491c9cf1d67c085ae2454ff2577955621e17360b1e7f266116856612bda1c5e883cbed1571df1207fa5d381b77093b1d49a8f990833eeb45c72fc12c29a6ea9aca6daea51e37c350ab2c69dba556764e665e114e51fc5414ac533b78c8af45db2404d89c1f3704d4691dec6c35f6d36cf086d772aabcdbbb66cdf8b1b2a40b66602d4829920e18a80ea04334402cb8bfda55c6ab71e12c682c07a3c74f7164525952bd51c2fbe051bb4b1a969d74631de27c7a2980fa548ae13aac9d02a93f23411c24f9119458ad6fca55a77919ea03d96fc74758f6a43382c3f3d5e30ca473b9bbd70db411401e7fa39de8fe94c5b947751727af243b5674220181a62d0ff0356c5f3f17eb4039b30bc5210e2741052eabbaa6af4062915d12b2d68572107c08a96eb2bbaba9b39fa96400b4b463403aece7bc1358a304f4df9497433c67c9d298785cf17da68e41e81547428353f67cd09219a58d78b10ef78f85f1f86b7523e05e817b4cab3b81f7d8936fdd5d9d4678b0dd4f81651f64b2875ab71a7b906089634dc70ec89fb8513b4cd60ad27d3d2ad58a53764ba93ca03527fc99b3f3320f7364c96eca5d4192c6aaa737003c1e3742d65d05f41ac605eebae82d8431942563d71bb516dbc99da65ab9712a9184d8bfef35d7a470cf24974d2045a491b36dc5b74f7beac846f6fa962eaa352ade237485f505409fba06a7e2193ecffd41fb7d3a2b766c9b9d52b08d350fbf138277c3b4d8528e4bdb7675c49e7801bb842aa78c2714ea9a724292c00d62691185c57d2b11f11367126fe70c5784a59015b1c94fe30263999d4340a16f45da7af64e254b427ddfe3def7c7cf24882dc1ae20f5f0bc4cd30901f62473ff0458427806d88eb78aa819d1f91aa7bcef960b5e863624df057892c3d07f59a23bdae40a03506e86591aa89953f957ddb2cae133acf5e0f6d21753c7f9f59a5ac9c421894beb7663e3d665a9078fc44213b383e5cc3c594e98386bd80bc7bc58a9a52fe5c2874d5c89f6236f54d5624d128bb35a33b60983a7e51ad5153e069cec7ed77683f1fb8ac81fcec023519d527cee728b19e4061416fa0310f9208772e19c0edb99f8a99dd2d2919ed4f0f76ce4de0c881cbc1aa144ee14d03be722f2157be1b8503c683720ac2746fa659044feb49cf53e26082d874786e09518584fea9e6b7806cdfad7f29c4dc9344b7418c848c0223e92c0ee79228ae5ef8050fbbfeb06ae7d3dae95b8d1ac14def76c75d948a2fbf3dad94aaca0ee3c06003ffed07886ebfde6fc2b71af208e2639bb3175aae4200829bff234190e81daf47635e8e6556a55ba08b1e75ece0ee371deb00d082098c059d89747a025cd034da7b1bdf1f26a178f8614324d16027c0ec185c49665758aff8b83308e8a3bb0da463fb18ab00dfb71d2843df6d355142295f5f755b26e8b9a1810a2aa5166cedc0e78bf4e40c541c21e1a697d9eb606300fc9a64e1d076a3fe41276dee799e8bccfb510fdb242d336de4ea96df0c780648ef3f0d6b7f44f7d0671a4accb754fdd831ab35ce929e465b6bbedeaa1e0de71aa66cbb6d23efe53c167eef5229f971eb1df17fa8085ee28947e9aa4a0eb910f1bfcbbfa00833267310a703c9c1cde9e038eddd1ff11cfc80ac8c683800df9a94d3604b7e9f26e8e91fe04e2fa58db70e64ff01d923e3cdff3c8546ccef5f20a208bfbc18d5786a90f175451dc23f87146589131ad5b758f0c3f810a6d1d748801015adc3bd5d0e63b1daf829568abc0ce452c438799b35a985a543ac661b9ec81f25f5a073153444de6cf2a093c1e4fef607f77d237fc795bff52a301e48fe6c9fcec0faf04bca490b71924d1f83d4cc773e78de0570aa086a21e3a224025fa90a4e7efa6dd154fa8c85dc7f90ff96c27e81349c1df8656a479964c525003f3d325aaed192df6f96b98407db5a93d862f8e2eb34c058999fbc6db65cc59579330aec94b52fd340a3a05ad28b5b798338ff84293dd85169b0554f42271e68dcdc2df3fe89246071f7aa5d964af3ec07b445775d07205fff7c68d93c335555a5d3da0fe80a37b80114bcaf91f963a10e419bbb094edb7ff44ac15c2f8c4dc422933ecd04673647e9a21fda48a461ed85e11e897becf698b69674b5a4456f6ef6f5ce537ea044a7e440cfd81cddebd41f15bcbde1a7d7c164e6ae20291512038f51e73a9dda2e8c60f4735ad1f46b1d93b31f51eb7e3ab1e8c6d1536c7b65380be9b39715757d6fc232b8df7bd5b233b38d88c295891a68a989ca370226c862ae12bd548857cbdc0f5fa23f0b976a4a5bb581243dc28c2e4d5206b7f9b607035d7cb7f1a4fade67c228df6d39ab6c0649a3a1e1d5afe9bf59976fdd86f70c0ef8cd02fd50b82b88c0c72203a18ed9514690b33571f48e33cb5ccdfa8af378e5e7f5c8c0dede726e9c6a3fecb781226911c4a0efa874e9a97a420bc7162bd67bf7359492bf38bb4a7f0e1209f22404d83001e094c51a3628a86e437d218e97c64ccdef15028a9d89abbafa7d8142e8eaf1a3d9901864e1e6adb895a38661ef5e4844c824bc331ba2ce6df4277ad940903cb5d706c756a141a7c28954ab72da71be9c4bf0b2d72ef85afd926bbef2e587e221a65da39a20a3ffce7eb235486c15d27fc1321a616e338fd7c254111e0f7664cdecfc1f670e25e307c9fcc87c59467946c410a594aabb5cf4899e19ca70f283aadd3d3fa82feeabffc922ab6f5669c20d247a692317d4db345dbdc5b5e98ec4aaabd578dc1f61056fdf36d38d24ecb67380b9daf71f4f8f6147ec983e5820f1332979761674c2479053ebfb4e1cae00b8d37bab932beb70a9e7073b96ab43001b982ef6c5aebfa9fe624fa72feb46844bd3e11e251c4fa75b93157e580c2560dc5771c15d08496add74591e6b81eadb6cc546cf7ef486cc4f5defa2020d00ad0650ef4c3283f90ed665b0308dc3c4b98e89528a45a3fcc35e536d14046acad4c06bb052f755c27b45ce47aeb8934385a687d7968aa724c9b252865489c8078d7233c8e391dc4cf2db6df6ed35c5edb5b7f6092007e77;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h75d7cde0609e2ec282bb59834d5b90c27abf374bf610d1fac9510514c8a9301ff9379a388bf7dc29c6107d407a3f83c110c2057b9ebd3428d92193944ab7773f1b59e321cd7fb836af26f1fb28fe1f73c3b2ad5dd1a58153b9619b13f14797303d8d3874a29fff460fd54ababa566e80fd8aba1daa06ef869701b54b0488de123bc9752797252a8dddf9ec137bdfb1131d426aa1c3b270bc7ee627aca8ee812062522f4ab343f11f796e19e31cc8e1d23f3a784dc944c04254607f17fadd056efc7acf6745d8a83d94bf03d918dcb3ad8ca0a18ea67ee4d736129613d0b14224a8e29c41a00c7a8218d4aa91f8de790ec9da8615caa0c59a318cd09d8403d7aed819f95e38a19fe753e23d207c68667a5764a0050be2c2a41869cc743db57d7d395bfe96b408816dbf1589ed31acd638062e9080e384cb3f6a9d5af1152e4c588df6f6aaa29fb2999dd9c58e0d1353e155f39287c6cf87693aa8685cbb0966ff7c226d29dfe1123a72a4bf48e963371e377b9f582f38de3666eb1f7c4c3eb4c035d626733aa5e6360a486e4919693dd212e7015fff887b7df3d9790ceae51ac9fbb0653b0196e0ce449bad7e35145682f30dac8d2d259c046bd6628ce29424d6d68c92e182748bde90e81b0cd1643c1a879e4e6e76662603bf315c391f3c9c5df2855c2d8f0d0ac5128aad0315496c2ba24be74df972d4c6ddfa94a90cb8f14e40e7df19a986384c1f7b5d57fb688b7f65c547357b9c4838f86eec114301ed5a8cb7d025daaedc1ec91fa355a2bf26668a2d588581ecfeee4cb19500b3e1c2aeec8aec90f6ecc7548045a4828a222996581e171a11fabbb45725e8fccc83358205423649f8452a1cd35e7923a7da8a978f7eaacef30e4477b90db0d9d0774b0e28f191f753c680ae26b74b9ca529f39befb9995675d84c4850071905539df75fc555f9a5186d80f43ed04aa2aa121c4994a794b69b44899f6d78822f1c744a90203405fbd6faa94cea82b4b5bdda2b19ef7d57463f98d7e878d9cef0b9492082b879ef976d5e6793cb1caf6ddd24ecbc7b7643e0b949b967d5793c2ab8aa672dc0f2fe917cee3a290256bc06464d67b1ce5ec8ec4b3b2982b765ed02479833244c4553cba85b0215494651d354e3e437631d4e980499fe16f00073c34ad3d8421843f5ef145c71bff88505c41e6235362de2bdbbcecfbca58dce4c641026cec338307f3d669039bb0d8def5ab827c7702cd000bd25bfed2ae8071c1c8e4cde7c2a7ba9c56530d29c33460a260e2d21fef8ab150f7509d836193c8c6cdf986de95d4723595f4e0c4ad900351838915ba4f44a094df23f6c5a34073a33f1f70f32f64fc48e6ee2fa3e8d4914b84b37642c079dc57fd92cba37ed4f6f7589c3bb9de1451135209bcf3846f2902f54e0d304f5406556161dfd1744dc713cd15db6543b5235461248cf767afc8960de663b7990511dde7a55ac5245df778e7d75013c5ab0702c31b20e43fd14d71e35c14caf803f588c895baf109081e4a413c3869c62fca30d5331ead3cc4280e86f6f0e3505f9f402cd687f585f79b20d5c21af5406091c89d9d37ffb90c4f5f8113773a5c094d2d6a06a9d04680f3e3fcdd42a8c813c9b8752d21a6488077b0f3c37f0517ea44dd7d70c8ef82d1de02ebd2d79e94286d14f5d243b7814e7a821703542001d634a15e2c071c9f383a758f083fd58aed86c631649801ffada7a8dd9730125e72a76681875d4838d2b1bd81966eb0589197fc1339f6580a2bd21094410b29f937a414e1e4af5e6fd1f7e5a2f36a4b46f4ad977088eaa4d32e5f8f7530ae2c9e8d6949b4f671d3750eac4cdc676aab32b095420f9a0b0c302b2b774c36ec3d9e949ae9c402ba219f3618e8ef05b8128545047ad7a40ab92c852ff4126e4c5d15cca2e156fcc5565986153aeb3918e72f02fb4d3a49382d655d5eb353473ae57e5e5a824b42c1b243ace3e4e4134eff99340fc7f6b2674c57e7e815159782080ebd6e976e041fc18aeb000b758a98facafa06aeaf4adb0b51a12ae9ccf41d432d68aea81897566eccdd5b49706e171e6da2541eaa798880eac55944a9722e77dd0023c03d4046c39e85a276de81fc68c9e53a534f2ab69b957d42926af674d7a71da82a6d129f2666011b341c7006a17825e550d0b4a9cacbd78856483dbbd3b1f91a83c97c9bdad273227a9f046124af0fa9bcac5007212235cf3157952ab8edc397bdb7ed69164b73dc09db3819b0ed4e6005c9281884f3aef92542dc2c631440699712cfb2f37a75cb5cee35641c77ee73968b6ad63dfd4b51403c8955031ff97a90ba3cffe2ea572ee6449d57b4b0a007e894c269a4d00367b7c58f270fb3f004975e3aca13c82742a62559306e01b25e1fada66e1985ba9d5463d3b2c02adcc5483c794b0686aa621bce68bd7ec42e7cc0fa7a26fb0bbe55579060742e1b305bb132d2b10c80c93f6f63e7a6a8bedb36892a2ad57a6c6408311f37c204d566207c8e85588d2c89a83058643749a68011302dcb565b1e4797ea1a22279c3fb329f767706dd77ab93848fa5dfc2689597f396c61c0dd7e5bd6397cf3377394d0982a5d2fec236cba2daf7dc7f077af9b07724f6971b7a02223ebcd0989646023b91f2cfe66147f2dcfa82c5a37f1e70a54d98cf5a20d3cae360c11bd589c5308139fa55f600580b41b8a3ee33bf71df4838515051404d95722113eb51aa99f86a1de4981f721cead31bb70329745a3813aacc15a6aadf669fce771153ebd0060ba64399a2dc5ccbd7a746ce43926e1ec277286e225c6f4fff5fb3d8b6269e9f1d751f3d3aae0d01f9b700a8cab553bf2d1f5b6862c7da2d88cf56a5394d8e55d493b6920ec333d99e20b840ccbc5e98660dcb008abdc688198e54239bc884739363d3dd0c11304047888865695eb5f3fc8eb775e3d51d7f0c07e0eba8a54adbec4ce8bf102674ddef605f41c98327c8e326c2578d27a4fc56234fb9333772896726687819f35ea35642e899045ade91ba42af7825777758ab0910d3f34357a3c924441f4b2104b53830abe4c0c3145c19cafebed25784e46b5c13c45ca12501bb26e231e5bcc8b89c70f31ef942828f251237e68f2dd765489df8d7e4a20394e450bb58f67c4c821d1d838094778bfa3d6f5cae9eb0cdcc4699536a4c83f7b61ad0b94051459214bef2a402432256b65ebd63f663eb587710bef2014679d6f84fb2eaff74e868869785ec2ea2dfe050d7607f1abf6775cf0dcf48f4301386d19a6ae87a77261d12e69d7d18d565da43f19b2385ce4768b312e1102f23df77e130a2039234a6ae76e13bcfbd6f1df883c74d33c2b5ee17f2d7e896fde61a8d9e571cd5028b67950ced4a948c6551b7210d3a1109342b4a4aa2fd5f0f02e6be5307972cdb30951c87f6ce310b1f0981f800d0dfd40ea4d54ddf60f769ce8952dab4841ca3083c124cf9009d9781a95e9aa70052d89292792a92a0c59a64515dfc354fd70d0c65584b20a7820772678ec13ecb4ebb6aec7b02bb4352de07d8c54c4ab26c25716afdca39bac69fedb511f542c0d433caa551b20d007bd7bd327596db6a82e5cceb46b9a0f2191f285074b9b7a31d77f998f0218b83249fea77c3746c1c35c9e36440a7588e32067548cb059e1e3ba03f1030decd0e1dfce649c1b04dc039febb01e2dd91ae2896fa7ad47b359ac20e667acdb06a44b295a931d8d030a9ac2fd645000343a5435cd27ab7c0d1322d0225eff41ba62aa0c349b00cdbb084ae9fe71f588eaf9268a8cdf21deed410dbf0697ae17a96f7b6d79bd9019cca2726eecf8783250f07c15c8ce693d04326f42a7283694202578ac19092c2f4d53dd27be390a4dadaaae5569b163ca98b9c819cf8026af5d0f3f47eada3575d3dc5384c6104a6e61aec043a651a8278b5fe69f0a8501a2027834d31d85f11cda4b3edf463ed2f77a02f394dd21fba7e844f0b36cd6ced4f82700f193f93935f1118ffb9ea2058b451d6b089cc58141374d6f8c50c8369e962796faa702a627adb8a1f35a3f838cc81f6b09d86776847622cba4d1905bedd1e792bf6ccabb1fe9ef25dd973717fafb7ac3c714d1cf9041a084dee4d8f16250bcb608c980947b7083539c0e751cf608f98ee45eeedaea16d6c12a2386b4fa319c13f2a2268a5165642024820429477036777207fcc91082fa93c9407901d860e128b18008d572633bff5eec4989504b672716b1113b945585b98c8e10e3ade0cd36d378f4067bc573a3dccc21c9962d7522370e6dfede5d9a3c899e4cdad194bbf85b1d868d65356d6ab1791e9fe49535a552cd6a2ba3306620a1eaef46f3e24c2c214c20f8e29df7931623f6ac34fe9f58aa844336532a340936514b56780317357c74835ccedaa0b36a9cecb3a87204189fde55266a00c5c0dd9048b0f7d5346bd379e1432797f394aaa18e42a5f2b3eace88389e6a1f786098b7895c2a066e7b5223f96ffc27ccc5b0d98f25a5f75d7981c88d65ff249f40483df6ccf045f43fb229c283010f2c191c5efbe9e9265e276676547e3a34ab595bd744ab3c07440871fe0ec7feb48b7b93daf3f0becfd4ec0379854a0a22eccc5e390326c1d7dc4f69d258db751e75787884cd726ba1d86da2f9e5e4a9db8fb88547b1a8154c59b055b2a947ae3299ed580ca2804d75f25ba01d019d8e68d85576eeeb875844cb4f8d6d4230a9c461553667f40b857222e5e176efd9db2bde0a3bcea68c6d393bdc26be0a4fe702c669651679fc9ed5b1f770b24957b199ddba062b236bc6a271834b550f4b25cbe3321e500c5347ad86cd93a0496fa84814f5d0909b861783a1da2f6876c470ec2290b3fbc45b425c78b15bc326077033b78a8028df9992050daaf6d33e411ccdbc12d08ec2ffce2b65c17f5b2425672e25a23594f8d3fc34f60df82da8153e64d44343f9b56d08d57674ca61e46abfb6bf46f0e702786c32b6b1f8bfae24af3b1f860ee2d6215b1158e273a971c2c2feec934b61581c9eac299facc821bc9f9591fea1781e8a732dad364b09298b433af1665d9d94b139b1df36617ca48c89e5b2f20132106f9fe6aaf4a5b8eaef49be093f2776c88a8d90724bd4d1d7768aa51df8d8ab0aa0fbf316f9a1760588c7ad7fde9755979bf7a04908aa25e12342472e8fab77700d60b71fd4c61e18df7bcd6a1713887ef713fcfd7b2270dadf3c2d08833c3047bada35ad381114cd2857a51a56de9c2e824471eebce8a479e7965d2c9581e104cddbde9a937334f139806189b2451983a86dd7b3123b371a335c99ee5fe5ec1aff917fbe19fe109edfe709a807085cad30d5e831d9f263d4c2a3c5702a7684d909494cff9a9f0d7b6842a65554a040193d30c56fe8b5c5c9245b0ea48a9b2c246c8c5d5049e7ea5d1135edf5d5fa46228ad7b460a1700c256f2ac33f5c8dfc0600f6002bbc1903d1db1feb5992978555f6d40ce1c3759ed6ec3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h234ef451dd3fdd550244a10cdeddd136a3224acb7ae4dec415923138133fdc3e5c20d54f9a127b39149965f6923774c875b0007dff7e85820bde2e39fe2a1fd794e0bb786b45ac37402e0c30712a0c0c430d91bbf835ac20b2d1e4070247c881df03cbc310d8f18c732293b7f1016999bd98b3a5e50b26e20125d5a671bcf69ced2595f3a66f4fdbed23aae37aa5620bd8dcff24e835a3fccc70496539eb7e7b2a8f1de73973b9aa148bb1f9a8c14ba375047016c9191ec52c3395121dcb2a97a04a3b8967e2ebeb38bd94c8275ae5537ee186658ea666c86dd41e53fe27e5e0ad88499bc831cbd2fd08af025d29b625990815759c552883ff7d12c3b5eddefd75e1481b573e357f2c0e187d6a0be1063eaa96b50f666c253d5fcd126007d0ecc9a39ffca3817654f62bca086cf7ad626b50b8114f2f6660d856ca7dad66569e0ca739d94edd66075b13437dc75a93a6fb19f7dbcfe7583a7cfe1a2379e579ca2012046d76fde76307343675abaaa94fae95aea3d30cd977c92560e257fb917983c47f411337e7f4088a11e75329e297e42abbfbd2aae86a573d558b836e0db4564ed0979a0d693804ee6853e9dda17958ec1e876edeff82bdd19421633e5a5764e9f21abc3a4ba31600aaa3e28a5eeaf6dd4084d6b054f27d10d8e5566fa0736ffde8f0eb26c44a3e49181e7ac13f62771e1ba19caae5e8a5ccfe3c5872b133074f5a76d8486c1f139d6b97a3db67d8c79785489dce08ff28e590135990cc285abd4c2494159bc161266f10db06eb4e87dfce2dca3ae43a0d04b0f1b6c21d665a4ded41b7d1f044858792e8e1fdc2a4f4722a86a743f352d0696dd29f3b9a3641ecf66f7d39f14e336c266197193060714858ea3d75399765b30224974330866cef45d51fd62b5d384b3f0cfbd038cdc057281dee6c6dc4cfc0d064a7df388f21146fc81bb24f8dbcab77d49fb576e2bc4a0642d5b8df9b98b6724322b56db78013d25131de81a66a594032e0be5e2ca34d2a19859a96f7de9e1baf9788811f7637fb9bd44d91a4681cb1e5c810e54a0ac5c45b74526ee4e53d6ee8774fcff2358756d38348dc10eab64bea42d2b62e3ae74040c23f573d2003cfa5f6c1ac1db7daed5c376c01c34efc5f12eda70b7838b3f15b7c1cb37db516def102ad14b9df6f4bc5c8f07446ba2f490c78430dbfb6c48fdd0633e5e8ebf9af7af633a7f58532d50c4a2dc4d65fd7d2efde2a1531352eb0af0f96d9483c46aaa0bae843c407db1c1a0c407a82201cf70a0a70ba204f3739750cae93dff0f1d9c00fbf5a1385b3b273db01b16bec5a6adbd9b3642fbcaefe1717432f6ad738faab671c8d58e234a5936f04bd9900acc517ae884f8f43b80b6a6379aea506afcdb16a21c3e4770def3c195c19dd785b85e523d7c1dbb6806889d232c3c3f6ee6cd61ce0cbaccc91c903f59bd8e3a6493aa54b714e32f1a03ccc0a62085eb30125e4d236f9ae642489169a83fb1a8d4f9bef4e1121ca242abb1c1809e517db1caba1442b87a9bf78f4ac1ceb16c02187f1b1fcadad038577b4eb93f4e7cb6f5afe5eebb971863a162ef383a292b991079a3c501ff422bd155a0bb36d57d8eba83464ebaa967190be1626bd0f2840a8666bacf9ff76dc38e3d2848c772e1ac01810ee08f956bf195b7ebd7fe9a95ceda2c2a169945d02450779c27d47afcf13ad710bdf72c84ab3c96c2e3d0ce52ce4ae2ec65c3fc8243124f76619343e909161491048c45c951e17a5e5125e57ff5357f7eac919f5e663f459fde9b43b26ce0a607d89c565d1b5defa53b17111612ef9f42cc2526d062e0e7ef8caf671322c0808fcb6893545980b1014a07cdbbc46d3566fc689ec4c857c78515875f6415c5f741a42f704d3e885a1f12170317833d99b3a478266fb8de1c51bc1d3cc510cb62f713a5802cb5242b7887ecf07da89d64553cc0442c288e9aa2c888e64b7fc9f130d39ac954ba522f686b7cabcfb7def70ac4fd4f018eeea92625fbc408b47f26ead7c2a97d51f9e364b3d0e2d0e3ad56a9e45e14f8adb8946d1b735cbdfabf302fea4116c2204a6d15afd424a6e29e4ebe4a293c4d3baad5430d8cae9a82152d4d33dc09ddcf76bb33e0c93a94f497ff89620387000cdefb7cdd2c3840de2841267ea0f288f1502b69766229d44aeaab618e9cf9a5a03f39871166b3382bf21ecb3f793047c66f0b65c521b6cfef196ac5f279ccbae4044ee866780c8816e126def62d1ef8980704bd658749cd62754d0c1058bb66a5bda889fa79c0fe1b5ce7c723b816d22a60c767e98c962880ce29eb2fcd3c72fa39361e97d94d580299b3a134bb844c95f26465c8a90bd7908b20642d46aa90108cc92fa1efc5c8b6099e5e55cb0b67e519e9803c3aa2581f39681413cc71eff35e803175b4c7cc27d21a5c7bc3630b24ecea49ab743972b7b1854ee924e640f155b44576e2c808c407aba193d508dc4ebf5f772e4b9c047d8176b994a6cfce35309d8f9126c544d55ed1f5d1706d161861307d869a6d790a12b5b8fe0793a97c0190172f9b3c599fe9b51dc2075f07402d5f79605c0c198339499cb847c848c6aab0c3375b4104066ce694fb8a3747d7491e3c9ad3d5f1862be2d05474e005419c51aa9675cb0f382d8c88d61d44b133afb4c9d68e95d3fcd7feb86914a3e3c521f28cd4507de5e57b85469ae3473b8379fd05ac3ff0ccd0e41f7eb91d777a998b28907ec7a6708b1e899e357618dc7a34323775a6ae3000af425d22771301c54088032d08076dcf33555ad47196e914fc4359539422217087e80c1759398a2bcd387064ebdc24d09399e66191eba694bedca1c2f98c731ea5ad899535761e9562e1011658234c9ec2af237a6ca9f3494d2b1456155b51f193177eabca05d294fcb321701ed2f12fba9fcab9c0cc8bb122a45cf8b691b18a7fe32a7191dc90eee8b70cfce7351e59d32bf6e8d6984c2e5ec652505bb700d0ade3b5eca7cee5369671de4498194ae1e089e0c0d2bae114a1d21ff6435c030728de646d9f3627ebf0d9539d07843c3256d606071d3062c32d418ff7738a82d942f958cd68f91212f886d530aaa350127580109c2a1f5286429efa408f4c2bc2b8342611f1f02f92b5f692d56e41f03cde8eaa4ef0c39edad9d8271d6d1acb7f301cdfa46af8411ae31e74ecc265b4ccf5e721f8a8a86159ba6c2bba43ba2a3b9ff5d1d4d8e08528459b2c35ef48bbe3fc48a934318edc784be350cb22e7be928ca7c1d3e0bdc63352b0dca4b25fee88fd4f2a88413f621e68ce7a07c4d120b6f47c4c4717e788144b303fb1d0a0031e16bfaf566cc021e786d28d8e21623ef3aef19902292946c02b16d1602d508657c08457fb99afdb716daf14b8b92181a2f53206a27b3ff81582f473df88d524d8a3b90eca69f7f090d53629998a0305052cac676c29a75bca55729709fdc0226805f0fc297f4c292b8f096d7a5553b51a1c0884c07942f2e98c9beae342a4a68aab761a1d591e40b67a459be4d9ffb27b284d3da43941c9a6a4bbdc48762562555d73f0d9890653fedfd237d820dbd44195b189764f0e3b2db95d870ae00cf3ebbb905ad8a2d3f51fb3a651945cf05f376f49e974808b22a77520ef1828337d2eb4d9d87af00e81bffb42ed8d610f565c2ca895b93d534c95074bf005e121d5054cb263b707ecb25e01d765d1ba8ba23c6d93ba9bd67742a548b8fed05b66ef86bc5b20a64a13a2f73b6f72de2e93e35d6a8de5399d8420cfd37a12eafb5d425acea51c21f0d37244acefcf9c9e5b349746be513103190e7aad6739b010b9d2d7c74c7b4be33f23428fae08c7c690a1d6a1047d4b3aad8a18f9b204aebed9657e1b5ef8a4238eb0ec634a207b7cd8b12c38c8d282a1a68a9f04be2ae102ded5f843a63c7c2cd965510eadb5410809218576ba9a4b7924442a68dd3df31d5c06816eefbef00cb9005513912f1079dd8bd2188cd01e2330efe2e23bbceef14e7ac952da453573ca84e5d3fb8f744a60f4e70b885080f14479a1394e1441bce4b5e0eb464878e8966f5e09235b33b1187c2c6f5f97a191520e8f1d6584bf6d65a6842ad1651f127848e05661d333e904edf9e103791e230d32833a5f130d274a26c9e3cbeb51abae6cb290ea6cc9fb483605c8ff0182593e2aba8e7ecb574e76aa96f8a176da618878cd0ddab0e5075cd3ec6e4d2c888335a8065082b5aabbd87702a3763fc8e1b1b977752c86d87324165180bfe6ecdbb5a9910e418f877658e173c3d90c1f8d7ac559e18aa7bf40eb786d613d79e27b1a414b009011e2d970c79eb343048e5783795ff03da96d27c7f38a6c15e9a326334f491b18d3288b08579f85c21f4d2a3129c889e454b138db3edf8b9437ce3da251f9f80d7c97077a3151e7495461db7b9624fefda30775611d92312a3d2a91f9af582c7e8cf6ebbc4760e76200a6d92f3ff629b85cb906e4f364e2a3d424a58245fc04f896d3541911a9f1e3649635f287e2ae3f6dbe15b00803bd662f13753a4d7e5b6e2a6e69c5ac3636699374da7c5608487405548b25322231a1ea31f900c6d9aefe0627705f7b429616d47c60397d2f6a26ebe85c1e504b9ad224bc4a2a6ec4bc674cf17aa0965c3b1826c096bc01343c8e5994baf848040539f28cc273a18b266c9bee62460966987ff06ee74c0185b7b803bddd42de787f8993cfbb3e407da956de1b0689c41728df2e884f02dcd23ed3da5ea6fd90334d5269d48c7e3aaa808c1f3a51bd244211c0e31b927921174570dca5c46e6e13b2602564ee284889410b92be956607d36114620d401b38a5ab0655ae33f021cfaf323d14197efb73c9417194c29576e6112883dee8a5802b0a3d9a9612fbb68dd505eea8dda5033097db26ebff4c1d0c22c02e14d98b0d6fdf6b87c84e060e0cb430a82818761cb8b78853aa66f4b3693ac3e353133243b345c324bf9456200b9666ca4595d1ca0b175ac8c040a21ec15a999f286b24a8059ff6ef980ff943ee946a68c8b141a54c20f4be0121dc7444f72c2a7e26556e21ebadfacd10656a4e1db47e45deedcca0f450660ec2ab2b44775a01342d8f0a3bc446894b65bdabff1467661d8a379394509bd2752db933e30af0f51f4c7d6320019ccd9166e0023cfefc4be5e0912183cbcd5abaafc32ebd76190f85ffbdaba3fc8dc77b014c8f7318973e8f1a05accd4944fb6294d63c764c36e4f4a7f3abf46b11808048d806581fa8cb5ed0ae7aa899214af96aadf530780cb711808eb543c954e017019d743591350f315a5884bee449012d0ba83056a7357d23480486cc2fe0fa78f6b0a293acc6d29651660a008fcaa6e06277c77a346ea9c30f321fee58bc0516baa61283fd637954207e5d2ce9eebb28463df046f8981cb59e9033c44b51860cea0a6a98c0e1d24cd6105624678d270d61868f6d7b47012edd281351561aa20f01208dc7765d59b4544687f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h6a01dbfeeec33639790c0c43a89cf4a54ba0ead0c2d8e6242542429b4258261af137d110b4e5d863e8f5fab44f172a3e2465e36a04dfd7db96e13578aaa087fb021f1ab1f5b7375c50baa4549531880176a534068ca74fe8e84f01eac3c731ac7dac1ead09e9f063ad131241ba7e24ef2f3ff0a59d26367778ec9b279241444a0380f10705ce691d8d9ae89a64cd032c32310200ef5c7199d009c062c7a4894e8191ae72e22e2d28abc4ce537654be4c6c2c381ea285b9d74de723ebf07cdbf61e98e7fb3db74c7d18334607556268187dd84847fb01a5ca264a92fdfbc393d9dcea8020c715577cca7e97c4fb401e96bdc66c322b73ce96716f5989129fc11341e1f6874a5c598e999c28526a5cb8d3125574493bd5290fe6850276b42b303446e9c126e98cbc7f52167debd96cbfc5d79069c53b020322c8066f08645a959bb6373395c50808a1d1427f83bea35cb49dd096840c468928f793510303962c5d08737d42b39ca8f37c878e10e4aad592aac90a1bd92d3b3368296ee4bcec0ed1903f432d933852a014916d2086c3a606745860d9932c6143b6a8f206d3b15148cfcb02e01886110499b5682337967b2da4c53e348c5e920950e8d3e74f44a42ba25fd1c9d36b74b354db9c0ce5e39822e1b0ffcfdd89ecf58b11c9901bd4c4be7da349092bb5e941348240103fe8ae54f71e4d95ee5dcdfa98c70256035161553997eecfc1af2792fe3a344d32e03c58a337a3d16b77078e8aca33c6934542ca0807582fd2bf38924b22019d79a77034a23976d3ca0b84baf08b3663aba9604204c33460f99a0f33f531ae44f4e4a6666d065dd1803a6b6f3c30945f6b59276453d23833ea78c713e5f4cb8b4d90dfa60a57476f1ce8117403cba7d9928a65d6bce7673b4f3158b3f32593c7b81edb4e51710ef94b3b1911f2b0d0ecab09813136b3bcb3ee1bdba1a3d7da9a4cf7910102c261e9d6374362d777e8c61ff8b41e3f293e5ea78db8bde1326b1288698e7feab4a6189f5c7b1941475bf7b20d00fde063024bb4a269d3f06cd01e9561db644713fc7add2d1f3c7dfb7025cce89436ee0722f650c64ba37953c9f516e88c332eb8ba7aaf331789a4f52ef4d1af5382fef87d33487163ad1cb8ccef8746a98e7d2f9877d9ebe936d00afcfc4bdb5b6f5d5f7b84c8128ce02d79539151d599bb7b5422295a47289074dd719b2b82071a8fafc02eb4bdebb668dfa4219b9649a616595141e504d14210339a8c95f0c195bcf14f34510029d9a83f7975712ffb63e740d670818aef19decf6a9b548a3a6228a1522b2e5a394f5e2e581b59f0dddd1ff98a72b29c644e25421fc688774d627314d8ae7fc9c48efed0f8758c34b4ceb484966d42bf6754adf0af566d64e587ba293d553818d2e0cb4887123e5583b82f3d0a1166894dbde6c5ad05686c417be32e0f8c2f41a8c84774104186ebda03ab337064d5c0365d706fb3747a0548fa8601ff9c98c5f0e6d4c14a3cf3382cbdc23f554f3fa81d664a806438c1db271457e86e25dcdd0b1400ba6e55dddfd8e3db836a405be6e14a5815a83cfc2e0e454e15168ddefcb5506e10dd085e4f3eb4e6dfaaf6ad28c9d37bb5ba50ce0be9b6355a1448c803c1de0bf0c7ad13cf4b5e944e2bfcd17eef643a922d19c83eb6b3d20cec4a30e1441ed0b2668d7fa86b0062f1e1e71c81d81ef9198901197899f22f8fc692af0a2fafc8cef8091674f4dc04d941087c0518c65fd6967b6cb6ca18d0cc8f787646fa1bfed98d85bf581951ca4507d46c947121023a163d22469acde13f6bbcbaf272fb47dda359b979290b8b83db5bc1a341e80c07e16615680df778052094b51ad1c1d4415a76bc9298c5eeffccf2010eab8fc75c404cb039fb6a9426313cfcdd497e0e86dcb39f3f9b475825c0907aea0db8dd67418b820eb2bd6192ce788f289364566cd818d583041a1c17d8894507ed6ca54bbeecfd310fcc01c18700f194d9c2a75a0eb3a8c068c48caddd1eedeaad996ee4a781c07ce332a9c3e06a565f3aeeca01e61c7dec2e79c83c2ebc102d04fd74b7fbd7ebf643bba479943c9d350a21cefe39b13c4e1f2c71ccb7bea27486c754def9d96bc55c14e34055f0a219fe1e20ac919c4a3d5491b5f7bc915d9ef74cfcb45b074c52e46a3bf1ba18415d601648a564a43aa7d0789eb18c2ab0f6d27b323c659cadf80f2179d8cb17110722c4fc953b9b11dbfc8e171f6fdca94f5e55e4eb1c1d80d7eb0707687ed95b827d68c58803101e7ec436fb7aec86c62460b7ec36d7497510533ef0e5fc4b2124485f2673c067cdeff0b3162412120217880c6e41a92f87f2409bbab4e096de37064c3d9ebf57dc38a3308ed0cf106f18bbbcdbf5769f5b00015bf191b37cf6b69c8a4adba5d3a1f23230658310884230db23764a421719dee160ca66cf4d3969c44c406cde8d79b8aaa65e4dd61715bb49724f00da26b3093d53a7bfc99728575e62f71681bd965d322f2a4dc0dc67e4cd618f8f6fd9dbd71d3f41ab491e29bf383321d2e3166e9b68f4a4dde0dae14dad5b67c7433e50e1c8f7e66aa36a0353290874c70b06de68d6f8de3a358ee16ec1bde30ab5e457a799e2c5a6d039d5fed66d47caa216c06f6ca535a7b0226807b68f7696d583a58defff1cf19b2aafa23d0663bb670a346f53a3a246a09ad9f454db39d57e0317564d2fe7fff4f414576e43424162a8bfb76c465bc9e41d02f1b8a98f7803f7f66960a412bc2a6b6446a4b32b0991e2d892c66f1ab1a60c57d8aaeaf519aab07f0b049baaff2346bd87cb082d35cd344c92c8ecbc7ad5f2127fc5e556cd9665f473f4cbbed26b08eac4e204bf216ce2bfbe16b609251bc5eeb232bf4d73dc53261c60498df991485c6fdb47c91d93793b564b2a18876c859594393de24b63b83ec9cc91ea5846241ffa4e5812e4bdf5ebe2ad659d4749a7e5be2cd0c984b9947bd934ad51366aa5588b75489bfc840a7269755bd1bf6cb9245577bc494724b56ed1354c77a09014c23399a867848fe6a1fa9a2ac61bf421d362b0187f3c2c19826e6d6c56c986df99ca006f5e85d30f0644f703a54eadb128589271567c0f1a127b837c919c3ab3f583225db39031981f3908797fc75eaedc67127260687c883cf8ae99988c06d710e4bf331571fc8b8a821b1dd708678fe323defc03e371b327ad6aa5befa6f56d7ba5764f8f5c5cc920d623adfcf385f11f0329e2299a03e0b2e0e53f042a7a9679990880c5decbeeabf5172de2e64919c470874732ff78536fd1632c3a68d34a3600b222d96a02edfb68848c41865063d126543507121520b186c64eacf4ff0a717c704cc2380377b6db39251f6fb37fe6a00a185c37f2824e51b3ca66ee3a5437fb81c201b8f0ee3d3c003ef50b112fbe1d6bff894edb732d248c099654f202df65e7843d02a5831fcddf946a297557393553a3d96d4cc0f1ce75b496a71fe39c8a8fa0661f9627aa060eb13e70c16b1a7f1490ac14ce1932a3a6678eb73e902d74143844eef5486fa945dfbd051c501b583db80d0ca8d3641dbfa87fd61403b741d8f35f5d935529a75adf5b37871b45d026fe7251d7f91834e8ad39baf9d09df8c759f6096974ca02f5876819a0ec6b20781ae0038a90b797289f24b989d12a9a70cc433cc05267e2019964ff3f3287e46172c488b9e8e886d1e8bc8857e34c2ae0011867d92215da9aa66bd638ab63a5be028a6cd6c1030ba549a7746481d14a20a0d3d684c85afd917cb67ce0a86576ae48a8fa30627e13c79146c8afad82482eb5d2368baecf16f5079d843e0a33c9bcfa606df4a569390de19fd158fa31d06d18d71512bbffe8d830b17e8ec64a17db1bf5e4f9c85c8424457950f9b088fa23f05b6180d2d04e013af556632b878b8fc6d0ffceff20265fee6ab673788ac7d1979523a6715eae8f2873ed07b5c58c55ff459e06b077f066dbc1e85bd716df7609e9950036e7c9b15a2763879ca80ae69eaa26fadc19afa558a4391b35597520fb0cf53a48e58546fcfae857c00ed1bfb67d41cef95c9758fb4a363827e34ac853b8bf75351a1ff3e83592cff667d975beae2ed3c44920c50ed8f933271f6366a20a5b69ced695a19d10bd5142dac9b5045b8283f399657c9c089edc2616f142bafa66fea5113c56dfc1b4c03d43c78fb7768ca4a11ba51d9f9606618364095b9ae7257bc5a5c45b2a363307033402c43a3b526b7a69137995c8e6f29314275827851df259bb1449d59e1716be282cd3b879c24facc4daed9c7fff9f0a88c2e651db33522dd34e2fa73ea10cebf84c8bb8ebc00e39ff086a36856d43636bc258af87783ed4ee181c086b7cfbd10c8d4a4faf89426b832a23f7e0d45d3e01844bcaa2593d8d99cb0fd0cea8f7d1a77c2c883e6368a3517736283ad9819961dac040b5f60e28fcfc795998d219eeeffef354766e5d1e942ca9ef85512ecd74eb3939d93f2d3ee22e74de915a28e0fea1ecf7f04edf63de43191bdacab676adb1d65073e208d8897cc3a029ce2cc0d31c73f06eea823c850b93151ebb1282d8e4afaf3c6a676845b61256c5b9f0f1435412a5c0362ea87f7f26f891f762b1cdbd0129012bfc1a26ccc166f0ec7ebc4fd966242525a9fa8c4da322d0822f01ca90e641de411de0bfb0abbe8d18417b33da28dd912d049b35107e2178a9b2240a5091d1205c74371e5cc3125de2f17240d4027eebcb939c9ea40125ab6dd80d0ef0834c18e8f91e1033c6915fd94919971a765cd2944ce3d2d10ecdc8fafcb330491b718907df93f0be18edcbdf42aefab419032688df59873b55fda9b6d0765a707047c6291979d2e2745e8d95044b74d46db8d16e26079c01d4853dd088a6fa765e54990cc2f773636ec9696f86c5652938e13e13c0dffbd25b3aac389f89a2feac6584c56b6f721ec9332ad2e02b0a4527f77817443e24a394a7865ad6532e7762ac427162953f289d02e4039c3392901c3c16412fcd990b9ca79a962972d94f8d7257064454037972cf36efbb05b78212fa64310a65db0a751edd5fdebec7fe41d33a5f57eac37f262b5c7c0ee868a64bab1d9cb2c3ca2a60b7361c99f849fa5190201e4d017de98faf36cb685e9448a1217e59afe0c9cdbe512b02fcacef26bbdfe69760634475e897a123b048f6e6ced43809b00d388facb9528b86b4fa5e447b5042beda2018e805f5d867b1bbd07b57f57dff555f9ec9f6707f8a4616601edb544e0891b2619c45562d9bcd953ae9217c5da072945e0fdaf56c68fe19026826eaba39ace3470682fa073a8c669995401273c3f85138a0725a99920d4114a048da9abd9cdef755ba10aa66b4263b0addf932e5559bd35b964d3ba05fa77409468c02c445a5451413d5921a72116ef74edd136805d20c4587a79350441384083b28897376cb72302f13e711aaa453932f3bfc7e370187f5f394e1144dfd92034b3c09ea63d33b964;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h460b2aaf95e37ce37839e36c89451f76c65632a3e97367a9a02aa29b4787f15b1b47a73bf66c5b4a1c9d587d12e291c18a46e8277a6b856d841d6465f8242a5a3d5ecf04d5a6d52c485430d3e3c86ace8de35e6f0a473b1bdf8100b1b409b5d6e82d06d59d920eb0d15651ba4b92c93d77b44da5929cb25dc03863e8ec5c11f0079ef98fb4df0c22fc38d2416dd9aaa0cec53783f9cee84805fd3e007a67fc00d2fb57a6997a8d164f3fe9a8ce4c23df0d0ca517f8b866532395fe895c4eea122f9e48856f111da0afffc2d9e6459841cc8e10e7a2901bbd7dfad7b0cbb840550cfe0b4349682cd6ff7d7cd5a33ab95a380fe9349426b6c4de7ef3d74707d3ab79d593da48fcf631b8e9e3c4ac6017a4744a9cb620257b3dcea19ae95c77c7426aa9cb791a8cf3d22d2fec932cd32898b7d5da84b677d1bfb5e026ee14777626bb8a3b09d3045334c4318dace1858d03b1ddb939af0147234dddfd03b741775a04158fa57d82ce807868a71c4affebaab4b5a9cc877108a830c855b0048a300241a4543265726d49fccc44c694cb058d4790a0b6b12949201ae6d65af43b3f6dc7a3e7fb893392b67c7c07c87cd9f77a9b590c5f35054b7a37a153e507db1f51fc22e1eaadef0cb8c610ef6c8d27522308fc175cf490cb566692bc9167c39c4dfd05b38f89da385f3ac9778fefbd139825b674296e9d0dce5779fe8379bb902be4a407de20e4985a3124e484c7b87931767e498bfa1a65d55a1e32ac864def2318dcf3b18c8ec629a1900463ac057aa57c3fa29a2a82d569b6c0b2270a8bd901af2cc5b69849943697922c8f87b8ba4ab429f4004f873b8452b0f8d2d8a1d0b44934c6716f86222263dc3c5d2e53a73d16f978765f060a0c9d24986f51d691cd9d490b8b2ef6623ad09dabbcadcbd19bcd7cc251fdf78bbc6f5e749a83902f15955c44ee23a18885fdeb1fce4e9edcbc27f470a955995b7ddd905382ce3372729c558745e41742e7398351d440b853eb4f55b0f0dee32dc5187809c5a6afe93fede8d16840bf5ba436988472aeb8c89403617918f0fb9b8df39e705ee8012229ccb5439c7ad0f99db36c9f003e4ff07b26aca9012eb1769f5f7de72785815c2f82b6d5f1c4b7511c9ab3bdd9790a5e55174310388f2440c0869032da31a2518caf7418f42b7cd88fe95188363604f0ea9bac260fa5bf5d804e3efc198dc7465aa405d17efa81b5a470b9bf45daa38f1e97051356520c30145cd7daf57f42d203aaea8599907b9bc49e87ff89746efb02dd7d13a59fbe7b2e16db790d7579023dc18cb754113239398819e62c97c7172832af8f0919dfc4c24b1efd52b9993fabf0b6d27a6a5f93a0ae65eac9f7f1a599c596c428b6dff6e7aac9cac1c2219fb2094468988f3746b1b1faf5695ceb272390a7da4c589befa5b9147e9164891c061d504f5e4ead1c87b0ec08c145180efbf4070d2258657dff5cd6ef8de250943051de6f65cb7573ff9bb8c741d36b67ffd48bad90eebbba5d49430623a94cf5f52391dd2cf1dce74c41d34bf46a696d1bd6085ce2d98f47bf764063e43e4eb894336b3e904a7bf403088fafb4ea2b53c09c846469352881f519c788dd8781f55f5b1ab56335d0a76c33406f9eed8348f0f33fdbba51997772419eccf5560f3f92f8aefdd2e9db42db06fa5aef1e62e272bc102703c2923205fd7e5317027fb81dba4199c6691d009174bbb554a222cb0dd0f662cb89a012487be82c97cbb0da3d96fca9eb302b61a6d8414e48529a7c16c8e5f167231b49fb9f721283467951443824972bee8f2dc3c88d85a283d596836f783ed408a1584725b7d4935dc30ac652ff63da6cff6fd012c5fb4dc9108fbf457c75d989a7c8b0bc7e7903d5176d656875aa03ea81c68915c77d1475f337df3a7192494a0901331d98623e5846ce42a79c4b7389afed885651dfed082a272f4c78f784370a2f82a3c15d8e895e9d93e57fa9a2a0b533a2af0de09137eff1b2c3941b1d11bd6eba7bb53ff979c688d3724858d3ae7f2bc94513db7faff28dda95b5c71cb9587bec334af8ac883d80ea4951d0fde11e5e2fdb4336e4f5b6608cab70b76e851c42abdd48a61ccd570f7d4d6708dd774a1ad67e61087bc3210946c86c383ce8f7a97f85907dc2dceac37801f56e415beedb730e2ccfda88f9d85ec7cb8f6838e325f1eb0fae86d0f30a1f4593fbb909a647343a7628b7cde9a63dc4e486fe5f8b22f138729607354b8eee1ff97f8013c4db738162e3251725182df1f4f9ff6bee11dea7302f6f4e7dff80bf597ed48a03165baf43cc4caa13476c543742cad674bebd41b48437997bca85cd45eb9d2a0932af38c225bcaafcefd3bdd011eab394d6e2a3ad64c3aa751c72ce9487a23fe77b5905459dd565173a6d93d55714e9086162228ef0860b9e1e8f5c2fbd9d7d016de29324bec9de7b08b4659e66a63d69445caf13d73c5f47df10ef56501fc601ff23a6e4f6c9553bde32962c07a8c01e6959f87d4eea738199e458c03310c7f446e8a5b617b9b7da037f9570f2423c74953920297b7b42f2965a8978fbb3c9a6e954e090e991f3412bcef392f7d8fe3e4f8e133552da54b3c316bbe77974c487ffc8e7930b3c2b23f1ce590e212f3ebf9b17da33e7e748450511e73f232ffb1b4540817b7976b2e8bd53189cbdcd6b605d6644e959ead3e1c13d512008dd8fd015904761e3284c28b4a794a93634ef8d525cadb07ef7e29f55ce07082b8ade9bd8c4bbd837d20435d59d328fefd10475a67d44f7bc03d0f935bb203090a863f4dfa7c53e9140ec888f042cafea7b2d571b957a1340b01f3e9b14578f970e4bd2098651db9fff27e14ba28c884fcfa20eec2dceaf3118356a1adbea30e40019814c595e80db30ec3ff2e3936d2994f0b7b64720174e8693b46671c20a4bc7fe1effc2eec38ccb02bfc8db379f08cea2e55091856e4c70402d917ace6c7531f5a4f0f0e9c42fb87ae28c66fcff18e99d0d07f29af4a7c2ac461379723bcbf92cf67017f4760b0d258ff1f30b0be699cee8f15316abbe3b9423b8d4fa7db945858466f3d4cb28d5b4c141eb7d6d63c635fd48d4ae19b0b2f68271867cb682ba1cf29ab59fd94b55d5c79de545de62d4fbc9081eaa69f8a282c63ad483ccc4c5c298cf599f6bf1b6061bd38a0b964bce662e4027f20bf5f20080efdf4c9eae5cfbc4b51cc221486f4e51a3ab2d0d4d0b22e25a813ad21a619a6830051cfd83a2641abf83b5e1baf03d1fcfbfa0f28fa6b816b00645ead1a82621f023d06d7aa6887e3de930512cfe9d1877d901dcd763c9a0b352611cd902c13c543f9b3a95ebc63e58d76ce5ec50d2c73dcb4b258ac03120499f32d3a7c5f36efaa372f061b82ec2185c30dae4de9c4820bd0c5b979f9144747d06c4e9c9a4a2cf714c3c8e999c83e8b6af2904fe85554084a1887d8fdc159f39472a61d5648744b028092c6a780c366ebf8530dbafb76c2f323ac786633ca6d42f900d13749ce67d341417cf77980789e1b6635c2b1caa70817215da2fe4f50340f10918856bb738f7a94f10575f3739b517b09da3e85f29fd6d05249df516fa87f0b2dc410a2113932346d1b29407907203780560d76550a303065ee83a876b7313ee786673312ab7c5b295a4b071e0e441af108a6f91754809e6cae9e503ff422254bcebc1e55fe3eed3b0622b84f8bc04a4e229dbf273514d2e101c66529b4ed06dcc0f4bd3bffa389046a1fff6759171dc329951d48c0bb4a9858bd1a85ac5cbc55e080a4bcb2078161ea40328e39fd1c982c4079092bcbe3d884040dcb0a5413f0400827a51aa1499175b4a71aa36a9b2f4389d6925f66a8476b72ed05d969eb6d00cff7678e1dc3fa13e3c0b6c17ebd48b735c8a837ca307858f12e00b1b65e9f69b8b4fb76618936e1655f76b5c82d9dcb3b78b1891490aa244c90289a2975e2ea3356c195b930dc08da8327b14dccb32b72bf7d45b5067b4cd559ddf738b8943a35034f0d165213659c5de010e145b0d7eb26fd46bd053780a62bd5c8eab06f20ff7768c1b1e34e5835433fddc813c9afb387e2bbadafb8f7e319f9f357ea6771accb1750986e3a7bab38aa8cd4f57ea4c785e44f3f5c999cd259f11bdce13c90dd11ac0df0ae8c0643613a9c817e2794c54797d3a8ffe43c7ba3c56d2ee2b3ebcb554f175e31017a3a1ee07c484fa1c922510bb7a0c4bb4c01649bdbc144c087b3a2ba07c24f828760eb8939a94b52e5aaa92fb4ca5fd0175ed2d8aff4e87e8718d2a1bd0687bc36d731023d615a631fa11c94d248853e3001e83e3a916cd6d41c91667b2c712ae8be7ced5f509c09f90980e6b52679b4a69a6cdb4f4ebe7cf31bc1e26f303c22d83b4af2cbfb3fedb81abf36830485bf85c72d25dd12e76b329fa6625ae7755b90ff23b5ddb638b9c6f35258e70fc01299fc492e6d47d478396b08d74f55b432df6637ecfe4ade611a490bce72bd2370e3ec75979a055543ed532c70d1598208fe527f9473971649b904173526661065cd6becbb79faf90c36f2fd51d8d1d53d2744311d6874fde2b2b7b78e3765d9b6c07d749e873275b84641d62a63f903dbfb6475717fc06109005c71cc4531c0f8713086d5cc87a48b8fb5c9b1de70ac67d154eecd4871bd8832932d94f06a073b5679ab36b35ace2a64b2733ea330247e7eb5da008c5969b6154cad44a22b81ef3fc1005775a41ba27943f03060103c33b9d29232fde8754142fb7c5ea8d7210397d85bac0a89a7d161d842c38689f43b5f7a6f9e39eaae57c5d24f25df8ecdc63270cb7faa0132dbaf2bfbcefc2011c03305d3d751f600e583ec00db2c16d1319586c15c85b6e71c3e01273905fa7735c01558383f4bc5e156ee39726375b0f880e408c661cbafb0ead454c2e29e1166edba81281d4cb84b47954103dc60f12861c55c35ce06bfe9b6e2d9de3aa686ae194b84e96e37d84859a7ad40ae309aabf4662d7125fe6cdcbe26d16afeaf8a605366c71207179f8618bb451b47453bfb8b24c2ad7953e832114a797d6fac9e2631376e360ca5551f9bb87bd98ae1dc4cac755cae18ae79bb84b6d5bd4e9b327a94e67b1f2dc9961f13d2a5fe1f75be1af0b4053e7095feb3382318d24957573eea7815bafaa14298c73f2ff2c5e60b732d786945001f792a4c9da144dd134be754c209cc8bea28f16f05a96e2c68a808584098393413902d3a6c1a2bfe7bcbacd87a2f87bda07836f28d43e38497bc4eeb340877edd0082d29e14f728aca688c612f7c9c5813257357845eb0dcb5fee25a0680d9ba175530c2b53e811786633e25bc1d2bb7f94856750dcae616cf755e422d3096ade7c4dafa9e254ae3a77393a9e5825b9d33ea354a1ebcc9cee0b377feb65810ac7f0a56af3d5e0ca391a557c6353534b57390a7239b1f102919448dea82d7e40e450f9436f096fb7bda95c2bfe2c4f07ae1e307c3f67ebd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc311aa1b5bd11be0ae61fc27dbda9f76866977af4aaae52d709e2fb89c1812fb19878ff9fb9d39a7e6e74d2598c18dcfbfe5c802fe42169a04234fbff5657c0f4c3f1ab16db7a05404dbef38e6e2307e2d0aa6bb1026a6a84175e82a8ec1861254bb6f8b7293100bee443f9be85a8bd8ce3657fa7660ff9e223730d2769e66c50444c3ddaed99ed11ee7e8843120f329cb20a3e36c8e3d972e3d28dfd7208061f0aeed6dbd0832a96e3aa4eebab8b8d68fb39ed8be423ab4040b91c80a975daedcb0ab34d314eee9e3c6e5383e82fb8f4cc3d9b172a462106c23abaace2c7905efc616a1c90fefb73ba8e3e1ba99cb02b72f29f16dd80d5d65b05c52fb817e0afabee6a918b6870a0a3c15d858f6ad00983ba448069880be9f9d192210a9a6d9ae069635bac483d57e3118915648067ede0f9f49221def0bc0b44f513da6b2647c87adbc836db0d57c2645868700edf54a2144c81dfef57801c20cb239c2cba40c3409abdaffe777b369cc35a3054fa88ce482ed40bb3f1b0c7bc07c0d9cc05db05e8c1a5d339e3467bbf3835966617718cfafed061fa1204c7456c04ddc4951c712b0759eabd1e8668e02f37745c413225e11fbd1323dc6b80f1231272152ed3d4ac62c6b0a9881dfc57ec24b3e0960db464112add4e831274bc08d2507ee734fca1dcc16eaceaaa8fdc27619286ac7525314cd5d3dae31a55f9179b63a2a744efc82aff67c0677eb0fe1d5a9ea73717bbbffac6ad9c3dfe538618bd9ad594e3fad435a08210c194cf539165cb043a20714ba88af217b03ea56f5db5dcb1af5e827856779fcf33bb7d75c0e3442bd8ff55ddbd0a43fa20374c8e836ce3f86eba7addc25a33a6bdabacfafaf13992468ef73e62fa615cc4264a64f7831a6c033525cd49e6c2464db9b22140a44bc7e96c955bed683fd03fa8548ca93d07d64c377469d0ba52008c324bb3b76e797c56da816f2a96783f65fa072cb430c4ba582f92ff8d433f27fbe391136421b2bd9c7df8f933b1144d35f79ed2d633a13395caea744a55148ec820d6488aab3a3d2d6285a5e53ff7cb9b8d9bd889e318b624f91506633e55c03f60201bbf8edbcffd5ab7ca3ab4ad609912d33f10fc5ffc8759d0238201c20d4385cd7ca2dbe5722c0be9d331a373ab327caffecde1a993db2ce220fa9fb9e7980900d55aa7b44c9d607ecd99e84bca63781414cf5206b31f0deb54b5f4a6e7c863d0279bfb64cda57eec8952c0b796220f4a4fe9d9dd16081a643f9c9bf1c701dcb2a708a51dbb6b0f3d44026c93037ba47b89a776628284e50e8aa75d6cd388311e663f504cea678ecfd07c5a204b20150e87cd4efcd96afde3ee7c4d9f44fa74aba2c118daac3eb8bd9aa3a33e03d42b49eacbc3be3bd07765297f8fc3f74f3e6ba7efdb9a3610c35b5836c473060471e5e04f72d95850697e3768a6be438565737ca8caf04431c84023325774b5a6dff8ff25c9f346013aa5e1cb1834f09a09af136d2a20a83ddb7e44b2de04c6a109e9b12f9b5fb22d0c7c02571dafe26cbd9bed50389e7688b866afef931af0a56f27c4f15da451388d335415f3fba06987c1ba797ed6f87d41c80f4789e0f0b8b11b87f2fc136ae6902207e4623a0ec383de7a660b98d61d1d25bcb18500ac676fda22de81a58a3e1da68058585ea0517dee58f2bbf4e01e77545610bffa15082b7536e0abd2e6ea38235a0997ca7138390d2d5d9bf20d0389ffadad9bb0e7574ab88c12e60047cfa6b582233df1d52d47015f4aa117ddf4c7952c6a440149b04f274a2daa9137e02cba3178082ebcf80b78bd974b59ba29c6a8104a38571dfd0315fe7fba9cd6db0ed2c59b7399685f99f0a64b24e38b88c3683b9cbb63dbeab2296a1797548de0f82f498d101bd84c840e77c27d3560d80658ecee9630b8e874084220f4f10c568b4f76c094e5dcb027a5b6bb337dbd828f2bb4d4058ced4b1e56ea919f67b5212b376786c9bb624cd8028dce805309c44a51d8c7213908440d4ad055defc0f6a141c570f1bbde2f2ddc0c4c5a910ab1b2d74e99d713092d583bdec4c9460b4ee1f27fc333bf7d701acbb7f00cba28212cb366e7c92a15d309e7f5bf1e67a7e26ca031b29ffa77c838afc6ed23f34380bb0b0d8517a228256049647f5b0511773e20af2dcb64118ea3dc475c8d86423ac6680bcb6789cb7551f9d6586b3c484c0325baa7a292d26379bc78e71fdc58e6bcdc252e08a6342e30eb8bcf799779d5840ab7d1dcac8ddc260d759d47d97680e6e8686f210ed4b05c2f8ee11192f56ff9d8d76a6331e685b67f751a3640c794ef499594b8f29ac617baf91961c9657b517decce8259bfe18a77af29f15d278be1dfc1faf0d1bc8339282b1a0ecc639f3c78eb9c6c50f0f65adf98e5b5cc23cae76097ac8973dc6df1d9b85a1f62cd1d2b4ef9ef78ded15260339d040b5db3549704fb2ae58471ddff3243b5a3fd1e83069205996e817d17c71bb9a2ee65fcc3f25fe0b3a98f06410c3e455f9aa44735f28aaeefde7ea70273fd40d0e9be87b46e1a16dc75ac6c1b5104bda911ce37335a74b2fd04e032a3cd247836850302799edd447812aaf3378802d9f2dd3e22765efdb6fab0fc87087eb372b47c6e28fdf333e906928fa244300339921cfe300b38d52e014fac9e8a15136b848f0d2e0cf1c5d02a6f61455d38c18a64259b910a06ee53a2ed777474d7faea5f6aa3abb65db30c369a9f89003426d1e2d75b30cc2ab2d540ab6d9abed1c280f0af7b4710ac2ba46c3aabdf7506e1b20c9cd168e5dd4d5e59fc8fefa9031e8307f940440b6dd0571918d306ffae75fca3770999ae9484f967a3c2c7b0432fafcfae66d133f782e89c4e1385ad563aff553c6bca1c74fc2c517a43f59f824a7a9bcba9f01066bd14aeffca69e1906256cbce3004cc8efd1ca1ba2c82b84e0d5f359b006afb53d4150bc8057a0be3b0c7a117217fff7b75c228b06392a6baafe36016416ca76bbe36e8a3c22764ae954897e86f68e63da5b602bed88a64353e47f51387794f7dfdff6e4a1f326fa431da765cc7417359c8c618eb9de8c8f316f485b2888e7faefb1e1ccab218a3b6ab29ab17505f9e4ff9631f0b9b6fd30e67a299f069781e11a3c2a894a1833561d6b9dcae8ef694a0b676fa2b603d77e5b513be81fc59e30a102c5e4597c13604cd6c965ae2cd50056c19a538a9ee1fa3e7d9d37e1df8a18fdac4a05fff09839f3909c8ad966b7212339cc8568902875b2b7225dcaafd172c260f9b8346c3a8c2110b852cc0090e6a08ec8b5a982a38f38d47773f243eca35399e74d665bb8bebd614bf6a8784bd07fcd69804eb1533b9e93d5b2e0c244cb340196392d376a594215c443d66126527c1bee66582b847a2fef18f7eb0ee1007df0e0ef8d275de84a5bc02734ae10073bf0bfaffc88c1c2bc20e50f83ddbdcfc66d7f195977956a39273e2f2a36e88cc139a449108624617ad814962e90a0edd870682c78431ab7fa8c1a3d0fb68d7e86c4fd80f35880362d8df88976b91c715d02f0c09f2bb09e3c57c643cbc834214d3eef90e24afcd13f32448792f92bdaab0491f11ce46b4ca4ef1e6fce9d5538af86c287019c46a0acc92990c11735943eca340a1c96b5ecdd9e0e189c2941aa64343bf0de65cd31431d0a03b6a27dea150d065cfc4f6f45ca3e5c33e90968295dd26585f309cbc304387cccf3ebdd3457615cd339526920f13b26ff07f5311f5c6667ce7770b2404a8b5cf63a758b5f179235f117152c4baf0b5a762dce570ed4dd1b1f9f3c37b99bd69011045823543afec96ad52f4d4873a7612b01f8d7f5d6a26ef502d8d0ae4cb300d15f0ca719cd150849e6db8d1a1077fa139d5d4c98f2695bee4515c5e02e2f231546762e63bc0a4b434ed55c5974448c451d28193212d5d932b4665516470248eecea21cacc883875bf2ae35c071abc7f6fc4712154d28647f3ae5c11e7534f413248e44c4f2e5f7cd294f9c40e73e3de9c0ba4f3116ce1525b06235f47166abe54177e1fe8d0acf9911bff655c2bb1ae26013c2c201648b3777710558786c2f9260c0a252b9e0e1b26a7b6177c9e59242995b6438a30cc21612c776b74bbc8d4cef60a5bf35858f4486785794a1a91b040ab70021809d0e067e88bf6ce998474e2cfb4f92039577a340532e8d8c38ce45f05635698b68da25f4e980d30cbd0e3f84c03fe38787d8e00e94a275df259d2a69527466a314b6869232c0daf333227b744f7b989c432484cc452182a92ed17d10c78130e5b2fc3e11b38302d967ecb6d8605c35c5b0bab0c127e4d9a8d08bc1c5b33bf5c95003969d67796f21a4612e89af21eb895c21dcf3aae28681180518da90c98099d9c0df4532e9cb5d6b2263550ce2932ee007b5cc7ca238c9b02c8de51a3795788f94c502681c0f0df06070e227d053aede00af901aa33616b8772da42cba1c02a64f18d98aa2c61f1babdc936ecae570142b3cc0ff471c87142e7c55392d42dd5dc80044d156f1adff02783569d521e369c20858ce50597f7898997b9f32b5948b50424ea69f90d9465d75ab951bedd5c9d410826b3e8167f9a1809aad2bf39e8cff471052033955582650f43bd69dd76ce3ec50e06924afd85d34180a9e6343c1658bc723d5eb3eaaed8e34e208043b9ef62b73a0a2b7a2634967d7b583b623da26e91a9f37a6911cd8b08df67bc0391774121faf431c7a8fffb6a96def1dbab11f65c7be9670c1ae90224e0a3a5d2a9157a538afa97f0ce1f2b9e7a8a1b8ecba871ad534599d64a279ceb46e2e931ba7f3f23f7af26c9437ad7e1cff64fcc757709a80f464e20bb6aa49a08b6a0f4e3fc5fc44b4a9c31e6f1c9575ded2a8d2abf3cd8f7450f0c4fc4245756fb15cfa221fa6698ec4ee88ac98cf519bfdf42c75cf3192b5757b2ac80be6679fb38393cf52c585f9dcaa106ee8e4fecb282b56ef298502a288bb77f52c1bb9b409745219c7e25ad56f345b7ad7349dc2bffafbed210f4eb96bedb3a0c794f3a18d033a6dfd3f4b3e813a7513678a325d06f8ec24dd072f092ef2228ea7addaea1be99a60b6bd178bce34d6ba980d3d9abbb5aab74a0ca4089737d2519cfdfbd587df98d3d3dae32a1de5540abacdb371337feb2e5ef7e9cbe4009886f72c99f5ad8d47a03ed00eb88f0ac38d112c3bbe08fc6f8aeab6bebc1f5ae35963a52278c060c62c807e6dcf74cbc2d2f7e54377120064a3305846b76f85af1daece2ab74ebdcadf7c8a679bb365969f8bc1e6204f68c5cf25d70dacd74bca6e3d24b23abc5181a0b1eb588060b1ca8574b061f4df40a9bda6c8bf5b30b337245c04da8c0ba1467589efa28e8cfc83255d823055eff31fcb4d0dd80966d461bb7e37bfef84bd34ad009110d41bdbdd94d6cf1fa99e5d43c5cb8575d66020c202160a0b3af6a93f98a959439259037e45102ce7fab9160c74f3536861ea864ef34ac2ec2861eec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4df15ddf796133154f6b50611ddefcb9b6bf6b346cf75fe2510bb37155939e88903572a0f473fbe97cbf48014f005ee75f2e999f55ac0d23a3978aef6e36ef3b28653b489e9749f933a0a1e06c05689c24afcab1b8ce46029c15dcbd41464d762abedc8513e807806482de7ea3694aec4a4e1b986315f6cd2eaa3ac63c6b7f9964426c265bb0250e2ed101a62548658aa77702b541c6a098e2700368b0b5c67edfa67dbb2a498808f713068a9e1fdba625d54fc9ef9541bfcc20895ab3863e1d0b09e22210aa97f85b66dd7c610afbf08992fd9d691bd731141e8c72b753d13a5d0d824356a9650ee328d95559975dd3e7ebac9d88e5461e80bc7b436babb70ad59800f6f6ff8901c59caf1dd7876cf620f07912e331fc674fa03f593da7002285d9da1ef9d6a88d9d3c0448ac0cf98a596f0ed4b01d020820b502c114fbcdaa95ff1631bbe9ce13cea75556a24a1e33d345d7c11e829968ca7f17ccea2fd953bed235363d25256149ea2a301ee79d65b851d54ac6977e2ab5238a2e12ef990eb9741a08017d803e68853bd471ed3de93802c673db722379ce0b22d62d417f1e48f436ed1931503c0dcbe8549df059da6897f64a4481f88542ac4928515799b8faa02aebd3c85e0771db60ca6dc36d4523e68c1910140784cdce9d0c9b4d45b0cf58e24ba20a9658f6343d45a77c229dd67d4c53d9cd1ab6e23a83debe6f187ce055499ce12703f292f163d476a97403d32ef5bec942be5ce1fa61b256b893c027ee57127f31a7fa67b26b2da76ef8d4ef2d0974bf3d2dd34df7bbb69d49a77b0a842409b64991d3db068fbc7f72b5a107ee83064e3c405b60f6905c7243fad8fb2f6ea529b88b4b960804897319b1679442e963ed90ff34d84449c8532914415e39203900c977ecdebb5c8c620184aba48c8d2868867caced249c9c05ae43662661de311ee138a366ce784d793794a459df75922ef2404bb1cfe578dd905bb7f737e6376312596a1017ba58608274a3f0380f5e08cd2c5a85241cc029e1de03d5e9707c839c260ae24b72c287ef09345a8640a53eae75a5c5b64833f0c9068d24303c3af6391a79553c4fd5c5336a5f27da304d7d3c8542ae19c4ff3aa76bc3d56662be93f29f1d5e095971630bba4eb549f18d5b90ba3b783b60c7b9aa6b221c80ee1352cc6fa53489221c05254715f5cc8dc69dfdf0f2ac3b0da411bd4189139c3e0d25d730f285ca5bb196a49a54e4b85419fd8d712c9d6dcd04e34d59e1d6a7a9947575ab165878e736b6e13f9143a699974c12b7db934705ddd08e71428dc2420722f74c0f4bbb29cce19752c4f2d078713e056f87bfd1a5b38d0211f9be0799a9e881bf2910e8f086a35022498d183a3fa431eef0b5c9ce7e58f3d21e03011e5fc635fa299bda10ab77949a76832758b1ed2aad982c3f63e86c06725005afa604f06fbad17fc589c93a05f8783403c17e609ff6ed85ce70b37e786c0941f9995c8eee5ef00ceb80104f53c7178830adbbf821605c803b9b40c6a137c198d6ec954b6f94f38f92899cde4aab3ae963ffc0534d6244c114fd9f850e94208948dd23c83866137cc27093a0d9967e2fc251a6adf606709975c5fc5fc52a461e21ac8a9040cedbbe859757be549a7a01d76d371b77ab72f81873b5ffa9c32a605ad751adfc6c835dec614c7429205f47e81f234b153e730c63ea81b3eddc49dfe3b66d08b693c496bbf6d4f9746b677dfd42c2803d5a654abcbe7404f2ae8ac6019de519af2cee2b88b15b9a54dc9937bdc4f8218406559c85dd6f6c573ba4ec85ea9e48640b38e7e83a49f7f42d7b9eb8ec55210b3a77533f2813bfcb7bd288242e8f4b0aff07ee1c680aa70247770e91fa7c6db017d21e8a525701a8a2abc316c1a26c77a926dc43c94b501c9af5533d51f96430a43e5b60048e77f3ad42cfef89bde2e4633bd0314ba7a84d42e0aa19de1ba0390807cff34d9a64e13a30524bc726f24792678c69afc7fcae1669fd2fbf6d68c6ba946bd23103374ebb61f9ddc190d80763a5ffe3a3d61aff5029d833b4cda6d301312001e6c24d07b23960d64c44ece0068cbe7faa2c3a8cab6ae5ea0924e3b4b750025e74cbf1dd98ab261fe2dfad94884e65e495fb987675a2457da0883b8c749126f0d377b1c7f41d68d357e4483e01020a739a1ddfbbf5ef7888953ff98d840366f73ad8319f172bc13f0525622f3496b825d73e288971adac5398779210473edc249010346ab0855b2ec461e498c275b7363d2653a93954dd5cfc2f79524cc2f48e9ebff874a94790e77377ede66f347e2739ab634eeac178370ddbd727549ad2c9d2c079b4c1487fb4a57953e0d9b8a1811fb8d990d4fc202e480ad4e05e84f86cd6e502cd589736bd019b66717fcda8621d38f9d287802cb4f1cc1cbe83a284a551bcda15659cba9c5d15de1e89ae133c94f11f2f1d005875b4f82fd46557480c5d633ea6e51e4854cc18c8abe40ac3ef78460db6235748e12cd28a232da7aa83c0de084039fac7e40f9f0ddd18d456ae3f770e952b25422d3ea8485aaddde7cc1a7c7dbbc52866afb6ca8e6be3533a303ed86f32bba38a3f3f2738faae604154977a4757afeed5d47fb5f5d9c656e6039e5d57574420e9c18f37fabbedb7ca48831a3c6fa1977b3fd7c772e3ccb0ace248c735b3e647ebceb64587d6f6788508303aab178473a06ee60cec442d4ddb43b8bffb41607d1c21a0fdef0ba9aa6cd333e213d2f5154e6cff1c48a41239c6e26ca36a6f1ea101fde251464f892f7ca7ad24ac0020415ab160285223468007ebfeea5aa0aeba445c73d6eb981807f8ee425cd60328040db82c5e805513ef2fe881a756b8f49a50f1c61994181295b9c4a2f5bb59054ef2fd75ba0ba70a23083b1588d131d4633e0d83eb900addcd5e9ba125ef6de94bba53428ffb75ceb2531c980b5f0229f3c3dfac1376addf2039f8854afa681a0ccbc541fad36329906c69a8fda2e9c92e4afb65fd19f729166f019cc01c987bb6cabed1dc0d1f5f0c6419afc711970ecf94715a72226ff517e83556addd185a0b9278ea02191c7b4f0e188348c65fd3a0431e344689faa4c6250f68fa91327261e8fbb7f2ff92e34e3a26419c7ee4677928cd7af84bfacd123eff2088c706672f14f9221321e86faf7b8443d2e568cf2ec12b72b51464471ba2b5af8cf791c82d1e9b14862b897afc9917e72265f958fb310ef94418b0aa57f6701ace72d96ce54808d6411c0e453db687971c3080d064c362cdd6a10d820baf805e6e5255bd9f901fde74a5692f9e6dde666a7eea517ce92d1baddf7939fc7a0ce5256e502cacc8a83a85c8e7f6ba34c9d7d96bfa2e268ee0a95926038740ea032374cfbff967b2ff64c3c53f20e3013438cef5133e6c5e73b82ef77ff82142966f070d198c6bed0893b5a9e518398c06499e4d97f898fb523e3eec1ae141af5db519a8938a4cd617aad3d29842a7fe20dfcd0481b3469e9623586b764c7e53abcda9a33a1bdabb79d5b885878f2863d60c62243cf47aada5ab2a4b09d4c06d88d36cfd8b2ce82ca05cda971c6316e210b55796f135e7fa946176536dbacef0455597c7b1ede6d84d1acb6ae55c422f093be01607d1630ba445b5acdb301d9c068bf520d892c5bbbcda6aebfb72f5346c49b965be83db00f6717263fdd5b3a210bde118014a1f08a80680584264b37b347cfda83783e03a9036327601c86c3a1025f79ad86987818df02ab50efd77fbd25babeacf890a960edd6414f407c928be98b59dfe976e63c8fee78e716bf840e347fb7ae1321ef23339938255f2454e089f0bf923434abce488dd545c7da1e6909999b26dad3be5ea65a2bcac0cf7174a3dfe9017dffbbaaa064186c17488226a81d278e9ef67e38ac7bb04b37d24f70dd428812915b1a6adb8e98b716fad53be724eb34e263b3e20a9af2d87bcead1298a85f83282e49e0d0daa89f00ad748043fe64ddf4b288a5d0d5fe8a6f78550ce4570ac6360857ecf624c67416cbec7b662483983d2bec2713c7d0229bf04fa59001b9cb63d0affd43240c7ebb5e8f8ee4ea7d1a2bcdd552e848c9d40ac61021c0c8094c9316e4b39e59e093836ecc956b7f3b08378ee556ce65e306c00f96d1a4e2a65a91d8923ab777fc3c939ee07a02a2e3e403d2c89e27164c45ac0ff6c5789965ea26ce674e44ab7ab5d49464ecdbae895cf33e8c5b93e0d7eec9676577359290738fbd90efd6d047360f951980f9b2d5991d9785537fa88f2e24ce9ef512c47be0ba76fd95153a9b775ba4637763bc65dd7737a6e5e5ecc1452b77801369179a266acc9e39dbbd9a31085c58add3ff507c2ec33a7dcb37db5ba31fa45300ed86dd52ec4af5fdba121232428b95fc990b737fd6165978ae44e377936a5eb13eff2736571c692e831716ffcdfb2607b96de918a2a6357bf08dbbc8a6ccfce1c1510501d4beb7d5aae4dfc57f72d02a0a0e9d69f92b125c7f33d823351e5939a07fd0993ca35dfca5a7a718c8be1345e6035b34f78e7110b181df414f5739642c572dc018cad9cba11032ad5cca2958cdf08a5b16b416b0bef133015e36506e08f001b05db62bf46d1363d2ed0edb456254ed0cb8ae43ccfefbe7a76dd3b23834f926808afda2bd7182d31e53131c1314297089b5d30d15bee814b4113c29c8b58783301fca3468b24fb51467e37e944918186966564a5e93ab04f4786e37ef9e8ca54d735b6e4ca636e5d7bddeed8933161cf8fda27d923b7d31d2f3fa788543e223a3b66581a2d448f82dda7569fb7f849668c2995d3eb9a34e98fb0036f38a2cf4aca70e679f2b9598f581aadbd7a73b32123b5bb77dac3cd45518c67a030b27849882911be2e7277f510250e268731571b0b2c7cbf91d4949320beebdb2c4cbd51743cd9e0aadd7c690cbad8e370ee8b6b45c78858d21dbe1ce9f16a068d6f06ff30ba17c59f9c078859c3f69049e9fbaf3dc6bc2ae211426300aa3d0cdadad535377dcba3ed22ce1a96aa826544972190901aabe7c8cb035390d9d68e5dc3d92902bc9768e61bc47e5abfc800db0c60ddb08eaf28bb8495409a034ca657d4c124cd42323c5bec6fb49b0ccd169edd7908375fbf998c64e8ac646fcfbbb59f58fc29e45acb9be712c23f43e62534c380a4ee1faebe7b555754d57eecf1b0b64cc1815941fcdddd0f0cb12968a0f4f99caeb8b5b59fc88f86b5990f59d841dc98b4672f68b17d78ee7d523cba52d372afc1a33862cbb380de802512bff38d0128606f9586c182f474ed43423d3ce90479610c6d0bf52bada38207feaa86f24c07c8eee2e0d0e3f5b518cfc27548442cc8b4b892adee4e1bd5cee48c52bdf0d6d6a69f255f8527fdabbeb0bf541d7595bb59423b5c9730106e033c5287884f15837abd790e6e4100c950f0f561c05857f6b7275379d63342e8aeb63a4b83cbc06d68cc4e21d6376c62e40c0ab5fe93bcfadbfdab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h89f495991d6ec5292662290e3d30492dd90fcd30af7a5637002ac55cd6fa9867a5d8ee83deb80b0a8fb22e4cbb0b46de8cd82c6632c3aeee36f767f7c5d694666195cafd80b6f899baf9b990cb62cda5f0cee78d87b0d7ac6639ffec0f92ad6c20e33775970ecb6317a2bdc6a12f141e052fc0d56c222f27d37dddcb98767eb3c87a6072618776c2d85332b0a8bddd0340bb97bf6edba57d14840b809be5a70ca1adabbe4058b672d11bc5445daead57b11e3b7fa80d3eeeeb09a82c65e21af2f1e4d87bb5366c5f9268484930c98fd92140b0ba143695ebf0b5a7fd82bd1f26ae2759434b4b1e792a0d46d7c5651707bb9eeb96f15d3ab8aebfa0918e8014b3a83d6232f31d0e0a290a83d81144eb16cbba8d352919694236003e15841adab8b597d5e64cbeb147daa54ee52c3e35207a0ed2e7812da4d5c030fe80e7c775332e1447a9981784577a45c071295238025b796e3782b87a6d7781c5f2a5c852608fba265acd97d87659c013bcaa4718a0fe0177f15c8bc2c5658310a22ae7154c556cb4d10dc2ba278f9515a3142942ee04d8b4ef4623e8e56650db3a276c262609cb9ed3eb2b7965591009721efb1496dae0f4290d8203c7964c30178357a37a98f947e443e86cec7016666569459a122975b6f47282cebdd7dbf5010c194f17f9ea9dad73c961ab325106a64f047abc485b7d36f287b19bd357c85e1900b0f1c977128cfe2d32454842be7f6f56b67f17cf8abe911c40895eb8bb0d01c3a40dc77b9941134caadd822e0881a671ee40d2522037d02eb786d301f5a4990806a5976d1c8cbd5bba4a766ccd91fa9ed46016a3bfac3b6b667ac4005f15a681a905adbb0a2a41b7209ce466f3803d2e40e31245f0088ae4f784a0f26310f3a769c13b56aa0f9ed99757c41111114496404ad93e7c234724e5a77ccd5895fda3d7ce5f4b1684c9beed84eb16a7b78330eb5a2ae68ab3fd7dd55824c317d205ac856e00d6b5720dd5d19da130fdc8c7533beff2876d216f123e07ddae00a3d547098e22d199be0ccea72acb6db30246850fb55d3613dcbd54fba8ee2b5fa2ccf2f93e1c12fed897e99728bcba6f72e61730ec80b240603350825d8609e6a8724aad5b0305f909eb7deb915780993d0a62bb44bf6ca92580a0684c1b0b64720a3525353174d2a0bd0a8380e91bded66977aaaba763e092396383692b6538db9a796d487722550948933a184ddce8fdddc3a04b7456e15d524ef9524d01ad122394d0a3be7f91353e11dfb9845d4b100d1abf9950468ff0ac0c4e959cb38299b5dc5af390c30e8ac21d951f431deab4d8a073569b8d73383c3413ed53aeb873c19c9d456ac34d3928be58d2cc1ecc8ebf6253a20ce4f9ea7613b4b8a24d6f3b6a056450f70eaf7bd3db93764888cf691552edbf19c742aaac9a4504f77ea3e4ae4cb671686b836e084bbef11e31d21844174cf714dec88692e3a4569b7d51df92bb078f56a09ee4c36b64477f095ef0e0295b7cef8cf503b74e1984373160d1ec979440b3188510fe612f707532300067ea59c3d95164120d0500b8100ba9455dde4cf36c1e929dfeed44879c54dfecd929b4d8e20016d1a2761cf1ca03d46b727a76a7b5439a9c989cd64fb2b80d56931c335f27d22c42d8da286348361a288cce473a22ef90f28875c53616226de2abbabdd82e9699c365f5d73a19fb3baa1224281ea59d9bd2a82ede4ec05fb1302813fd785483696c8434cdbfd83acab4a90b36f84e4869f3ad3cb35db3a5b1e8dfeff8448a47223a49d6227190b4abefab0fb408a4b9c0dbdbaf681131a735ea9e29c1225d6871a55e62b6480232d17f71ce793103fb3409f455bb054400eea1ed71aaebaed39bab991564e6d41c465b6a67ecda9168bad4f20026a9f37ecca86596963ebc958bc8d539e1d52c80146988a48e9623ffc3b8bd2b90b02bb64f6f341307b5292b6ff716e78c487fd275e040b18ca92f1c4eaba0d1b49fa95a542451612a9b1b44315ce12aa0bcdb824882d2b08637227aea0dde2828480fa63b8959c623b0f184ca629e883c1323a9ffcf0be6f4e4a732c8f4a136a24e61bcc429f7cefae53c459fc3148ba6706a064c5e4fab2291a660c185c737754a6f5de4decd222bf502fc26d4ae03af01bb9e2761865fd47cb297e6146293dce653ec486f44e1ce357bde29e31e6c2e586a84dd5315476bbcdda1c61dae371812b25866294b950f965514474178cc3c3125d39eccce61cc10a8be0fc1c9c5e4d4bcd8c25f9449d8afbbcf191fd7ce6da09c5dac04631a36c6cf323027892c31ad0f34f2d0c5f5851b7e43012abd1126fb6a22bc3e5055c3e1cc4214bb1ef79c9429c7ac7909a92febd904f45c0c9b38a600ff01939e451da3ba29286bf0c8b71266fe4c571b7ff37fd5e90c3069433964d4c26a4b1bb61349cd7c07930fe5cebd82cbcc8a3790b00e5ce77084d83b54b0812383eba34b0c5f7a27d8855ee2fb683b7bc36ff6b1916e53c76d35682eefb81f1fdcf952857a1b97db27837939c3ec51d506c6e3085078d1b951741d79a55746239c02823644ccde50fe857c247e4717dc6eacd08179bf9e75001efc6475d895f4ae4b85ffc6130926217b1365ad19527d1e012dfcde44dece05fd792fde350f827fa3866855134ced27e3dbc1c794ea1a1e3a63606530b1ecb529a2d5fa6136fa75455d336641dfed02a0dfd49e7f589f5e94d47f2d3f9ebcb09701e8353c90a6d31f0d710f68c2d96df1901c476443fb1211a89af3561dfd6f9e4499eea31e1c543768789e19d7dfae3f199dd9779342fdc84e216212f68bffa41d8f66efde374f03128c48d0c75c4c6c57aba872b350953eb5d264ec46c0c58cf27e157ef133af33ee37a2e531a8161e87c6af90a5b1f97bdfc96640b85e18f027150d02d658074c2699c870a618c1a06c54b2560eedde81c9f198402c4f17a901594030d665d457f952cd5b5583353043d645946bd1d01f68f8c139eaf9b25dc8d8dd5018c06c0c0ef301f940ecde6f62330ad35a2e49c63f795dc05197f69277754c5fe048b22bdacffbab12d88396e63bab2f9f17b0fc962d1e953303ee5c530f4943f05f1f5da0eee8c4598b0876b53dbf58422a9f78a8d217aa274bb402ccc63ffe6f71a13a893b0d6c17c242a4cd1f14defe70ee3c783bbc722802fdd6a1483524a725025d299c4538e47f693b628d3907f2d434605fa6584438d913f6ca93b2ef44c7bac1dc8bf616ebd5a0a9ce58f613f685938b81ca5d4a61625ddd36f9d44147704df9e7a26475b178085ed3a1e89cce83aa48eaf43a394eeb432b92099b81c485cd8dacaf0cad1cc19e1306871a6ce9a5bb13285f28e23f09794f69b0962edfb83de91d41065e6a742bd5e9a90f204384a9ee6fd4c5c7264924c7c73f7fca5f0d2d33b2204b559659ccdfd9f59da9e168798932b147945e8e04c433d59dd55a155cf5d34eb6745050fc3ea1160b57c137bb6dbe7cc7847b9afb29f497f9c453967572c8f5fcd90525c27c1ac88c338277373577961499ad1335f1681011985f23710edb7f38c96233526153fb156dbcf8452597fb131a8100fbfd023042e2cece1c067f99a0a37956b91a04450c2663ff38d4dd7d960085f3731e2a7108ca3f61c8cc19650b157b9ad2036429bd12ac3a6640e1799bb5e6dedb930baada850c22406f5a80939cc826053e146b470f6dcd33aaeed2a1c76af711a0bec2a349e64bfb1c8c0ca2d7373f3fd4232f53e0084c6ec3ce18f92f6691d853832445574e968c29ebb7c91a45de675e16b0f1f80f0b950856b4da626cbb32c5d43a7f441487fb405831aebcb21ff060a56d82b910bad757b1465953d528979ef07498b1e34d1d97e1c6a6ba7f44caa6586b7284bb24e19f57fb70dbef01045a881652eb54d6818e9549a8aad5c93c7da5acadef45b30e085150c5a1323da8ca4a902eb749a5e8a31dc842c12094cd8bc67764ab2cd97e6f07121a62f225bcde303a8c0e607d47396875058ae3dd57065ce3d73ac3113822f7b0498b674273f468008c70b70170bebacc82f75f0d0012fff98253dcf188125de3ad4e4c0c7124e0a76846f885c618e6d5528a5b8141013979c76718feb6d79d9fffd0edbacd2f4a0024da192e39fbdbdc89674c82ba4462425df49936714ad9b00440b2b444198318575d673b7a7abdc11f3dc9d4e3bd4eef57bcaf20c41a2392adbd35d2ac4ae92cda8a6777cbda29dd47c11670b21ac238403d95a54a78d83ffc3180f2969571c19b334713b0feadd6285b134c3d48aef277ca931c3cb47c576069e22faf7324fc7c70436aab0abc047190c776f0c0d815eb2717be06cc7f289127316c57b3e41cfe2369804d3856297ceafc8c88969d82a3508c9de6688366503da5be9e7702d974ebadca800ae57bfee3ef8b45895c5fb5a8ce0a64ab99566e57d190a5d3f70c6c30fc4be2a1d978af143e681cd639910005519c863b3368715f244fff40bbcf7d7d7a23c7c249971a03eef692a66c2b53a4304126c1524e6b12403874df802e4257700626966ad75bffdda9612c655c0809233ddb8b41f03424d74f81fe914d5bd0e8a78b2ef2ef4d800b24a8d6172e2a73c34060db0db0cd1115081e81c33fc149eddd5235344b1e50fdae8cf1f0c869f31c508ac8700c0325e1270a0aeb1ef6bdf90a4ad0ca3a672103b20e0143bc552184cfb50b0500fa5cc6e37d509909496701348c90e1c173f7c8030a620f8bc583cf6c2a501d52b322e2f834440af756cf61e49f01a5fb95df2640a34c33e0f576c775e164f8d561754de82ae6c542a0347bda7c4862d7146df3f8c05a0436b17a12f1d0ad27a03c1497b5eb5a22ce5a03c60ca5e8483da56bc7b5a098d6235a7523ebd21a34434ba405b9da2707c6c7fbfb050089a01ec53514afc91d5e3013b275b64edf5c29cd343d2240bac3e06e9a1c841f115e7945368f102f727fc10c54e653ac1cbe8fada9341afc476604d2c64309fa4de478a5e7aff3481742703d6020efc8a4246affd4653e3e6223f5e56620421dea453fe956c23c1c409a891c314108522c6ed9f5cf2a33d71b149e7f99f03392d0169b8723f3d801e544eec899e0b87275e5208d2905844551f3f4676893e97a27f6d8e8d8e2a8dd26cdb0c2120d096854ab14e116ae3334eb61e738347012be71206bfe627c329a3da3ca70eaacc63ec1eb34119ea3fc04c29faac780f4c389c8501f16f1ff7f0701d00d4a13dea34da96aaf0c2be075fc4353a7a823c26fa766262bc1e6e641ce492ec0f2a51b480fde8cc78b5702794e573788d4242d72ea39f2009145ea2f20478ce6683f191c0c905d695bdbd0b78b24035e671f27a96c0bb129b40adc5c801624a385f460f09f1f13bee086b92856252392e06eae9807e1249082c01b58c5baec7e030e25cd0b6c4e3176e8e5a06805054576985dcb3527325e8cd108cb7c466564b8d88549a2516ba95a79;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3e49cd4567a987b2dc4c7371e034f8a03e013088e44884e6b6b6354a150b3051b4eb6a4ddcd2636e148a57c7c39630c830d8588aeed064d95c4e4138cf96bd1254fcd96aa30afec211db95b2c88bd3b3a129ba9dfa04c3409b7c7465d33bfdd673127c65e83336c00745fbc8d8e3f9cbc74763335b331c73019627a0a78721b1f2bf02161e5804da869cce78168a020f5ea7fc0458afabeceb4fb409e664d9735fca1b25cd848af4afda78cfd4dbb695c042543442262f0f7ff0af541ed88c10474bd5710e41fbe8680483a4d0e7330e7582ad06c243ca40078471995a77175f7eafd91b38ea7f4d4ea45eb6d50339e80b5bb39c7830ef1d466927fb9e7711d298048cbc3cb3d9c2953dd13a10162b1f6b66f5ff9c65f0658f04792028964ad0d5c7acabe516c6b64a962742114e1b28519496ac29acd3e336685cffa5bbd057fec5b71e0780db7557849f76d92e96dabeb8f155a46d4ebb2ccd8d35494df79d355b3b407b38499198d917cc927d6ed770629b93de6f9875bc60831532b9d1ed885a53652e5f9445bd5e6761a77b31dd31504c81b0f07e270f62173a33c8645076b00c5a2e82b40c3a07e8d0fc8f2f383182a536f16921dd823e5c7cf742ffa5b990db76bcb8055825d3da74dbaa1d13dad64af713641ab80de984ff4dd0814ebda2b02e465b14c9074c2d83da8b039d768ffe497654298945b89873e2a77aa717c6075d270a84ac1aa6a9bb0cf4b178c77e519a33adb7100b94e6298541b8886b8d1299b3108d5d9bbb71400840484aaff6889d6b91503b7eb906ab9db42fb92b4f8dfe0886d782dd5553e5f14752b33dbb09fa2feca3853a6cda05586b8431ea61e3a19c6577faac2f2cd0ff7791217d25899ad32cc17df2ce5161c34d410cbfdfa74d0e6d8c68981de3b18e2ea94ceb63558de2c5b7af94cc36ffd5930137485036563ff032e6e6ce874c3c98051e62e4c3cea1af7f3940b1c0c38b201d46c609708d6861702af6177431f2cc986a6282d3d484446cd66e2c5e871b89b802c141cbad0d7bd455d5c4689d31d5d742ce8e37376bc692e532dbbfc9300a5f5512a6b3bf9ce5b06a85585ab968d6a651a95afc17b2b86e18e84cb4687e62c67af440678914903fea0e02ae7030b79ed37415e661ee2f9ac52c15e13d39947d4c216530c75ca115ecf51708d086c9817cd873a1775b1554d73c58c58384ffef8f20593b1a46b7796c360101083dd5858540df69ba536f57e1f894d2cbfd5fc57c7aac18570b5b7eaa0f2a83d75b89279e2d48fb64541c4a3aea25b1b0274f990ae6ce9f8a391e91b049fd059f22163abb2c16d392eca409a7ab6dee1deccea4546012cae18eb732ff5d20f421418272799da52b0e8bbc7c4f23d9c3651e64956218e3561068ce5a60070eded3f791bf4da324d861fd1b341679c4f6ad1f7195d0f55ae3ae67f300d3357028fac03d8fbda04a33201e3a1b84274e5cd670067d84d12fe87743fc20034525712f5e44e3190d3ad31c68197f76a7bb65465653807bbfdf4b594e5f644079a529477609b8372ae82077aed9b72e6a686eb0ae65c5af2fbde9b507f62a122d7cab734f607d759462e629f3128c65da7255487f1d0b02fb366c332ca6ab8a33adb0af6b2052aca15a72ed6ad601a36409dbf636da5afed22c634b356752b7be4bb9562d07c89231b787f14489d23e17c89b564e8a5c6040a82dea8f5394dede4f0910e1554019062ac5905023486e1811f41b256b2670f3f846e56c967a828697d4e2f3410838fac96a516fb763ef31b88e930a9953e688c7a5a8ca8c684272667700d3eff74ff5d9cf82b69fc876468a5ddcb50a2e0a98d5c690251def4defa5bad82549bd435a16ed2627cfeabd04a626a4f3c0211502e652df5871c829afed98a71d887c145dbec0235cb2ea5f293a7cef5e7334a06f17d5918296db77945e4dd5879baba8e8f44fe21b8f7400f2f86abb10144832d1379374b3cd1a98052ec5eae527323c6f9d013caf06ef7910f41170da486f5514aebf49f5e239de698fc4803adddc7fb6e5994fc6c9b2e11d904b71dc5dce86a3ff517eeae4d6bf688395cc98a62263e8953651930d33dab5c88435ed58393bca7ece1d3849a8233c8119dc55b89d48e2a64dbaf170c33877b8193f01a7f902e08928dc6f0cce43f88bd10f73c0e8bea5c084d4ebba4c98f4b2e36a873ac5e2643553937a34cfb8e7b43aa1717b88fa863dc8678656951fc68c18c6b8da2e04a6dc662ef88c6f57db97fa6abb0bbc1fd01eaefcc1aa6a3df0d64b4f1e326bcfce9afa603df5cf0a7a21c159a4f9446e88e26b77385ef3589c3533099c29f928118d0cf7be96adcf943cb7b9f9108944a946bacb01d988e10c8701fa404bbc78bf5a5f76916e1a1143c32d5f0fd4981e207fa45c12136e42df6b7b2ff033f474eff80597485d73033c6096735376752d003d75e337db87627d3e63dc53369013115cdf27a4410299037c8ecbb7076fe2ae2a6c55efe81e39287beab383ccc0798abe273e1effd082846e3dc3dd9b1b4c4202916db44d223265689eb78da66d86f87fe95303765b4c04d53de320439e954215846745fa850be696a31d08596b525a11fc219a1d6f1e29b45d67e4abdedd6ef30edd4655f3914ec537b785fe66e531d994f9a243826c936afc15349967877e150054ac124a8365139446360dd5f8401a189b954ece39cf27dd37ffb7a2c309ab764edb0d05578d55fa397adee8dbb18068298878740dc0bfe2aeefe4ef5912609b25a28fd95c58f471430ffd08436db938986dc11674d341535866a1909776bd44382944a34eec5e6b0a350374d5d6d60e5e9d18f54379fbd125cdb57fe1d278475296c364c223e4a26000349456a9da8e89af85dd27272ca8099ad24872449a9af7758bc2232400e417c1fd4de5a12de98171c09b71659980468d7c6798c512194efb8b9602535321f08064d46ecd001ccf869524915befa12713c010b4d3438d195c9b3e445445fbb43c06dd41a3e3adff34786ee1a57a46d1f9b8c9fbad6b179377669877207dacb0a97b69fd6f313d822ff5a6f1258b85881db11ac61318966cfc905929c8c974a8719cee40d86cd70c395a7061bfa310a047e855767ca45e5158e6c811f7d2e84ac0abfec91fa9eb191c248ae1c27678cb4f2499669e00e8848fe61ead875c25d5026ab06449c6ad768b9a9c3e2d747d4f2f8529d196912df3908a47c8572d1003891db697683da66a971351336bc8fe3548fb80cc89cada209d47628940287dcbd77d182f24f5cf29c29ace182e27651ce4c5ed83ca675278d6e5b8f24aced19dac443a429fde92edd3c960e2de898f69f37d120013653f68dfbc6d158d4e4c39cbf9d53b08566248a9b5b8852e5d56aaf3d340a8ee4936c9a0446eeb10e76a81e72ffd5212372b77a283c90e8109b3f10a11b9284163774ee85252b1c4670af2c33f473231d232f119694cb64da8683db440df8fa7db7d949fb7633d7b5c1945527fd8c9115fd198cd99bdcb5195705eba9e4397373710c535f2704f165e33f0d05217074341404a1fb22c3afb7ddc09b91481e0f39daf7666dd0dd76ea1390682c534a8addd7c381f2c9a91f1866a65f1d614ac6cc04a70fdb873bc178542638a6bee8a2f1b930e22012393a6b4ccf37f84172e0ca20bb59ce0b0ece588900f046ceb1e438d398da5ed9fd13fd40224704f2043b2ae945dc7e60ca625cf806b50145c290a69f107f6c9fbb28b1b3751148dadb5eefea56ea5723f303793fcf46111abfad034c3746895cacd0a451e390e3d8cbd8255f8139f91e0d90e29aa562263c1a240d455aa2207497c19caa08a4d27535781146f09012e8cdc346b920ce802c5205c07de2a9b867834a2f27a73081718d9f7cf848bb40cac1df2d84246255c34c4d15f541ba862df7c2083501ffdb72e7bf4c6de339add01e812a3315d8c64c24d3e9e3938389bd245f66012840c57b136b7a02d9e01e48d280fcf4873c52aceb64a59ce7c2627016aec1b9bed45ca94f76045d8ec93e121a1f572e97a01d926793e6af7d69b827dbc186a5761286894202cc2b7dea924448a9829e62c0fb248312c056b0cd80aa7bd8274dd303773573be62da45ad25ad0886ee250eae492267e5b80b506bc93e35073cf9dd1bb50ea280b90701cecbf73926931173d4f9d5265009902b40df7ee08706f83fdc0df368d1717828fde9d3b4bc73e7482601e52b504fb1fd5a4c937759a8e03a0410ee1474f7d6a7ffb9394b194a1734d77b31a88f7d79f3808dab1df62ddbcbbd0c6f0d32da237d4dc4d5e944790440607e68724d4e5d5160efbaeff24dba77c28f9195e336c5d233043a1dc40134aaa256c30e41ea2bc482a41c0eed2c4aaf8973c42bf62639a082e404a27263ca578c11a392f9b5fd26ab07f8b9fc9fc9a7d9d3fc8bd6f4273c3fd3dc33c98b4d313aa65a955052a393c0fe0e6939033d8a5ecfd4c34928f3d2654e50d0ff438399e8be0344f65a4d269795f39033fa78b2e1ac7fb5ef9ced462ef69caad890732b17b1e790fbe8030ba7a201fdd34f04349d51d32aa9797a4644d9d83df66edfb797a2e0c26e0de7e243288f141f4ae18462edc54600aa6740488a5f34b9a4c449b726becff5417319e18c2d94f0c84572494705b2471cee22ec6dd0f6e02db9632fa9f856827a7ac2b5d7de85da4c02b1803bd7596aa66194eb9f89755ccb17177db527f0b730058fc7d8be5664ba01f52f802ec9c9b28801d726438bef832e378064c863f0f47e9f357873318e477453f71d25b54bde0ad8909fb0baf80389082d8c18c5b9121c0f0958f3349c633e2015e7d27399de53c2f8d6be2e44639685411447c75aff9f38bd391bcacd8b34201bd2ac1b09a01015fca9a1bf9b8bbe9d44e486f80f15762c3e5df57d820395f4b8c474225533939c63816bbe8fb8a3587597f2061b10a7d546a4b67e57b4d6afd165385a902511080799969d8fa13580d927dceb4c39daf657f7e46fefe73ea707581403deae156a7764f55d8d17050811afeaf0fd7a029687c4792f2c120100b8c9add17941efbf28d1bc4184390bb3ea990c6db7a396edbf1a6c74775fac6053551aa120c6d12b4d75e6ee042d5f93a590735a3f3fd7b89c21b141e5510cf30a45da5c7c2bb5d16aab1b355a1dfdc264f95d579178e0a2bb753120e4b1f8c29dffbc0ba9d528e61dbab914b9a42af3e40b0c324171138d0b93c600c584e31d26be50fdf93417712ab748a0e2115cb9df12ccec5b1f0fca0f8b9d56ed34cb44eb797207693f3b3f6b52e0328013f111b712f9b2ddab76dbadf5fdf6d91b067a2ac5879b03f07a7df0f1cae5582c13ba35134960c11b25b9b3ba94acb2dd8e328881e088752a35140d752e38cf4faa5d90d19fbd4dd32a42ecda844690d2beeb15ace6b56065f966c8b3a282f5204945cad01938835afebe00b535f16e06ba5970bca28ff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h273593e49957d56b21db0204bc2d6c239288476e7cf386930f6c2da6c80539bea48d3051de1fc045c8f162c81414167e0c28961f64b95e2b6d3d3aa26ab33837cd6c6e9845503587654daf77b51dc3bbbc78e3531b98ffc29b155356c30ca219d9a00991437d7e973f3c4aaf29b940ee56062e27149701d9caa5600e657588e33dc28f06aefa641a555dc7d7eb073f396ef5ba0604f6a323b914027ce82504df9e51c86765fe63cec552df82e523ec0f780cedea4a2908743dc3ec3f8564ca5cda949d97de7bbcc6c9a310b5cda1bd1a882c52471cb0e4bec9577595fb4132ad20d938fbde9ca1e69a8bb21a695b8c50b1f29c01e515e7a17740bf57d2b5025912c4da5a8364b101f1ca7dc629b0cf92f58bfacd3404af53f7f3244ec4051460605004680725ad2e45e9042f1ebde7411bb73c9e4f39a61ff080fff00fd3ac63a19cedd060ea2fc854fef3f7d6ecffd94e82cba8ad9411bdf4934c1f8e9f505f2d4644639094572f14fa09117e182434602bc1b2d5c941b6383cf0aa4cf13d0d1c5fb194ef785f916c128f578b7a5ce36261fe1e0d0d01635a6e8ca567b0e6814803b5138ac2d331c852cd007a88c3d8465d9f9826f06d31921a6735aa63288b73b8df2b0ee407c7fa8b049abb4c2abdf758234ae41485f3f4e91689328bfe5a71fe4677a11e36fde94e9650c5a3f32d1b8dfc8f51cbe0c49803bcd375a1cb644d29131633b2f1764ddf98d2014f6c9849e96a1376b62135f6368fba88d5fc5fa0cc70b985ceb6d94887a73248f739ca2822bf2d5372d1b50fbfce45f60ee8288d9f2d8c16f9eb5aabc1238ad309ca1df4662a587c7ac3a96be1107e115f5db59cbe945f855500dac0b9c1e1c9141e542f5236b320d53bda43aa911288ceaf2df4e9e367e6e21df2da3024a05f5aee64a6eb1e7861464738ed5c0ab56763550e0f2bc9d44dfa664998c70db199d603598508d5ecdac43e2d1ce6a01fe2a7c826f29cdbb00b5ef3cb1fdf3c81a9fdbe60daec2abd0b16dfe1cf0ca62daffe44e958c718142ce04547f9b6057f16514e59b308f1e3f8ad1c8bed27e438bbb34aa87a0c0079617b119b8d7ce949dbafef6346eef4780daa11f5f95d730984a491bc196fa6dd638880fcdac412ec7d77f16ca223f3e65dad742d50b6f1afc6081a5d57ee1166a9f1202975f39a64ffc13a5e6f98db40ffe8c16533dd176d4256d1413af75f4419c293be2443e90b8ac536123010dcaa405d9435e14905ceb499919cd49eed14bbdd8c783b110f5712bfb03deb7d10018faa19be2128800e23d57c9390f68715d2bfdc2c4ce590eefd27a423992c6f4cc2cbdc0c02156bd05ebc2798039c2ae1d1c991732dc7f0d7fb6df633eeb589dd2f7406f58d2e5c1b0e9ead86dc05b1c7df706393a9f2ea5601e1f1ea6646bc383f91b9137e386a1d573592dff786cacbf4775d3333e50f40f31b34b759abf6562279e251fc81c96538ecfd414fea3c9713bfa0fc77fce9698d3ed0f18ea187ea62a0aa3929d5bd26ca4c22af2b1c5608997f5f4b862c33590c13824efc8f4771e9c4fa55da5fc4986dc102bcaf0af25f67ae66fb277e2f211c5b5357bf1bbea6249fa80bbeca6681c1b3b6d1a7bf7c688a716e23a0b8d5fafd206d7cc1ee538a46e5662548786c7a528507bb5639d6a9a3afee99ef0071925cc607b2c1c5ed32f759dfacc3a2e4f712fb5becc3bb885d891020e07979f93c9583754cecc78f78d81aefa6572054b0cc2b91862e4178bb2659ec5e6abadaef69fadc3afb3df167cf8ac1fd74489586b4afa7f94e07f2398bdd6c36922f7444272d47c6290400bf798b5da6d44f9c8252878a500eda6f5dabda52070c66fc06717ba0c4eea5b6c03d85b63611856b97ccc63818b9501bfd17cf891d8a2fe289a2ee5dd3b3f3303648bf9e88af41cd195227d3bc6328e3d1b9ee61c532f7bbcce09e329195b908065a811605aa17014419f598663aa6b696b1a429596c26edbf23f9c64793194c197fb5c9ade9e686a8248bd0ca5a232a95df8da3b12c4d131e57a241d5c5ea3c153269d3ed33e01c4e2e1b47daeb3da502aeefb8556366510deab287e63078fbb956205ca618130bb94e1672f6d0219184fe5767296d4e5f232b760de23c0ff48000740efb16e5d1b386537d822fb64b254d5b446724a41c275ffee5104407127cf7ce87418c6bc9e8516b4bbbf1ffd44145e4282b7ba42ed78093a6bcda355eafbfb4e59864e6acea36ff019ae702821c80ebb088dd7a28add298bf5d443e0ef11597b6e44e8b7313f76c723427de5749adfcdc27fcdab10588f5f842041a8567fb435ded1a56e5e52d008ac924ed86d254891f9fdeb774021ce41c96ff23bdb0517a70335ec7cbfca259189a4d12d822c646a57b8936243488527b617459eb18fbe94536412d009a75ac16206b9f6b5e2a6968e511502a66d463a5bdb7a510ecd3e10f63dda8cae4e58adf271ec15fd80c0f6d22a490e158ac27f3527552606630860c367bc515a0bc883ce1edd0b1c872c84917c0dd9fb074052dffa260bfb35cc559de713a557cdaa45db62cf2f59af33b1246a52bb2330378b79e60a0ee860cc6b1ea90fc80f099a8af555125b89cd3da094a25235cd29726d9079f9b038d21283f62132acd137a1cf194d389cd1ce42f1b8ce5b97975420fec3cb0f23ac9bf1ed8c3f2331615504775d11e46efbe564f0166189b01ff5096c4019ee71e860d1a3163f281deb390b3d38ad75942f346606092729fa2c2edec99cf4922c64ac1f8fa808fa7888fe8cb6d410385ed9dbac190afbe9892043190af6d9e39955d0c8abe926fcbf70ea1f92bd17e68870f84919011e7f13cf900efcc18bad7a0c0087f34257705f1bd6e32854674102f605192143df8affd2b3cd7dde0ff9ca8fbeea3be1a72bfa24fbe32ad69cfa811c39c4fbb43180d02f7352bf79cc1a0affdbd2629a3dd9f245c6db4bac3c648a7233577f216b2cf1f4820f167ffc40de00ec01e4baaa4be673a184ef5f490f9cd258d259e0271f288d9a945432033700c626f763b76525d5da546ba61fdd4f9e237f2a374cb021762e27ec92db5381bf4eb4f01cd627393da792d605432425a45e4a8f67f0781c452450208cbfdea886fbadc7c00a9d29e7decb944da66e47488d6511445a08cb90425a04e694f717b7cd400ffcb0bbbef41ea0d5ebd0aa70e3c83754941e1695afd1708dd299d690065dfb48a1139b1387eda11d547f50feefd6a3476f8f86fa663a3a4392ebdd1106011d5f46f15f9b41be401e5a70493540292e268a3f1f6a71a0a55e02a4403d21555f8dc53d848ebfdf30b1bb2fd6bd33aa0bf8b1d663d4ff308ac76aafa6376c3bdce79b0f7f24fbf4fed5ad1232de59e056b005673c43fa615d1119195a4ac820a8977b9331563df092a291b2a7d52c7aab081dd7b6d7919b3e7d94f56e39f06b081d368817f4acb946a6473a2a0699df7ec4b6b5e144616c8d76b402606c03d6a795a8bd23e152d27b4b08046b5b936bcfac476e2271306290e6f75f55a8723ab7f7edb11719a5584595e0a6119a8b3f46a4adb343c69d74d260823ca2e46d98f117d5caa22ca8ad1165076f62569841ba37f9ed7fdf0451336ae217f81a20e9e6a34f81fb5614981eddc7e91ce99c46084e1ef320e75d49f07b7b9be38aff98cc512e573d5136072678c30c25c52e115c3313961b1a533181ab42b353b5eec2f8808e37c258ca4c20ea7820dbd1962a432dd8d1321e39c55cf4fac646e4727f8927f0823ab128179bc1ab2c073ee7af83552c190caeec3706a524993bd4d2270007269a1e7c595d356f0ad80fd592835ca92b8ba67069fb12f72176ed37d821abe35f2d69e0520fd974f6c7d3c01ba749b3ce296a164fe45bdc24f328d1051a0de33080c245b564e39bc16b590131e62a9765522d593ec85a989b113445ed2f2f43f3ed0d9822ea0dec33da7e7b7469f6792b6190fd8c5d48cebef17027bd2485b78872e30e3db526b2e810f0f8eab93b3f511a9b8f01157dd6b7193e18353bf9ed1164aff68c30eed5c73778f28bf929ecda1b9f1f8ca1a3beec600b727785cf1ef71e0788526d1690e5462f0575cf0b7de18547cadc30791544e138f21618b9a9e593ee4a2142fcb3f0ebadcbe077f1de4b24fb9bb833f6957c91665ab8797723c25b35c0de52a9a69bfe2a686561a9d42e73d85d7834ee5adf0bdb111f54940a3c7f1c595b922113c00a203122259703ccfdbfb5ec6ea7c06541b4aacdbb1d45019dfc567eca39478cc7f6df057d78fc726082d16ccfa451253a1cc01df6af7af89739d83debabaf8e9fbaa0cd80059bd3fea76525b56998d721dfea584ee8243b4fc24a7220424e15894c9ce3f50d2f1e2e4eed1eaa92b2a303b69e79424cb239f485de38e76b0b87c6379a6200fa73928e83623ab0ed61b7ce2124b4b01d0a2647a0d27da8782cf409ae69d938a804fd3f79abace6a1424740db3f83354b494520c179c6b0a9995668f092a379c6e77ba7a427f60f684951fcef86b901e2b4dffb6142c6f54d358bd4faeb7679f64814965ac99bb7c2fb912ab5e8b853b329e672f3eafa878ecac10b6d862a85f816d0cb5a267da3759ac7de4a2a61a7675d41e1c93b7d00068de51ca70e05010c5a9276037686937970b5caba78f7411b4676bd7085169d0b3048590a994e5fe9ea8deaab1fafc3d71c4b1b3748899e5334e9fa0f35436b5817b6225daf5266104b9b01276d7a36dbc50c1c4beee1bb39252bdd4b6e6b3cf31ba95f5fead0dc64efd8c6d10e19f73bc0555a0aa5e9b6352e31933b0be2a19153a4d828b230fbd4b3701fe185859521920b62bf2fadc7ad53ab09f369da6e79781f9557b86743afc56a61d8fe6d9841348af26e232493bf8c15d8f6c69b77fe84287daac9f27641ffb49b471ad2a64f5572cbb111858d0babf754630afbc995e2511940f65a1fe8376dbe20a68cf7c2088863eb8a935ec9fb0104cafe329c7c4fecbad2f75bbf8b7514833958075f11ecfa8f3bbd6481eb95685f8f62a7eb813d1fb770733677a2c15ccece225e2d05b39680192f865da24f03f5f87ebd87f8d10c10f50a4a7d73986e7fbd99db6027ace10c9431e7e51d3ea7705d7e47fa17cdb4197f203daf5bd5bb780cfcd4b6088c749308b76b1ab87041db026b30e736fc318165c8235d11eea6edc616c1613f53f9da1d2e6952d7c9ba0a54af392dcd38d932730eef25b32067d1425283c0797c1fb8ec75d518c2c2d436655e2e804644cb5a91e0f0449124b1c79ab2ecc3747ae961ba59a82707a0c1e5a2ce35b623d73102adddbce0c6b36ae153dc9ff6b22007bb6977d8981dcde26672b3e2a65872936f64a3e58744eac93d90803b9a94ef38025a556d1531c24ab2209e74315b0a18ce0c904ca8bdec551d54a20566692d4f98f1d8f5cb78f77273d39d53683967045c2d0fafc684bd72c25906774531b33331;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha7d4cc3aa6cf494697e56210770237b4c7e9b56f46922cf79a563aeb821a0dfa259039f45923cb224503e2b30b87fbcc66d4db7eee6353f6439e2b78c363ab4959514504e1eacdd723429f89b5b9d4f11e5145db654b57c55107eaac7f6a8b55e0f80448a51ce0e5fc7964e4bff8b6a3d37a8fd316b2f76ae632a2d18de2a2934149c6d4e9d8550664aa220c1268ab59a374c813512249cdcd1cd914257cc2202c742891b8ee35f62c569be6fdc31a0bf15e5a55f8e3385885489c139b3ada3464c990ebe6ceac0d05b799bf2e2d712a9212b9a97a2f5c41fcac3cd1949f4847cb893cd4a41d51e6f54da54a919e9968bb57186ced9e8fe42ec4f97ade05e2733f4abca1b5e03b01ab9c1ddd8ab1816f5794230c96b26f5fef23156ceab92db3a3441e60427525708dc75480f31b553dc5b4d2ab2d4dd161699a6f238f89c6741933fb0038aff0b3588070330164052d7f10d445eef0b7fc21d62b2d8ed3a703bf125d9939a8889f39217750cfa9c57131325ed06195e45ad56d17c5f698b9eb365734fedec86b14d8c3a140094587d1ead98a645b76d4aa3b249a875eabb431c49ab96ffefc2a40217f804fc36f8df182fd71dde294b0a207e6aa0bb996500803ba7eea638b4b2500c63f209424489f406e5343192696f0dd1426e08d73ca541a705235384eb5d553fc31589ac4c67f420a4c549e20d6487e047f2ee5aa65bbc23d93be38ad5068845388981bb629b05a7598fb8d86a1dc62f37bff99e0fabfed40ebea35d3c6516c6b2bdf16aab655b193215ddbc849e7a195651713c67d250dd4daa60dbea945b0c3e1bd9a6900172dd712d94618486f24ec6f36adb515d12bdc024e4e280e934dca76e60a75876996efa902f6fded37f322f31908f81cc974441953d3678667a280fe5c25a27da618fe2eafd359b15fd9b0695a6b1e2cd97ed5d11be21d91cf1e6af644cfca69b17c298398a5166d3e49324662686d99d530dc545bbd77c42aca5d9642299a04f5024d54ee2d062eb8a601a22b4c6b4b5584e6770756895f287dae93b5d3405e56722d57e1bcc57f87ed82011145fcaebe58c996c1f2dd171619d16532aeacbf8eecaf6176860108cf8c47ca054aee99df0e880adbfb1566473b708b459aaff9bc949fe88bd34105df8c4148e3cac425a141a9ae6a0193283bf70f9ec084cf5299f2428b479bc63701de2ab2908c735f384e05fd56d08d32acc11576ae7e4caa143d6ae75ea3ba640cb3c9543158a2fc09bdfdc11a6bcb11375ea8db6366dcb3529913b4daeccdde520727a6d17f1e39d8021e8f1f9a401c51ca1484c1396e86853b4ce2313be2c607d0776715f545e9e8c4fdd171d03769e20981ecead16f280c17e28f39c804747cbdc1d6dd0f55ccb5fcc8f7c2870c60e0b7b37f24f104ce9ff12922c627b8726d81e6821629e66026500d6272349988673c310467745ede7e4d399af3f7c176e065bf41b2e013345483a626b283facb226077384061bc74bdef5cd5b1d9474e8525972a495108956b933bbb0c1fa70fec846bc368db935a083725b00645278a52d504a68ff42646882cf18f19d3019965c8cde73ed1c378c6ee151292b94cba0d7c36f4a618d53a95c8029a7aaba4b85cd48d5818fdc4d3b798828b3a2e203655c7e98937253343c799345332720e270fd6fa12365249b712bb80d16774de7efb0de8341b333c4a6852ece1b3315e1d24ee726eca3f1c5a6e6c9acd56daa16910710283b2b3df43191382634820d4709bbbb3150a8e35773713b4c57a6c96c7d96c33530f39afff1b1aaae273fd008464650a8d1b23e0fce9f3ccd810376e075cc6a913e2c7d6ef4d2e74d7c3b1163bd4fa58fde9b0ad5643a28fcfb6a2b081518bdce5e696ae8138268405f18858a38ae199e6f1a666ec89ba27a3af37de501df26f19683754780eaff127cd03a847108deab2ecc3cc69ca1902a1b6c967f09ecf30120d7da817773f6c0cadb689f1adc001d55f93a6c9ee6633613ac0cc9d52d04beaae2220530ceab5d0e082af3c9f995100a724cbdb99111291a04f77585f5de869a547ce930de2b78d2070ec7b8d41239105574c6bd7a927288c1f28e4780f97224fabc0bbcfc17359a4c708d47b8c3f1435681338a3adf09d04143fcd83dccd6ec147e6bd344adf59282b683eaec61c25201c2e0a5aabb5993ae3ccaec3ba003d11522bc0169fc0c324eb8fb9f586a8ecce6e6a791e682c9ab503059c0959cf2ca91e95364bf13f966cfeca2598726df5ba183441192ab9a16aeb0d351b01b01d6edd8fe5f944fe33ed8a3161386665e9fbe987e0fee07cf74a42ac016afe4df2e0eb5aab6bfa0b67514ba7361f8e5da6a183114f72ad19478995b8976d8125cd652c2da9992bd77a89d09ac8001b639459d3165324f26668cec48f5b08fb857cc75cce6461d08cddee83c962b1bbe70b71ac76c7b8aafa5edcd715f40505fbddc30d3a21f01a6f48de254fb8ed98399a848f256fb98876ca7fcdc8677ba7f630b284950329ef01eb0f3eca8305297efd674516af42e15664c0dd8768875c530199e3cb7106010647dd9bf63c2820766006b9192ea43e4bec3fa183b013ce4e0972549f80cfe44a1c573ef67e23c50bedfe0ae00c962539ddc34899f5f4b9954878ed7675383263028124b8b0a1a9cc77c10594ad97b94be98c3f087b7200331e09f90c8cb6c131e2715687a422186eedcf9451ec365a7f352ebc183bafa630508fec1eebd4fe0d74b9242ff9aafe79385921f2cd29c742197575ae33e1d3afd05533543a8fbe364dc70eb42109eaa6911f70d9c79a716176479cd6ea11b554e507bf0ced392aa65db73504294a58645ab1ffcbe6492310c373785c13684ffded51b0a2d18875871f21237b7e070c63cc40a19ac26c2309b74b869f7e9c89a81f1b29fbf0ae4083562873bbacb63208cea93a483a3d545207e0f60b8c2b946ee225180ba867b0f298a368d9ec2457e433d2053b6733a9566d0c0ace4d6e7588bd57b00ac7f0af2b8f66983d2b5964cc525c5115033cac5315cc828e5536112919f7067b880a682e461d16963e9222d011b9a2c47970c1ee62168dda7a30f86fff7e6aa63ffa547f81adc758d7d82e29d6b97471eb879fd93ce5f6392b2373d7adbe4ada716bcd609095db6d0469e039d962a2724d325f6ac1f1f7ae3d8f9d51ca84aefb5df41d9763f6b4a0da6bf618c98430eb0a45a70be090d067cd67f4ff412617466ee6ea8a4251486a7c5fe624dedf8616ed7e1989d5e69f7d3fd9e1ed4f904a2c3d4c60c6dc07c9e176647779fe1ff360398e1bbde17f11a34e5377eca430646e66759d42578d414027a382d63891151e9371947a417fe3eca9f153e0688a366bc8b8601942012a83ba62296e43f4bdbd11814af9dfd5d0206f065e23e085eb1cf8ebf08e1772a2b8460a0e7e756929cc12e6c1988d78b65a1404c077867f1d4cea6407b9ec3ecf91f0673368dd8a7a656dc27d2173a16e588946c30a0eba25addeadaa1725d21e6dca0a63536a8d1fd1c8611e004a84a7213ca50a510c6500933ab833e2e76960490519d901c30a9f2479acd58a66312636b5ec462e603c79ea037458dfe37dea9db86e39a23c8d4983a3bff391d32a5acac0bc733553c24bb1273d3c86e86e5c99cdc74f0e57a762dc8b81ab5e73aa1aa941000e10f51656f45563427b94041c13b67b792289e6cea57014dcb13902b842260e8435d5c8967d82b1149fc5718c91506afd8983df2da00d2da014dad388bb08a6491dc4c51e517c7f6c66bafb2b1b27c698bd1ff18a11475da2d0adf81de180c6441988dc769418a56df52982de84ec2f2954071d21d8854479473db08b09fbac09bd3a7cbdd8a11c07d0f72100fa76710f495c5c7728878fc724c65005a560abcb8121d99568dd2b53b5eab801aa919103bc275a8f02eb11f19f3b81b449b46d1260c60b6f48488a63a1c2aa18fc5e693b28dad57d65bc061c9938f6ff467a3d3e25a0aa441f5cda5b999931ee1b90cf111de1f6fcb0f3e7867cf2530262ea7e37243de103d2831328f9bb354d8d5b8d5146f0d27864a84c9e2bd14a9dab7bd420c6297835382b9e403e7cc888956b6d4d6f3f3e9303be224bb7c94334b550e2de218c7cf999584e013abf1e478eaf15abe13821777510c81400d782e8552e39775c766a736c977a587b7dec9e13894444771803ccded1a1b5ab7a06c86feb5bb779d44385d7ec0abb3f71b7a6512a5d80fcc1ee8e1a09d0a3f16a8e91a94a1634b4aa56f221ca385406e9831f7d514230d1b6744e3d4f8091e329486f65ed421ed08c14be97338acd2a6a063b3ce9b1e4ddf7eb040a6037fd36ce6f8999950eaca1d9b62d5726fba1e6fc29ba836c113a67b414217238b4a5978c4bac25fdc29dd8635795a1c75d398f86a2e494703c5449633e0693f13d5a8e0d98777b851f48139e712b157810d8f7f4c292f8ec1321e6d04b65f65817a57badeee9f4a6f413beba31c76f14b90ab9d35a86ea9db362942e0694a428751a3aa3d8bd58477b14e1fc627747259361c62b5d0928c0e6d5af0b000a7de431cd4cc018f6cc03bd2b476fad7905014aba75a9d341f41065a2fe532cbe0cf60e8a9940d3a75b52201a6d37425114517597326d663f7e01a81cd18cd7eec9bccf7fd96c7251879493116af9eb6e3e9f44a10a29b963d69ef261dfd5d88669e2489661c86009fecbb669cb31af09a364a7344fb9c9cdf8f43bffeacd79f254c3174e18e1cf2184f39a1197c4c5c963938f0a899f115ac19b6fe677294de2188741522b28f12cfc5ab63263f30256e2125fdd1bed9e956fa9261dffd880cb7fa9d87a3b7f7b9f30f061880cb38837b8d23dc3f823292c9b2204468aafb7bb6d07125dcee7bb3007cd5697c6b1c7f7def7f3515760af325e38e6e8c5b8875b54d43481caaa1d5f29bb80e868519ef91f93e113b9b98f7eb381ba1d047a8678b7a5631c714eda0d1d2b3e1ba16154e140d75fc30a2c2385346f62c92b4a130e4d8beb18eca98697edcd797445303ceeced96f52e2ca8c19bb69d19b02b62ecff67c9792705e04d8027b18009ba4e6d33e157262f3a58bfd61fd3da8f6351e234ef12f8b3a77e1069d49c2df1128345b60e2b9188507cb1e04638175bcee12b2e849af48e6b49366837a996b80c8b302e8539bc4841b5018778bdec03443f0bd446e95558f68c502f171db297b20d4f0c8884a011a8693f0f6022be9b62a46eef1a1ab7f35f964873fa48705d249f73adebe9497bfb810b01b20f3770d6fde63ab68ff603ff35a409da55c5f033e3aeea5491891865ce0163b04b0a89d535d5232447e31f78117a30281de7fc770f43d5d78ce37c896f6c2322a3be9370f8a95e3e469dba0128893628f0ce353abb8623552623545f2ad9c1e8a7337e9ff699385ba39ab99c207d82840792e1551b6918d196d060fb4d37a2627d8eff532ae941dfd85;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd1f88f8496d9f801f661c598046ec7e172e5b09cce2a4b7f23bd704588e2f3e5355db21d441abec5df1cfc0082d8533cb3719799b81d5b7c056ff56162cc6032d94fed52b6fb3e45848d7af9d6d67cd8267229189fd6de55c041f8421131a86313d54508e48fba26e2cb6063753edcc3a9b58ad100c9c5a05e9a1fccb1b1ccf39d27eeff9ee22d643b6ec9a655d0d21ff0961f8a0c78de75059059987c9f4363b8423faeba15cb371e5fd8e554fcd646980efcc0c46611bdb52634728e1a9ac94d46cc9185e062fd737e7dc2f5c9816bed57564718a7ee3ba3612ee14115b67660b1836372acd38952515c0955eb767c5cbb2f221eb520953c8eea1f6c0b7e62f48d13b4f55bae3206d719a228642ee658b28dc987b4825c4b807e4131e8ab340971f8489042956a7bc6059fb48b9bdb2966e7f11934a207a87dca198588658a563eabc006581252bfa6ebfab8f84151d6db52ddadada3506f9029a653ac98e4ea6bb7cd7955b2085f4bc23d791e34e731e47dae86ecb511df73b569426c7f0d2d48444bebc2f0ff64ba11439b1db8c0879e774c026b91124732922630c1835b9fe5f48c1a0cb9242a3443aee74596f7441b5ddc38cb8a8d73fdcf8bb067d197fc5be42e9bce2f7ca929b7efd21deb03e46ee3d03a53c581fbcfeb0c8360afc549294a84f142c0967782077153e429de37c04d972d578775b4f53bf30fb40f88e2024f798ff6711d2548573166758f119cb358afa3ef90b6dd20ece8a302555620f1c09216f6f599b205f059e4a2b9d7b26fcb2f5cd6bea7280adb6f604041e8ab9e289bdfdd44065f79232ed41bed8d6819cdf898fd8853df0f54d5d5ede7cf9c75e010e6f55dbe60954124f743ef031289d350b836c284af193ffc9eb8fc3441c3075aef2e45f18ee9b26a2df422a2b2fd05f5351e95b6279c204ebb1f2532870a6a947b1d93ab000f9ba7b63ddacb2c525f946356bf4085bcaad3be95f6510fc6ae59b70a8e40fe78d6ad965591cc155e35682dc02436dd0f2345c3cfbddf8f5343c9eabe8e2e9f8c82215b41e3b8b81e5f68ce03d50781a86601c63300301be329b73943549cfcc299374c9a4be10ae8c350967a231c040bf39496ea9181f824b08717bf34efdc8062e7c62e8b90dacefdce08b33921580ab6a94bbfb92a5549c2bdd1ca4149c6b485c52e480bba30ca830ffd3eba231a54bb2c0b1007eef1101346bfaf9539a82b03c7f6e8cf31a9216b9a8eb9f4afdbe7794673efe166c803e9967d2cfb88bc9fe26d0067e7cf8fa5b88e650e2703b1fa7d628141360bd16ec334c3867d08374fcfe31121d8ed23825a99ca062bbe2f5993f1e8fe7540b453f1a12d90a08a22a0aeabfdb7e6a0e6df71b205a2dd6b6e01fee31d4427e39e18d7df6c63fe201b26082801e86b048a19a68e6523047956b6533d4f5eb189ed9c79c20803f5a0feeb78ed11f8b051662a09223d11ef5198ce67e6e25b3e183ab1c6459a0e04139517b0ecf9e249bb5434c5694eefb4e39908666b15d6879ebbfd71133fa64c275ad0a1c0ba1e6bc82006891dc32fc9ba6d5081a7de4367970844371a9c1f74d2b834ba0f167a6f6f41aca26dff842219091c14675f8f3216e4f836838459bdd789d6a86275e7273cd00c7cb8d80997e59f7a0fcf08d372aa17567066a04a3359b02bad4010c504097c5d0f41710eedfe34747132d169dbfb35b11fc8ae78b845984b6a2c4da53948ef29ad60b3e70470d4aa272e4e4774c16255bbf5c3b84b590d00fc824653d0d0611c0194d5893da1d1f5f240dde71d3622116f90f7469f367304a2ab8aaf89a747f887d6fe98d663812a224ccc9eba84d04d1bdc340ab6f833d675cf06208d638120f5fd0c8cd383780ec4400952fc7296ee15011b4fe2dec85310445fc2a09120dc2df8970e49a50dd61078c9158ccd9fd55068f550ffc3aa56e89e3dfe4f427909dc6576f8837de5379b1ee921dec8c3bafb867e8a5c7ac53cb2336a06095d18776911c4e970243dab51048542cdf3d8bc7fc67cb57bbb63f68e839d3957b8f45e70b80e5aa6f51956bacd591b205016069369195e4c3d802ba57a027ba5412ba17403237314f03ade21e220ccf4162f1a81264157209ea0058c98014cf85832fc28977cd66e3dc42e6b52122a1c4767aad7453c1bcef42ec966f720d17c2f446746fac94a7bda49e95ee03d0a928572c5598af63154ff169bb2e62da82360229e84302ed0fad2dc06b584db5a41315e00343e9abcd819d3c1f6ad660819142832fe7edfe3cb8e16f13f7543b26a8e4da1b5bdf4a280b2885cd3f9f254e345e6240372ab0803ea880e804d4b06713ee43a751606d68bab1fd16eefe1044330f0b17d9a76a86ce2fdde74f77331827c8096fd727797c9e0714a4f1753944b640cd698fb9979c794e9027cb7973eba57255c09e31ec1f16d05b75bbb56049933aeed510d97e5b13c60f73fce74822fcec4dac595cda364a1b3ac486c39b8fce2ba9f96c14e0217657ab271c33aa6cc7b46d9f201092fa1c6399aaf528c11dcbf7d2c52d80e75079e1b32c27b92868795a166a90bc7354c7c3b59bf7a53ef302a63eb48b14489a28321e60d3433bfd8ec6e7a92d15d0c6a240f61f363543d4a190dce81a90850010c2792765ab8573bb331b50b19c9f0e9087ba67be95d02386a8ab38fe434d33f50314a563a9f8b430a1f2d7670a83e4f457d5951898eb9de90293bcda283516f84a74e890b64476db80520acc5e6a9ad344fb438ae9b832be7b2020bd961cf498dd75083ce4eaca9619e2bef9b3aa85925564bcb8677d6fa035a238b5cc02d6fef994f4a44df44eb206c37929a14d18b2976ae1293b072ac6114aa7353e846c7bfbfd2f36be1fcd9323b4d672028570783a04545fac4fcc80887d1c6ee2bb4002db80a906a817207b1eb9e3b816b76d93c344c7cd772c469fd427ddaea3b4813185df77fee7efd26210548f882a2fffbd6e36d9e3b1d15e7a9abebb7cef47d3b9b0eca9c8c3dc5b6f325b57f88969c2200dbc99f2c3e6616c4f7fc19772b3f70caccf3c4abf4425ab4d6918df2fb23c9eb30defc2d597293d6936d2eacbef8ce27a1b0549ed6faccf1ac519c2516b62afbe5851abde079e6e1f1468be083ad733ab7e5024ca8716aa2d20b48e3ab740204c45251f40c7dae722f61e192ca4e957f9a13ffa2bd92f6d3b5f1cc86be14cb65828963631f38f60987cdad70de59640fddc9e9fd646407a2ad58a8e4d34a6d3c1433c03ad74f4fa6348f9daf04bed8754ab3c40e70e63c880c24cfa45d0e152c64adfb767afcfde8290cb7dadc9e9f5aad34acb2922b745f6345ea28a33b897175ff1a52e7e4f801b0ea3c420afccd29b65567faa624ade3efa8370856980e332c5ff0e1cf061b724162aa21fec8e86f53caed6127800aa50d077784aa19ac9952531991d8f76ef690a6e2e606494b7216813b71626221c1c7b116829a72e6c9508aad6c20ecc590e72d8c447cd9b0962f88170b1091f7eef6ac600b033cafdd3c2fc2c7d4373bf15f9392519837ec196a313745cf069f9e38ac2c4c529e2ac5d648a8db2b92bb0271a385f480ba4f867b7842c9abbce7f6f3167139076034f8d185667d5999479829006033ff7e0f8af811b198ac887da5bb03ca48c7945a254fbe66c42fc4ec3536dad3cbf9490bc6f66ad99888b1a38c4d7734a6a9616f1a7d90cb8aead9b2e79773efcb05a7fea25f3a8e076b5f4cbf8c83f91e144edfc6954e1061affcb3af405ea6068967852144a9d5ce717f22c04d518fe7dd180c0cd3eff0bdbcdcc41dd60f1630a8530a5e03b2d58e975e1f39f064e6512c2e40408f6f88059c470671d59d067ec012bafe0bba4c92f335a4fbd096bb884fcd90922f66f8844c3d3ef9b074e18b84fe24eb2af2463583e29f32f553578dbad4cb81434a34ec97d2a8e625d6ed3bb111f1edf7c4fedc0f6d4107d8e95667760e3da485f953bbde41eff5d0b9da0a7ed0fd5e23b4a6f6375165e16ab9fb33ab3adb04fc3fff35075a2e6717d558897eef6e8d308d57db08dc380e2f5573887e6974ca67fba07daa099c13f5bb8261f8a73d9b599b2b456b375ce2958d8054f0b30cabed95533de1bfa597295880ce8bccb501a3634de5006d62bafab745bf62edb83d900fb490b2a7443c9b92b46628d12ff751ddffc9db7c74398f223f8b81a37accda141bff1d924eb9fa759b1e08e8ba9771899bd176fc7474586a8543be6d8b72dcff44fb000465d38f9760ad7bea3104698525b16fbd33ded20c270768e7b15c2aa9f2f6abbb2b2b8a6d457c1b8cd07fb5287fc8df6d5b9dcb0551679438acb60be13744111408728801800b2c9b968f3b9f282faee334a760dc33e0f77ae4ccaec5b0246d9d3e98180a604e5eea17395a5920a9a2233cf9d9995f46baaca589878e2ae800a003a0fb4a2c556db323cb6b5a312ed538ab779b3f3dab9d7b53c9cf9299e70de2a6371d37a49aad9da8e1c2742e4ef8003d6f6c8327d312a2ef22415d9df66714547f6ea6781d3ad0a61ecba76aff69504fdd3e7f696ba853d94112d888fa1497d397d06a19374629786026069bcf6984881d8caa6fdec54f544c3d4aea5ded4fbc751749e3784ade4c104c6ba7e62658439b70bd83327aac9ca2a46138412924c202c8627c6a9d80f98cedb34a4afd06507a5d2162c00be909323963797c9d370f6a6436b112ae68ec6957c4ff2ae60b081fca87e4dac13a429f4606a95aaab84fbdebe6e1142a4083e78785d2a0c89cd3fc8c6121b823195354d1fdf02fee43fb2515e7695d4e8100e9753042305f4d0a2e18cc9ff6712ceee812835ff12c617d6dde4e04e14328f959be0b900aedb87cbae88c584bb41bfc30fa1ae2f200c6987790ed61d5b3f3a040a475736af1a3710f435793a7cef928a778366ea0614539911d813767943eb8bb67ebc1f85c1610a1700c349b3c11ff19f20d057ecbc918e3179d65452a556b82f0c14d380b6f63867cc05da202375ba2750ea4635a5e694a69700dce9c56aad81f57a6b984ce2814f9a6fbcf748b5c83439e1ad6e25ceacc0ff5632223efa8b5a3002d3fcfac481474b59d66ecc8406ae07b3e43392e635cf1385f58bc33c9f2dacabc8ebf842be6b2be80194fe022c4d413945ea38aa4cf4a38319fa8790dfe57304df9601d016bd071ace1c9c38bf1bddad5a1c93ca95e2000f1daa38657ff0cd850b4c792fee6ad5b3e9b3b6221acf235cdb32db07dbdb0fcf866314d670660a06c274ddbde8db30229beca1e191a24a6378ff9ad5217b4915d0ee0c2408d0f5405ed345e3138a737e8eda099875220c23edfe515671958313876af0c21e23c2ec3e6dc09e562cb52e1c3ce180d506f0264eea23989193c0c7413fdcb4046cd17ccc981a148470b3dbed36333ab35c7b34df08a42c1f28600c1abdddad23ec56661d88f7616fbc4c9de099e1d96229a69a97f43245263;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd00bab67923c8b67ed8fea349bca0cdd54b7454e1e70e5047aa7383eeb329186a74e57c4106e34b5e29d97ac9353273f28a9089f2845a3dc91391f3ad5aa86da50b4d59991618ae5394fa2ca3334d08b00c0391960dcc45be23323b43876ad212c4368e6b9e0c361b629887850324d93ccb7e706877f56b0e380aa0b9aba0476aff00cbeacf85cfdf986ef7ed146a85e58cc0c4c18a151d45ddd364a7ec16c2e24e80ff57616f2545a4171bf6347da6389daf7c883ab4a8e9c7e2becd0f5734dee9dc9530aa4d63ab23617514c174c0d118bbf377fecb72279d8909cd623c9dc5d52baa22f7ee9487260ca11af9ac84971e81d742f06813dc472194b1fcd2f4e25c56fd5ab126360a2ff5342cb383a7530c5f2be2a3940c3eb37bfab4ea99f84656d63f393a8c376cb75574db507a7efb8562d4aaaa45cd42ecf0472c41c50998472f618ffbc326baadb922fe2adbcb29c797252f2c5dd50bb755fbcde62b626854c52cc0c6f888208a19f5a807a43f23f4face5bbb49183589db49baef749a2d7bf356ce7fcb49f865fc5bbb7b45651d4886e207c111d2551778d01b037559412115e5d25a17e9104afee2aa741747e9bde17b223a081ef32cb76a4e3103dd5321a2dc844dd97787bbf683eda2fbdc11173844be2edf36a31fab62258249d3e301ac5244466d23b12e799ee1a3ef6c4975dfbffaa210edb3dcf8d561f3bdb767d34118cd1ab7922023235b3ef50026346f3c42285a9e7c49c708f99e8afa085d78f93214511903a80ed89222a2d23a3ea9eb74ded2c31a50b357c1ed11ce3d7324792a9863edefe419fddb6611ca0435e8db1120b97d15d0f9e5bf672a34979b50112b37f09537472db714f02f3a72c073365b0a91ada1b1d67b912cbe36e875f02a7a9afe7addec4368740a6490e0a6f4d9f6bee839284f6dafdc8ac112efc3d88db01ac42cb3ffb0c3f2e4745f25d52f257df8cb883ee01a23f0a3d86f1a923f6614b88e499de888b5efc21fa6d704c52d9263deba640f20b80f08b62a05011cf1e28f69297eb2f567740e84c11136b75c847f910fd20ba8e17705bca592df356f0f5cbad014c197437f4c5c925fb06cd0538faca4aaa010d63c0fab04e7004b51a1c96693654e746e0123eaabc5411bd2e71d9df0797d87fccebcbef481a2ddb0ea5f75f07330848fb77ba10f823826e8405630e7185441a419bd9e494ed59a5175d31bde3d5e592f5a688000cb1a76604305d7089f5119f3542d40596733bda3e3ae5ca97266aba30da90b7bd115e33e43cdf331c72527f9a6b78913927c2852a7bbd26cdca57447f812350e853c34444f7874257f0c9e68e6490982aa301ba35e604bdca0e211d4bcbf48a1095badd99b10caa1cc0c735b6e1c4e7ea3d23ec2bda793c743872bfd8b2b948d28ad8295b7eaf0b08a8a6f18e6db5e698a651ef39703da3b0a2e874ac332b42816b81044d34e9dddc02071c2b2938b03252a65df13803c88bf48bd12cdcc057ed2751655975b76db5d5c1a4bbfae6448c91c7b5689c1a08089d23504dae5cc0c0c2ee3622645d5fe55d0039eca76aec51e77d80076648f7d23b61a607f218f9c734997e9e3a44ad96103dcafb4bc79f750aac0ccded32b42e2266a6391cae6b9aa6d98b55207ee3dd63bbcefe3c0a637cc2495211785fe21d05858192cd0c2a05e5607f3fce03050991d9a8c07bcaf22543df4b52aa22daa33dc8deef80fb2327061e2be241da105d66de3cc15d09f9f0807739fd610bee6cead28dccfdb0b0331ad10e60f272ebabccdc20011c50e3a8628d4cef1fc11fe308b6945462de5affed58581e2eeacd235f94ce82550fe7316cef22a3b112e46049e74bf233f979b57eb62fede922ab42818256af83d331b51853ca4606cffceb06b8784bd4fe332b6355a6fb3474daa6c5900eebe91f388c4c6d8efff9c461eac06aa375087a0ce49a2bd9c2af7ae5ede783fdbceb8c7ca4bf0feabfff932a6049a6cf8f4d79a3ab46d3c71214eddbfc5b934bfc7c5a4b7bda7e4412abd927dc3bf1f83af527d48cc094b92e32b3e5d5264c579c135c762001019c992c872b1dd92e92cc720e3ee4ac4a7560fc465c6f7b0089df2fa2626cef74a3e64f840134a70412e057963f92bf611cccee08696883b291616cc81db8545639f37e25c396e9d8b1779a4ca6e27be5443a25fd189e817cbb61e945d6f90865302efd0ecb71c3e6f4f50e1c08384167db35cf5752d6754efdb9306bd600e8b5f84e812b49919b6aea0bd3fa312953cfe64e35c9c061d40eea60df6d5d02e2bc820f1bd035722dbc6a67c397c29a4ac55e17a206d7c0839804d52931095f7af6174f361e5fd6545a5fe368fad61b9232ba00bf9841205ec0773faf2797c12a47104c951bb9fab107ca861806cf5ad1ba0eaea5dbe30235747c9d4b4eab5a2681a34952ef6b12b1a37b0a0ff7fbc173ce6bfc7fbb742b82575790fc16a6c0494cfcdc85273377e59a754c8c089a6e589fa6a738a80f891e3db0590469a95542955ea82f63cf3189e3c059f798fcfe0e44b608fe82d395161abc1d3fe1b6bae002bd6a836bbbe0259b335294420399633539080aa7497c24d6d32eb02af512927487c151cc345b74de3cef6508586f229f673380b7ccce1a4b96bbf34ee5040f7967ba8878ba99dcddc0019711d1d676f64be8b81b2d82c17052b25d4974087a3b99b8a39ad79c4c0b3b9a40c1abe82855ccddc450fe79e00e9ed64d3dfc58efc3d0d7c0abd75ff04c1791522ac3f31f7da874fc71420b9bb69c9e7762b7516b1be9dbbeb12ee0cdafde54c980e35279720f04e9bbad756249d63f8281ab80925c6a696462a95c8093a88e7d339e514969580d400636e10883ef61be5703a1f3cca40e2e19bc774a4ece9e9ec533b58a49ba0913aa898049f159c5deb8cbf8c786e116fcbca3a303384de2768c2c85433bbc793cde53e407f900c6bb28967c071a07d68e70b464aa8b441ee9a9671f1b4cd104c8a180a4fb2ab5f33415606ed2a057fa49186cf61db3a897d2a1d972b96c5d3475825d137b6a5c1c26309fa7e90595c61f4b8bc7513daa80b1e91a195d18fbb29e6aa9887ef2f8bb89ac724d360b66173e06962b037bbc9b0910c424e6ed5a5a39923a75920e1575310f2dec3c77c86c5e7a40117dff1edc0b209d878a1c133f0a93c81ff3588d6be7cf5ca83d2ffb678a4f8894155ce62bedb79df3510eeb043baec2a48cc9a5fb3d27f8d40c7d5b753a42d917cfa8c8d1ca0f1f6214e645e3c236d079835841a43dcd802876cfd77337f84308ddf6a402d7cb61346f548ef4e19a5b5e9c2584585041f07d2d9707b5d6c93b2fab8a134766a1784f119dae87c1c19f534376c14fa72120a1b625d092fc614db7fc774614e1c474fcc5162f0cb9366efcc1b3f50e617666d671ee56db2d544442837fe2237c7c58b4f3b538746a10ffd224aacfd09c7c5e17c3f617cdff9a3df24c6774f12d4321ad92120989bbbd5e4a69e2673c6d6f57ad7409f1815e7f22e0883d667e7dce28bdcb29d9b8f2244791397ff38749f8def0044eab71289bd65c3165baf7105d763f3d2a3bf3857f4e4d6adc53efed83cb7bf46c51707135cefb86f6bb8269cf543d9cfa6e6a93681750097c7670debe1d3bdb02a88a637aaae8895b5ac3d83b755e26b1d79b2fd145ac8190abbfc62fcd2b80821dc4f8386b69dd34a66279a6fb872e143fc8287cc5f04717e12f06f21491ed65bc4686085a3e47a8a17af830e514d7de3ba336e0a0d571cb543cc1c07b1b80c67fd1ea10d145190ebd456c2bc400f0398057cd21e11e324b02fd4d666e38e2995261b0bb2f5cbc5541cb6f408f9b7783c589c62527a7ea5f6d6cd869052df089f7f623830b708e59edd69371dd4c5c8bf132aceb965dc089513d4182381b8100842a29f623471beb039bad314c859234b9c93796f6443a459aa3a6984e129489365a4111ae3a0fc99c9cf160d086430e11280b5e3259ed6afe09fe41b7832c2f8b9db2d213039fc84b02f147e724b35e35b0da8251d3e0452d9d6952877d5173414ee18db67b7f91ff474a948b861fb38c23407a1f4ddf929538556e1dc1f490b7501be9335a18156318a9863f512c5f57d333de91197abd99d64209f6483f0e33a2bb16cdbd767fe155ab1906006b52dbe23388b10237635ea1ea4bc2cf86b5a0c01fb6ac78b9fdcb5fdfc35e0bc7f5623ce7bbdd01bb68caacbe9191383b2e74f54667a1efcc13db5f45e4e4f9869e3c433584dbb44a436b8990e2f36f4124e41c6f154266dc47381400b054c8eae9065f99f4cb1ba1c25e521ba6eb239f9d644eeb54cca95a2c352f0c1f5a63c85d961ddb5dcf5d8d97e2ad6ecdef617c46f5ba83f730530ce41ed625dd00238c479e153cb47abcba907c568dc0616a7dff81e6c72fb1cdebea9d300af235c71422e324922acde5ad5fb22d69cf21c509b165a675d4a1f9b074156f91c906fa3cbbf87012b72dce9d867ddf5c62c16e71cf38778b84fc05cb97eac2adf42afa964da4e3785f4fb17702d1451689af08280434c1eb67e5413e5ccd8f6371abbd2e0aed3215c483f18138bc397c74a34c262a48c7feb62b4257da45d8754416aa9e1fbfff6ec761d6604174afa3c5c10144ad24870b5b21c6d4c2c2fde4dbb900d9e9a651dd5b40c9fd69289aaba32f80f6a47a210f5f13d5b00ed02e298abe9a531fcdb20ba966c7b02204fb1922f3fb3b12dc316139c08a4f7f8cb7d0b26ea898847b342e318984cf805b55fc4eb1bbd7d54f595da695c48877ecd3b088f679c6f6b94f9904325272148a7894f576c13c3e2ee016327cd1d3ff12a850142d378be6fb3d1e99068d9ac2d377eb657f7334a1edee0a44e4d3617aed367882a6b2da39c2a01539a7b6c6b21ef7d33a2e2c5fc757966f90115439a8a49e8a761c20a05a08f44ec8a343ea141e8ea5f6d67d342d761c26c542d4203b3c63ec45e766211b6da6cb4f5cc780901092453f1c4dc7b4a17c89c1430385a11774132ceee86ed6f596bbab775665b67b83e2263b0cfd8d8afe88ab9b0713d28d41a90e9be0050b98091de893682257279d5f588356635c4ba9b3d2bcb301fbb3f5721c0b2ebd2f7f4726e4a52b907d542fc6f542d1810d7e823a92b60902d09376def17764b2e308ab6ed7290f113b74f231a699036ed186e4bcb46db474d4c6ba8babf79908452c1b67397f8173a2ce3cbcf156a6a0a216c0786457f05ee6df2a19d903ebc22e46a1fec4038fbb9047168e19e11239875333a0ee147df20e1a33099f6e4136d867bd930fa5e7a7e1953d7403ac6ed73c62abc6723e3a3bf7fb8875c5d59cc3059c92716a02a21310b6fad80ee3d8655aa606167d3f53b5be5a27ad545738ad3c9318b857a36f9ffdc580d397c02551a1daf98be2face280ec27ae686e59a4524d5a5baffd0364f129b388b83ed1f31e3dd59454958287dbe19e38e223f6b4b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5d62561df88ef17e4a777f535782efd956effb048d73acac7cd6daf86ab8ff09ac3c483c5aa82ef8da009b6ecbbcf29908a16ea0f7d158ac3d1764aa1514b4a14bc92358096f13153d11cbaf1f9b4a1fe67761a52f9c5b1a9f5f67698a91fdf5f538e16cf0e01b273dfc655f0f97cf5b512a09b4bff85e79556ff99af9ba16a4c2a3b769d8169dd1219f2afee47f3870aae76c0158fb140e5e9c9a9c5a0c5d7788d9397a794a21a8cd244a2deb7e04a9babba91892f917d07ef2f53bd4032b1b1d62248c96e5439049364fac65ce8a1715a429fe2e9241e032bd0d48962ffe66b32563bda8bc314568344f9d3bf216cac602a91c4a13d0148373afd3e6d3bf6e09ab9feac2888177df93ec31b06154f03646ba5d7b1c6548bf0a556f24cfe5bfb330afe0e1dc965dd799669ac4619b7d7e0904106a2eccb2901650c0a3126254f5a14021e60af854b60a396518eec882003051b9230f110ee943192fc8e2fc5e9d89662cbba0b06ac41d280988b868eb5201876ac747379660f614d6dd9661ae53e0efed44222eaf914852d36ca8a7d86789d4fbfb7ccaae86ee0975f6ac4277646d13aa80d71caa903f168f9cd5bc5737456e931d8eeed192b7016e096f9fbb33140956cf56d39431c351d189022989b769eeeacace113ba5895b8f57f2dde93cff04e9de0db17ae3382fc2650175551c1c5b5a351376c9c7a0e6c1670f6dc29a8996d5944064ed76a5b1c03bdfd9d551e21e6ece0ec1942c65b62bd19d27754ed88f4e0afedabd1f1c7f23365fb36e8a517ccbbd6ae0923057d84912793be218df4c05c699e8f733b898816994db99265d18904bf5aaa7afee25794c7f40ab6ffdf9db40fb45a5584a2aebf05b0f4c001e2467c2ef1b9c481d493f35a8ce61c1c75370e657a8672288bab901c2cd3d309b8f182180c12d767aa7a046290a43803a9ea5a1da4695b5f00bc7c0abf43450da00538a8e9c460e3a836f6a1d35a3cf136016fb7abd309d26e088817239da892d028b54c601dc708ff1ffbbfa412da5d83e23a6dd8bb38c319d741d4cc746c6cc94d7c7ad4344e206966fc7136d8fbca0e11c77448674b27b504de92cb348156cfea232bc32ff6900ac81e280a5f61dc315127d2d9846860dba468f7ba1824250aede3f5d433459c636b8c215ec60949ecf501fb9b7c5d0657b8c8233851a4ea9a4cf8f8147803e43e696c1f6458ca690637fd4d54de929ce3d8eaa0ca93932eb13dce2480e3b7998caaaf79446cf6d9541ecaafe145f8706eb6882940595586e3b665b570733f8af6f213c5eb3b3d01dfb19eff0304571b3958d114044c993c71d2ef1c0c56111b9d0281a792dff3de82329d6e7feec7b42cbac3b154a4bf5792b3b744032bd9aa1561d03c114d2589dedee8cea369d458b2a9beeac7babd0aef13284034e57059f507a9ae51436e97920abc9ef1b8d18a1087210154d1836eef4ff2a5778116737fd62260d138c01d8bd04c65a1f914c3339a827884c63168a06e1a92ef28fd875a996b84eb15ad2d52f87bf838e4268ac8cc087e9c3289e0ef2959219cea533896b2e4f265242b06147efc333a47b839b9d3bad404617e2182ca051db4c01b7765106686cf753cdb21a39e790859b1b19107223bcb22e6add3ec3717d05568ba10f6f75fad34bcd337984f02db4a6f6d29e7a53d5affd650a087c5cf598b9fa4b76f38ab56e0e20073497f3b70c638f23f2c455ce3bce99d7e39f239d33a320085e675f25fe23eb7b6019d11c9378ad86ce0f5270ee673cf89182412de37d4854df2eff282f33bb893d9c25fdf6633f023eadbd50cb731fe0e4a9e67413dd3b2d63816a9dbe68d8423eb941e9fef6a51bf2888c86f5111fd39a3b5068924a854150fcebd45999dcc3be371c2ffab71cbce5046630eca76f8bded151ea9168d68232d026b3462ebc33fbf572e6de85f4da142d81e62952086de22621fd8ecd9bd57b910cc6cffdf7e1e5d45608613f3bfceb349791a880a0a57a25068b6e392e84d7966124b7618535a9af8620c1c22ce285fa1741d84f9732792be627d7f6b63bda9d2b2ff36a1078b159ae7f97ae7cf4ca19e3a06b58a5e9950cf9262a986e2e4261050e8db61e89dfc081baee14e6be68f3511e5d6afd7edb8bed5db41af7f9f8c501bed9d9c9776cc4d2ecc66e20d2b86aded2069ca678808b5bc546a675cd640946afa603fcfbcc4e6a2946f168fa39eb81c3790a17c926a1de40f921985b84663abf8540c150678c9e3b158cafd40c6520d0d2945b5832acf5c46a1b35b3212115a3bc4bb37817d346f030bdc3ed5f407e3f55d2f21a617fd1c06baaf11a3219486e6dd0a249290bc0468bad598bdb5679a5884cfabadc4b96a09ae88a8cf8c21381dfa02c031139cc207bba102149883e2d628f1cb895b7d94483f65f4bd1a283484c11dd1e06b7cfcc3c72085352025fabf8b37b7f4927ef6335e60ac62b25c00a8bf5069d0c29d90f151ef55020de1ad6573859d1bfeeb0c765011ab1483bd47b6afe803dcce90146437bb23f8df501d3808c452c7f83146a7ec680b934850a1c456056eadac11310e343c4272d99f2285394eb876efba074915f6f5d0748f04d8f2a63505e9c889ec3c5b77b2c15ebf334c3d24f4f67fdb4799f19b1be45e9de61345aef67fb572215a8c34494d2e01b870c942ff923bd16be725350c969ad51e18052697e21c531ecc24507d60ff7ee7c75418f6099acdd960e6272a1d627810230d956c6f60f20faf5b8cfe73a4f1421ec1b1574417d39edb1528e4caf8de63b70638c7eaef26795e3fae44c363e26662bd9bde5b7eb9cd6efaa4de6500e4bf4473a10adf662c75f92b4bbc96f6cfb370e9b04260edc2549da828874ea713db5fd5c696042661ff1a9e0dde64885adc23e1d0eb0dd9da06246c7514c03da279f2e343d0788de19a2908290aefde97a6662d6fd2df2290313473cccf644e9b0dae74605ea1240da5181a2058369a1b05b50d5332061139b6efae7ac00ebb49b5306867ccc7a0759c95bbb5adac1f68e89a17d823304544c0e7285dd9708aa3fbb228c130c2e5120d0e78b2c0c769a5f4311773a504fcf57426cd34302e1515b82e0354618dcb41d8d4d2fbe17e0d50be2992776722e8116f429d931b9b479c5d7378c616b1d1e03a8e830e976fe9bbe9d2f2908da7c42322c34712f68570d5a3ed7b382cf155647d32882570bf4ce38d573a40c6d7c2f1f5957bcb86f0d9a324430ca82bf15586bfd8c74cafe0a0454911b3da9924976f8bdcd07add9c3c61bf501a96795aecd7320e923e296079f0118675efefb89ea9b387ea66071a1803e691bcaf13c5285f30efc2f90285b4159771dd301221bfa114a3dd8f512bb48e9ba99232fd5cd0ce296a94d4758218d56800733cb7ece6e9a5d667060974211feb11e4f2b6ca22ad659e6592d71953bc6886e972b6d912b7c5f3703303253368b596919c08a68924f9a0765a558203a9a27810e4e9231d9d212feab1a0ac753182d2ce1b1dc2c148fb6603eb9eac82dfc34497535158284aeae519a20bc0415718b9a35f56474445ac369215e10b627cf8cb3f8ec272db6cfd646b0231e2b7d6bb6019501e384bcd1bb39be4c1d8a4281f187c92354205ab2251f76ba1feda4c850e4cf08965c1d8f9d1f09c71ab6769dd1568170843972d7255a03e5becae5757c64adb01ecd455c28ec4ea518a886f5c84104313d8895e15b812b4e9873c3cda7fb618f3b02088282f267bb239517344f33a893418fef856f3918f884cd151585c86979c7a1628ed6b5dba777b9313ccef635b31e9857be0cdd875cdd365038e3681f5051cdfb184608bff08fa72a1f523c0a44f70878516b66c28b7aff393de2de4d7f199c919179dc8c5a62c89d33ce2c30fcadb1a93fce4f269bb631d81d05dd31d962df4ed152c5d68292bb95fc3a1db04ab1de8fd860e10dc8cfd89f7913a472054fea0b7f1d0b0181e959c632f9219df6abe857bb5def4ae44ca982b405558f597a3824fa86dcec64adf61a8193860da3f3883052fb68a0f926e0e066347d48243a77dc0bac127a570564d14a35feb4550c248aae8f3ca3fe11c8ccf4e8ad3a791c3efd3ce5fcf2a040a6b1cb65bc8d2ad3a1e2bf73d0954c91447cd225574d8c2b065626f4fc313f4f2e4654d9e2180f19e1916f1478e7d8927853090baacc035d9bf962c43783efd08b31925f5585b224bcc121e76043a9f9ff4d719969744a4b712f4f7eb64d81f7d8c4a741550161e7a145d2d30501abeb4bd347360c17ba0eb6ca0a67264b21080f8d60f5b74d7d8e525aac2f71743791bdacbc9a2b0556681b7ac4c6deb0806d9e1216ae720c7398fe30b5755c9639ab4d18ccbab30db5aaf3b70ffa2a771673147c3736a1e40a687e10b85de75a5421bee1515694b25b5dca5da79bf13e4eb7ee91f9bcc0c75afc2d7903134be27d333508b0ff1ca1d56087f8f887b8baca886e8c81963475f61595324669446482b8c979c57e952071d7b560ec717e79783ec882cf70758d089c03cfc09059d7325d9da4969b3518778066fb915f215150a15200db9ee97e1da8f875866544eeafe255592d547a0b6bd3496192efd0f642f95482c13bd1fac69f63350061b53df61f4356ba89e3bed9f78d30135152a23888d6b04ae31338d70481a8db5fb5bf1b45a1b8200ed56e3b8728d9d29e2239fd147bd1e7dccf5bb14ca22da0274c08054ae4c1de54db8ffca0e1074dd6db000450c90e220084949239a92e0ca55c3447e9b1a24d6d716f4ff09072ceec4a9a433db563da57c280a38412ca97563e71340fb743ac337998cfd9e79d3c6509ce6c89978a57d5d8d1c99341c5cd99a91d7af80aafad64a199b166af58f3bba17c58a6ca3bffd521ecd6efef2051db2cdcbbf6edf68af7249b55becb9b05b95d4396710d70c12938c67bb155a2cb22942786c0f1cd171d2186dc9b2e354b88949ada768a7d0809f88636e551a26881be0c97a7a8d6f493990058ba101d8b6c55f0236d01a52136cf890a35c24e800fc3e03321808a865700d312aab11165f18cb3ece158aedf4e22bdd26cd6a585602d91f6c67b30a2c0a6277759acba73a201086efb05556ffef2f68ec8fdb91776af6b80cf8e3988f9f0d54b208377cb43d5c7ddad5ae623712ef369f2d535260ef94698f9ff1131bab715f1c43da20f14903cbc7050ab229bb1ecf12301b1d78e4b326c6a9f63934e2268fe72f8ad114de5541c03fc23b7b579da47ba52915c921551765626b80fb208980488a40488152fc44e281bce5abcb4822580b1f8a8bd02722c20829f63513b18737aa78d4d11e86c25ada48f37c891986b73129a65bc18dfd0e56784328efb935296b8a84c9757fa9526267003df805f875aca40360e17edc1c3b2b848081d8acf982506cbaf944abda3403b262ebec581fc3c0407cb93ce99faf25d3673454cb4bf392f64f7cf50e08e28ab2f2ec9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5bd69a4040b89372dda7c5e6bccbb2e9aaabb566e4f673837ea5933f1e80e10cdc105027ff21f9b6afb507f935afd5a02b1d9521fb6d837ed2269066aa7a4ca7bd6d48aae68704b27c78d4f56604f4c89455c476cb2ac6c8aa160f3b885973ec589aca33b8cbc4f9b0bcc7f95f0a05e363434c3ef3a84cea8dbc156b5f0d3a7711006bc778483f4bb90edd9c8c68a0755f79b0f0c2b465c077ff4a8203c6a5007155b93986465ca69849216490dd9291964e9d937a7ca9e81acb443318c928230b6b4cafef61c4c4e5191f15dbc17554ec181a173712483a271ea2937088ca5cb501b85cbc7cb563fd14b36f62a47150ce0afe5e4ca5574342e13943e1f8744ab250b5dbc767e643469e4d166635b5859f162eac5e8a451d6de5351da98724fb0b9f57c0423c9f3dce24e3fdfb5904670d4547448528a032269100762924c28b94e7d8bf0f37d697933624cb99d2bb5757bdd9dbd45682870bf9b3666c29a2b105715128c93a94cdf6faec46438524689f2298346b45d6ed24136f4334ee1a281eb23fe0688157295e40cf0347d6e8c7d3a0ed9ed44a5068e9bd05b61c8248da6c5b5c34360d42087426db1ac788b007830172f68ae486c7831387ec77e62a1f0a3b19a7e0779080fb463507ac8facab6b0dbc9687a764cc2adf32b747edcc742ee69a475781641fbe010f9e6d740946daea4900803365332c4f1fe956158fc01c381eb11a52df917b81916bd771c17c13f16bed8cbb84f5a284664fa52cf8397f5c79d4ef64d7597839cf44fee3d1d77c586ee4e89d2156af1f2e153808b0282b14aee1e919424f7a2268dad63239193e3d5c1b74faa03a7dea22712003c411d6a21dcccb1938e832f6d87c3dcbcce08fda9cd5a23906fe0a416bf3250ecad877e701f956312d3d7bbe5e8b80122e23edc94ffbac788ed1e888b4c1a225fea3057431133b3f2cbb21217c4079dd3ddeb517ff7725395a8fc6e089d63984a3f1971d1a772187c223f90caeef2390bbcf4a3ed07669fb0ccd71260d23b7e2a07d5fe9b5188063107030934eb2f94a3aa1afdc931f126b8c2a2024015ae337785d73da26f62cd1b68a7183e2a085a40c676871a59a7ac878de6d18b8fff5e1349a445e7db10fcc624ca2b82681bcfede439eea56e537905159caa62d6c8e657a0b284b919873597124c52a5b916a5a380981231ffda60242ab94c6d8b0d1a92c2c77bfdc6163e514591ecd0882fc071f48c3d207dd7222539ae845007bb18516786c21379e77cf25ad87ebe0ab087a068bd555b18c0c3f7e67c58e26bb9347304f9ba0ce2005abde9c44029ab4e73e75a620956362c8c7a1269812b268397bea1a79e18f99366e4752def346e44d14bbaecda90b47c70e2323a65e51ea3be4d7f33543b45add14adbb187f0395d09ff4ea87fd78cec27682a722ffa69a04d36a4c685461d1d3c190fd99dbb69f8deb3b94704ecf2107d3a069088b6db08e58adfbcf288023df65c81b0ccfa0d10f62552062922eb5c5cd0ac7b497fb16c13e9a09d3e07c60561ca972aa64e1c73dc38d14f638693de8fed447a40b6f96ab0c8b156f897bb192930c1ddfc21de57a43851de7d9365c877359451d9a5c4af19105eeaed22a04f19d871c1206c66a1e2d784d1ec3eda779b6dbeb3f7c3cb2ea52dabe5bf854bc49924b61f5e43afb665b8bb1e03802841a3c364ac6d885b218e90ce0683e17815e36df728feb9673f974fad57b48d2db08edfe750248b7d3f08b37ed03d285264e765c1a6fa96691475a7976055ae0e288e222e861119fba78eba3245b9ad827a8af048d188f361791ab95049632b287a486a229289e63fba0db50d4ae5c1af6cb31b9de9cf1db5276daca538b0b572ec2a7f5b87e88c78c851c9c0703db8b5ea8fc555b04d58ad09882a524672c1d988657e812af9490289b7371d1ee8c62d01cea2ec1360d6e69dd27bc0490e254b59c8afc24bb061829f21deab08d15ca4be7c87f930fd63459bdfe431b1fec0fd307174821c85bb24cff4e3dee996d076ad884d79d93c48e14ca9939e91c084bb9eab8cf786f3205afa9209a79b0114155eea9916c85523c81457a5206e1bf9631a53292e5ed14896a14cf1a83b6665d351d8d3eccca0cb43049768d4e1a1e07069e7b6ccdc1d53bbed961672b1c35de36ee4aa6a39d4f495520e9b3311279ff2279f00d6547f0f6a76f2d391518fa7e8cef29549d459019a6f9bf38c53a7f55e9caea66be89528ec82cfa26b7a02474e74bcc3ddfc01d71d3b84184c7c0403968e010141fa9e86d92c61ea6a4235cb7b1d20b529533dc88571a9bfdf69568148d197afbfe5d04a6a9b0593c2b82143024ab871801fb8453e0372142425f56faf9aaf148a05f56b1e54cc441404570c70d67b72f21cd72081956096c8269b035ba026df99e785a692418202015a7146ac1c3fc3fd99685b5c12ce076c0f456e93ecf6eb499c30cf037d6c9b9a9b0684e3d6519ceca56da57e9af28f712126dd618dc4cca76196a2dfb571e3eeeeca3d2209899d2d40f0cd5aaebbcac635474df55e4f948ddc8e6752738adb6cdcd9aaaf4f8b94f5325f2c0908b59d61d46b094609b4c7b0f04669d8b9d08067842451e9af57fd3c711cc477a5b5b7958dc92401bf486ca34fb3e1445f0c3b08cd0eaa776755873af904742868c98d37c4eb4c74f77bd7996eaf3a8f51cdfde0e1b0ec7feba5fec54358e6a23486a1c75c8e298c0cb458b74b9cd328a2699ce3966cc22779e740061528bae8fae70d2b11a6f89c3977f28753be72871971a6be2fbb63008aae9315f72c523551715f8dbbd88e850857e704ce76ea7d43ea3f7d0b3fbaad609b2111edc43b82668b18d73d2b0aeadd314b517af8ec0642ef197fb6d276b7ea2a12d9579046b5e4a78150aecb386b5043441c1e565cec413f5c8d34beb5dae59d4cf840f7cf40022ff71ad513a8a10012b28880db748d8a3ce1cb5e3f6b2c108d3ada69382591e8be18b322f9650e79010d97d35541389fc43a144571893d28bc4fa0af7a65cd39d9a1ebda55f1e35db5046f801a5136153ff5435d4887bdeacf42fec9c9d03f1f6ee07c8f1a7b5ce8aaeb893283888a28c36e83605f3dec7ed44ce750915c314eb92352f160042fad5ee63223785de59e1cd0ddc283df5c1bc862f453f0c94d3fc78fbb49ec424daa20937728bfa23dfabc26ed55922824cab222a9fb5b1124988669afeef18dc31e3a7024186108885e8381fdc1a8d7c09192770395316cdf8ee1255c9cde8c8e6c1a3f531888793de8215101902a28d6e6e04f9ff6701f5d0e826abf7e1dfedb666ff6b92d2e576e6cd279cb1985d00e5a2a85fb1d702033dc29b56f3f2f0a2795bed1304fc6ea07ab994df71901d5a8b4188260d6fbe9dd27cf25fdc1ece2178f9d640f9a5a79d93b40ed196d1d41b537cfabd72fcf8a4de7a8347df0a6df2d639e42d523e66f80c10b02c98f65064a63e1caabd6130dcb78cc22f234600c5ef39e206d601e651f305ae52b986e94ca384a75d6618bef2bbf2cb78977bcf281f62fbbdec319badc4d7954a62d791d696b3e4b26dd9ec8cb4f7ae682e873c39c645508c0b3086c3e36e1efca071b14f8287d47bf01a567f6f0039fa4ef18aae727a9643b71e08dfe34952f365a3a4d68f91987f3f6a78018592f1aa83dde8e0f2e96797ca7fe2dfd04a7e15cccfb33cbbeb4fbfc50c6fa3e1ec57c98077ea3360767c14737473e129211f7feee81dedd9c089e8b5c824e2a2bf552acb60d38c6ba89ba6ce0156625981d52957944d59cc73e644bcf5c0079121fb4af0922925c3c6303cc483c85037904028b3cbbaa8d0ca69e87d4adc269cc7018b6c80531232b81ee8146cd03e187fb4b8ec2b071b49a193a90aed07e48ba1dc5ae2989f1dce35bd61be9fda2dc677dd93f7fa860fc2a226bb797cc733da8a759710933bcf221e644fd095d377f16748614f126ce53d80cf9022385638d169e7ee8fb1cf6be07102186de5a2137a53d1d64ff9e16005c46dbb4bb2dbb9d90fc0e4b544326d77335f9f0630c382ec98867576e3258ecdc8f5ed18058fcabf0f97d0cda9117a61d0e316ae732088f387d1437a0949f60ee7b75efae79ec171a4aae6d5520899af6e93e3bd9276bc09f058c6dee06ac814914412e07382a56a7e81a59146107b28f2030765bf92d1bcf3103aa204d47150d0dcb91487121b22daf40fb470f9f5dda367f5fcb6d87c77f6c1ee947d56771c1e500359457e022a7016ee5d66409dd67b8071d65222f0a648e280218b67d92e649dab8d38cfe62b8363e05e27dba6a503594efef1ac63075242c17bce3c2f32bbebce8d0f80a78759e0aeb14f9643a6877deb05960c12c7400f8ded22d0346babfae4c91aa14f9ba8a4c51b21f32deaf086e596dd8c164a6b10bc404a5d1d0c72a720c183b98a9750a90897176a2533ce84235b967370cd0a15ec5e9515b6d3745d369d8a6ceee28321e4beea07ec4d8da82cfddc07af89012fc985ef76e4ba81cf6a9c8fb0eaf8c3fd22d936586cae334578b9421bc0dffdb63e882ad83249c5e57d159727d47e3e5c6c2ef198fe570b0325343ec24592539c7572b3ab7cdd42edf10398fb0a42cb8d9a8c85ddf88ce22c80f34994542b5a5ffcc88ec735f1df36900b0ce426379435aa9a3980081221764a9bf4c35c550996df1395a30f5b9c21e5bb15132a1356ebd86788d8382eaa42f78a73dd52d601286867bec730763e73bbb5a396d7b4bb6b7548978e10c42b166ce65837beedb745436475b288531517d6a02ce6872faead8bc66dd64b13d56dba83dd3dff2af7c3e5643068826e20c5cc60df3fed391a1108ec0bba43c5a1fa2d1714c782ab3a687ad68e9eaacab9d488fc8472a7cd6061603a69d5b1ac58efd8204abf7414f4e6ff18a908ae7a7c66af7e8a98072f16ee6eb861027dcf5e262c456ba23a987d21bc0db12523b02d001159addab0d93a816de911b3e9de8da0d9352835411f2e473d0a7bdd065119fe717dd6cdc6c1171727bc2f12b0e77dab56c635f184b9fd7ab5c06ccaaf3d0aa9ff3045d0c2a2157a74db177a85ff8124698505babcae36be88a4f9cc80911ae87127b553a453888d6cf93fe6b4a503454ee03059e72fe150141c5fad9bbd6f10df99330fc775fe23a9e9a4e9ee1f8b6d6fe3543f28f6697e3cfff26c0abfeaba24afac2c69bdeff4ee65e529353962a3de162fe2c531c82c5911733a21277a511ce62ce68c82778a60d92533c46a7885184605eaa5906a8e8823c1f2a0b60593ab58dc750b5e0b253a35be2bf8c1dff2f9303ab1f5bd8fdf7893fae5f1bbab7f76c703f3c6ea0c4c8b73d4dbccc2df4a95b06a9839d3d20180469ddcb4b4503a90f24766c0e2b8f90eab488a3c1d1f13fd507c040320fbe7c16f392d1ec73b7db7f5ee96fdfcbe79be61a4cbf2a67253f121d95fad1485b572c4e91acd4d9ee1b42f19b569e6886e53a5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h9a4e4d7119299b171fb61336fdd0e8a0f1aee9a5827d420374cf0cf6d0d20ee03b0371ed9a44ae85fb16c01764e0487ec9808d76e20bc625d54cbf876ced803398cafb7064d7e1d4d831075d925979e5d7445b6635e0a47127993da99c64c55df64dc27613d12836104eb5c6d3664cc0d11c29d2d3d94d09083fcf9d159b12e67a20adb3c3a5bc60e7097b98ee2b86222b092177c55c3576739b3096782ada88b21f28277edfd1d414e40598cab5901efe44e32cfc8e080e0b67c8aa423752d5eba2db1c283444cbb9e61c84d06ce435f9fab948424b5ef0f36a4b0e1c44385bf3ab517dc1b997a0a6f050067fb6e1c32321ee3d7e5579548589a3249e45092bad729fe33dddc853624fff415e71d6194ee70f3e198642cd535311a8abd6553df49161a5a26bb4f3782de81d4f9192b6c831188f5b3a5edc4a6bd1c12a5337476042ba814549b7579e64d3888fd2d5587a80f5f3785dbb87034b2666dc215f1bbdf7c5499a8009aca98b78345cc8ab58ad32f7c7882fc40341eb63484c80398a04082554c7c2d11f559f1b50178883a03f1557ec76e11b0c6d7e418b3156cb33d93369ab3050971120a53892ec6620937758447ee38e13feacc9ab3643ec7b11b1c4338ab524aa2551d8670fa2a9414fcaefedb07cf0461fb736af655fea505e4c3a104195544ef2e8c11b92eab6835fa750bc173eb1fe4e5441612a231c453e06c7698fb32ec9c13d13437f794de248a6e9c0a3703d4e12ae13864d0126f65bfa7eb7b3cae8f0873b3f552b56df3d4b743789711ebdddf22274f1c15bc154edcb291cfc4b77037cc7e54f31a6525b9bc15fac13da3ed3900bc93966309e955e6ee8d30af9df602c039827673a23714e61708b46fe13e975155ab1d743576c73fb6e6b2a9656650cea1ab6312e51165c44d6572052794bd9be45a34256cc10923d4c40a40b4cef2c01f6d2efbdff24b45105e3d5d023d9978be34b56d2055d7f5f2b2a3b031b00edc99b75d688f637b58ddf72f539b2d88469e27a2c3a22e4afb7a02aa79d37b194cfebcc20916d0e3fb1b34fb81a3db71c571cdeb11aabdcac455e60f89b49acab4d8d188893c2f2704848a09ca51619833ab92ebc3e4dd991d9a07ca6f84d8dcfbf90640a5f44116d0946b08ac6ab4c4760b4e2c20c37476e688925716e2b1605f5452e6c94f0f5e0d516cfefb5c9c1a7e89f08faa6f7e90ef99d2e5024147d0ab42643e7539a8990aaaa46e736149c9d10ff0417c9e207363867e9c79a4691b89babc02359ca92b4781943ed4eddd3d6a5bf42b66ae97c566d2cecbc26a192a5a9f1ce188e0b59782a67ac1bfeeea3ad1e8050f9609718963af6ae6cc4102c315760205e51057269049873fc2acb15be11dc248362074a723444d2e003a450cfad21f61740c79390b2be533613e99caa27583bc8ec4618d2f048536c89233600cd49a31eef513cf1f975ae4c25c3dd7eacaa406fb38f8bf0f2d39183ee2a76a38e20d110e177b65bf5c774c7953eda002cf0d493b9eb2c8650eadd7e9744ac71e34852a7ce62f9135c78a4287ad8407fe2b3376af5f295ba998d08aa6a080d6bd0c8af721ed30cdd2e7a81acb9466cee3a994e6b36bb1365ca827ab0db9e75cde165fc52ec528d66a134847629c822447bfc1b5e98c55d2639ff5e95f736e60c058a36078fc26b631ab863d218490d88fc290c3395d4140c2ff70db4fdc26171d7d0e1f8a97b178531f44e35ea063e1dd6e21e2d2d33f5634a37486186519706a3107368986ddf10850b4a23116f5c60c2b5f9d4b74f21363fa81527500615b1606a56e4896381b41efdc7a1f95f2a99d0fa4ebd85984ae442391434d0134278b8fb394b7511a83fbc0599b61f6c1d17bda447cd6f4a1139126f173fa115e9e8dddea12fa5b0356beb4c0184c82a6fc5df7b84301b632ce48ed99c6d465075c44124f3a9ab762d736d0822b5a26912fc964683a47fe9843bb40103efad2c4f1ef49ccd4a1b42ecfad4993b76e639c7767a266dd40111ca8d272598246b1e34a7c845dda93d8cd09c5fdbbf54518e76eb700b5abe8a6a692362c8484447ad697c9c12e96021324aa722dea8608bf59aaa64c35a3e1b5c3e552b599eca0ce74f41ec199375b302df6ee4073c042cd0c6820ec783819fe021c21a416c2f56ac5c57ca2744f90632510b5a3e31b9c51435d0a30a0a96336662a3b2f710515a12470f4115d1cd9de2f5ba2037820cc6d66459a68f167690170c82ca456766170f6f556616651541b0973a0696ef7aa3e6f2f85ccafea6b00beb02a4b4ec3a254f7acbd9bf6bc20d336e640608b6f91315e3ba388863b60e9b74e5ec6b97513bc718cdc76c0f6f9e3f85b477664870558aa80ace3f771e12ee386dd7b56efae8cbe4ba3298e2d91045dfb410b786f91970f30c77a62bca671b00a31eaede77c0b1831813574227d2761ef349cc7ae0c0682b65ea5a2c2ae350eaffd2625de69f93a8b363daeeae5d68668c92debdf0191e626f111534c35c0ae50548f5b6477bc8a7ae1e509a9c45ea8b0900bd29b75ee68cae6feed2a93e5a231c2794320a35df18e6e0591546f93140d86802ae1da56e06161b2bff44d1542e00811cb95640f40c3c9537921478b9b8efe7bafc58dabafa83edb81e9bb885275a19763db463b6729692faa18cde45c62a18b2c4c42feaf683989d5aead00b8c69cd6b336f45fa26c5835e241a5755ce8620c38bb9f12c69a82d4586d8756be7758fc9518ad709f5e5bb476e3e8de04aa986ced4f4f53f8ff0b3b73b8c7a2859de228608cc6cd7c3eb17b18e2c6ef85488ecd1dd005f633cf4832d5fdfe5a2acea3392c60b92e88a923f4b248b83d637e01259e2d73368eaa1fd143dbbec6d22cef20e3f4dc40e49b299b67c51fa4be0f5f995dcdead823cd4c92c192d302cfcbf1043c303075f5982096b2c9c8d7652c64f08425defc5850cf257e94af29823d1557f55f3044692ed244c5afc4256db90a061860af0a2f515c1b2c345c00d9aed8f1c8ccf10abf18c855ed87df04be0704b8ae2b023762aa297c4ae4eda22b31d63725c302922e981d79859b5cb3dc63661d50ac6891484d273d7d21291ab81d03acd49b6d33d95b7dd421a571e8a3659b66ebd0efc56a55853675e91ffcbc77bb87a61a50a0a4c0114f183cd2ff8f678a397fe9da36b365e22d228c7a4cd20979e1c34b100020eee01a54dcde834cc9164e5cac291f3b05902b7da177a29771d6dbe2083bb22c3e7f690b2cb9403f368998fd81b9d5269dfc249072e399ce3fc98e757de50f9e97be7fc0d89406fc7b54284172d2398512daa3962e32001eb15cf374e19231e748a11f7b58d64ae74e845856f12b5586b43dc5f0f7df1b736acf2bd5085db293e8e91ebf95dd348a0a5df6d8fba80591b9212cecf1dafd834f1bd691936d5a31612d6d05762641b5f96e9e14bf3e66500b721f6de45094cf39bdbe4e99d531e686ce415d16d3e01381e1d25a4115298892e51a9e0d3857ddf17a93319a1522a646c4b9080ed820a07d50ccea177c691ecb58d432e304b2129f486d78d0b63677ec3371a9af8e3cb66390bbccc82963d6bccb531fad183165f8320f6c458a14cade99decdf75f505665bff602aa9a7756b9d30878a855397cf7e16b71b0806ae532001ae17e4ef9215c95c415880733775f879fdd966b8895c9f01a8a1db3d8173499c7c8057d2fcece0473d51e350296cabd5892045e324ec9634a55302dc6841d5dd05b6ebd49b48a4a0713d4f1ad4d213a9f5b0b5ae89e54f30bd074e2658e17f9c4013d3f683f15332d585f0f26845e0b6840ca639da390b3849ce78c78cc6e9b8b930e8b4fc84506a1a16a5b384a52ad2b1d0ce822b0f03ff6c72e57cac0371eee8f0e1ecd70706dab45c21db13b2bef67485c7ee5762230c17602f1016148fb438c14a4933bc2a015047e2f9fe3d59d50edeee0669758f0ed302afd879de85c41e51e73e7e5de6724af9791b37048164cc454dbaeab3c4dece566919a39820e04c41358aa5e8f4540cce9af50f39d5d1b0ac45d22ae2ed9dce17106d1c573412a6dfb9cb431d14eafe34229115b606ed2e6bff1469482258ccff57916083373afac2e24be6777f7cc934533dc3c6316b5353b04ea4ecd0c13bf338546599e7a6cc753756482f6e07dc57958cf5164c31a90463ea0c52c0ece8cf1be340cf58ee3647039fc35ae7e90e6ecb8414ea5af3d2b4cf3c1b1b2e4d119f7185e7077e80361f920577f5ee466166780fc72d22ccd8aae33432f32b8ed8ed096a1e005fef2bc4596f2fe541d875084beb3d72d8407ff16c71ce9c48ebd6498bb3abba555c82f4a35c319c80bc2c4e8c72641bc08dd728f32c5d04382609862d3384089c12af0947efc252225768445575f27d147de2d8d457090ebcb19dab2a5d0f25074f9ef45ea08e937c4c559c5051509576063ba15d936ecc23bc6b7974055b752b2d9a79db5df33adb04067ac29dd41905d86c76c70185562fc02f1d626fd872879201c4b806efaebf85251e25eca1b7221b11e3513b635a05d00cd5470b9b713e968e5a43cf716ae1bee4cc8847fde1ea55f96e9bc7246573030b6f62045e0c83648ccf123f454be0e841dfa1f9383ae8e206b17b6db2b1284bd878e6381caa68406a6a249c72a973fdffc61dc884fa97160011232836997762a6ca916a5848935f01fb81c49b0237673a5a0ab594bfe336e00befc44a93d0c3eda2eab562fad4ee2b906a785b6803cf035817e75f3bbe0a47109cea158b4d8a732efe50e0358484eb4901d776361facfd56a234f8b9aef1cb701960f9e97918d52b06d05468d5a0515e7dc8367bb0bcc5c5ad9e138aa6b8ccc8f4897d5dedd087862786ec9afedea6e992632dad1b4a395957e3fdc573d688b8b2d2cf41346333f7502db4692104dd976e893d5fabe3728a846dc0313af7ad1ae41993c7bfc9a23ff9fe119fdae4d2e77f1142ea2cd5330b215965221cd3f9030636216644e81043cb3abc2de1f0e48e65773f819958f0a9eae52da53b5a5e5f7d57336ba99c4e68bab13d14ee262579b73177922609646b878a3ee840bffd33c1433dd8648b780a1c12ba455945bb7253324a2b4f7ce70fc864021179d89cccc9b9b29291efb769cf0d519fabf04e7528170dd44f144419c92eb523561f2f9efb00e2b35bf12372f43d74e77e42c4013a0dee7c6d133ea0a35d6f17508812752876fcac34eb022a749060affb3d85600425817aad0615c62c5ae27a4c975eaa5c3114e84af2051293136ea47dc43264e5d12719a156bc7f8096a9a358a72b39b5ea4fd6fb1134a1ca3ab6546cb6251f0d72c8777b1caaebbc1d01cbb69bc7c9e8ea9291a74153b4862ab44b4f1f5b4ab02e86ad5c3bba5781005d8ccbd38a55447149e2163f3712f51627ccb032a00440054774a486f4c54f2960134b5ba441d9074850dd518150b71eadca326cd7b11d9752e514;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h683f1e17ad91e7e105ea770b96bacc1f06dc5daffc1cf688fe6f1f113a321a573ee81cbcca6215c5084a4711989a8d4eb69a15ea5ec6ab27571e1b48ff0a40301f1b9f1851c068b0b56d11b5901e9bb544f0009383ceac8ac6ad222ead3d74e306df75c47ae2e5a8bd58a15d88775010f0000e27fc2c3ae1b2e26c72c93775bf3d43eb20b9ce6718e3a5486d6179cba85e8120625984b65b4d6034e1bf19e2dedffca167f9bcbf237df245729e6dad6c9e20f61d57275a2763405755b56c1964f14d63beca957e4ea2ab6116ff5a35a6f6160d1036f5db6141857404bb7267e53025045f63da65c7c32ad23e949b42a190312df99e8d9ad774440655ad631c480c1981421fd00b5256688490178dcdefc3e820d07c74e31cb1774ad2d329daee1b2d697c18c98430ed85e44f6de5c81ca73e0898ffe42a34f3811c719ccf46dd37128ea7c833a589561913ff9209515bf99450236b1e8b8feeff50ac4b3d884b9cb618df22291bc4f764e4a13de22329a25595af6134f9724bdf3442ee3954168060810cb9aeb9e08282da2514d7aa1184b6c742a0fee3bc9b0346081048c4c06b1de985fdcd71282b95f7285fe7f7ed9a052ef2c9fcc976a5c4f873bcf9bf77db2e4d5c859679a9ae4105b431074ac001d699b2e599a3bdcafdf0b0182d75ea41ca4decc06775109356bcc4e1a1a0b8ef175160b00054ca9fa8feea7c4d0d7bca522db3d77dcfcc13a9388675b9913c977643b71cbe4f23ab777b54d9e0acb91960b437998e9accb0a611b2151726ae83d1e164c39b48322e60b5507787c085173fb69ba67be4a1cd603d845c35cb04b7a17083608b55076bec23282926aa1f5ebda0acec6d723016a3777a916ae20b698b3b27e8032a35d9d75b35320ed171e029f2d7e6b8cbf32f08bc2c9c77d1141496238d9c219bd6f937b2ab1f57d8898cc70f52829d1cb155eb84e6d7b466cce42951996ac4164f620ae9e4c0a3c4d90f686c891dd6ae1899fb585e096df94f8f8bb17c1d44e1bf160a181049333a60b033c0f35c311cd634cf1f2e82b3fe4788c6f11a36fdec8431b03025b44403e7f09500e0d4583995738d70b52fcf31e7c33fa33a40bf5a707eb518a52a177c5da4e4b133d27a58d3592e5304390de500c09fe3927c886a2a3c15f9bb01bacc94f7cc49034a52a07cc085e7b9951af4f24ab6bf80a9f34fd1d75e8cdf79fd3d4a36a0440671cf63345016cb373e110331ba46b0439a9006ceb1590d06b24761cd0867eec5b92e67373d6a81dbc27cce18c7334d507cf54972c0826a307e702df44052556733530e9b9a47e8accb72dac4bd08db8e06d7d4468cfbd474c36240e4f28f86d6c63110034506c3dcb7032f3da658c46ea9038bba627b1efb237178bb7076d021eac608fd00db20f7b0015a9fc727835e7f5f27b6fbae1cc0b446d09ad9f30d2d63bedec0808ce5a6023c8da98ccf398ece753cb3a8d0a53866d504e584aff637d5a52fd6972d1977342590baaccbf6ba4cc6575b12a1ba6ceeaaffa5ddde3233029aadc4c1ad8288499a547ae25d1b067fd5cae23447906b734a21d10cd44246bcfe4f76882c7e3c607a11c7e59a4fb806fdcfd8e4feb0d31044137e186f230827546f93dffc4b535fc33d13c3e9631d0b88933c2c4618a4e34e2900bdf8da79d3b4809acf5d1c19f326bd0c11c73cda78d5bb86eec2d6091b8afbdfe2d1fa82814ea1c3915e28c6a81fbca8df3e1f72dc758f6cb964ee60dc89f2c4e28a402c5dd46d9b8201873720380d901af91679f7d684b87e48684ecea9a8647e5f4133de8eba2df7a9bb33e9e494d7f5613ce532de618ce86e86ad9dd3afc0020aff6576b5209bd0dfb5ca5250fd34e3be8d8a775e0ac4fa99d015c2b250fc870b1f9e7a5201674aa1beb7bb7d330301f086e9fe722724d262579dd283deddac8fb30fc7c897c099de0b24618d7d06ba4840e263ece9709c97856d5ab4939d866690cfb69a7aa9ce7f3729a12a2ecf7663a30d5971a18fe5f014c293b5ba80f8820a0dbf14b6afd57c095d25ab0739022f40e1590033b8efd9076f67c35c4bf655a5852a016125c647a6b839db80c4658d68f213e65b4dd9cf4266df56f8e14d4f5591a50f0a447bb0f49ce69a96959d4181c4889e4dfcb761f3cc31c04e811002239de10430e5e6be49b074f1137ce1cd06e315512ea98d33b2586b08fc8012e9639279efefe760c92866ccf20c7cb914afd852d93b3a399bac2866472aa29b4a38d7aeaa1d1e8857fd4cbe1ec77bbff4ee3803da9ae22c619f28d371ba2412ce0254a614870ffe40ecb9cb7ef5e9ad166c21c7ae458e6f3ab3309d9e1b80c2ddbccf4af1446f56ba90bfd12e9e1c031be7e901de0a55d18049fd2607cb622951a09478b0cc7303c02c7377867cdcbe053a406497a6a06ab0cfb9716ace7e7d33e5b2d800a89bcf75292a119c9275f87c3d138ee4caf864c7def0111d3ffdd6b95ba30f4d19218c933ea7f6d3789ab66f2c3a8e67d92a05c1771f0c869bcb83596032c58a050fdf99f0780a4cefc6f4589bb9e074c82b96a54c7419e5c8a5dc3967b4d1b63cbc8af82834743a42393e7a0a88410294ede24cba067ce88bfe04df5d2a0c4d48f7062e65e5900adcce85ad33927d0a6a504b1f5bd3eba7e34290dc6da10fd39468a95826bd9ae8316fb2a9ac6715bb8ff88a1def8960d0a1704ffb0df1d3a349f3bcf85352b742bd30383441b9a2b43aa401087c3f7989eca7a4b040b7f26a241a52e32ef0e90f92bc8e1fafdca724b36ac9588b6a9113e7aab688922a2f641bd6b27ab2c12a9de17ef43ba4dbb928d24be744abfd6c6b08e3c068105dac76ddc7caf2061a8a0bff97f449d6de1f3d4375a3827e2982ee1a77c699f2817c73425fb6db39144db774300f44db0f677bbf6e8a8311affc169a9897dca69575d4c368a8b7f6b0ed3faab54498eb6f8307e233fec304be3bc2bba7cf74395134a05dbdbd5215d3b9e6c550c6f3e2b42645ed49a2673f625232e4d64803eff375eff3d21ba05410bb4eefc16b7f0df310beeeb9c5d95ff8eed45fb8041af645698c46fecf0ccdbf3564242d98b1d15763d5a1504911b5b14d4a2da4a415021a400a9a9e4cc5c38f34a00d8c40bf316a0098fc1711c0272c35e62b1ed09cbbacf3094753993c90fc785148bcfa5a37feff997620d9e249d9527dd3cfa5db53536e3f838a5bc14c32485d82596fe8016be3c7dfcfb726305c3b50a05b2aefb3531bcd3c83381f30d91159abadb07765f8a0fee2a7bc31bdc7df3a85b0ca38787e80f2db548cb0fc4b01cf7fb7ddaa026a624cebd3a1ea05f35e09f2cb1e54afe9ca4e302b813281c744c6b080b0fc40aa3592a0d6a586465e098f0d5c6672f34314f2d79b6953a6c8dc7aa93f3ba5e0eb9b865252bb0960cef9981abb487c434d9b9a18e6bb8f7f5fbedabd862c83b5507282616c874705c1a11949a795139931ff1bd1cb621af47ca524933885f10d79c8fc6175a2bbb0714ade9f9a2d5e91f756506f693e362a5d7b8bd190ba72acf6bcd82b3d12e953f7f4ecb214feb2ea9dc2dc82c53e63f64e454792a27aa313fc2bcd37e01ff3b6a325b39eab7f6d052a08d9281e5cde540b063e0a9eaf4709c9732a1658a1d35c3ca9a0c7b0590886cd9265224d5717f41b4a3246c7f1147a33842d4d40f152a8a9f6dcbd1b905051b82e8a5ef64dff33193b2daa7d8260ec55015b1bc884ae01f1b36c918dfbba4766728b23794ec9abc798a9f48cf34b60956247bedea87c9c35c0d911c7f65dfaf1038071240221249c6b49f0edc42e56c75119578cf1017f4f26d76239a9b93522a95860f10861354fd207f0a6fae08e65b9e1b56fac6204e100a011756f01075151c0c5d8485b9c644d370aac82bd53b03c2c316975a774bd7631b36822563755bc4cc3295f76b265cac483760c56b4f02a2fc908df6f7536e942d9499594000604a175b983bfabae01bc94bddafc4420fd3d06a6e3cef11461200411fbdb5376c994438e1bd8b86d178cb88aa02d4cbce65dd4e1fd764fccba128b718dc93d9f9d14d1ab2b97dcd238c7eb94f38c342b0a7643e0c5f018a3207fbc4908d9cecbfda93057e1dd652afb8c4d24d28c0c1a35b9e18c7b9634c808fb66bbd8e23018d91ec37f21eec3f25ac44b44bffe591157350725775771a25a201cff3d05c321ae5a62a20ae78c1b46e3df1384c12a0817af92f5956ed2e70115f2128f6a28579a6f0a64c108f88977820dfd126b3ecb0e55f1531628689e4e0830e9a0b79026aa799a4b442d3e7d23afab3cad5a49cddb4b75890d1c5e5c8419db587687cefd2310c21487d969cea521d677f2ed2b6662719e278e89f67c49a97198c314b7a8eda2887a9371b6c4d1b64305ab9d8e25323544d78fd911ad0b299271a7d49a7c82d2e881ce87078818236d5d60743ee23e7decf977a2a86adcb8b26843a960fc9ae6298aa0a121f67c2b6bd8d4826b5758174ba1f373a01e4d8054ac8a685bca1dd09c8ecacbafe9a4a273e4fdf976ed54f6089fbb17594efd81426000a340c6effa8f0eaa51342c666e6d1087115b51105b28b06c5f2f581171bbf9c3eb4f234582ad885b169056db95e5da7cd4a6997a8d678c2120677f7b275f260b651ad205ba5de91d0c29ef4c8d62936d86951f212d1a124aa054a18dd304b0b2dacc6da17a0c6db689935b0d665e641a23d25ad2098976915d88a94d55e9c7782601c53d464553228e2796e5980d165b4b3e5c9289d44a1a58b280a7da23e49bbcc9dba17d852219f972caa16a6fc965bb061616f8e13c1ed5f7e3f6d049bd796daafa779a18c6fac0e22babfce26e49b888a17ab0aee3b78e57c668d6a64712ed7344d7b371f278a4e0fbcfbfebdbd2838c78c13a09afc99d20ed4d06ae802d980cf667c4fd4c463e14be47cb36c6c67217c1e95eb4379cff4770588370c3b8db26813e392817712046edc216fb6658d9894fe78afde9e6046f3046b68deacf21fe81281ebeabfc107d9bce110edaad485d85f9c64bf4af47ace36b3fde747543242d111c7b02e3f9a09ea210205460a8c118f7b5293fdf17661d35a9572738bf18a439fe36e49943ebe24d59fae08a3b1b1d0d26e2856a15378d2a19a70986aea70942e4df92f63b8545e1d5ae814443ef7bf53d0e1f3b4ebd5c0ed1d0dcad128d38148de7daa99277e19f53c4ad8b0ea4ae220a39488cbb165a5ec0de0ff8d16017299b13751446342b836c918747fa18fade62fab836ae5a05e9f5d1450b301b48cc5d6b466eb2dd8c9c60040d449287b9c778a6dd4f7c6abbe51206e495dea19d907741772924c37ea6ec9c2d0675cec645a257bd93d5fdf21aa33b2e3135a4b8f9e60de16b9a148c3da32b6cb37ee6fc88d049e2223ca55a3ad42f5d919a12506ac9880008823f5b2a6dab831cfedb84633c8d5d2b6b50256ef66979cf500a8191083a0a50d176468318b92b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'haf8489a5ecc07b4d2e462d1d88322ca01ec5f77a1e56282951f4df5fb248dc30da2c1f1925fcb6fedd9021f4a6fbbf9377e21836d5732867034ea8640c8e5cec79ef7d5066cf19134a5afe2916c81515324074f44a36f9322e99609c4c3c9a17f115e6751b41cf504bbd65bb6b8ab891abc32ca142505e9e506ff2803de0d4da50a68ac8de24e15f6b12453c9b31c11d1fc88cf25f460fdd1bb4c0cfa5b2343d01617d643fe192fe3a2f40ef53ca9bdbb08afde33444b13673d2c01c2bb06f43040747ad7f63d1cbca0fe845de40e9f49e00850639ef6c4b2c25f0a47f2a85e04c452a8c1245ae096a6e2d76aca6a91f3322f874f62777f7b4548ea2d0f8e590de5944352468ee69db4ebfcdb84a353c388ebd8874d09939bf9b5df6e5d00c8c67ce231e89a03eaa4689ca7865407b5d1a18c8b22f3fca55777f4ac034c1be8551f7f565d6c8259e17ad02dfd505fa60228dd18e6e52cb986209e38d7c57d66ca3b62536363a3f62a1c829a5ce305a505c3b4ddb6effc5583f89ddc9ad77967e3c551991af8bb6be6fb0a42a3c43ab7b3e8e97d44adc802b697116f94712b8c2984aa5b72d705e4e146de697ce273458ad4f2d1db08a65e296790f752cbf7cb6c4f1616a383b92d34e908e5f6388cff399213fb261d39f63af50b60f4efd555c3cbe6cbc3e66e55e98f9a64457948b7b7bd960567d2eb45ef9f434c5d64c9763f90f8038cfa36852344bf9c3f526f2f0eb01330477f91802477b2052a3401ec22bd1f627b608a6ad469e288b9949405858c2ac61da3093d232360d4801a5dfa01ce60b5a35826e8374b8c2f508282abd8fb390dd7ff83dacc0662718b0783b23c3f6cbfb0fcfe245d10c39090b9e47ebc022814098be9dc71c496286e12de184b3e4da32878a36192fb40d2d2ddfac1b1198c82c67d9d1dca48728e9c1a466631271a8189827ca3dc3a6bea50564c020b001a5e5eb7240bc213f89ac0e9b0f0fe179a97b38bf4c70acbd483ddc16958f025b00776ae103250dee10647a45c1f24dd69f8aa282027d792173ebc4960563327513fb35b5aebe65238a67d1cc01de3638f8c52d08b3a85de07c8fb4520e0aa91d57e6a4f67fa9eefa098a09fc162a155add76eec9d3c232886958a9e4a35b2d08e8f6673967f184a4d1ad0222ec087dc1f2f584e55f5e822e875c85fe4fc6dd86becb6894bdf633fc0de2fbb08f8dadae8d582fd44617cfd35ed369e278f17992cb3c1bcf60eb35d6308357923ac3fbab295a9e90b49a69e284f1afa4af811d76c775231a794d77a3be1d7de5fd56150af89b3b0f60047e96307a749bb49a0245bf91f0f334337789ec820f6dcd2fadb88eba236f2178f36b5c9bfa757a5f9281dcee0d9b0f47246a10e6b529bbdac655b1ecbc49dafb287592cae4038f085cbcaa6087a1fe1885f62491001f1045e5a03c2fb7f884463f5580307849b80f2c91a41ef82f960619ab4473fb49a07a6de2d6f33e9140257a3b16a75237eb22acd7ee047c40ae97603a4afc172390ffe32a4e62f24fbc930e20f3d51d7a3cca76ee932299717fa89e06f536f027b400369bc9ebcdabf6c8172a7269f88772ae135466b42f107aa8f26e9bcd4a1ae2ac26bf583f2ca7a2f58fc08a2999e468e42d904dcae650095680b83fc84cf5cb98734648aa0a4fa45b5efd932e0c511a353c90cdabb7a84855505a3d8ea6b00c26adc00513552192acf443cfdc39d1988db807a72f6abe95c66ef9b47911a5ecd4e4640d500f8b87cbb65408848cc6447f6fed13eb86495d5151d4d62f3266bb73f2fc2856493f3741ffce59103119cf6f2b709d60e750239b9fa0cd007177962ede8fbbbaf752b5e916921aa3e503cffc50ef88609125e98253bc3756e341cfca00a6c7d7fe684c062d6f23fe5cef2a22ffccf6fde0bf01f4b75ebec4f2a06f1022fddbfbce60ab4549dd49a8fa1eb0d8be3fb27860f77a2ddc261995fb8bf747779cd819037b695b5d0a02fb4d9ec81b2cc91b169e3661876679f491d65e7e38d85a590af38c6fc8975b50d6bb7cc365dd5dcf15a4edfa47d574bb615d9bb1c35d30a993c0e5021147303a455c4b39347a4559399adec246892d6e0abfdbb28ed5c6e30c7b2b2115ddafa0d1070578a83bbbf4bddf43f1211c8f3c0e8945ef0070f1865e4b9e982c9cef682aa7a2a89538b082d6c365f3112120db4fc78f99d20de619a97e27cb14d37840b4310ee0e84abb10f54906f4340444b93b8cd3a8e841157f408eed1c5a140251d3620a8116b83d5a68a502b456c06931546617fa1cc069664e4f3a988128bb147416f1c54049f5680de3ae4a64277fe153f6316d3243cb83455c29515b5804adfa308bef34d2d9b38915d7efa34f67cd423d3f2c2b99f78916d2fffbd78782cf1670e8f95be5e1471aaa279b35b8c63f71b5cd24e02285e145925001a4389fcd0a11c22d370aae739e6e2bf427ec2ba727248152a299906d34d61c3f2a1681a57e26e87b5bd757bcf68c6efb42c792a6d185ba035fa8addd7e2e2643f2b63c26bd7a1ce915c04c9d1ad3c788eac631773df09b50c3b538cc0c66508718da747133be89e440d0a2ea8e3a59ec48754178b9982399ed0ce341b705e31306b9d142e7bf1dcb635fba3ba213df905c9b9546bbc60775ee934297be63894678922bf434f5fa4ae806d9763cd92c423259c66cd141325c9221d7ca397f0372b9bd960dd5528337ad2723933c2fd7b83ecf10da08b920799a613bf674a6851d9b0882aab15201eaebcbb40a1b9b19b1fdffb492c748aab1a832aacf0482edb167523a30d87e233d585ca22c3389625ff3d587c4e751a52da5914fceda49b500eb862b54cfb30cb93a731888eb88e1c86693400ae4900c372083b562c59d1987a4cf0ad5d32657e0834921fea2357d0a82b3ba9a91b72e629fdd39758a7e8b3ded5bb06fc4a2ff611aca97390a4bb89af97ed7d430655b16045b4fce94dc48d9ca2924b6921068b95be86d9b011d9340606186a237e6672a9897f3234967336e21162e69968faa74249e9fef5a53190b7011a361442d6236b4f9c1be13ca508a5248be0d2926b59b4cf8dc71ff91582838f5f6be9dcc40dfefe350bc5ab2ab03cca430eb3be18bb5dbf58500092eaee6545e7193758bed40d8daaa3cca5809fa76a17d6c237ea876a6346d3ac16b9fb2f02e784ca857f64ce3731257e6d1baa1764ba1c2cd619bb934bb091fc00727c5048dcfaace6440326f3b35942ea8bd82bf16cffe5d75eddffdd92fb21f5d7228e96a5c31a51906a6a01ec35f17b7db5db384fa0c7fbebf02f2e5fcb2a9f60290ef62575bad1ba62d653e869fa4442666da1cce7abfba62e2f9b4342c7c7ebea07838858f326c3a9424ef6b19fd4f8ed95bef1c9f37e78f5d127599baffd76147f87ffcc9aa7f22f57e28abc6ebf8053e5dc2ff74d2f49deb4e87673f697b486feb8304fd2109b304431248b09f4ccaaf795578acc931cc3a243f5603f3b87577fd357e3f838a2846530fedd25147d95f6a187ce63fb6e78b62eace1c6af6a47470e1757fa77161360466a2192becab7e8640eb7432d9e6f91eef8e42af63130a6d070797ce8ddc05a53304748fef5a0378803d8a2b6300563bfe43498e10276a2e7a0c769ca804caf01be7c7745219e54fd9a401c520d9d403092c5dd18f5f7d035bac7d650205eaeb94a15de33328f1b2675d9ac6b80aadd3f868f586ea990a610ced32d8ab885fd75fae1404948eda7758dc95920d1478a925e4f4f578c52cf21080bed70382c290d7543e4083187730a9ad035fdce06926dae6e0509811b288dcb9e5bd72f2e49887afc91906cfee23bda40528b976b5f07c89a1ed5f28e89d49c2111f1fa72407391d14fd08b6ca86914b86d1c4c8edaf18d8b74897f1544c2900e20038a5e2a23cf97a25b700d398c6b4b70634c8035d0e47a563d1848d84eb98419546a89fe9479d21e3b7abe4501a7d46c114979516722e7612ce62efd4b1d8ff34fab799944825fce252d19d8fd4bbe022be114efa1eeefab4bb6e0282f0634b1924018bdb66f6ec7d138e2563c3e7cd6da4b20da53fd5506d75a8ef49fbe5d3fb8b3a51fc9a141e856d3684c3b84e0ec3206dba3249a457872ee04a563f0fea297b616c553928f66dd1dc3f240eea89bed9f7836bd98a4dc46166105538180cffeb6929c31361b9ab5d94daa286b0203ad051db1e1aceb0659a453a79e0759f0e096328c4297d6470e2b26509e29ccf4a1c20685f32c15ae247ab94b74883e5965496de7689162d1e43d79455b209ceeedf019d3b10275118f6ad50e33ab8c53d445df78ef3d3dcf0c5550e12c42c0a66aecfdd320330200094a4ae955f2d15c5e38eb4affa6868d1b4e6e25c59612888cb9130449c478d16e5e25fd522dfff8a5f5d292920b5bf2f70bb9ebfef543882e07368f988961ec2ef95404f2b7f4d0c226023c6ec746fd0534b1eb375455f65937899aca10ae30960c366b5ab9b830129362aae319b3b05a0ecb7a1fddfb8ff6602c46351d8c2653df96fde41d64814d66f4d8e49d5f9bd26b17ce7997e3659e8d07d84d8dc367e61e8ab14bc9761087ceeea81e2b17594dfaf94a945dfebfc1c90fb2fc60ada6fc37392e5a5a89c3f9d909c672f4735f58509cb4f35475f14d33943801ef3738b514a6c29742508c1ba016585b29060815804fcf5a48b5c0a4ff4fcbee3efe2fd8537e53e60ec0045e32c20fd7024b79833e67f970e99505f80e927691e09ec998d08c158a7e8f051a51dcb03665ed6f91a8fb294d4108aa578730e07b68945307ee9ff5b6c6032888f0b9726884cc0c2ca5b2915ed96115d32fb0fe63430180c4f5cac79a86ceec60afd934c5760750636e46dffa1b8f956794ea402c35985c925278617e70e9f1e7152fb99b4f3ca7b0c99707ab8347c4e25adfbc89603c5eb5cadb4120b6095bdc6db54b0ba3d6385942e7757e336f66fdca84de9f5ee029429fa45383e99b946a4f6aefd160b7b7ff5431174ea969e2ee6eba44e4f785e8ce356f79a7bd39db7a9ed991927c28754c393d9081b1ee3f0b584f1d84626ede1cca702cad4d6e43fdc99475d6df8b3e100f821d75970e82a3fd2aff16e7a3d97115dd8ad710de8a7f404ad1e6cedc044f65f619f8d68538dd632dcf944a0f72469292b8a03d0297cdd68d6e66e17a24bc27bc881bbba48b5be5fedac0850e2f798868bb247f9f2ddc0a457ff9df29001a3d98be792b335e1635f87083197c7dd2ccb916666f4d3eed23ef0004a8b3898fa9f0bfab6c84bf7fad1cede09d238a6cd745ee4993afc85232c6fc887e436f45f67a8d0a4a58229b1657a4db62232989a1d279b2179bb4498bfe6fd7abcc61686a25f4b0cf35504886da66ab18588b6bcf3f9a6bb4b2a9f972b8a2e90ab8db5cca3804c9dd078ab6a252a2832a690da0aa5e6ac73786176bbbed8c3469a7a0ba2e3049cad13a5934b97f7f5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1b3c7e1313aecb618ba796386fc6525304e949b61b9e8c306d9d6ad70900d7f687d0ed48926e7a45e79f8fe4e56f378e3feef2f9d4b31274feb85dcaefad50c5983de212a4173d3e1cd32b561dc8bc698ac75662da0e816f3a663f9b1f0a171698b1bc2e35361dddfdfc41e2497a35b738276d35597c5eee4fe9fccf2cbfa8e7087fdad462a1277cb1d3b08caa838660e077d126d8b10f11287998d2e2bd3ce69688ebf45a9f3911c2eabcffe04fc08f8fb5c56543bae8f31423e75d5baa86e08bbf2be60bff2353999a5bffffa9e9e105c61c01d0e0089b3cef672e8492739a502ac24d69d92d40dfcfdf220b442342a2d46a031eac9854699b6cc4e00e0bafeef59f6ae6560a662e860502e61c71684b44b3daaa4f1a07383a6670496bd2b9ae806344e446d248349d6c132bded6754ec27d084890bda0ab2dc77595f33cc5d9832066525850e5c9215b456bc2e30e2e8c986acc476ac096f83fbca031dc1385c60c40ab36a8bacef5252e0fd7607a1f3ff6a5398909834aae4bcfde6647a9a5d40b59b9cd2e3db0b34ad0daf8f854793804b4e134ff50770de64b07372fc62351c41e70d98e29e1f442bc40d0ebe738b24969fd6202bab3a8c7cc84321e6374988a5f85d24bb1c776816a99151e2a2338e4ac35cdb81661373c9e86a4b31e1caa86dfda5f6e66615527ea2a8d04791ff9e3b760b14ef739015dd1a707165e13d8b8149a7cf7118b8df27c211300a44dc93b8614037d1536460655a7b2ab37e0fcd28c95730fbd216030196a853fe0f956e2c21b83c7746b10f9ef132c856a02974d3e389b61f54f03a6feafadd52d2964cee8cabbe992505a3dc975e1739076e430f6d2afc86bb2a830a9460bfc65061b19a51cd798c606cc8cc111910e2372fa048c125aea2fedd1a8fd233d0ecb23f2f321d9d5997d02e6f99be9615c3d8e3c25da9df22c4701dc7d2b4a1c680e900ba2eb8ec8bc0bf83aebdebc5b9a03bd0fd977e7145abc4b09f8a1c04075b9241915bd885135894ebc2ed6db7961c153e4c6d7a55d607dc43dea7b5dba3105a6c7e1ac66101d19affc760a08315255a34c797e2bc817b7cfbf39127697ac98bc2ef8bb1171e13a0716680f3b8a65f0a435dfe1cfd04c13ffbe81c1e27f82c6942da30c722786333d6e4beedccbe2999b288437d502af486212e9ba6b26ed57a117d03a5cdadc6d0d8af46eb75c75ca6bed5585bee3b7f4511bff4c3eeeaba1b5714c72d18c6aa59cd4b8d7b51083b458f10054aa21edf5cc8171f76440de5cdad7b9e6468c053073afed14365bb7efc18153d640d25dcf00e073c27651ac897c036be64aed62a6830372203cf41bdade66f567467eb59ceeba4abd97dfc7aee2d2394968751b57ee066b2b2b5aaf304c99c0aef9d6c0c56c8ee2f894e5f81290c2ec381e80ec11cb04dbaac103054d964ab6448fb2c4221e11df0dc243884d8b8ec85b172b13e6595fe1143c5d619e787e97075e277a6248cafeb3f7a8c931e11f65003870230847e76465f12f5033e9ac8f31e4981425c048a9e9678239f6d30f095320e8bd39798b20567e8bf702f38e5a7a339ea1296f4b6ec724319b9b79104e5c50f9d13a8be3efa7c4c960a2ea73f4886b10e5121452f481fc33fd88605af2d39264f6fe2f532c8a111327635f5c42d18c65e5d866bed339b0856c40d2987b9d047994dbd96d37beae7bb4437cd3ccf4ecd5f7767a4508631996a7c105f71bea80cc8591bc71befd63a74ed1da23038f769670e6836b97e3076f06d948b9d97345da1137b785badbc04b715f7cbf69dfe4fb0c0721598dea64e985b9fcea6412f1f172bdce6599a6724573e092b2d3f055c937778d5263f5a0eaaf87c1a49ee3ce4372fc8c58b289655c32cb6625efbe9ee252fb2b3948de0bb959395a2be3195a02b787e4c4ca2bce5c3c88ddf7fa8e1b8a45232442341136211eab502d02870c9e5cc506538377263651e37c2981d4e0756b80fc3933d56c7907b39ca84ca1195ee27c7df360083ebbc77b43c75c1b5e43908d0923be85f36ec28f42327d8492060491e9730f9d3166b054206ac69f2b1230fe6b1c427d3d9cf3b32bdd6b03f11ff330b4f905463663afb83a5d8f8780b1f99a1d5b3b8187744c84aab9185e9902066a091472439c2a01002444dbaa3bbbb1392736693a2a1e5b52d5b75b4a3b24373d5167f003c3057179a960c8000011155b6387595d2844b7b1d52159d40338c0f90a505f8ea9f795c6dab61db7977b033d4f15664bdaba39f539cfd6fd9cb9b8911615292444485f6ec17376fb24632c4e3c90e27c21168bdaf258f94c88b9caf50e40360ad56ddcc108eb105f2aece66486477ef3efbe013617defcbeae316440c65a546afafe7c498971c540f2e91aa08c2b953d5630738b2a7016ff2f0aebda998ee11d9e6f24509d373721c08f7e387999a56c3b23c804132c8785a45593d08b7f3698d176db62f96b5b593a2a7578dcbbf5739e47d0520248bea2df76543c8a47e0f408b944a423341d8f9ebc20bcadc98a3f947b2d06b0a9fa1951f253f824b3de5d600cb25a24b8feb7a930562190016215db9a5ff5657c8bcd03e87f9b739c6e9eafd8a8e0de7adc33312f8f6ff854cb05da7e75bf00640a3e6cb53c830e86eecbb25111f9d1e35dd42d98ba32b54555b2eec6deed95b9772c948f76802adf38072450e064850a83532c8b9d483c34b67ebf7774eeed1b46f59e23551c6a116c1b51998348b9ff0efde5e72c1656adcb232fc50c54fe945bcb6dbcc65deaf95b6ff2b7cd368c9d2d55bc0042d16e18a21e4338d4e8184708be14670bed4b7d1395c5b153bc082f01d58c1986abc9a0e7063f9648fc64a79e2d484875c3179d286b2a523a438040f9c3d3706b9db17d53169f6d26a3d921e4c866e65747a49e121753a1f85b359e55461b90680103cf230376671ea0d65d45aa7a71b04ab25f542d95e11bf60307940bf43e8b7d487e7cc7b6038aa328374f1e4c95b74eb1dff57926721ee8b29c3fd8d973d14f715b8a542469a505ef4ee753331a3557bc6fcd242bda1a6c267dbd8662ab053550b75d35a983584797f215114d82806a2ca3be6a5756c4bd0b822f9510f6da3da7afc7a0c35aa4fba3393718015ecdaa25e41380ff8291f5aa22da7a93c0b6debff141c1bacd5cbad91d36f1f627247ef7d706b330d6b8b9bed8669a623ad596a9eb22a33c00946071b9d0916bf80350a0094ab945ebcf756abcd0b710b8c6efd95b734667bbb57636d7707e9f9416d2b4729e26d6287310de328376ec933419c047e74443aca6005a8f73e81f2bc860159ecc278d5a17c5c72dbab5394ce2c747b105b15f90a2fe9880c8c0372770414fc702733c5842b608b0189e24d2151d3456febca896459f0d1f6241922eaf34e60e735f20cd18074c27e33b875ad3a984ea8c92bb63af9f543f0d70dff852899236785e8b152773406b53067fc808362b9ec45c527b9dbd67d9f634975a5ccad4822a1a8eddcc16b999954630650e1cef3f92f47772ea2575684d8ba2d3f8b0b34e4bd97c51a6455f5118b7d918c3693ceb65432872db4473dd753a941b4a497945f038bfa02360538cfd6f618309a2653dffac94ab3640000aa8ca60c0564784e778a6568751e03be527c972167d4f655c6540047b7f6f4d48250eac8f22479ffc10fc330adeee65f0b8b7a1568eee5c9dc0b371e4c28f1c2fc6c01ffc3923352477ca5e4b089bcd47c4219fd5b4d6e34522d1bb75cbbc3f1d35db4786bedfb3e32d883073a6b00fa80313975c4df0cb4c3abea3bf13ced765d83f3e79df28f7085994833279ed210f8f8db688270868770b04d08f537c7587b6a4a2f029472c7536eeea2a25ad3f0b8f2f2726135293dda98639e322a188507bb1cab237c11c6ae2713f8a1fe8e82c735dfd2da72839b157a238646e41d705ee5a2d1c31bdbce6faaf56eabbed7cbd21f413a6d5a4616f3076332495b9cd195bf9348f41b26fb6bf2063179cb06d50a3006aaf869d6ae6a1c0cbac92b6dc8c448015e567d0a1b028e61a26334538ebb9e544cf9b5a0e8e9b09a200c89699ec8778fde2e671561701434be47796794e7679c4750c543d9bf0ed31748cefbf4fe9f80e11de4e805b42fb12ae54652b12057be6a8aaca947342f6343532f78fa12356d95ceaf22cfbe6d38d45d47cd06c51609a2a3fb13992cc84a379f39075066f581e536c9f024c269a3f0ae7ce5709e04974d2c45c6be465d12c056ac2b8723ce2fb641d78e35456781c152e59a74acf811efb850f5b0bd4d1dbe90edd38f1e28cd42275390dff2a4906b9a830cf4a8c9c2c8436326b046eaeb9faf25cf9d0a2ad509c7ee62a5d76fac295c11b5269b8faa1bcf93da70c1093cb3d848e766ecf8ae5b91eb62c890dd090fdb7e2c9c5a9cc6617b4fe472cec649af8d067ca899b9066e05bd039c37b50f0f659459150c81a546384cea7c91646486d512d35ec242eac961d5043e4e9dc373277012be26d05d7ff65d52dc6d16158c7932d094a9aa7afc7d3bc1bc6d26cfd83ce116f0ff22326f6456237c338806c01389cac499df1bb4f6606d591f3019773e0277c05df988dc81891f40fd581bc10241a191e7832a21d043418c71d7b58955c72013047c5b0d9c1c82bf330a1d4cdf62a1973c1713f7bd310c440cd52a15532a51fe914e40610ed726bb8e74ff98650e1e64b3da3805bc3eacccf473277f955845ad941dc94155fd30bf8358139e4e131819754ff185146773c8d4a4a25b7261f04a90a24d020ed2f5acdec5b553b3649ebf0957a55ceff447a7aedd4b9b61a271b72329c093d636a84dbc77ffe3443ffda3fb16eb2494f9b0ae3b256c1988ac9aae63563b321db20de649afff662d4b83a4e3d5fca030bfd65fb22f53b2dd07092a98fcf77885280d138936beb0800b3fbb36ebfbe4d3303f0d23d5a734c8f0a3838a066e4d9f48ddd148ad24c587abb882586c7d9eab9b0ad01ca42881865ee64a60ba2d50e65a422a928bee979bbe6c7f815b304b59b25e92b718ae314a23dbe65a3d27e22d985fe2546221f28f9cb446725a37de931c930dbdeb95ab7b63f60abe42c1df1816696b3c09a0d9deaeab51324f9a16916e7cbd036c7e275cec440b37b933e74f958ea3b7967651704bac850070acf489ba400cd318ea00b5ceeee59ae6e9ebaaf2e10bd4d0b37b5bc94c9d5d8f9e0f62781391c0e5e26a1e07d0fd541d4d7fa2a5eacec70ee679c61a0f64909281b957a93a8e790ccead91007aa530a12af0cfd80160e15ea70f28ba1f2c06f92003a57d6cb78f374a719107ba7a1915321f097109cc356a15dce2061b7213932458c421d826c7bfc437027bf5aa15d1db2516e2cba09548bd9d22c4a32fdf50237a03b8a38dea4f49a9b145b1a0a9ce9a1499f0ed63ce5adbb7437e3a65b5241147d1808a98f847dd7cfe847f02d18f61c2906c6f6cb2591001f9280;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8b83a6073476c70736bd2c18d89d30fa20dfb14ea595b1874b083516ba7ced663defcee9aeafaf2a948e4c017ffaf87e23f0bf125089d2961ba8aa0c8c806ed00a5c147712b0a454b7ce3f6fdb50d5ed86db6c648672c4f78ef019f53b19e0f9131c5574b82b434be03aeb681199e401ed534ae7f1c2329e9fc102c353faa895da1df2bd2f728d296c469e7b81d7fa9c12a2efa987b89ccc0d49f1c110fe3ad43a196afee58b989fcbe4562e704cc29c50dc562efa7f67f8dbab615a2bf4996da0da22836d7ba0ada429a1f14ed2082368227714d95d5ac69f44ca5ac93997bf4be576c897c854d9f2fce94a78efe15bde6e7960ea93b70ef3c17584fb5f778827704095f2db79b4cbf295327d3b03d248ae346ce065c726f557ed913e553ebd852ba15b237d849524f08600dcb82bee86604016c0394624c276aaa40056bf6c8a4f60069af6c22ae7d6fbd2cd605eeda6647baba071b66e1090092c17fcc2379c68e8dae11a65b5d7a35635819a7134af23484fca19cefab08696f65d194c20c518155147db8cd1a20d1db0a8cbfbe4c7e60a6bde32e7422ebc7960a5147c39b74b03ae23a843c37bd64aec0d3a6bb69e6f58e4e5d31598bd6db172661fcb98e9e00c5df0b6e107703cb74377cdb53ce05d8dfad7e40cb9eaf24ae4da03a030c7e8b9a664b81fc5167f714cf495e88d1f889cbdac1199b844055530aca5699f1aefaa792f71be78c2fcc137f0e4f2a66662a8a4ddc8e64d86869848132d5faaa3c34ccd1947b215860e4f036ad977e448cd4242585cae733eb84ed7f404ce8d2c0044c40e29bde40ba6d8d49e8f8d7c3fc0bd0860c89d54503a55eb9363500f9c4abe5d4f6a3bdcb3bbdd92165cf979f03a3fcc97e6d49bf6de8c3f240a2d3dfc6ec0dae92568c15300aac077c2859362c28eecc06d32aaa7d124cd899f4736f79daaae00e5dd762688c387840426abf355fa9a92e7dd6bca5d8cbf38b2da7443ff53193acd955c3c89c9ca03aaf311ed9ae6066f824131d5e42525de586eaf1387a39222780301ed6509f08b43ea110485545cbd605ae85b599031b6b58515548519e11f0378fcfa9d0725db2823fcee8794d4b0989062234f2f1b11f7c2bd4eac5d948edc52fd64ee8e65fc62871ce85655ad78ba023b974c0eab71f9e388d56c18ecf88e82ac77c4937e6e54f6ddee90bd00ed6eef419604566422a30d746975b22c94db1c784e7b12a886da74476ac7d897615fc95751bc364cd4abfa7408b1c62378d66148a164f10e5bcd0d1a8f0cfb112bbd42826b8c7823ee682472433244341af31308b4671a1315e5f8a559e0688e9b2ca3dde78db86317391629f24ceb1b1fcfffce5806621c3a3bc32cb3bf879cc77f4d31415999fbc9f49f5ab3bea767dad56ccc47ec3cc9d514365c9fe4000bae5c4d2139cd56cded6977b96be7787c507563496033a37f1c621aef733837207a32a7017498fc934070a4e5e796911cf3efab9eba1abdbb29033a81d9e619aab3d56aff818d9397f6e92ae459b982b309fa4e301d3bd8bf9013850ecca20116a0d7d1163b9e977e8575b27de687978bd1ab2f3bab63b47f3dd36688e77149584797b021f2fdd7935d520b2f291e87ec9a6adffe32f2b77a9e71dd064069b07849320b854073a2e3ab38f6732660eff28b4fe2a31427868bdaf6ba9dad8ea2deb3513ed2d41324199192fbed679c3ee6c2234c12a4d281da868490d2593190b50705807d4f7589b01d17cd80f21c6d80633abb782de5a1d0f669b3bdb9e00a74027b3b15720aed48da0876abc94984215aaad545ffdbdd17eb4e2529af9dcef69f3fa87785b8df6c28f8e63e707a78dde73be41027990b88d9712d7b7dab7a309aafd4884e3238c3277c1510fd06e17e8b66ab33bf9cece4d5f00b682f2f8aa79dc3609c8b6a9eb84a745b397e0b086be4a1dde1460ca0fcd02d47ad38fb97ae20ac23f5a29a6c47fd6b1ec0bfe992617ca3bb8656c5542ae9a0d57d26f5bb0f9571137916bef8e0973a257fb73103979edf49a24d3268084178f73755f4fef051e67060d35c79f4f46128460d41eeaabf00b476be89363e626858f68b998618bf469ff431d89bf7e5b7752e2722ecdfbc8037ccff95d78ff8abca568ee9b166fbc0b8644ec38e27ca5c60b928cceebb3a3f9718c2a45c99dbe4a840e39cf2663bdce8c4db40a882548b42fdecc19e9b68f4b9089ecc9d8fdf12253f97ac00d4289dafb31bd48817a0c480ddce27c06e5d91e8cfe0ab6ed3c38bbc9561196ed9094ed42bfbbd3abf29ecc5a891ed66d34838eaa43653f3f9f78183dedcd8e6397656c78eafa4976e3d7ada06ecd951044ecc458b1e4fa4a5425ac1d5e513ca676fe690e69465e059ab17d65359f4a2542f4aa30d85a2a832716e5fbac7fa50ba11d7664d7bb9edb0dcda07f6437f82e9e8c8fd20f5cb7e29c43240894a9a8fd4afc474b9d1d3e44c0336eb9a409240794fb574c443cb7d3be2f69a4e2899a531ba0795cb075394281b582fb6e4eca6f51965518041a875b1e341ace8ba60e14709ad9df04a17484b05d2ee309a5f4d25310bc7fb50cf802acf337c47b8d9f3ca85dbed40712f62e3087d99fbc6f2be1bd8a413e6b6f664bf0a146ea27519328d8d3f1f3a657667016be88bea0d862ef17553c4fcc0991c04e95dda46b959c612f3439d4a1f41285e6e9b4642e349f421e293882d55638e1728bfcb3597cf6417a407f4d3d47dcdb82a4e5e93b5f25a9bed0c7066c2aff2c2eb53794afed88ee27397b58bbf4e05921209ded80d0fa9f911a42b11e57d2e3f988e8cc349a381e20a4a945a7627d95286f83822c3b70a5fb908e21fdcf09cf9cc58f985a1a093b224a74746b86857c353256f0e8a944f7b001e95c52e051b8c2f9bfbef188b5c55565339824caac7133f3b58489d391bf8bc7a198f017601d69f89e8b682523f1afa79feea0fb1532d0d724fdbe204fcf861a75aeef5a95e55e8a3a337889875e022a053661affdc40efa9058f7a345aa1a71d8554def4dda57406deaeb1e68b80361c829118e47e571e03ee84cce2b839861570712aece3387d6b61dbe1ba767ea11a40a1c9fd410228195746e23bf0889bffb81d8633beaa88a0bbf8daad76086162b58412a34bf0e7c37fcc4042c69b7945e2f1dce8c14fa1d4d898c43db2ed7b7221a9c76f2586566f92acc18bcd7b2a142caa897c8e861bb15f5e18da6aad16a4a72211c690be7027936959bcd730e8237787537632026bb6695e83351d7b78050f95823f4a78838093c30d2be77d7bce7dab3f75c0cab7992d3564cfe50cfa3f7bca4ca533ec3eb1cc13a5fc643831f053585a21704254e2767331057bf39089465ec369870913f52d4b94e17d3e847dae56900f914146ebcea3470a97d3db132230c62bedeefcade264e598cb5fd72654fb0e3bbb4ac42cf2b6bee4504ea1e6095d59a3790f3ab93c49fa0dbf9db3ec154b4333bd482c980ca6fdcb90406b81a6d1606853af3187387d04a8ec3b7d9975400d8a525812cb5890cdb2d24b98c6227026919342cd7e01c3b67d2a71b1d6a78f9fdaeb77aa9c882758616ff23654ff23bb075789586a818dc2774f19e5049724d32271e093ef9411ca2e8c4d879db2949cc04b39554e1a866d1cbda0c80eea31c0051832bca7669a54f0266bc0fa77716c3d6e2c3d23f553fd889dc695b95cb3fbb210d5dbec710bd57126781a8d5c5c1eaf8e8694acb5d8582643c751396be725cf4b96981b2c9b0e3041eb7aacd357061a78c54dca1c9e643f4314752745ea67607456c387f418d6cce8d661424c765b6151676ce44922c3ec18a5b962773aaecb2839f89f78b5603dfa9f4a8001122ee7f70a62e12c1e6711b38558c08a2d1f27b80f94132a71557d95670c87f1db27cbc627566ebcf99d205fa611ae678d1e7926b65243eb1f3963641d8c4dcd5554794aa2c1e535b523b0a630eb68a6ec53e4405ae0d219486da817930a2fe5f73b31569cdec0d7ffac1aa379be55aeaba75df0e708cf8cfd43c96c7e6ed3b256fa802dbdcea74ee1cb09933ce76c24de9525c973016b3dff8639c015da4c9aa2b3fbf3c90569d3ff5807daf4429966532f25dc359bb1329f0549b775dc27381da8fd73959ca086cba134d2c190db5d76c49631fe21eb3969d28123608f631b7bbe5348197502732664eabf5e383e39157b83f572fac069a8ead1e46854f3cf83bcebe3f26a5cceb81ee97804888384fb3463d92a52ea1d324820ef52c95c06bc73399e16ced0068eac59be9789eb4d5b9c5df5671e82267f76874f8eb4afd334942be1ab5a2fc2c8d597f356c5ecfdca4c6350b78e05e5f7ed740a3eafe810e8e9353ab687d32b817f9ed34061797c1cfe8204d3289041fc07e9a33d75cbb5dea6655194ed3881bec248ea12083a0168b177f22cceb6d039de8400079f84106bd9c802bb3f49b6b69944c5231dcee91193bd7efea963b70d5710b02f820aa0053b144994007d8ebc9d3aeebd1e29d5386685dd76b58958960da5a9097a7c5e605b946bdf1a379e04890107e1f0055fe4df1ffed93e3faec57dd3c1e23f02966d9ceabaa797799dd813bb8751bb5b52ec827e91e112f2c0fb3ab394e4787af023e2075ea6b8798c30a5f560727ab2f5f28b0f8d64fbe79b9b95faf92b5cd4c6731e2a344291eaae1eea9400de23d3e8fb642a136bd21dfff33688a5be407af1868c3062a7f3a3c87e20fa9e1ed0325be748cf1ba8c1fac760cf6c64c6cb7f40380fa757e3a6955959fa1ffdc3b2da692ee891787948caef1ec09d4f8adeb39c5efecf59d0c66797edea09e293d3e29912e3622d23af5df3f3338b4b93b64ecd1e5a4ec2d8cde80cb6221c36f98d89b820c8a5afd54a5c85d0250bb22cb0940d2fd7bcd5f610dda9971b52b8bda8a0f86b34fb2482da8cd08f71db897ddf0f54ad280d0d5b2ff83452fd40e2b1acdcc7f43dbcf6dccbd627a8187c9359f9ae98d972da611759de40aafdcac291e3f89fd95f2dc159a027ca1b1bd16f15fdbced64206632e47396d99f7500015ac37e1bad422be9ba5386e124c611a7a6fb8f36f9224d7b4a5216e476c2f97a29638571f0d811d45da96aff5db40dafb6134b709cceb859c37fcb25246f86add43807f1208b505c13a69126edc8fc8340d8ee37f4ef7cd0a0f5fc550360615de431ee7997311bd4844e04c0e6547142e29cc179173ee6a7478e154538b81a20be3432a85fff7d03d43b5de7ef9b773dfd895dd6b8a49d528ef4ced3706272db833faf1c0782546614c09fa237c55dda43c4414bed0a409856af4748b4534c173e39267b566b77a3417fe9bed9bfa57986f3ee1d3bc703961e8e434a372142a838e166b6afe67e6a619545620fd8b2d77c50d2b3f91cf00bdade92b80099fa3aef121cedf94c25ed88335adbe12e610f72308692294e4e437a065925b2f4521c225340c338e2c87cf24f1bad35;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hcfc72edbc0848f7182ecd0dbf0c4dffb4a90a7484aef7477f1b81ba45b48671eb04366f50bc65f474dbc937f8e4e20b7e5e4a2b13b3a17bb3275839f46f0df87223abaac43b8f64cb9f4625eb9f1860c515f622840743409480bf25959a499bb0872ae08dc2a6eff54f6b221c2d541daee7bdbf5aa3c4c19bc6d67f5bb8052fc962c2741914645e761f854cbd5c7b6712440729de73022973c9c40f7d6ca8ebd601f22a7b5188008b967dd64e13f4f40091086b5e5a9d0b19f75ec1d53a52193a419caf7b8272179827681f3ce08a474d0b7cdd9edc4cad9868669f9e0b942459fd54b8ad130690ca762960c674b00247ee02573556687cd695afef8be50d8598afd5683d318197ebec53b54e3307c43dc4e6c6213b3675d802866e0ec8bce5e35e75fd7b23553062d7a3383cd9ab815ff87c10ad36688ebc36be6dd1667253a768ab03c1cfa67959e0d7bcb2706e463d2ec8898c78fffe70ec53bad618633efddbbc09967c469fdd7d2ba3b3fb64a9a808f43bd17e245f94819536bf39fe633ec8b11260a285bb56257bb04b89567eefc92bc7180228bd1e97d24bfada7ab2f1e8327aef9ef3df86c45239ea7dae0e5dc700623ff21b436ab4228accb24df41fb28f1cfd931c1c6b9250ee3e427b00811de45f49c58c1e74eee100e606f2a66542c6de3d13b62b7a0def1941aa090e3c786afdbee4097851fd95bf711a651a5e120b8c0906a9b206f9551fae129b3e0c6110be73b9a5ec03c86dfeebc74fad5a33d9d0a7c98e8ee81e7c1246d6cf95a3fbfe8d568721bc2bed59216b79ece0b842ac8fc257233e55587eaca8e788d0b8b040118c2b7eeec8561dd0d7e0160cc1598a8628ff1c5c9f65de4fc2bee22646b507e22f9ae8037da91e6e805bf9e00578ea227aae16122e796311b3a45e6b12fb393ec3eae99341df170a5bee7131fa955b8904d5beb0e8871ce52802041df0dec9e17b8462690d53ab4b2dae2c67dbe7d6c88d6f0ae4975f893a658d76e38fa940669682f03a9bb877c19fbbce050fc9bd702132d37f420ba1a7b06c3c8b8b7511c3dc7808dd3ed91aa072565876ca55b426ea69432ea7751b2b6c6359df381936f0c8e79c249bdcd36c4756d2835ba52fc01b6ca6edad2401f0d834e313d685cadb42ba961018a68fcb6b947ae7085da884a70aa8f675508f634d251269530b38a466b2ed9837185adbf726120d4f90ad23ec2a92249c26986b74bffa2820b3f85c88a83fe321330b656f4626adad3412486fae48e87165ca7948eb518ab8f61adf19610d0f9a391cc2fcc3e778051f628107f7b96118fb1d075d8d15d4c4ec868ec3d4abd68c0137c815ab6ccb1d33ff6d4ea19f2046429943aed53214aed4337a51994585ac31b6a605ca6ee19868c557baa99af37b80a2c02c24ca9fc057c1ec2d11b2e91fea4b806dcd6e54ec82f45dab36f3da233bedd5ff5656dd369617f9cfdf7d7b8f1478fb6e9f65e7a528023b49aad2d1d3dbe4ce275058afdae27670fd9e53155f341719209792d0466a7e72eea87e6302b0ad2536d30d1e1c259cfc1daeb86ffefa044bf622fe3433309fdf29c2b41ce76f92228b932bfcdca9a0b2db34f146c1e7026397b9f50f5cef1135401a193edf268d0dccf42d51348fb4cbc15b4bb1099a3fcdaa42bd5d5127ca050851d0bc818931afa1a6886dcf2225571922de4bc36a23a5b33d91f586c242e48872200ef5b989321826c1429978f031662032c471e7722399d45a2937856dd12471a06a967914911d3d8293ea8ea49d5376d1c229d64d350e2071b11f8493cf7d76d24a6a27f665824160431025af47a5b372fc7e3ff10aacce9af2f61b7f43d3ed438073f9150263a2f3886aaff133c3ac960671cfff829c3e1ca1cdb1f6575e14bb07b00a2ed9518557951c5d6d447f6ea7bd5cc3e4ac2d38ff2efb2cfb38170ebd9f608e9dc8d31d2baf6dd6f50ed3a88b4885d066618bb8c2487bde1c71d60586f975c56d4198996af1f96e65dcf0187426929eced3285e6282ace5ad3e0362da890baa446b78ec20171302fd59440aaecd611d0074b80dfb4eed8456d7b0a69bd475e521a2b348685262d6031a12d8d4aae0610dadd49726fb0a3184efdb9c38bd6341e317ed07d671aa2af90249a0c737fd6214b003f649e270e5cf7701b4786d1eb637f2d1a6f56dd6ef537d2ed638ce9996c5638e7b103bb18a6a03ef406adf0f5179c8677bfec627157e83c2674bed783224a728094bdb5199962cf328d6868b0a4a57a3c323b278ddce92ffc43407a611688b0f8e5b51104164ca5a2cdbc53b57de8b32b8e21a2813ceab3a9466c9f7d5571a9a9fc6b568e799373756cf902ccc9bb3abdcf648520cf35cbe06c383cc7305a5f6addec526f264e1ea874dfa131d1fb21e8ee091109cc1e8055ba77e620206ccc3bb8630dac47d923692e8a54c8af2ecd150a07c8deacc9463d1bf2899fe20c68a2889a1b3275713ee331f5c06ed59414b10089d7509d7991a29cb75c1c841467b21f854928f9f67e5c5dd08446f29c9d75152455e3df317f78e76c5700e3fc211f64cb0faeb1cfeddab5ad9c732721e5452fcdaf1a91c3af910993640bc4d3cd0cef7283ddc58ed1dd1922e4edb21d6cb51b9c16a5e70bd55391d0342070cb305ccde4500cb06fbbcdf2a05f6d7322d8647b6abbee40e1e5bf94d34eedf558effeb5528edbdce160b15aa78332911e0a75ab37560bb8486fb0b2b4ed016180f13599712837f0c8c2a3aa9692128e7306c3286af35c5e8b01662fcad20187fa53096b17b3513fe735d4da2c44c4641d52bc4a7fa4e15c0f784d9bc94d05497f1d97ead9d287acf5b9f75966be518f637f852b06a86c88f7ea5a2993ab5308eb54c892a24b91bbcff8642af101a55e63c307a62c41d9c5b3e9fbde975ff6bf5074111749ba1d5ccbec57f044c44b07d29653f5d25a79c044d370ce3074c58f367743bf62471f034b58055fa2264b22e7cffc6ed2a76bf47a98f00098c91181450b40a72aa16ef7d9a9cfb4b48d6163fee1f75a54e40e508fd46e99afdc0a47017ac631964438474e77076ef895b29879cfa61a714d5b799c8d81a0531d87b2c53bc4fe2ae23972d23477d659898105a18e7a5e870119702bb69446a9d1c871b53173e2c0963da80288836512bdcf656c2595b27ac73012b88d88fa5903fc739a0e74f4c0ac662ca55cd53afa0fe795563e610c27f0c55a9f976d1f174fe8c9f8989f1e3d59c85c46cdad8aa10127585b61fedd866a26e0dcd2a8b0f2796019da69648cdb6e9ad9abe3dad6156e88190b5a0e70766c617f814ff0b5b34ec321e33cf85a58baf6cceec6f0b30819ed64bcd34d64ccd7022b62975f1268717994b130923e1ca95332f8f0c9b528abf00fafe40d5a665fda62d89118bdef5e5823feedd9e1ab6083064ef8618e4f3a255eaf9c6b12d9ed8c5bb052e4d2e0c478f13bf70885224654b2d9c938669db8b339cd7fd9a8be5823d1f072333779c0e18e4a414fb60e976894b1e6ff8294ffb7afe3ea754a66b71aebe2cbf1be194535bad9c0a2de42b295c8f19ceefececab22222f2eb5898440e17ac6cb96d906f52b7dab38ec332e506b7850f2f8d7fcffb5e8b768cfbb5a9f744ed671dd7b5d4e1e882e73262274a7bbc031f0c53b89bc711ad744a576ea59e15f436d4c5161a1ca7cd5dc8e46f98851728908076d0e6b8a0efe2ece0843291594de627309821a064110db374aee522fa0b39657e1856dcc17283f4390a450224cf1bd8d879a40bc3c01831277fd7169f0df118697d7d1a8a0ec10429cc48b655bcbf5fda9ad8916c97a0d12cf7bdf190b5e3d24a6b6b420281147843de9199063ab135d50335a9f8556c6ba23e3e66d876f6855755423f038bb1c768168257c59a2e2635c0752a9d31fa02cbb4414333f5039d44369aef8ef3d269f748ed80a64add76c022cf5cd8b5eb37d566976591fce9bed7b6a444ac81234cbe08f2438c33c052adcb728d395c8eced766e4c9fd35b8872914876cc901c4ad229a73e084e4c084a7910d23fec1e2f0267b47cf62b875b33378d0b76ac7de36f8bb2795abe2790b21394dd5e54260eb1a96c6302ff8058155dcf25008701841a41fdbd870c69d9625d012cc67037953fb34782e57a7dbf95a3bcc4ac5420652601b91ace298b8c0648cfe9ff0cf480fd43f31469d8215202b0f0d4971bd4a7b28175cb92b9ebf57b83bca21531cf9d98ddd872e18c50d0460c1302167f98182b20fee45cc61dd35ae07f7f2621737adf8cd6feb5807483b06aca85513ef392e218c4c0c8a86454c61dedbfe9dbb15f9f00d9c4a5423272d4eaeb27e21c53c2b8a8e9b9a79ae60cdd389b1d91048326a846eb8961c20f2c621b8aa5ee59aa1592ebc422e721fc6b0ae84b1c67fdcaa937652f9e680064585e517e0c25a001dd73e905da2e6309c338ee2ad38fbedd1d3a50b448f4a329a1d42315d9e18e86ed05d8de8c1d1c02b6747abacd90b556934c62a75eec9c1d112ab2eeac827d3e9ac709de1c144e17dbbdef2d53385625ea17cbfacd1a947e82a35bbbf98c319d33c9a26bf8c70eab6d8966454c143b51fc5e830f8af69678e51417bef35aaeabe575166dd3dc91e5a1f7ed7cfe152cc3f48d1a9495eff49a79dc754655d8b2c1c88b62f8ba92cf8dd58e8f2488968aae8ab064daba4d4ab5b75f4e122a2e1cb9dbdff16d63c68ebfabba84f5fbbcea12489ca28933e6ba139b55b9fc36cef147676cdc8251a7d173852edc791ebfc5e08d796d65599d625139c1367c9edd75c7af1d1b8a8a11803096eef1c4a14ae6f4a17057de3616970e156db6cdcd662c11792e5d965a3ed56fc2b3a1090270f61e14a4d341057e0d086ef98003d2622c3f545e80779b19c1007176d6ff08632a9c421f687a5ec1c6cda0c90d6783aa3726a6e7b46e4b1c5b6f27aee0f7f5d3077decea4a86b9809e9f0383f2ce7571f64b2274e0be12ae9a94da16fda5a3c65396e90385e4def407c8ecdee0aceee8ae8b0fdf6adbc28fcf29d6a2ffbc169447d4f678b84bff164a21f46cf6cc43967febe083e8dc3348395001ddd770a84b191aea5ce94d2eb3e97e1d441b8650404340c59c95485a588e73ff21dcfcafa403799a5a273ecd887821b3fbfdd0524cefe2b05c46eb5ba263a3d8c69fc0a93e76ccf7232b844fedefff96043180176c74b0e9d7f01f003c4809af8492e387b63cab45f779e2442dd2b1c0771c3dec626f3055d0266894126a5fdc641bc0666246775a84d3f41c1bd6e3351d315651921e32a70a505549eeaadbe125816068ad3774897bf888b1a05d0cde46b03443dd5cd85185c9159d89ea5c27709dca6175da663f217170bea38ef10ebda2dcc8caad84712dc2f7b1fd808b696168777fe71948bb2186cb00829ea7e6a010eac470fb56013eb5dad561fa1d8deff63933ac4bc22a007e114db6868cce404a474db24c7a02288daf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hac9899e4ba124e7641395d0e217055321e3eeb84166828faa6c1217dec2b75c33919819b7a3a36d329eb2cba6cddeb359b1d7b38429a749d3e0c3564c751b24e771b77c305bf907b327db1fbe3403bfeea4bdf53e2d714b96e3da0bfebedf57bdcac6819a79ce8316aa6dc24720989b394de02a80f78cde73f14ad31afda5b2ccaf7e762292974825e983e57673e2626741f60d4017cd1eb49463f1b9b9dc7c1c47428064a7c39dbbe59e8e124b470ae95851bd9ece8bb29dc65b69d1ba6a11d8b3fc524a85316053256f5fdd0bc3de1af6928d47a852d69545d5b71f22486f5852a58291310562888ab9eebb3b4bb2e910c23337011cecb03db700d80c7d9415e1afe775b585bf521be0c563d010e2c080521606f507e0ef40dc4c3c00e540a9988242803ddfaf62e0a4b1a82d697f4df4b55a6b8797d73001cfe3afcac32e687644fbf9eb2227efd2313eb90320b11718e0f24cfcb9ca5dd874bc6a19183b862ed73e2514a581f565d30081b6bbbf2fb0991266ab68ac236061bb76b30ae38b33fab1aa97567662c0105db7e8a41aa7a8f09d900a024e7205b188091498630ed011568c38905cb743730175de452c98bfc3a422db5104ffb3d5682168101253df9d1c356fc29d42299bbf6e9ba94a42f40ec2fc9bdd4b1dccb962bd67faa7b8caa16fd0d7a670af684fd17d6d38e2c457b71dadc9dac3e78829a57d3ef32c3d3a0721593d426686d44a38c397efbd1e2e1b4926919660faad893b64bccd5496b33f63630d901833597d49df47b8994285f1be02b57667b876aefed23c864d2c9fad8090392fbad12c80d53d0b9d1f90d9e9627fcd3fafc7d8deb174ee8e939dacde35ae431e5045db324503d605ab6631f74e7db7c1a0c300c809547e313265d334a3a565d7cc18e7d0aae0c10d7a9a885df63b16772071dbf9d273043d69525cdb85fb8d11f3595575e341adbbade33c9145f0d59993070b66dfa50b925c50acfe79c5e27163d69a90e928b9547beb0e04b60d76b399b676c81b5ee3f2a3578660cce13468380ce870376185fd6a943f1d7ff7601a0c17701b3fa88107db60e8dab10db0f3be20f175a11fc05133e1ff36dcbf68c6666e1a0ee54a40a360cf8a246bc9380d580b1f65b8044caa0398853a9aa61010d4716b131a5f16607c00007d896bb4ad331d074ae9eb76d0e759ad75d2906582afe8c62984a6968b9e9d18c00272bb33d89076b128d8552063436d0f683c7b1c2c66a0efc99397ee250e3931ee84471ec15bc315f9a901766ea6c4fbc016e78dd1935e928d35d07dd343d6391c45873ee8fd0fec69c021ae1eaa9cd7e6d91fc391052d766cfdadc4e212c5a4562e7f4fd1d393c6eb9d0867982076bd1661ba65447d81226f444c8e80714fe1a1d6777541d75687d9f04b94a7f9edbdc2ad49d55e76cefe5d99d6edc620c642b3ad3ba96e63c6916d53beadab5d91026327321a760aae400be0418d2a080730280cbc659f2bfc5435063b18762dd6a98954a50a3965d643c341a5cfcd240222b4d52f07df168ab8beef929c3929a85ef95cb14f31b63372183a2649472e3e2775f60b1ad214c100763305abef96e32bb2fec41fc3e3364488ef810033b68903cc4b3ad53f730c341ad7b383efe8ff665e21ac93348740452e4846355e91a2a56e95764fe536bf377772d4670471a962cf96153ff89f359a3ebba6167b093d77de4ab6c83c63b767315c28e076cc32736d0a4211fb65bd666c2d97cff459345ce2e17f6bf8d0921c357907d111d32f41bf27ee8af60995b859b0501c346dfc1f57b8adc208161cb13ce4c4516b74715606ed34a196420e2932a204b3ffe8372471e67ad3ca1b3c6215d11c108259b9ad82e726a99e91853c56ceccefbb870b8989b73401156b6e28ab05e9f1d2110c97e2985a81c3e809994543d86239daf2aa33c256b6482d90ce17729667d99c7a758cebebbef97a68aeb2ba6e8398b3b77c4589e29e5685928be94956de5f278432e40aff68844b10973bebaed9f7d160b5bd197eb9d10ed9480e28111c1af5470b63789a4e40128a0bbf7d596a8410ac7ec605e82d87cfe09265848a18e80382152d73f655f1c7aae697043c24cdd8c2f411263de1e67af77a110b57ef11a8b5eafe3c7f3b1e109a8d0cff53fee9d7a8951523a588133bceb2830eed69b526f216cc17daf72635bb0fdddba01dacb378ea180d7b13c42fe4916ccbb8519c5b5fd100523142357436410665856494d67761669af47d11719e3f71ba3b1ca2b3e29f5285eb0a71f9bc7218d520ced421a5326acbfe712bc4bbcf7a3509498c58e5638f20587b2da26991737a517b59e1f09e4f7d8734c141cbb1b9a41355e0c821408ba0e406e859dcb5008f069827669da77b24a31e0f044904f87e27f369503d79d50c0c3a4df27a3f8c6f7e17b7b82c4dbaf0ad74f03cbae806287fbc1107275acfc19e5389f9f671118e40d919be8770ebef3aab84f9e83efa036abf5830555f647d059d6578f4c1928c6157a518d57e2bc8177aa1937445fe0d877c9c861cbb5759c320ea80311768d7e99b289a8fd213a0bae143946c7dcfd46471ad5ae8d4355ffd5f3a9a0ae0110766d88cf4c06f5a939c6d4caf27409be97e979a694115638c2fa176328f092d1703dd5e3baf350ed1f7ed4ed126f67511c5479c818bc32a582672b851655ccc613930dac175d95b893ce507cb1de38b1b95da711b6b3c114c86afabbba4dab01db4b288ae0d3c4c6f924e0915bf42389cc74e0136f57c24d0d12d7179fe21c13fa0a7c898b09ea7e6da2b14c346d27ba3ef73d24cc3c9204895d015694fc1191e7e6dc3153ed7dfdd848fd12493f8137a63f5b2011f54663f4c580aaefa8e2b66e603ab6d69cf6ad606228d27b49a7423425a2a026f2f1387833d2d1b8bce035ee2a26f2902390a078d3456d9c9b943ac9e29f0a6543d8b53988771a9d352031d16051dabc3cecd070b2c59c95a668c698ac2c3ef2d2ffc71b5eefd614101a5df195a6224131506f9ad83095c312816622e3a07cd75b2f7ddb40f2b1384d8b52ade0a53b960d6c00620deed9fef594731d3b744880b490c302865f1f483c49b92fc7d519fd8283b01490fc7e95deecad63d559475ee51b311bc2743584f9328d1d5018ad5a394a61ad9da4c86f999b7e0b9e28eba50d4a4f835904b41a4c0d891f30bc911b15b6cf53ecae7a04fc0f636418853021b1cd3835cae2726e9e389446449878125bc209b58990e86af43ab3c7b90c4506b28c77b5e9d5c44dd273582815230617eba0ecdac3d314247ca26757020ce42b5f9c536447a01802228677c17b4edf1e54e2151e604e9b401eed701b289a3b1b632812f5ce2b5c8e0304fdad4d1e2ae749daa8ef29224c22160dcbed7c700396b81b466fce19c3d074f07dd1f872a30a54f0b528dbea064279bf14b9d89534a74c40175fa8cbde375dcd13b4b9993f8d0bde6cc6a94dd05ac32ac6c9e3ec337bb027d12f4f65340ffb8d2706442b594b081e907051489a17d0b7fb24583f6b258cf58866bcc081eb664b1ef1e2d01add080cc4c2670f55de194bf7e27a9bcd3a2e9115ec57441b7ba7b0b083fbaea141f43bac9dcd32e727aaf4568002e9e8f66c71c7c2064ef35eaf8821e4acf2ede8a0043d3f78e957be7eab396c7700510b13d471bfb7b58768213ab00d9df3d5ae084c7f28189426cafef3e201abad8097d488b66dd85ee4cdd048e84af86d06a31049c1b3b631868a190ec8946bd56144e73595bc87b7b351c92b809faea00c11494f99afa6e8043c36ee8c01af1e2040c3607c1a9078611583c2568ced3c2303ab2f74de9dc8ebd106607a2b31d641c3a973b4692a6684fef13f66ecc5e9b381400e28c2fb73aab125dbc9e47f652cf80c6cf0de9c59339d0fd554db17ff6ec31b49fdf507b2cbe23210f5663817365710793c4c53fec6f7145ccf9d58bd8515132a40ced89e8c0c35f44a8d394ef475b35d2f3635d3a2d4c2a3b690ea438c5e99c0b126bfe2a410033bd93b8154b6b7fe68b6ebe0127920685d181d77f0bba253a2261f2aa810bd8bbf56780daebd45cf7dfbd173e4f725759c40998bf88b355098046fa0c129e477fc8d5990f71b20cd249c9450a582c3cc1dfa31171fb2292ef62ae3d047ef8d4aaea3660f0c85c4a1a6eadf95efe6db5114e6841a3628553cfca93e47669c97b525dcd43186f4b7c816cace65cc217f0ec31c20383734ca821ebb916472103add28d2c8c7c27b5ffd2a599a9face132184dfc92d0af17259ead48a772867d7822c5a255b23c588a18be6bb20e4455695f68b0b25c9aa81de6b9c74abde3f443d45f7f7c82076847aa6c5be5d73cbdfdb7f6e29a7a9d4743d28a0de421fecba2ec8ebff127b12c8f084605738dca173eb3b717d4c8bc820bc5865c2f9b59875b8f92c8c9d4b9675e6f4ae1c94ff71ead1cf4e2b489293271659cbcfcf38e480b89284cd80dabfaa219d1a3f223bbaad0f93dafb4e4cae9d398b35886c9a2a543b114b17d013bf35ed8b644f10abe8691865c1f06d4ed49afd0420abc0d415abeb07be11d270bea46a3be53cf54ca232bb3edf376072265920c74bf17bd4eff3b5c795d264819376858f7145cb17c3ee34ff19ac9272666010a98c8c4be8618a7a56b31911a64ae2e234eba8162e8a7f1813e405f049eb2f868271ef88797eb81dee1284712d45ec6d445a26a8175dc4b9395918d703114184f757c9f07d7ed0511426175691f9caa6e0c9cd8d8b48a8ba80704c5a2b848d8cdffbdfe04bf64736ad79647c7df98cd4d2ad60897fcc05f18a03580e6b09a93ca862be84b5f7e06fb4291161fcd9224f0dea1d3c32472d573fca44edd7cf4b8f3998438062b574750925bdcec559bc04012eec16c164d3581439e18aabe55cb0fe944cf05de600a2c671d40e1259016c8acff13289a82decb934ca9c389ba0df14d8ef019f4dab425b42100ac36770ceed78f1c7bb52152bf0b0b663d68abf37a217a157ae5281103ad8a20b513a57cdc56caadb683ec0f634291b6a6e611bedbfdbb75fa5a665b4e95ad3feeae03fc9fb6166281b6bdf2e7130dba825cb0976f587c1830cee79016c06380692a817afe3676b813bdac04292354da008e80c710c56619f1447d8c84b6e7b2dd1a6a1ed75790e601cb6a9b79c00453757f7e24b0b6733620576e746becdddc41113ebcf8653a0e0e8799db483c5d0d11c65fba1290d950c97421eea99b14f87f5c22d098c09d04cfbe086c5731768cd21c422db511db2c7f18718b64e24c26c2503a202723bbc36a88f497843e7197ee2cf24e0acda0f2cc96b79df68bdcb603b0066c7438c2e298b4b7f3ea91856e3a276e9555d74380e037eadd36ea00ef3548af074c49796a0ad02c482c012d76021a60ce1707826929769e6a5de2bcb7468e4ebdc60c5fae3c4569122382dbe697b3b7cdd9ea6eeb1b19bdbc819654691e72c8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he157c7a8203e277b1e4cf436742e585895829325c7da5f624889ab6394f509cd424cad7b35a83ee39c0a7b199cbebd44cdc95991edf7367ade503238ffdfa3527379623b81bf14ab92b7de55c5f6b0b785a50d9244cb781ce2be0d7922313cb80b5e1abec5e63bee76e3b4ea29aa59ae872057693474d817df833f82710ed3d7bfe8f35020a79a78275c53364a8dcc4af881df306480b371d165262591216fa0016743e5220985927eac0a8f009c4e8a717426f1c12e8f90a9d23fdf2553299bdee5111801c646d7688fb9ddd8a7a0b24e44c40db6bf977c4031732070e3d98328768d7f7cb96a233c3a95b86a447d6fb4d046b599fa35272825635eb99c3572ca09b2d96bae54828c99d3e8a185541d0e0ba27cbf16652bd95ca5ab99b8307f76285deae801367ddcf0417b93ef9cc6186aa5f30450e1f50906449ff778a0b5b6614bead2d2ab63e9035b266322fdcc8d54627b7d6574c4f6a1d4642ac995c86d9fbef9332b9f41f5e2d9b62399d03eebac395ca8f042a30760c4c53de9731e693524d6e04d3332cf4165847d6899cf47b4ba418beec0ed07e4b4fdb7aa66ab4380778e51e17e913996197cb699c552db2c5a446b83c1e8136910dc5009e2a025cd21a506bb5624a6281e294d9b1d9ee98df1bf1b9028559084955b534dad3233105318893871fa112f01d884efc52afb7a51a693e13bce0bef711d7e2ecd0b0d0a23964777656fd1470c12b2e18e40630550cdc2b3aa1ad7779bf2fe2597f05dbfe1d27f1657c62cbb42d79282e611093cf1110ec404fa1eb9a77457f5a5191cd4b66c73c41ec2cdd5e19935fb8c6db296461790972baae8559eeb00d61fc15bb64fd247c013fc22e05c75a89144a0467cfb2a4f8a34d8f8bd4c81a5fe17a936b9a2a00dc3ffed980b569ba55c90c6485a0e1e1e314cc6bd9ac145bbb067326dda4d30a64bbe99f95f475b0a1dd4295e7b637d0a778bac6261b85f38fb5c8bbee8d245aed17695dac4ebc28c9a91ebb15f12b38e6ddef2fc293e1d1a56668262ac307e22f6cf0aed770af34a712826916b00e89a1e39acebff215a0f2dc7ea51b03d27cc4f9d910064b8a154c41cbf71cbdd76851d7c59ec975a9652e843199c96380a5881ef85329eb77e80d2ad49f07c9dbba51edd0cbedbfac134f0ab93721976652492e0700583702bb77602e14340e35d2d65d86c5c8867cd3ee069d4018f9f394021a2ae0bd2d4043a24b429884288f9e22b56c472828e0575330ba19051239a5da82b542088a3caa197d725abf9a425704414e7771265847c013b7f086d2b96f5e3d29cb14b8a1317648a961378a066c8d26aba185e82e6ba362c21dc4eca4a91d1cebf855d1f3faa3b06c41901ae832cd151b28039bcde71a05034590b6535d4068a69be9f0ec6b574d2ea76a1d0f707d298574ee0f9e170a7a860d4d7ebb90ff667b85e23bec66969440424a3e0fa200f52ff215c3a6db87d123c10c6f9e8b6a6c3989daee0255edfc35aa4967d7e75d47bc3974ef6e2247e1d3a0c1929442f533b4b72689780eaf50ba8ced72c62e05ff2ddabbad3a4aab1aa4765414beba471fd65a6508604cecb405f34bfa951cdafe62074ac78c6dae44ac7670d3ecba792798674579d9c5e34ebe9876c1deb75c84212d6bb08c3d8256439b14ccd699fce44ea621cd2508cfdea15ecf1c586e0f322d87754fe3a4a74395535c0ad9307ba0a7e47ee4fb8f80f537d3b0d0fabe957e918594c87cfb1fbedfde6a6117e509eeeeb5bd79c2af2f16b18fe61a4bf99398445f52874fb4d03c3ac133a3cb38dd291e9610ea88fc4e2a336bb4ccecb97af8f32b3a91936422027506b6c08561b100c228c751db5c7c8ba9e337de7cc5ee4acc9752e0dff525f9b12b58342d1d2c5da5755d6de755bcfd384fd15b4a0acda0e920ab1521153376237d09ef3ee336bd832763e96caaaec663bef5cfa78de02ea7ea3d6e71b7d18aaae9e34892fe5e65c4650b13d7dd3a9e9fffc4ad7934a92090c4eeed90cc2ae9ce0c3ec066c6b50487ae71bf11921fed5402db58eb9b056b4216bee4ecab4eb85ff01ac4c673697bce3f5a69e5c1a1bf8b7024fc6158ea4828c6ecdf9323a4669d63e53fe456dff6affa0957106cc69d655dc1740fffc773f877282a6b2a8daf195fcaa7ccab9126bd67c4ed6ad5ca019ebc7ed53a7bb14e030862c0ed0eb473d01f5e076957283fbfc2ea6513b3d7211216cec03ea4b63a91c1cbf17abaa1f51798261309092c3d00218721e5dda541948a84548dc3f6885076e1d7d34bda42a7800d39892cf4486578c746f0f4bae7b0c68820992360a8bbead4774d279484299812e72bd769fdd436400595bb00d2b07b8c30d15aa34243d496d3a7414b44a790d42c5b3e02f389d5ffa5ed1334893acd677b4e23af17dbd7f1fbf6046470f54bd2505e172dd98faa1b98587685d743939b77695e182091d2c30ed811cb65287a56a1c7c4ee243617677a196c497dac0d4508a0718d2a9a75e614d4a11341cf13975d03685b5703600945556e4365d93bd1f415ccfbf5ff1ee2c2887394ae7159b6484e3590b05e1c1925ad815fdcf10b46f8285382865292a0900307e93f0583d3f12fd76fab94b7e25c1f01438b113cb9d8427c7e898725b534eae502358bffbf16730dfd7d36c60178e154291615f230a6d743498e829520c7ce50801be9073182379a0ab8e1f47fb91b0ce675cffcc2beba340bc31f5be66d6eb843ca36354eeff0c4a810b3eb2800ccce4ae4dfc1e5a288471faaedb9b12d8dfaf9f8718e0939c738c50a8ab7f36ee3f3b37637e730cc42d94081507d195ea7c703f76ddeb3b0b81b9aa103bbee8b9ef7e16028e2d17e732aed8b7a5ddba17485c00e0fd28fae66a821370838ca3f0e6a2bb804bb26ee8758d8b929c42244f1e4d0927a6ee992a93f880532016f35b9001fe01de5e1191a76c6759afccc717289fc449c6b84490e2452c4ee6138a11ed49a6e3d495af44725db0bb92e29e769a3a56b92d81a39f11c591a670ff1f8831d7b84900753ff991bba6943a1098e2daeebccc5864bebdd99f32bff4a7c27b5a60cdbfe5029edeaebc0ff248269cfa82796d1a2ac5d77b562deab22ef594f9e033c266780a1030aadaef55259f8651258af6edf0f8874d35b4e6c5be18422d0113ada578aa00eaee808176b0cf8f4cac6fe74039a6887a4286b3b8bf497cb11363b8d51f5394503ec52c8c94a53e294898d645e7cc30d0341ab2b5f7d297bd19b2eee79d42968bab1a05b2bb661d1b8c7d2a407ac95c651f4fe51dda0c386ed35127eee933883787f5cc9bd5ac87c30a84b2fc7d973733d599792d2736e6c8006b117e642d4143f2537b9a49668de64a96671e7b6ed0d9b79f7de7629193065789a0bb9aeec6055504c27f7dd7c10c834f6ee2355ee27cdfe9756f5f8cc4e6ebda3c41e1805c0ab08eb660fc664e85f158efe9e5b8f262bb80a75ad2cabb42a7e796536dc073082316e1fe39ce8e538b81eb7b92b9c625bd03444664757997eac3fe4d19f201482068f7f5e5e30a7f323305291dbfd2d385a9c351c85c8ab01687003a5e73bac5c051a52926ff1e50cf81edcd366a5cc20bdb046f2e1b3345eb640f98df6f0cf6712a7fa562472f89f31d6f12660b70265fdbc2269370ce159b82a42eeb87a3d7f768eb026730d778136653ecfd130d9357676a80e07b059467f87f3779b6840ab1926f1501fbeee6a44fb5ecce7d06054547926441dbad9552060b3683ada719daacc132ca896047609264bbf1614538a09780c7094d39feff972c78252726d28bb882f299e3c847a479269f44e5780babea55bffdf6b5c998cbf26683a8adf01b6429b973e6cb968af8271ee5019f5e47363e9b4188ac3188d13319d0f272d8a6b5d5ad3eaea83335d5a56d7c1243a21ef6e0c7fe1f7462f8c40ae3d24895f3b3b4c59ebe45d6dc36b6675092c32536b757e0b9bd280318a2de647cd0372fa24cfb2e184a745f74cf01f3de89fec886ea5832da8654bfde7c9b915b528671014bcde73f6a5a972774f0ec178359581ab60125f0536688d523393d4626d2ebce8c6a28e4dc42f1f1fc0f50bac30037f9f9885d93c5145fb597b26e831d860e12e2f9ce4821d36f8e8cf046a54026d75aea4e81d7bd5290692eeae401e63e86c64209f85b5ab1318a172da475d11be0da5ccd976abfe08c14dd70325abece2ca3316f7d0c7eec78fe2ea814f3152c5ae3e2bb04029630a01737290662dccbfca8aec14cabc375a91db4b4b0f8a98b2689f50ca08a20a46ae788cbc7fdd453e522e58c4098a9ff76497f8471b45e4ac3aada15b9c86ef3b90a58b72447a2e454fc3b325fdc6b4aa7af143c8b0743692f6035c9a84945646122b5c2992318877a32eb9c9112cea1eecdb8579f1ffc0c3e1c9e55f062b737fbea6a1736ea7ddd20150650acfdd59c972a2fc4de1a417755d861a8256799ae1f8dd3a8b7ce04eae1b1cab3371634ace52dc2d68cd0f47f408889340208ddd155e62824560f7e9261c715f37f44fd4a47a809f9168ea068ca502b4acdef160233106c251d63a610f8c684ecf62f2d525166e10377f450e86861c6ec895f32b2b24e6fc1bb7cceab94078d592716916e3cae1693da96c66e823014d3837d501d47e577bb93b1a78c069e55274291a48e77140298f705b4efe0d33268a7cbd716aac45ad24bdb5df6e9621da5b65b8061ed4fb5933d952385d1680d79556c806e4ecae56cfacd876a0ddb482231757085e75f56cd198675be19495e9a295b661a5f960fe6b90d04902db912f8c08a777717a050f243195484b1b8cbb491d5617ff40e957461a883e4828b58d19f17fd1da3efc2324bbd09e5020a56783fd14e52e4cc589896fd5f2da924ed4d202ada1884992b5f689ac295074a7c9845c44c54820891ec19f00a431a27ed51dee42eb15ec759ec1fb252fcc3ae69d698d71c83374695a3f72613d38a7d671c9af0ef6f70e8424fdf0beb368c4f77e7f5dab9eb5ffea9eb8408baa7e8aeaa65c541ff1d379fe34a3f8ffff34f1d31b9c8a0ded20e8188a77442d7a69ebcbe671c6fe2501fe0e9fdfa109f03f27ae0aa152d901c8b8826c50bf6571054ed2b31e3eebf655c95240142151875b1bc7406edf3c73b64592c757dbfe45b8138d8870d0b0a170366ebcacbe8050595f190f377cd1f4d64192c5b405dd9d77e8d63d9970ce1020a3e0c4592e9592761b6d92af6b5d4ddd0b273f19381c4f16bb7a0de15d107eb3c2725b4a43c5b7de3524fd1793f55f5bf07df622972b8dec6434b644ed01277c15b7cd525219efe4b1528b4f4f533034269866deb3a29cd8f08975928e4c811953bdf61ac69e0549bcfa518628e744012204771cb6ddde1c7c8b9f6237eeedb5fefff4deccead30a2d9b9d9eb9d5a9cfd6bce5f92753c2637c616dffc6d3166666367c4401d601f3d94a93d1ef8f230d5f52807a9bc10;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h70b985b757aee7279d7e27cc25c74b04c86c35a3d85e4d23ffffe12d973246b4b3e40675d4ab4fda6277d27266d3d9f83a98020b7f4b52713a3acf8acc4edd8de2dd0cb124c73df78c7245a60feb16cdb9824d70ff07c074a190505f6ec7d7d0faf6db9020324ccf6be2ff913b1f9d90c40a56b7b373358b00bbb7c8ac9081132e958f243b75368d3c4caf4f8eca7803a6242f11321d7270e43fad9bcc2b077d48191b25da9f056f158b0c033663e8c078164b1e6260bb0014f3d14d6de007de237eeeb6b93d30a8e124a73b5b67948df7ca35092114cb2937d159f8e46a37ce0889817ce6dc175f7ef4f73a995d304150e25ea0496144abb1ee00944c1ec937f068c66650c2aa60a64cb1b72c833e64d4035bf411f3d0a36540b1ad193cd7a6e9fc8324f10c10e560c93561eb7ffad4e15a16f82d587fc455c2a5a8614c41150f5ea904e24545423869e5bbe870f171fb35f89174a872f20ba1095df90cc049532ac6fbd85b5fd6234362814b548fcfb0adc8ca13a2a092c72e97021efd697c84f6b6903e40be9796680f420967cb7480022b943fb16e6066e6ce041732726a290f8eed31c0b8721f8f9f1b9437c9e276eb3fabca0a7cceca9d662fc7c5bab564ecd2a2eab23c1c09490cb848b5c95055dac4fee87bd426ee6e9ec3858915dab6fcb212ff54ec41e3de4dda9de58bb41f9c42c2933260a7200a7edc4c5dc74e2e493393dd2f9779bf1d8201332920cd26e720f0b8c8ae97d07623389528f151b8287591365a52378f7c5cef4076d903a15308959b27968c6a7a35400c47e0f9fb7a292e5fc0a0bf6ff86b16128d3284840839c4f1c23a9f1be50c2a7c287330d888c4a513d98f91adcbfd6c164b8dfc6214d1ab69fe2c2d4087c3fdd8b6477dbd7b23474f34d5b9887d44c95e4b3403f5506e411dc538274bbdf3b04e805622be90c3e6299dd1b7cee0546a73c7ca6e8e30ac378d582842e4eff518e92a24cd0e07f3695851aedd2deec533384958328701919337876ff891ab083b6d86e0a9da98c070360f20b60afd5d2f5c9238c491c72be280f508ca9b4dd06c8b1f9743687198a157ad6ad550433d5869195a4103440fe019916cbd2ca0819fa2a685b243b97013b6eac98731936f27af259791ca937dfa9eed7a4be33824aca68e4c61b7136a35f5fabc59576fd53725d43adb495f55f776065551c955618ca21e2bdac3972d6366c74f962400a31a03eec5a77bb3d938a90870ac7b1eb80b2dafc4faaf517cc623cc7a4819bd0f086bb98b985cfb7fc52319dd5a04cb8215b6b876199de119ca80efb3c5a11593e45131056186950999b8a738e1ced1dc44002f8bcb03a7d5859ba005908dd6f16490d2aeff91639a3907aa1eccc8ae3ecc506282acd7ef52c301222d4e6d3cf0214693b149c0739adaa2fcd85bfbd23095b4775e6f536cc247b09b6a8691e3ab80999200d4fe407323bf7b30634aae5eff15bbf6d4a63af1f770ccf3f732380008cbed8854e13531bb4107e9ad6e8d99622b630485b12629dd69208efaa919e2d0649e2899c12a2f0e6d192678e3ccce3b69e051a7a10d19bde4920da548d5bd62b16c3630efc421be8e455394fe343b04cb659115a6b12cb2e048afa47d1d283d3fad8a3b3f6fb007abee22d7a174abe7be20b1f1ebc8359e29268133838ddb33758661294598af526cbba24cfba8d2d56b4248f478d9e41450aad648eaac2f47191f4af6c2ea450863d6f9697d20459952a8b0ba1875721875853ac7dd517d8ed5b94d21ea1ca6dc11920bc8f94f9fa25fcfb01ba36cbed136aa8088db37657de4d2f91a7550c84da99810808ba260cfd6b505c6c8ec4794d1347d322ae4b20d021b60a418d094ea92d2cf8b76c707e8905fa8f2a62b5ad84961a3d913e2a6043950dde9cc9f66df5d2c30b55c91cb207b23fa0c27a80ef9ed871a19180ee8f428df9ac1c00fcf251f428d1170ff1658be20d4021bfbecc26c57b314b36e984faf562bfbb1e53c7f74369264ba166701db17e79fb0bcbdcb00e02e21bfcb3fdcadaf7ad268caea0837b8a03878482d36483abb22946f16ab5a991f0fc9da0233992db3387e9d9b18123df7f5ee8e71191b178a6d9c9c65678038790e7ff6fee22a839faaaf61f58170fb6c3545edfcbf3f412776e597120e9b7145a527ae12d080c83839140372bdfe325e25a159cf6eb9522a52b04fe854bc683b946f9cbd9eae47c10cda08db810de6d07812d06b72d2ee8d5e18882f1993efe27acf1f8fd0a49dddf4a5b4e4aac9a547b63f3bda7961f6f10b9725a2c8e9ef6d89cafc98d483e32f0a9baad31bfe5261913d84266fbd28b00cbed81b4318a82b547544158f79cba488793d6131d33093466db80144a16df8db120d64eee432c90c2c497763b8fb935853e941acab6a20b29acf2192d01d03f573013db78fbab463e4a223d660e48b462e8661de0b68df9b85d7c87a7f7140ebbfc0989b5bc8e9957970f35316e0acd6da3dae7de743bea46c745941da9d7f87ed26f662fa80b9d4711c8b98a3bfaab96e475630cd992c49e3a8e1d9429683af16105e3bd16f33fba76407373b268502457f7bde4e32fd9ec5576de7dfe7be09ca20ea1156c62aabc64086e270005cb17145014a1f9f34f27d71bf42905bbe7fd2cee2bd833338f78cd517fd4c2de2c572b3721baed6467ed4ea0bf1a2054633b657bbb67cedff6f4be8a9124dbe2907817946ae441109cf20004c65d72240ccf62c1f6cb08e36c816f276d701b799fdbffed1cff7e10e3772a82a3aefdc69a82f6bd752bac262aced16dd189d63db210076aefa2aa45b30fce3b97b1806ef31fd741f48934bd22d3a38350745c4c68e419045335f810653a01229e35c0178efad7bb54b85f140231e7021d8c24c6fe01df39d1b89c0fb68614d83723fd243644db7b834c6e5a9898794d33172378a14df999b41d7ea14c1b5d36015f43de611df889375f3bc974bbb647408ec6732dd05d20732d8d204da1b82f65cd16a01fd8355ab58a33759a02361096e9895ac399bc68776dd44dc3a11b496beffc4fdc235718986041f70c507bb8102ae88cdbd74be44be0fb125c87b5da52b57ea14f447898696835b4d13f222459141d1d39cb05fe25b6082de7faab5a72a4573267f845c019c43912d58309e3859d2080caea8415d199572e4044aa205f8f1fad145fd0c3d94a146b25fc1a9ca9bfc5299dadb7ec53aa6905b8e1fdbe28cb733ffb5d8700823f3c39429f22f58f2915b2bb1d1131f6585812adf2b83cdcdf09380c244e5e16142bdaa96f8ebb6e4e877a13485457abd885d9f88911847f5a4dbb2da4adc7873d2c7a1a763c3cff79eb2d56090b21de0a0f1478d97934d8086a01f35cd28572a4e2cb80c3f0b83e1d403f76906d3d51f7456cf1a6c5e715131f59bdce8fb48fff6c443e91c390789680b04590fb242e825daa6c5f1b6450e182b30c0dc888b7f954f0eb577e74e3e2c108cd1038aef3320824f4607813519119e7e38e439bee18815039a45eca24da485792cef7832d25838a4d75793fdd77ebd2afe7a97102eea7721529c3cc0f698e7c1e368a003a5e9aee580348a7f3c7df72be7408b26ed6b6b1270557d956d8342088be5ea62733b0b7e2aedab9d67bd8e64e3a76774528eb401b7997a4da07e3c7501cae5e6ae7b63be54525c148823189e36143bec5a3f3c721e94bb08f77159d412c69295abbec68911e1615ba971d5f3ec626a56e6b552a65d1724d3fb14f8f1b28002070b7bc3bfe498e7bed83ea09094feac1fed3f17035d203e79b6bc0489497aa60a9e2ddda07ed52a16de280b8968a9c660be3531be487c5c212994d8c40ccd2cfd91fb16f2e5c6cac2b466152dce12e1ec32a9590246c7c5a60de75cb25f6ab59ecb1f89207eda79b87e5b630ffe943b92abc8d6c8c58a7d2965ebbd2ae8cce0fd4b53fe4b8bf29a0f7384a58fed2adefb757c45d1f95a5aeefdf6b1d227e081350895eeeedcbf38f57d0bae4f85fa35ce3ac64a83e9f86b4fdfb4582204fd5b48a5e01167407e85f554df69f84e9d0af5ff4cfe094307627e5e9580299e10cbec67b8b3d1a8da5cd9a030014d183aeff89126ffcea3947019638daaed10ce28533743115357c9c5ba93093812877116f254abba6847c677a57c6eca39abf95947812ed723f5cb914dfb5adcd301ba77a6ea21e67cb2990fc196588340ffff35b06380c6a51dfd2dd4435077ac5061b548051ef869e03cc8c7b526136a23e478da9c9be70f1336e457c0210c3e071a3c21aa846c05c44b53dc21dd1f4d9db6e638402120b7273640e0d9489a7733356df9291d3ef1f96daefbd080c201ff7591dca8a378dcf965cec12aef099e4aea2aaaf6d0c5e99a68267bdcd7d77e64c51ab234230d4808b929720ec3d769c28b246b48a854df6ade1af446cbc20f5725a56e4bd0b8ed9f6797a513057457e3f38c02c49b1c7ff3b324e46826615c37604ef74d0302b705210bdd6236bebe5845a0f17476821a9d2f371f62bc2e3cc06b2dc8fbeb9d8d33df91d4b10797d3ad004b711bc49e238c8776c6804ef800864eeb4aadbe4bd910606a5bbd7c71cf81fd607fd86206a497fc694153db70db2cff8ff9198496e7caa126830f4bb8d14a38a987fc714c6505379ee1874d604a816ac9832efe3c20c3b620ebf0591256cab422c02a2b217b8177878922dd9e15c88827e6feeda6bb8735ab834ffdc7bea15d21db63884b71dddfd65a6728ae84511e2e0a12c7f7a99e0f9f9ae92d89e16ba52c4d7fbc504b0575452fc82d6b8db88472fd490e686a87f5f76ddc30c0fc50d6285fe6c8d8aad1a3a1cbc5f83ed605843c0f3f448639677c4fb7e572c76e8a078bfdb62d04aadb76e6199200bf23ad2ad5b0644ac5809b16b45a46ec2487f64405c4f125e646209ae538f560a9e043a9b0a463cfdb5e9cbd6124ed7981370941f4005cf063a1ff5173e364459132980a73413b653dec222f535b7648219bc9ee74e875fe4a88811811a5fb804ebec0780b57d9a3f08fd4ad8bfb6263378217aa5c8fbc55e5ace68f5335af242d9562f010ad520f3bd3321cc2b51d2ad02424836631755e2ae9517af0a12598590ec46efeb40d331b76f84d84f3e3189138edf4b2778e4b2acf1d23a327199cb0ea26af539cbfb9dbf0715980e63a28d82b4e4a6167b098a69b6ddd56fc0745979222711535bc3715fa61aa7b29e65c5f125a20f5a0f4e3da74f25e93e63f6590084ea6b66c8fffe5b392a342a28f552970f93743a092af3c3abe6b675760bff8fbafcdc5571c2b3319aabedc61bf4d2862e1b9efb41dd7df2d4d67cb5f4534f336129855ef315584a824437cf0ba462add9680519df30f76950bfb5ea70f1aef34c067aa5d91660837c9756d77ec4418fd7ba0ae4ea9e5a73d32cdcab0bbc269029da21fa8c65f03f24601c08d1a9f193d7cf4c8e29a4f52107d10206710adc2aace;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h725e13cc96aa632199ba5856721acea9a78266986fbcecc60f7762014b4e10e8720979a33cd49c0bd8dea1f3745ded667630b259105a31686d663da95391165123c3e94ce0ef0f60bf355227481d3df467d4ae44763fb9715efc82a88890e4f3f314f227063ea072e3b54733d03828cd54f13e19ca9aa239bd947394bd073aa28ede0aefedcf57596368dddb8fa5fd838c59c533b06d1bacdec46a1c6d97ec3e17658c6d2e521621bcbaa5737c0dc9c88864d4bf310e3e93ce8b165c6ddf0323f39ec6cb61c81612db6f45fea327f24fb7b9e1c9877924b6f642c758e70f3fa78b3a461ad18a71ff30d686f83ea07496e9bd5d8bd7e83f1269433612d9d7585df872d14c397233d3cfa9a2a42fc73a5d2caf82a373e6db3a0d2c233220452fc21f07813ad9b6449fe440fdd616ea2e73fc310d4b3286eedd42be82b608ba0ffdd54ccbd23d5c5c5f351bf2ac0d6f94bab361d376566eaa6b0f7463d70170599e7b9c2d2789919dcf507ea53a9530b4d0398cd7d994627cdaa982f2039d79ae6158384f9a4f07ae4d78e107a5425d3338eb264bf0f44900eec2a0b042ed158ddff848984fda50b035c5cbf4276d148c2f39463fa0b971bc86e4aea4e8e61905a43a9aeb8a120e8067f70071d6f24d2be710106560d0f75307c447800d5360cc429efa03a21903ae499ce16b73155043d167fd8ff86c32bf50127c7fb6bc82444d4ca944826421cf2e7825ec1ded73a9c2be1fa572533a9e1f0cffaa0194385167fdd43387af911159b657aba920bccf43f49f626dc6bc623226f62a3da23f0190baca86fdebca266a1d5207cf54c3ab70eb687c8b85034d982b6a1e31f42bf5adc8ac3b5b3e811e618afa96371ffd917c2c81d1f2f1a64604fda6fddd9c72902d02cd674ee3f30a5d8d6cda47a594f1ddedac6f0fa6b41d4533e2051a24289304bb77d9d01c64cb5aa833d8121e0c7df9e6349f2898b2eb1b1844f863de8bfceb2ad22424473a39ebb451fa0a5118706b634e02dc153693a1c0bafcbfcb613a6f026af4f55d6b4a001809965810aaf8bf08aa6521e94c9c4415c3d6c6438b238150789d3ba67df741014d9291a719aa5610ab06393b1a109f7b381171c38e45d25b9407a319b8af9c300df27d25774a42b6f67bbbb1ef86290c27523ed7a1d1842d38465223d1d40382865e081904681276b91402c23ffbafc8e42d4ec59034e53850f7530f109f69ab0f1a0abecd1801493782df308c774d2cc245a48e4eb1f94a63d92c0c80d57ade3f65dddc24909dbc904104efccc18c024457dd2784fa162657851a5ad36c94ff0245b0de6766ec0b528befa7029cf667c124178da132502be18aa64a5d1d04d4ca19cdf0fb55ed23c3ddb0d86b88f38f9fe3a8b156ef82898b4ec29c4cfc0411f2389ad58dd85fdc3b28b9ba6f6e05ca1dc1cd3eb78a9cf1d6627798cdc2e9c494195f24d8f7c748d79fe24e890b183828b9ae7513e3e5c8c5704279bd5d8d8bfc6f5b5f019d6dddda6ae8309b7fa801e832f86726b25106541fde048da65189370be84283704ab2368e56ba5afa81deacdd5bffcc62ee258492bcf10b10dcb191e4b4d007517583ff108b5672f817d7dcb11ed51dfbcd495e94e05174d0766d0b2959b3724f6ba98f8c099fa6ce78630c7cb9a6b139b77aa146cee014d300059dd984d3201f2428db9f5ab34f0cff586083ff6ee6e485893864358addf8b7d873d93438d14472fc54a3c91d7a029cb375e510c567dfbfb5ce64f74b771d841be4a76a780dabc992fc8fea6b8437ab213915adbfa874a875534e36bb243a7fbf45bd18f7038afe021962e07af96e6e63bf9049c0f895ee85e0fabebbe0b9a18895ad107a15a52aad031f3f4713267d61053b4b273f28b832bb2656819d058d415d829ed53f749f0c31fc50483d0c2a5611a88e0e4a54282214de3672eada106bff2640deb15baa05127d53608f4bcb173225ec37bc276efed84b3f699c936dd90e3b9cad7927087f61ea7bfaa80b5fb1d636518e58b64cdd06766a2be0fff447ee04c9d23d94d999efcc1a6df9d495e9980c9cf57944b2b70f30241f14fe2bd9693f348df36b129c24709f7ef0f60db5e41b9d36885e1de5c85779257dd5ffbd189aa4078c4df86bdb6e9c5b6920983f7583a6b9b66a4495549bfe9b14c5b80fa85647c2edd13efc5032094a76eb85647ce1005b4106c45ff57e628a1bc2c13fbeb7566a2ffd57b7718229d871ddc35c3c977451f6dd521373d3a1058236dd2eb0bf7bd53a55fccc7916ea9e81750873f33fb6e0b4cbbd054d0319c38042718a2b245a823037fbd604a27a49669a2d3b8b08c950455b525f88bb2fe2485a1e62d20e4f439e7fe2d71c8256084067231a38a6b8f15ed596c5eb29e06de13c151c9c37efcee12c50c34fb97fb6c7897b4460d0c7e478ca2a2bb206f52d1f8a639d6045fbe4fc173e948bc4513da58e7207573162b36b3c60032ed417d9ca7e492d0f6c6b7fea20370bc1d5ca73a4baacd88ffe8bca3519225bdf99b5ebe86e0f633b86a8afa8619f0443518762127e5fb0e79eaafd001ca70ac1a903290f90107472918673d8976d6e663edba1aaea835177fc7c744dfd3cf9ee74e1d689d8846750ff69a5461c2dc5fd2b35c7696461daa770f8ac27128c52b4459edd223be175ade9d123441a8860f2e995c01fa142d95e838f21574015f16a923b03f22b56d87969878b2b9f33903423d82d10202f402d1c8244e9f6c64fbd9d0684feb570e717a48747d7e832b1ff8f9f9f7398ef9d2a28bafb57a83221a1c84f750eefbe3c292e0ef579aa7f97307d8106fb32c5752f0b8209b80006893fba8535d6e1950782437e9078ab3b2e32f3d3f0227cc3f60c5d61ff870cb556324749c1da39b6a9d13bd2acc9ebc101f4da6fbf860a547148d0ef5c170135a7e1959d0c4bab6d63fa816d5ddd281874ac4bcec96ecc88fb3ca6235dd013b68949c0a93d9c14ca4fbcc338557d2f7e3f133776e5e84d268f4878de3e0ce6e76f35ea819897af21ec8e26771c493fca40ef522e2c53f90263c9f97021b6fd6056ce73d8fdb15e53f18ad9e4d3fb7b11225af413d7abe77025ef8941077bf06360dc297b68984ecf482e5cecc8a90b31c0008789c2a903e9f511c2f4849909a9fba01fff3e8f369b410429db27236fceb0797459b9ba99b603c3fe22e09cac64ae57fa45344991e09567dd772c5c194e21f06285b9c41293b53bcd71ba15a39f02c6357da7f75418267dbe31cf14968c32f219cc5b0c74c0e9c146bc60c7e332c4ad69625f88ecc961a30cca77e6a0656fafca887016d3681c62495f3643c673688e524ebf2857fa64e3cb37a8d2280e6c3405b87f34632b2278272392a263e33daeede3e63614bf2a696b84339968192998bfe475a8d6121d7d676627c00aa0805e6e8e7d375136300ac003a5c807beadcfa996b4118aace503af37e34d0fcd12218f22212a1c04bc2903b3bcaaba45c809a1a08de600c4f40bef12f3ac4566516d0d1e892be945ad9ca1b233101dc94d03259e5bb3ba863b8156e4ee1f603c9f9c926c9ada91d36c7f12b2626c6f5266f430ee8a63f04d826b551d4b188a8a41402c75838846f7698a1e091e85ee7e5680bc8e8974bedc6c255eea25bbf7c12ec65e36a72774db95a3f37afe4e10295eb6f0051e5ddcc1462910ab6832ffcc6a3ac367470991b4a52430540e94b22c09934aff3acf9a3e7a8e734e5ee3eb1826ce226484f1819a9673248feb9eba1ac90e7075f041b108f3d74d85badebaa92ea00a4cc4ea2e4deb6428352e4270f7766f11f11485fb8d67ce5709fb3a9d8ebbf5cf3cca2ebe86c11f9c685c984ce95e50b73913933d36b2d94442b197562aba6b78d11217cd286b3700f38faf03cd09fc7fa7fc3dd176dfc5f991f8f9f791a6061f2f62d25873a2881ded4dd2119192dbef3975fd775e0b8adf074d8d396c6c15542cedffe7aec02ca4d258b71f2fd535a92444077f35edd91ad40d9e66604a77a27280d890fbac7eab736015e5748732948c8d89eb49376ac8361aaa126c6bd02c33482b6a0227ceb573c175f00e498e8704e3562432fcee67e454acdccf1c2edba4d53a5b0483b04bbee6b09aa0a21019d3bf6c951b4dd446b0986397e06de5371a02b8174941205d264769c5f47ccc1632337c51b3966c2f43aed8a1820239b233c1ed4f2e26d7866df6f5c6b19fe2b441ae336c4bae7e547abcae6256968700b802288d5b73f2d41a9004b1de5d377ab976dff4c0eaa5408d3250964e30a175909edee7194f9c0159e6fad673c56cd7afc68befff985c97742f836a23eed2a729686be2cf09a8d031ca6d9054e1e30dcd7ea144bf6792226e5fda76a1290eea94030e2dc717abab09324229f480b36ba0ed2f52ca456e2ff100497463c899964d062401818a952379489eea468414686a5403e74a128e72cd1270743ebabf38d054f304add236221d08ae573fa39c56f238a4b5a4b6bb2b00f071e1ca311246673c50d56b8d104e8aa24be02dfa46d64f9af639aec702ce0e006ebd389fb8f0bf92d03ee8086d4d6712b21c3c2c96c491d5796dab8b9af157835eaf058e9b592b2508f4b39a97a0faabc92fd77f833275c377d0eb365b9cf66a17ceca91903ed859841309856fe45a00dc1bc152f6f0b9b1147cf135ee28f6757442e632d0f7bca2c606c6c1b26d251ea62785d7dd919d1e54e10dded2dbe66e987f20ad97ccd9eab8fca553bff05ad84e9a7a4f9fd33e70c4c9f3f9a22ef160475a93385f4a8de5b259ffabf7e0e084a6f9a73d0664589a1d27b9d744228a2ced7681d13ce80a21ed604982f66106771edf6e67a14e31fa51de976e47f51a09ce29248fc851c13276be151f69b9cd9f8adcfa5fd51241ef3d4003daf9d27766669dea9852c9e9a1ca332766512b4fcd0eef2c34e1ab4740df417695665b9bf905823651fa3a73353ff9ffdc97ab545bc269a6f7afc2cc7cb5506981fa8439c0a294d21bb7c4683dbdf9c0e5cfeac9ac9744563a6e23daac0350fe55e4fb52ecb220eb7f3639214c96fc99bafe61f9da0827f74fe5b05074e00118e9fd65eb1fe0d60805108a54c75ed9732ee7f1865a07535397fb11624422c1c843818639c63afd06d73fd32fd310b11901b837e8720f26b6073d39b59f4b3e596ddb80668a1065177fb2e7be12d278d46ebe1ebc9249adce7b68abe6c2e366ad4ff9443b08e0a00d84af564fccc016cb5d8b1c647e3f2fec9202248ff508f551091634b36c95c28e1178d647f009f91b2967895b78ccfa0236b359fdef781a66ca96ecbffb880e797ba81e1e94e9150e395b034d1bac194e53560fedcec540ae781f7b69392f92f13d47fde2adb84291db3546e08d30eaac239beca922b16ddb530d2f0a4c7a70e25120c6129ccd9f8334df71331be44bc7e811d46fa49c92d757c8b9487dcb7ca641839bc645aac851b19d8d9489542add;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h495fbb160314aa4aa79f307fb9c66c56c9d6ef26fa6059c0bebc60bcc15a42fbc1ba73db73fd0b3ff2012b28ccdf2868e5aae6b237abff0b1575455b53e1cc3f6b6d364fedaa991dfde8f0aac5476b9cc11299e99110e97649db2ef418a98a4d2961f2c814add193ff2c631fe5daf09d11dc3fb8c926acf754726e672aad1b9a4ff3cb4bb734ec61c82066df9ad9368774e29d3bd99e3182ff7f313ec3465b46a5d0a8f30c5624c40db1f98f8f238d05cb46e7607e9ded2ea20f7f125086960d676f00b7414de1cdaccc17950aac5f1cb31cf1b0b26f4c491db23cdd4aff2d851fb957fbd2c6125de47b08217487c4bff03723073367c593b93a662efa9e04a3378bbc060075e000ea4c8d8e17c37e86cd7657b0c7d5cb94334e35fb5f5f418301d7a6e6e3f18f9caf480ab4f7a5e6ae423bb031a88bab8e2e0cb44faff38e95ab8c851dfb9f889f893ba8ac82c0095e87e0bae854a4557df4b3ae121549ec65fdb42e8d5a80b1b49af6ddb30685a95d13121ac93b72c217bb97e0a9ebc9a8c9397add124412163b0868fd8bcf9167c073e0e8e13d12ea9ff5d2452082567a660bc3119f4b3221ecd1befc78ec2fa8e4eec8976b1efc9047259382cd692ec48443c3cab1bdd0b51f75520546042595cc447c41cc18dec557b6374bc7b427edbd6048380492e0c0a790a801c35ebfbd8b70c38d090e184da9135230131413e9a1e79f0448d9864b3c18371650279c0b400bc2c364038894836cf5f399f571feb9f972b6442807b8fac700c2d4ccafa55280b51dbf7b002bfa20fdab1d246ae394c0c70d67c485dda7639ce2f1d620b0a176c098cfdaa23fd071b62d42b652250a944ce11c0c65535072e5b8d287ccc2268a6e5c3eff39b8922612af4d8754be307ded10d144ac434ddb4b991435fe16a7cf3819b42346956624bda024f3bca115057c33ccb8671d24d2179396ef5e0ca566a0c90e6f6bb3f26c582269e3ee2497e8a97ee466071cbd2d61e317fa93c457f4fa19cba8366c3b30deaede76a4ece0a552bf51767096947cff4923e17ced89c531fd9ba0b61ee7b1e706322e20e8cd5ec09af4213ff1f0fab44ec35b49e41433445043d3d01d32759ebe85b200b1ce2a4866a05e9ff8ee6a3fab542c3c4a5bd24d0427a43be6b525d3d70b8d723486b0ee9a99ec9bd949e5e6298fcebaefeb99387c8493ed0d0f3fc8e9184127fdc84f2d5b57cc0e8c3e4fb26b49bf05e3f8d9948909c6b840fa66c89597c01667689392b6209c67faac1d7ae6fb9a659927e4ecd161c121135609efdee80fe8109e2f59521a93c7d360987e0b462f432b6453f320a51e1bf10bcdde7d35a20e3977fc83fe04dacbf30d2d3ae51e18d25069c79eddf00b6074d26446427613e112e7882e45b0ac2191ce7e2e0aed59a4bf351ed1e21975e960a1c6a8ea9cfa96392fe06fd808f5a726a3e9678b5a77efe3cc5b5359d8bc54a8675b46027f551f25379e79e0ee2fd4237b5fb101c09827f77baba77509f593355a146a700ec02a24e0b2c3637321759da36fe0da89d31ea4a25aa2736d1b0f9a1fa4c0f48ab89ec40a22d7588cd8a6111d14908b0450e0868c54c81c97b06b51c636f0623a9400d8017b39b2af50a53e825eb239234b5b8dc4510cc4afac40f069ecf12adb38767bb8a4ee52936ef96e4012cbdd39ae5ee74df61a9926b5ffc9afc8b66c15fdb1b95e145c27cee4d80ccdc8b8a2d1efbcd4706b0afb666b738991263fd20327c40bef8e3005225950a981d6569e201ddba6a7715e0ac26979dd06461a4627f367c5a326ecd4ad60c5c6cac027240e7555755901c7e22380fbe63729a06a086a96c349e656002ffd850d2a3dc351f3d2bfc66ce63a155b3b3e672feef2979afecc28a0404253f977cf10721fa9e52ee5be073c8a2fbf3a608f6cb4ebc74a6801ccfe57230381d4dc1f28f4171ebdb0352e1f30b2fd1b9755d5cd04a81cbaba8495a7e4067f75979c706e46234843798b27cfc4d5c85c5ef049599a44a634b188bb7365cf1b0cae16f08859db75712c9da9871e71f090a5c36f8cf9196b24c8448c33a792e27b4ca36d411d53179c420bb2ebed632579b5111fbe97b8958f2f249864046557e5dcdce53ca78e48ce088659153f57f2f5356aa787fab640c09a1c8b5e07e6d1718c60ea1169093dee1de4ec6cbf3b984f0a603ea33763edf8cd7a985113858bc8cb56b017426be81a9ee51a51f74dc825919f2d3122df303bd38ac3f415e2182d8d5d31896afb5473f94d3c6aabeb0ffdec8b63ce33f63d3e2ad4fc39d158c487ebcfbeecc9104bf5e0bd8e5057d5eb9cb38d017146c8a2ec301e067c9937cfb0c2190071c076b41973cfa52f9730c8d55bd235a8d6acc4b55892d7310596acb80550d8b96d3958ad3b1fa7effd58c1ae034a31f97f7011422578746e529f56b6326c35658625aa0a2bbb7ed890c9232305dc249493cd77a0324fa7c5e9f8d08914e0048f3d13644c01b39925fad4c0f6f3185cfae71df5e1424501334414eb40a139a5ecb19f09e228bd2060ad02ecbd738222a22e46b7e2e3202d47dce485bf88bc7914734d78982cc12634e8aaf647a0f1c0828e2d7b4d409a6149c5f7ce346310a8ac3e3c4afff8bd66980dbd996d0041d31f1401b87ebd282bb0540edd0eb2ffeace2277c41cc53f7b011e21a1513f7495813193d2565da4258977e8f1c045fa3dde13b4837a2738daaef16cd346903bfdb79fee7c83cb693073180bd9ce7cb3cbb1d2d00f177259e5619fea5babedc5a9f5afc9f8f0fbdfdc77d3ab37e10179eb5f3acde36c1c4a737ccdd0ff75d57a20d249d90c99af0ec154e724461ca1874668abc2192c712404302f41edaa9cf4ed37d176678356217e4452b074190107569a09a342978b0a4938253006f421a879a798c90ec1f76bd745ea719e750b6c5cc26a0a48e0328c0661b40123e6574d7ccf43d690868ffcb85261a97edae25a62e21ddc7401b4b7514676c3922958dde5325704f21e9e1bdffa604b6f9a72fff15b8e508425f9a037af9d4f04b2d1b00c0e607e08e87ba7beb02b2423a30f4742d08ef5059d415ed7b2f3c2e6ccf0bda8987982b5e2da4660ac61788bdd6132d52f5918eb442b50b349ff317efb6060a3973fab03b18e72d1c2130d6a09878d1436debce67786845ac5917e361b93617c4cafcc259f3555a095c3edbb005c166de3e58cfc75048b7d3b91fba43d1574420350cba8215ce23c922dcecf8d6f2801a1a93d33ec731f09f9adf03de73c058138669ef360e1eafdd8625c4149a86b02b62229a3775a1b5ae17e67c49f34ab94a7f9fd2940d17a3196bf3510d17cf96dd29ead0b9ef0fedafa23131f696ad3e4f1a57e50fcaf740d40f98f11e1ef602eb1b45fa7b33352b411ff217e76fcefe141cd6346220ee81059ccdae632c1055a9665b06978fdd0f2ad4fd46ccee4789e0d9199d894fef64fc7ed6919a3e47650a9de9815847a86ef7eb2fd213f6b66017cbc71ea51e13549383e6570cdf6b6b9b9b13f57823c6dfb3410d7e1bb42a632b99be2bb145516a5213966e0470bb2322cd5532d44e287a6f6a2acf00d37b3027d20cd504dfb7482a133769b82f41a98cc0128ebc07ddbc1fb153276339c49163ddebe9f9c241e866cb8e8afaa12d9d39c795e386b342a30b306cd2ae79144ad82dba61038f3beeb81a99bdb9b377e2999c00d1372699f59b4308a1fb2ad634bdc1f01a3a30dc66ee17118b524dde8b98615231fe67551a02ecd83d71061458c1dae3a10513e257f92cc43f28059e5b9031b1a558f0e0ed954111a296f4f9a5b7d0eaaf152883594cab56443ed1025a6f3af993031ee04762d1875a11f2dff27d24c7f255e4d9e86884d9b5236b7249bd2fdd884f2035a1c7c96471c3846fb387562b2440b3c9abe3bbc58c6f1b15bde4c88b6fddcc0dd1b104f16f8d1c67c9cdbdb9ef0de90c8f0537fd6624220db4e2e0cdfddb133f35704c9785229e0756c2f0cc29b54b1bd989d17e91d5845f59f745950d7338f2e1d36698d173a6d27361ba3fb850a1829c85f6046e45170c4edb918fdb174f798bf6fd6c60d68c0586019a758890d50fe7237d7e494774edef3075214423382d390ea63414e4a622a164dc6b7a4de7e60ddc29289e4f7cd22e9b3a357ed8543ae206675fceadb53e0ecf2c85067c58c763090d7140e737e512414ebfaea5288bc539b76e83ced41a2bcca95cc3a1401a0232bcdccaf89da4eafca932f8efe9d1c2d7db556dbcaa4330964d2d8fa4d84c63d6ac521c8563608d8aedb3e630d4ebe7403b1bc1d5388e1714d9421e12679402d6ba5aa4bcb668ff30363b36ba40ee8ba500660a8e15a67a13e997841d418520957ce62b89a3c045f28f542653534c2599c0417229892e23c9ea8a630fde28efbdef1a366854c80f0f3c07809035fe25ddb1a591787ebed5c6e8e43a3b1555939e3190de3b1d7c90bab373a87f2e912508b13ec41e2d721ccfcd201c381e3f1b70f2a513460782ef7c1e6887f82b30945aa74b1ed6b226bddc97a634022a659097520c671560d4e1162229aa2fb3402d524aa2a3d667961f38bf93634ba299c625c7f67dc8a5b36e764526da0e9b7ed248b8c34666e5bcaa375c9c9e18e2d47d93bba1be6d28c725080c44139bc36f4bcc7584dc2f7c8d54ae7a9429d418295bccdb5f203f8c463a916b32527de8fe5c28976ad2fc662c26d2224c77fa2ec9f8f477160e61bc5c9ae885348352793807372ccb45c0f89b56289a2a80a6f1f294672007cba265555a5337cdfa05e89223b4e94ccef4b55ace07dd71894471a85667202257fb4c66eaf1f64cfbd3729a593fcfeaab42e843d3cf2713bf7d6c19419da7466ca2c137a148ff6dd4d8fdd82e245abd1d4496b34f763431c808276a4b363481106b1f11b6566bca47deff5d2998f92d9c0f827a154f50123e6a0e3f4dd0f0d9de2c1a4eaf6c9fad3173891c559467406066ef039e2f4777007d891dabca611184867ebacade7f915cb328f1da2f861f2fc2ac942914b9ed5cc28ee9aa5949ed3518cfccd63fb2ba29c5eb5d013a03353380d849119cdc629d25ed3ebb318d1041169232ce1c8ac87d4c28205242298eb6e6b5b7467afad672da46c130098fed96efbdfae7be48cec6b23c45986191565aa8fd2614513653a5ec20f2dcb83da67c23c211bf81ed0cb38bc2c309bf47962dad9ed8df22c94ff75456aac23216ca185d0fc1f3f7dec226151639bcbcc871a68d1d34040f67e1f55c1cb7ac6055f962c598001f7c150fcbebbfe4915dd6655f977d3b3cc191eb12d872d6756b975a624deed5c882219a888e64615949133fb5d1dd159f61965f58010898872034fb0a3d6414091238d59c4cceab3f5ba190a447d6a55d63c1c62ab4c6009ec45b4b7cb46dfc8780de4811e8c8aa504097510ecbaf0e02415d47768b5764fa3695c13bcb7f103f89c83db271fc1d73ee749;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h61834161b0beb1a2d9902a9fcf7076939389706d4ada1c0db39ebc0d28a193cf2afa5ebe3d9eabc8dc04271199b210d5c198c2ece6c441c5354f7a9fffafe26e9501cd057e6b8c84aaba0e743629f5b23efb7ca711bb4cf721597660e90c6e08b4727340915301df63131237a405e9e0a08303a0f4f23e032efae0fdc0965c6ca94d6df5aee74128407333e3c4c45fed6ec7a1f25ef3de7c356edbee445a4afa8581ffd862729905b85de36ced41ca4465edc8b58870109f72bbf1dbb8914f9ff6f915e3e29217c9f74267f0a8e1164a35141b7e939e0afc05e0f8a40feeee45e22fdfe2973cf78c01cfd568924c48e4db397a0234fc9459d4c4c472ba0f6cd91c3e6276db9fdfd5de7b74d8f893e9abe0ab1380f87e10ffa5418324c659bc84536daf5b41967a2445b5a5ec857089f1acbbee64f58e17420fe66ae690ee7b0fd78431e10eff2888e7d4a76cbb604e24280957c3e742cc8b0500a888ab28357b51b0ff4f58da173cbfcc8a0c967be6cb2a73c06e626eebc4d6bfb248cae8f1093cded5005188d644feb3b43d43252dbb6514cc3464749f3b2885345b47d0ef9a9abb2f0c7428da5743dae17fbbcf18f3305ab14a41f305e56935a3c6fa869ed2e1d53540b0f30016f0d9baeac10d53f94d517a34773fbebfded6f6705ba78475a69c0b12442a969c20d27d713135f076ee03a14b75310833b499d0376c405134587b53c81d3788a410c2ef0ea308bb4cc8240aae0df5e8deb6063cdd4f02edd8460b988aa221b282b01ea0d692330e3663c2591bb13eeb9c6d988577c91919570e8ea9b31e5e107bd6c0050a7d7dddd0f97cd0e785f1b82ad073467112400d8ae2de2331857176b99d361e4936039bb76ad942179ddff72e08b1b6937b0547f0230e6355e3d33016f656772dce4e87ae234a5316f6b9647cd854e96484ae6a14b990ae119b88041c2a2348d3f46995f4609244931f4c195a9f1cd797278dd04cdd224cd78e1a89706bfdae053a2118f141237414cdf78a1d3ad53d004d4fb577f4f7d67df129404c54b514b7af1d537e6ecec9bc648b3c3255b1d99d12970020046133db4531806918b1dc02137d72ea1225b8c1489c72fcc737df8858423bbcab255b6e72ed3ea065e52c7eb7271ff65d345c8c7942105e744f740049517e4f4188937917943cdd53b23bf4cf23e7474c071ed190700e19811ce878476b6d4717f997499d094e8c37b5c19e56a1ea0918f7b3ec8048f3be946bfd24cce5a3f413648eb594c317b09896af9080ddfe443c0d5896c6a2edf7b7ca762ee7fb8c067673ce46dffddb9a2426b98163b274d891a29500b5b1208256d8f2a36c33d256eabbc57c7b7c83c4f5aa5f4969bf52231d056a724a5ca87d56a94515e959c3360b6935b2415fdac7d03c1d9c543be279aa7f92f6a6429698a3c8dc76e1c508e486f02c3530371ab7197083d9e76aefa571139b919892467e26659af81a02153a2a15234375d6de2046a835ce6c7c5c5409a27bea6a817477a8150ad5107cfd74815aa35bc45ced222750da19603eb69420cdd5ffa9d769fa185fc7a8d15d5b81ebb086f386bbabc0915d87618aed5677181b12937ec92d6deabe0b4cb60c26544ed3e48601d4579837f500487440e4a768057284b1a027384d30dd58af67488de41fee6a13bc26c3c28f423c57103b80b1872213bae9cbc67eaeaa39d83ae4f5f87eb9cdb532cdfc8025cf84702657f1bd49468e11485c514b33022a6097b52e7e4b7a9603ef04e89646035ff2e1cd5ce3cfae3497f88d8907429f152ebf5f3fa3ff8f76d6c3fcebae1344e104736188b41c6ddae7472aaa01bb8797cabd557eb84b99c05b0fde71b0b150796a8131113733e6ad3fc2c5b276a1942aab4ca2adffa1cb6c6933f1a664b8b502e33b13fa7f3a7ec3a71b22cb30f94691107aa7c38a6daf17d8bee2cae97f42d485d5ba310d0332b77c82c15941a19fcf23271756bfd1c72968d4009a95183ec4bc0ea55d92103a6fc6e034e91ec712aaaec012eddc832ad7372b696fb4ddefb51f63c2cd52110438378d2ef11087a3caea57164dc4c38b693d95bf39a244699ee8e17d3514d0f4ca2e940f5ea1be9f366a9c833c321272e6f9abb75e3c05791ebfe5e43237a067c230caa646c24e64bef1a31a6e8f9fdbbd2117c591cf1921c2bca34f2326b01123595a1056ffcb155b3998e308f67c314ea252510ad362ae5389bb20995300872d3491c9835cbe8043900197692bc5d904318682e28362a2ae73cc42d72b40ce69df0f8c500c81f9ccc913136a853910a20b75265ff993a286f48b3758ec511bfedd66abc9e2b52365620bfcd18e82f01de3365614dbfe03cc1db857756648b4501b1dd7f2a55e58728dc69f516f76200c02545089741c21f8c4f2563ba58e7d37d77b6630dc93bb11416f760eb7c79960d12b4e788bf2e0352acb48095c72b077bfbc6b59940f0cf1fb944be7e8b515733f816c1053437b84222d0bd1d9d1b984fb9f1ff9a867df29c2395a114eabd1eb717bf8d642f77886e77b0a6234cc414085c44f640a09fdfc08f97886c0270766f5ec21651661a06993bb84dfbb3b858fa564b2d9a368a25e25cd81f957f9760ad66c1422236aa98accea4a4b346c45b76ddd7883b87557364823c43849b2463ba1c36adeb9a2b26b4d3c456b3c9bb6bdbbb7eae1968830c8213bda87bebd0f8ea632daa1d01131f954fe586aa829378cb96a4628f62fee979316a94ba18529bded4062485e9cc81799e2985bbe2035179671b97654a4664494da8c62b3054443d7e9598fb5d754891d15354723a418c2c84fa6edab76361eedc95e9360ffd91c5a82dfeba1585b860df0357f61f996d9baf501c0280a7a3d36a89d20418daca19ba54c262b81dc54ffd018d2a65f9f30c598ed4ba5908f5d71e2971f2aca510972acb48cdf27d62f080abc4953e8d44e4a71252f804d51e269cdc9468cd2caef7c36f4c7530a3f50245ac438be68b25c9e713e4ecb3e27996808b7b63f0e7e703c6361e69a15f66f60e028a8be911cb38fcd287c9ce0fa0b626745e25dc21892f7060bcbb85edea41bddaa459e23b22ab41bb4e51b2c09201e9f7d648a3e137e8e2985a740b1bca0e64b03bfb8f044a392e8f19fc9bf60ce897492cb9f81d5ce29051fb77bb646c560c737ea6e16b4673c9afe5bb5633afd4478dec4330f8a37a0f7001817531b9e274b8a4b0eeec957a3fcdbcdec0c02e97dee1759732a6b672923f446c179ae0f9ba026f933f61e81638acc405cb52f96f90063e24763f1d658af6faabe0eed3e2e2420e3900c6d80ac8ef24d062625ac276d6dad052edffa5399d50e64e88c50b9ae529344851d5b42d19964ef8083bd8358baa06fb3e0e4569fafff1a598c18c7a354e03794b8e4d5800f5808a9ab3e01c8fe6c3a1795607668a82c36a7f730a3faef0fbc67469525987ba36dcd21ca95ada2d48206568ab7fdd31ca680562f4f612ff14fd77904bbca47a87eede448e5bb450b1e7b8b2fd48277fa4ee23d9e8947133e2e30335d668b88af7b17c40824a0494047be7961abc7881ee6c932ea8ed1e70754f9b8f318d5809bc4ca8f6d97c1ec6396357056f17e532cec140a184199fd150b008c22956bee1604ef4119046df84d85b89b3810ee77de7289f67bf20c9b2803e5cc868ec4c2d15bb10d7403937a56373af4d43a02a8caf80c9f6a6a8053c04cafd1277924d508db8c417241ce3307a0e8209e697296177cf97cb64e3500d469dc90f958595704a7465c2e633eb4501b0fc20027f41122fb72ef55f589c4abc6aa763076232bffda2e231a4bb277b5da19692ab239238705e02a50bc1759a1fd3ab367610bff9fb4d9bafba1e7dbe5e6b709c373b49e40ddc81f44fc9654588f7fd944e4b7719d93a2b160ffafd4e288d459d2ea8383498e36a272f0c622d2bca064dd767725429a7b7e6d894c4522c0b2de7b20331f38f87fa73844a4592fe09dc399277509eaa195c209fac72b2cc354355c1830951c55d15d47ba3813d879346560e2b01d558f26cbf769a94cad64100460c0008846bed351232623ccc8655e8abf37ca4b71a65d966089319679ab0e4abbe73966cae1fbc5fb0bfd292996ee1d13fedc7a75df41977de378f55d51542d9a091148678baf82d2b56ce2b3947be37434c4077188b40610db73343ec110de1416dd6b4e17447a6816aa3c114a5028c356a160d423156a9a2b047e43200d288641ef27247e4b0339a096d150bc3ef0351545f4b0a594cad0dc1836bdad94ef1a0b267ddde71a91f6797b14aa33907d714945e459dcd4f9098d2760f2126bdabe0eabc93be1b0014174c13365cee3cd510f0d2cf0add937eeebab5370f9ef6df6455e2425c672ccbb89e59fa56122cbcf20a211fe281f4e7e9e614ab1f9ad94239e1006f4104fa93be68ffe7657fb5f6a7b405b1df1992f0e20b2ec3bca04a035d7daa31d8bc8dff627fa6f51ee5bd9efe025f5bc7202f2b35226647e85e955f785cbb5b3c1429be8bb91b59271d1856cb271d260107dd00125d7f180e4e868638dad137ff3e00b9b845576bec7bbf53542637c4968b0cb40f839402cfaa347754ed69e02c7422ff0bc9a47f6d27deb195fc8d1530dd99142a0faa57ede7c1080c163f718461367117f65b7e227f5674214bfe17e4b219ded9f20679be6acb59fb1725181c4e13243b1540ff1bfe79ddd7f9503faba2b230bd5357f168a9bd45bf65a6dde75ab7a5b2cd7ff28041a4bdc1ff1af83cbf0520311e8c4487ab89048da763a4fdb54fdcf81a7b0208c2bc5eb430a5d469b5fecd67089f3e7676fd4802cf855afe17626af304bfec541aad6df6d865dab9adcfca34c753ddaadf7b313bc6c7f345a6697d65b1880d32735edb7b4049823c30019062b8680798e764e0a53add454c67c0fb6fc0f29506090ec652b8b4f22fd775e9ecab70887307022e5ef24f0346e0cf2458e238f2d1e1c468bdf975a17a080d9a6fa3b7044c6142b02fd7aa75148613bc6634408ef7d8cc2c97d6ca79069226bf4ec61d206421cf1a8124f5a678c0a7c204252aaddd04d99cac6fad0d7f25c061ac06a5fb0eeeb183b386cbe9ec9bf2b9a970ad5ef9eb6c105ddcdca38c12a0a1ed1a0e7d26d3993da91d71f457caa2a3655fd303a07bda8ab92ce5b540324d43f58bf85f1ee62053a9f13e68f17d9e88f47a40bf5c25769c813df83d56a9d017578a310c3a935c1b2eb430d6ea92a3d16216c8b191c0b87f07a88fa13c3a0aa2a46e54982647f1404de05cf105ab41c826d4d342b94c17b1ae32722d64565fa9ebd7de1bba558e9a447677e54f4e37bd563cf155db87b8298ff54acfcfc321324117c07b22243e54bcb64732afeabbe996efbbcc255aa0d33250d41ab9250b52be5b437c08312a0d46c3713bc90444cb27b2310e70a46037045d53df392422fad106feaa35028a199987c6bff11cdeb2f527a36b5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hae4f9a3b666b6445a73868930e29bef527cabee8c3ce04846329e5afab88d22a72a08317e6403d696e3ce29004e0016533420b0161fe3733f96694580f8ee9ef83dfabb698185ed33d6ffd425ef6d9380448045565ce73660a4d76caec1f7fd59495ba6de5050566cf164fcf87eb251825b5f5445662d2cbc36e773b87f9dcd5ef7bf92439700a6703da897966c005ad7b19b42ba12b924b61d9bf68988052b08b80fb2a2cc8c3c50d16b650289e2852cb474bc4f5973af1681732bb4b25034044641d7f67342313047397e3c50ccfceff126ad37d501f273252c10d36207e0303adb86f8e5f7e6a3f51ecfdaaba4e01d4c7c70491d4aacd3ce087c49bf18307ade159cfd5b820c92c5a3acc7512e830742b4c80293236f682b461c579f74fbce90d88a058a64e85a247151b6c8ea32de18f5114efb4d50c166810dfe350daec479fa2bd7ee7a66a930a82aa4f0a73d70247a0baee9e7cce27efcfe5f24c2847aba7378ee9aed3240596a38f5a851358189954376f5ef5883e71b51d44ad641a7a497e9cf54d2171e5e5a83f48089107736683d15034d79a0732c3374cc36310edff52ea978fc4f15c682c4f786911f1d25d65f71fc1747832ae26c76067cb3aad286a320a4c90d0109db233981a20c94f179fbd4a578bdb199dae513fa2b6db3db08db968436c0b44dc4f705a12c2cbd47397b4bb502a1203fea8af73d1a9cabe487599f5fb8aecf995c0131e34b37945b4c1fa2c9e39f2bae6434456cb1cdc37d80255e2a9430955fa6427c62aad4226faa3929a774b72f0a85a931d4c93f24521eda8002c076b787adeade568c2191a1982ea84b78751ef2f2a0c9fd5d514beaabddf73953cea74182ed63455058ecf6c14989583cab5a7a3587eae60bf1a50cb9612d9b24e011588e6a0216578a1468c38f33a9525c2d77a81aab69984649615e2b4be74c92cd7f4eb662f43d924178198b81dfc62940aaa38631bc2cfe5b5263516cbfdbb6dfb87fe8803044635d2ef66c6636b75cf37d51810558e418169bf74b79d518135f3e6922296dab4445c144b02a52ebb70d99bc506a0d8b74ae1d41ee8620a38a8066fe37ca37168b75ee141a817a07752cb56809f2337d0b44a63701c72cd84e9b8616f74007b28f31befe676d9540b3ceaaaa6ae0d0d292ef4b4abb01cf2a0b8d465dacd40f6244db8b57c6058e299cd56e5ab2bbfb56b8b0c7b761fb00470578be25a92f6e1d1a0e7d91ed9ddad0c5988252aa66eff3087813e61981fd3c6e6a0baa4f444dcbcc976a5aad94b664b3b935438c88636a676c0b2d00e917c58da49faf281cab75c3eca998af8c3636651e7ee5c38ff9f3b8cb6e44262b8fac2e52fac3baccc0c88438945dee0e67d592aaf258f6910f40668139c8d8c222384b53581650d07cf3276e7f8858b939f6076c27324e5fb964eb2e29459dc6a17eaf84213071ca9b2e40648cdb073234d45df3b3b41f06a0fdad398af22ccdd8a2bc1fe43374930fb13d9eb7d4baeba16bcbc59e76564f14735dddc5297f1f6a62900713c596c565661aee28ed78ac348ecfdfc80255c3e3422610ab9db6930b97296c237f965ac9daa4309445e486f95f730abaa6dc642ee643e92af0d83daae941725f74bca46ef9b3db2f355d9b00c8530f0be0d3968cfd2986a8b6a5a7772073dfdb31f560f05c02242e71bc4d1f7d3e8e7e4bade4c1a352a8f3cd4d424927cc1c6552868672a15c02b97b0d0793630f126a7c7ffa1c1600fa5b03a4f158c5d596bbac3bf4945c273a0fb68f51303a21505fa8eef7d28339adc0cbeb52b224f0eb222584acf48d7221ccc5066849b76f78e8b9ad34933dfdc8f0870fbe4a6ed7e82b98a34c27ca4237d453df68c439ff33781412caea45c8194870ce4f62ee592c2ec565c3ba93bfb7aa8c4d7a7c60b54eee4e087a02be2b119b42be74a8d3f9297ce903c356e8ca7351f69817175e088fbf756e01ef11b9bd2e3d3518c616f311bbba127e687c41a8ed35caa7430e1c08be0c1af3cc7b211b6d7399a53c7b2129bacb4961cd3b5c478be48527d040fa9c42a219a3356c07f8ced6fcba5120b7877a2634a1fbe19719eddc869bb2bac173119a9f601a9afc37fab7c46239a9b50fe8ef456ffb98c270aa7a475605ee10b69f98fa325eacaca5ecdc03d5108e946829b2c25ac61eef9a9cd8a3be9395159c2cfbea43bf6bfa1b18b5504efb3fa1ba0224a9ec1c9bb9323cae9253fc82ea2da392b4503ac2d4b417b350d1303ffd3cba2233d1b90d554ed232db72df29fa5edf9a8ef075fdc431958567cf648718fcdc5f3a3f3865644cba3b8198ec39d4706c2744e67a801f07da2453514bc70c7404a7d8f9c94bf62e1dae0d6150cb67cf0605d352c1057c085979918208350f02a19ad0b5e62ccae34d263018186961e453b99488a0b0a57d02c937dca15c3240c5d0516c8330df365b51852af244c149f825ce9fa9461b8e3d01ab09f006fdb371b89ca7d55737d0a0eb10a931c04f8efde8857eda7880ba15d95f26f776c5703a16708c9113ad9e3d3fdc0a242ce7d1f670cf1d634b22cc50a027dd323a520aac1568d63a785351f5d6cea4c3fd2a9f4435bd0ecb44ffd187063309349f6c398e2749aafba5db376ea78c36693d680de2b67bd88270ed881002e14d3fa2fd7727f16a1deb9a393997d9237367ea752e6b92f6d528ca24a47eba9cc7f04005b5325c85b0bc925687020793f9e9c39783888ec10944e410fa22f70fa19ab19e40c30f06c78303ad095a3bd5d7af5e988f21d2669735f09da01f2091035b0d06ce01f33cb5ecbe2fe43b0a0dbce73c57ac9f555897ab37f8b825dac4d83dc0d6d3f00dd29787869fa2fefddb6a3f521cbcc1b7bae111ac48e69036b41c131ee1b13760478eafa032f0bfb6b1df71b6ab163e404fdd12c844a58ed20811d9e319411fec35f4d65292124f6f9665a5f7fd12ba5185a040b86aca7e227eaf2dc8ae425f641fd5cf355b966d6d2d355c59b172f7a3f0f7b0934b808601f0300fdbc549ad985e9c4e6b03644508099ad98a00bf4ccec1466adc04431d348b29a86ebda4eeb9e26d3a4726c386a33008709b6e832cdc3aa853dec0e37184c63c45c9824d9c97e2daa559d107d59b74683e915a6477bc2e2c21b409e799ec3a920e4c6bcf36e4526a7d30e575eea74574587a5b0f0ed997f61779bd6302c2c90ce8f688bac752948455b0392fe69225ac526896ec377758b0c49928ba315e15678b4baf04db2d584dad216a906901eead30e388d0104f6677353c67627bcb559a09a3438fec1d9079dd93f5104bab0d148b70cdc6da688a3d2b0a837d8df5c141f81d212011195a8b2d393e0dcaf30424353b3ba2d4a6089c32e6d8ee97a772fa3b7b7739e7f8f7aed5314087e88742417753be8f015e393c0a746dd1597fa1d0c365c83682768b1a186e699ded21d971d9d334c040d854b9c7034070f28e96242015dcbd3d4546cbc5419478bb18bd86e9de05675065a68693070610af4dff04bc57b1d147e46497f481f91d03d4da5a9ebc93b9b81c69de543f308ef55611a92d9e99a2b365bf17f53c1b387b6b3426e724c28179b7a70c6a1b3388f18289cc4cedf788e0656cb06d97e81cf2cec24c8eda2f31a8664df225d180d034e31e58f5b2a7298597fb2384d6c6eec303eca43bc0547ac37cd6b6271f2af2d66dfbc6ff991f8c934378aa2c0c4ca8288dc7d4ffc3e171a7e370d172f20107509ec4ecc385556dbaefcbae4ecc1093c98d3d7c173b8e0ae8f4be458983f9cbaa3f6c74bc134c2551aceb71315eda1923444777490b97512dd93f08a40b15045d1912e63c0ff892b924ee267e0c70aedd3e4d5444b6681d865b000ae1a09f78a175a930a215adbae0fc1c6690989002334d2c8d9508846b781d6055e8796332542ff73924868bfe078e7cd33e0494e140eccf7a5232b9a71ebaa71781f30a7c345b60e3669cc32990ada56677d99f6a146cac551c308383369965183a61870db3c8655c3b08313bda353b85c31c81c4c4cb540fcb66131497b01ab2059fb6b37670b24476b8f7512c1634ba1e615c863c0f03eb930ab95e15c54302a083ac37515abaee2f6e643fea5797558da122764b70725d95640acbc33848474fa1cec6871d3f2757305bfd59e9c17f9199352fea396a145e798773ac0ef487760b28a86833e880986b656710a55f5a8af5c35196e081658d727c743e12584fc4ca360905d3d0fd7548a2094d9ca63d640dd7f5e4fc3f5d6fada10caaaf49faa06e03454549428f5bbac1fa05968a6eed917a964dac0082957e1cd9e2f700c1901b8bcf17a34310e0b8e4d1e93aad0136771c11a3d5daefe4ca962f7965fcd4b5ae9aefb0403744a262c83201f708b7abba448ef85f34421f6e0cb0637b08f5127b9599398563efc541c2dd848c3df445e4a1c40ac3529ebd3b1e18867e4b1cd0b19703c8d00fc41c3a4e68d98658a7790e786765224657b1d4773f6762f8ff4a3c17797c291b8d1ee2d1b88980aff254e1c130a2ba0e770813442a16453ab5d4d85ba4167baeb47f17ab72219c81f11a015d3324bfedf57b0f3eff972d90c87fb86cb7acf6526ff3d276c26e76a26805586ae8e5a960bb7d56240ea383566f6869f5750c513efa569547c89986b220395c8d4c7d8fd5a626d814304d831eef36d0c1f5425637f934fbdc174d7195583b1095f726615e8ae23cf9a3e13e5d130d097e7d9ffb240617c7974c93635bce875db87da7728b338e732e1b0f46d8d3210d491fb5614184212776bf5a6c157d8d206969c83c808838c291aa1cd1d7e145004e84fbde78c6626823b946ae6bca6013a1d078647abb59ef351f9c5b9f0c109e2dcf384ee37609905e044ed345430c5ccf145b9ce3ec8a027298b98d930001c68ab865c80bc68bf3fee678a116ea8f4a7849b4ffc1c72cb0be67c9307aed62cdb4da2754888f9dcef780efb609cbaf89994fa4ced699d20362851b9219c8577b93852458f3cf1552b0cc304b3d33adbdd5d8549c6f81917c3fe02f0443c34ba8ffdaf17f878eb6f1c51a788457c9a213015175db6af8329ce155a6a0a83a965d51f34fa4ec7282c3225a1017359088e09135539fee603a9c91c31f3a72f67d162144a823c8cd32bbcd83841a1144effe1f66eac4e2bd0845aebdc1f4083af3b5d5c4e777c68ef33b2a6f941ccf08c0f69a56e89cb2d90143eed1307120bf902acee3fc812663c1c58228d1e0970fcb3d4b2df1e738936ff33577a11e8455ef11b65882b82e51c589bef9082a7ab961a54ddaea41f9c79011287eebb31b772c731d7f0bc1516013b2f9efab600fe0604463b561249edabec487faac809beaf3439a6c1af68f6d710ab5bcfed5f69c9c5cf1c04566acec1b09e6c171049ef47190c98294eee29169593c9cafea0874ffc52130c7d5e706a326b3279a3653589e41664d7cf468349d8e1a624392a5aadf079d1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7aa87d5c53d29a120fa5fbbec46c0f4c5084d997f933ccbce3b5c3df874de5972d5e8fe5d8afc0920460751956b01fdd67fe816aa1841d086a08e44f51d5068f011755467e552d02845d9eed695264d2f575a08b47695f3e8c8d31e1041273c3324181c7a40335d7b18efe39e7ee821cdfd60d1a1b84982adb637f910a5eeebe5c5cef0543d1d3d70728c9bc433af35a2235b1eabefed187df17c8f74a11efd491f34d2eaa4e4754fc78884d0bf19a26cd5e0cf114da3416066d6a062f7fca704d913a9767ee00e5e3027a7d73845c37c45739b0ab2339871488432d157a62b434c36f21d87161e8e6b44e14875735a26fe45a65a9dadb064852fd18f0f0166ded602969dc2c891d7bc302992401f3f9c210faa41012ba905f4394a45f6650ca68a000375cb20ffa1a7fcd2d094bf78c1fc3fd7649e118d41ad8a43b9e66719b642e480c08e233d7b61a4d69f461c3c80615a74da0e5b426c4ea31967cfeaff110deb5ebcb33b11c8acd73874e7cd99b67806f101598a80f62941b9e53e7fab15d150b540bee1f781c58ac2a6a9c0d4124292d1ed696847455e9077604997037a2838d6f92ea671168af4b60785a98347fa3ee89dea0130c822e31e34b409fc1ff0d99ad308332603c43daac042f9a3f3d3aafd44722125ef6ab622059639004607b2666395290259ef196ab531b051931827e2cba03b2d255ef20e3a21a28b88e94d3405a09013b589882550bc7b8e2ca5aaa5eeef31da45621c2cf034bbccf47e9498ddfeaffe44111afc558644f5b6f1d0644d254b19e6f51317266959b7030515eaa22dfb92f10c37fe56ba6aedc6e5a8d27e289faeceeb7bf9a61324340c91596bf019b79bbb7857f7fae19267693a2b3d8740122bec0af62086d63f9558adebbaf44932c90d3f75b24cd9b9b5eaafadb1423a310c7b30aba0b03115782589d4d3de0b3dbc482c0224cbaf6c8f3223a21da6b3e255ca6080b881a931386a419c078b411b04904c9c9cdad2e5bfea387adc703c26486fbdb1390b5169f9b11312e596b58513375975dd2d415e287dac727b3a7fc0f4d794bbd5a05f386a069ec2f048b07ace12b5c133b70e69379d4bb858653e6f4535e3ddd25f95dc49f13e15cc48a639263171cfd94f5448d837964213e241e2180c6d0b1f70066b22cdd4e4a7a321943a3e629185cfc77657631b27c2d717e83e1d527af7222091ff35e1111e6a049ca929a9f242e3062fafae4923e5e95dfe3bfcb28a886f276c7f373fec41c2d4bd04c4996fb0107230da754d21345e3898af949b33fdab96d5f5d0ea50067f70d956cb8c41e1e0461e844385be6a358ee4e8a13709251f736b2747ec3857c31103a34697a3ac8c0e50c874f23349b3412732dfb357c64799c54babd2db2c8592dd5f12f3230b12f89cc4960efcf79d04f2305490d7e5a2b2d3487f9400e9e08ae2a753bb4aa372a118f4b0c419479eb0c2d5a59197ac9db460f10598fccc9ad20a3c6bf533894b736e84e059da27410ee038eeb6d86e44a49e6445d2763c5e469641848774cd4665edda3da66957f3a871caca67851401a7905f0365d4c263c6a3afbe604a28a159544a573920bc8f0ed56ea46f36b6ce2114b98762c99a1373856604b0e7c4c605e4b991ef25ed093ef2ff08d56de299f27299c85f5e63b9bc5b09b600a96de4630e9040f9965a2699667757ec4c5d79198d376b80595b9d4d970cca7579126f2a769666bc7e21f6d3764ba7dc1ce2475c5ad2605c23bb74634155b41a3f53cc96857a45a0fe82f58d63799e805efdb94587226bc371db94aeca647d3d7a531d24fed604f65aedc454b90e1e3c346ea18962500142290ab28085100112f79109e87a4402a35da9dbfafacb2d2d072006d766106b67da90120322fe69e3a7202d4bfe4647934952e2798b6bc1bf56a69d61a05fce792b0e4ec4b15503ead7f3332851fa431e6046cf031293724123ad67e735dadd720be712d7eb9609113dc051320408d74aa24250b80dfb6da54047b322c69d63b0dd8307ce9ec29e1cdd008cfdb0d73e8a92a0231988ec15ed8565a6fd5f9b16050b0aa5fa4e56eff6cb905d795dffe7dd98d033d14ad7ce7b9aba9034087f96e3280cd77b72e5686960ccf5ce3c3762f5e9c3a961bcfd712b23261cd59853ed10ffad469e393d3cc7f977c4b8b495f00d30da894224eeb6c6cea15ccb8bbc1b76baaa2c082e0f8f7d7bf1439ac9e729bb32cfa7fa32c5897f713a5f7b247abaea0011e908d36072755478da40bdd56edc4b2649414b5ed0c510f897aa0e0152c4be8bfeb6da89695a2be11890b416bc2ba9c62110a3257e555beba119f41219718fa8a8e7722b49e8e2099e3c6877a9523655787fb4571c98493faa67af1b0220be9c2b9c4e241aefa1a489f63495106d75b1095bdb0d8f082e3c973abaa81974e8da6cc8d702d58f3aad77a9f0eb7c2f510ad0698a5c3122bf1fc456e4d6484d3313e5afcfce1aa2f5e6beb400540ddf8fafb5504595ea9b00b806e1c7f0603a9d149a972335df07b9836b824f5fa4e8b2fd3083822f0306a5702c53ca931294d0ff84d910787bb77bf943a374d38744facd4d743cc143edfad1cdc3e9291f1b4366e1bb9cb8abcf256737166dca5f65cae4b9c33bd3663e345f9826ea541090b60e8ccb41f4753696eb7bb07a0a1627abf0c0c930d98260f19d517804bb759efe45993b4544d7fcb6d86ab555e7955dbf54bfb7af7a62cda65b686706c5b019fdde382921d6100649e7ae330dd315a01c9bc390d87b8a6034391dec5bde72e9470970969a9ca27a8cb85052ff6a25dd9a20978672e7b7695d65ed41e771119e03b410da015ae2059b51d0cf6ef80a7a2e7329aa476a8dda6ae5badf513bbb183912ce16a8fa8954b6ac3d3b96865a9230a0ef170ac7bfd5287d4d6f1ecc012bcdd241aa30a1823a95b8b7f1b81f0df80d7ecfae81b9921dc27fa8edbfe05f9f10f58b81ef8b5f4be8bca1fe1ebed49b204f34be39eb39d8017d0758c222c5c4d9140c75a0e525798e47db61bef79c399c7d55a39d197b556535593a0a62c90885be9aceb43b360287e43eb2ea47b7f1554935f2686ab21bed5ff4f25e5fc1fddf2a580d6e3a5bfe9a9eada0227a23043d0ed541458ee351093358482ae89179dcf8a15832b2d1f8ec95f85d3e8b405e2d353daa1a8ceba68b967637f053efe7dde5198dfd27d2d41d84424fe20a9910995f8c752dd7a343feacbd66a3ff09df3dc82d010c388ebc95cd027cb1c8639ebb036ff170b5ba1a2f4a059e911c04e6a85b33375e066643881926d73b906d9cba44cd6f767974bf699ffc8804832b08f7d51f87800f7c9a1321def31a29cd96516f6904bfe12c86318544a84c7d5d29c1b6660529f085685413fdd8fee87a70e5565c620f5d3f82f9964ab9416647dd673020f5bf354f5af98e9afea16c614f0be8da5201dbcf5a8cf1437bed01d669753d58c73014adf409ef10d248a9100a51bd612a6c5d562c836217caed9980183024e70a3a3222ed92e67a44083e2f243e4ec33ecb24027e90a2c3a543fc871174bcff9dfb404ddd9f60fb92f4b001f7b791598ed8e41c4323dd42748e329941fad1decfa880adc34e4536bae5c6f01ec26a6930dfeb231e9461d5f3b19a409aee7524a7cb395076a37b4c1d7792005cabf6b412841644456f3f3df7295e784cda0356964ad94f82ad82fb012ec5ba46391ae390659b86cb5df8cc6885a92b2a361812ee8ebe4cf9c1bac0fc886807e155f4f7105096c7bb021b2ff29a7440d8aed81e4bd4b5c3bc476e1b52512cc651525aaaa1d44487eaee4fb46fb640f9c8a7e92134d3510a8eed4f4668afca2a271fb3b05e3cabdbaf67d8097e29d072070df7acd0e7f875f7a1955f7bb440451fc355a96b17683dd17ef5ad683e30ff860513c1552a9822c36ecfc78e09714770e0c7956b528c27d30d03c644ad803278b1a6187120775fd74e0d47e9d4a8a8fd0d55722f67a49a6a0189caedcc26132e7ed52dded2dd93af8eb020fc080f14ac7748ae307144fd4bf21a5ff0435974b92b27a946f1897d9257e23bc5df3e72ab95359777be65020765a085f327190e761252f95b4f0db9eb057932df527887f62063e114eeb57b669852107c04eba6f7eb10b79734a834f763f0f2e51ca548c84c71ecdac18fb1ba92be36554baaf872d6d037d1e1c0c25eec461ceb9c9c648cc5664f15273883a1a66eacf4dfa123960e1b5e8b009660c1c086fc2eeb903b6a4c4ed55036e7a52adbd7479b5429ada95b448d7746d10dcd1cffabe37930346ec7b50928c5673f19fdc62f79e0ebeb2a002f32aa351f19e1819e3a878912ee5f800606829fd93582e98467f9c4e0e5ceffb5b58344f01065dad7f1e8a1d123646255108725e9ecd72d5012f8ccc3b30fc44ee03b03298590bf53d90641793fcb0b1912fd41656deecdce6ac165d91393f2732491d5bcceaa6eb1778354838fff8b4b453745e00ea35956a1d99742186e25108f98f7e5e7196cc350a578d31fd6e08fe5287c1f7403d03d336dfc45d992d41983d5c4092981c6f5c8603aa1b90104eeb882ea45ad8f9d5f27845fbf95793321b290f70965d6e116c8bb071e08784c8b407b896daa5f6e693a1e0749390a0c906609140ffea813cc516747c172ff3f89979803268f1d7985b20bd084ea9cb260b61e5201f9ca68381606559f6a2e8e44044e173e1341bb8371c77e56b14d6dabe53701b718808e58c3805d1e451d1b2b18e8e8f2a1cbb98b115a4134986dc677ae85333209414786af0a0e82541fdcf1fd4f49697cd8b387d801d38633a3f37cd57268e0cd659b26ba00019d781a6370d041edfd5c2184cf80cbde45cc216b04f3748b399cbf2ca82bf77634e6ee4213e4113edd1223dbafc9fd663b2fb21bd0a76b6372f87d5f78ebf1f8ced3bd2970e08ba02dda923e92b2a8b837572696fdd6afa637b49390f51626d07c71a4c683b2d18e3d2dd63da9da73fe7f39e543af19d80420540fabe88dae7c6a1c152cadb51257304c89d05c7fad1d9ff9f3a6d27673d8c0b055c55c97cd12c55cd5d3e2c512fb3e9aab5b7e6fa880f28c0c81ed6fee8c03c44d23142f6e4886d961593bf69c2c12750bb0727701cefd7630a079324323fceb977f24199a0555b531052d758973dbd43fff98447ccd313341be0d9183b2af0bbea62e39dc0408da1ca809b4317ba7eec6baae3d110b21eeb567d9e27a7bb8a32f43dc215f4c82c3c223fd2ba1323a52ba641f0f878957d964cc04a5f889a780395ae8b007690cde13a6701d08cfe1732abf4ca8bf019663d3e3989d917f61a05938930ae37ee7f012feb9a9e01d615a1ecb083be624489105d70e97ba1ac9ba46a823a46a697db5683d4db290aa2b054b07cf1c4e1929779b2d7fded8e252599e81997cc76ff0ac2697ea17b0bf5ffde999b7a630ca8fcae7a8ffcc14e592c9d26ec590086ffdf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h6d809f5f2b876b8ba09b819a2adad9cdc6306e08e74ab47374d7b24de7caad0f8524706551e3f13559ddf823d61e22e32e86388c64321bfefa4721d8f882439b3481bb28ac129451c7cfaf16794a87ff05c1feb63df0c572d5801af505888acb53b5c61050a7b69a4348c53da2d4f435850fd72f6b718e8138505253cfa10200f684a982ab00918e088250b8bcec9de4427a8e54651d0c0cc3e44e7e17ac210da37f5869d77bc1555458f711b6fd27ede6dfc6d504cf0721d6fb7de32d3ae47cf8f14ef88e2cb8899b5ee496d83361619f34b3b38048e8af05b85c14bfd8a0bae3d0afbd8dd00b8df98d7b2deaa2efd48a4425b4e7968ee88ee6be36097765c9e376156f412e610c78e136ee0fa5a184434995fe3b207624a2ee118be6755e7f94f52cfc8a4dfdcf2111fc7a2fd81322f9bd11999ae17d100e4a464bf9a2669c7b8b4a2972f279122618e3152870ebf396890fb72e041a9313dfa699250400a578a22a711808225067538cf35bcd5747e1d5b6d8448ad78afd7a642d8f68b147f396af1ec7710bd677e9288d581d63912cdd9c6fc9aa89a1b986205591c58f5ce3c190b2612a3b7c302e4122047feff414352edc9fa8be056335cba82555fc21e2982f73132732c025c488c62a57f8acccaf5efc41af0c1cbda8753c28258a1fb80521b122bd8ffc2df2344e1beea8116d0e75fb20f6bf425f2844a8c8431456633eeaea1230529f3c1732330b9a1c35af06a0b346b75e5378dd737c9d1dd4aeac9e289fb79de9d09b67c95723a0013f3fdb6b24d0d7ef441134b8119cc2c89bbec1e9e9abc0d664e3112d49bd4cf0c12fc5de0cebb55db02e8962aab95e29fe29dc31047c8a3c726a0188ca58c395ea0f8d7f341bca093b62faaee5b2733366a51a29ef4ab2f2b764c88128a4e8e1af76241c50836704138ec31ebd6c9a1499834605ec57f36bd84e96b89bef224fe5e37ab76af7e7459d52c91a1a7c68c901096a044987023154187cf3622fce16c3e0de1dad8471af87786d192e7e8a85805c74e500a9ca348c10ed4a9a2d7dedb3bf058bca8b0caaa1a0341873cfc4f21a06b15897ad9ebca6c4e488c910253d4fd9a4b32b73aa62bcffde5dbad8c64acbda5fadab409708b6125216e347385f9d85d246409a17fd889e38f05861311029cc55c71032a13add5a30ce102df03bf9774a6bc4c2a924e5bf7ac1e1a37c2a3c347a81eccacb290892a70ef8e284bee52d1b9494f3be114b6007796f65c032a17cdd0d3a5b6befebd32401ff44a4ef0ef07bf40f48ae21211c2270d7620e5b736357f6a0218d58160e990534a070548d7ad448b76791511b8899708f1dc2ecb3af54a4c0c4277a4f53b686dd53ff6b7892ad8cc8e815edc5e8409c966624af809e318a5844bfda96a4983b4ced70cfee3b8b421282e9364d0439ddd3c180ab65fe5d325ef7cf7cc3d85cf29ec76d60fa415b5e5d8238b84426343916d481542f47094a31057d5278c2206803d10d3cf35d0ccc53293b051c156ce9e4161ce5e93dd01b18c2e298408d70910d88b5cd53d91cc4c2422b1f3c293cf716422fcb3ca8ffabf66e6f39140b5c7cdd93794320516a4ef8fceb89f567551a9f26a8013a5e2b0907af714fc3fa0c6987bc589954679487e506ae93e7de5887b5113c8f88b39cbf7c6b10d14eb4e6b7a651541ff8cb26777e76d6ad24793f2ada8e6969a7975623d14b305caf95e3a2b9d09b44d239dd7d982668663cb5c2df1a7113754b673c17f8ae87bdffe05654b89e9a624605aa069c549f58b7adca2b45e5dee412c0ede4ee5f2c2e886b561d1e348390ab09663d90e6fe36144eafce7d226ad9cf57e2a88fc75e232b38d601cb0b93f9dc74fa9dff2ccb2ad18e1a73435381997557c48bbb5c0f3508ec194bed5b71153e8f1cad26c28a95ecf67fa3a8de0e9a644e0e6b46b61ce2849be69b9471b1c0cdf98f581c1c2ee1cdb0f314cc78691a597227a32604aa66122c2c7bf2c960c18ca1700a890caaf22b238fd7216f2d0d328e69f623c8024058189c8aa27a789a61a89fb081740c91376addb31253a2acb9775dcaadfc198cc868ec62cca39364ecac2379fa6fe2c814008c3050b28fe012fccbdbcdb63ce2f605072f46e6bbb93d713da5865b339519f58c45f088afa5a9661203c8360a994d7a2b56dafaae4994d59c5d3663ae391401b3f830ad60eb36eaa70e5764c4c7536069eb593441146314751922e3feedd6631082d84d52d081e2a33f4d0b6ad5d03a85f4a982fec24f438aa516ff63baa1077191d1606c6fe94ce93ffbc77dfeeac472345efbe2780cc54efc59d081dc6df137494c6f5041c1fc4fe7222d712a9d09053953266503557ee3d1543fc0573f3e48b9ec5b079502c3905f26c9de7d2363babb99464b634fdf2f3a01fb6feb18459128d9864192756c40efbf1f365f8fa9dbe71b0cd54f7af25ae7cc28b2277c79d9383207e6a610e4c55ce9699a430a2ce039c2d1f443cefcb561df69db2d5c7eb15d8b6e3a31e78f5a8e480e71255db6b4575e44bcbd8a92cbab93c2f26598120a02b441f332cd43eb50af82ee0e70034e5559d2782ba52d65ff1e8235a9911fa9417ad25f637149dce3fe685b09b9bd15d1b51d8bd6899506e5cf558a48d3a7b7080ed3a20bda33f852b1305ec2e1081de4c76f9078fc97664bf9fb5ade4a4291a96e5133964832c533356dc9cb2a19ecf7b71c8125e4d585c3ab32a1c5e7c027f6542b3188d7d8b070e7f9d5fc3c3d5883ecc2ce0949ed623ea39850d92a18472f76f211f35a4d60fe691cce73caecc6587132b4e62d4d24963c1271eaaed10e7ff1565c7fad8a9214b95cd1a0958ed1cf625fc39682e45cf66016ac2faf3812556902cc2175f8e90ee549906455cb18d9b8447e35bfe50b36d6ed802b9a306673b5276f6352a07dba16895037882673afcb2b4d71feea3059eb12808eaf5919415e632fd71ce819903d1f4dc5c62d4a2d670d760ce5c02d32377aae683c91c08a5d3a4e40447de46b7655f4bbf17a788e73e4df70d70b50e029cc62d8299e902d19ec3cfc87c292ea02afd1fa037972e5318b50e04e2d043247ffd80be9d6bacf9d77ee500fe5aa35bb969263c6b1f64a6ff3c1f96e91f14aa2e82a77d78b60d01d7d15f9842a5ae948ccfe63eb66d08ad1c19fa51b95be953de9c22465a836de921a52d9a545cc8aa6f28d8150103f29e433bc773f61bf3bc6174268b5ba8cd988a64241f6596041e1555db495e4cc96ca659a6f228a54ba0f602963a8c9ead19f904362953aaad9c032f4bda60fe6e21c4259df6f2e4c40b3adeceef430353f4fa71f080e52922d6da7019f6d9b72d74f6ab2bbe2adcc5337c49627f0e79b3ed54d822d3a6b1ae1891c4c514287fea3ac3af097ee6300d38aab0f00730eac09d48e919bc02929028295d4256f4b2f1c18846697a7418d452f4b42fff3286f0e38ba7e209ecd076d5fae9c33d28eb484e066e7022e13f5f73b56aa45f33e3393266a74f62cfe0796f68a29a5e68d62a982529f3f5cc75a267e5e0d60998229ef54e0105a7e8036ee01d39431a03271ad9415875e3c9f0b5f0c85ad61e7f5248a4c4dd4e8f941780c329193743df5bee8b8e7a382e487f8344a05a08223f7f34d7a137083c3b7bf32698a4fbc2228a1b00042f6236f7abede944d0fb9be5a1f1d4563d590708d13084fb8d08b831d4620cab2b4f1b50e9745c64056eb55f3474e18d196c6691614413217230e62e67cfed77e294a814c972e4ba393c82f3f0256879334c22b8192f06a902dcc64cb2f56a33f59bad67ad99f4decadd6d25e7bb793d3a1e686402d4cae368a88b387e9bf1771eb510310bcb43cb2a82c999d86d64146fab54d2a347410a446a5363703004fa4705f4bf07c7a63c4c36e4472787c770ab90d651c0959d48304821e6e2a828940f5f339e2362b54474ddf3505e06d80972db527699af76540c2c8c8091347dc6c6a872ece43cf48cac46a504aeb723bfe6b867ad324d381540b97edc03bd39af9ad3269ffb58185c02ba7f8df9c2c582f2e67aab01f0713d302997889e2516a70b619b6dc3fe1e5a1f8d96f58810c07c11d8fa0aae47d44db4746d78eb175712baa657134eb406365acf2251fb474c0a954b1ba6dbce12d4ad341559f3af5d226a4dada5f646cbde1adc340917ca528650e4df31659ef4f91e967924a2124bca820847f6a45b8a32c7e39ab5ea3e2c5727c6e7dbf0167de03fd2b91171c75f6342a5e8e406fe7141b68abfcb6ddd8fdc80bff0d8a67eda8164f1bf436d93fd346d2c8202229f80e9a4cab36fc55492c76c2bb802106559eda335b4ed582e8b106987bbfeb08fc957628c3fabc6bb555c758c50528e3260ad95d6d7a8b847ee178425a28e96410d24380c5c841ba153a6ae90485b7a4146e34da7c6ed11a1c5593acf717c190200c12164ac9e6685bf07cd34ebb6a4526358d764c7354761b6c1a231c59ba7cd09d4fb2613a67dbb142b29f86618b826bb2d9a9b5f09210e4edb18f8321181f1832d231a40d61b546ad5372771d2f595c3e4c56d5de08194c5dba91c81996f335090c541beaba98c1475e6ac3f5dd662c033b5014b97d9339952ed207b63293dc9fa0a8eb996c31ad16126ed5cbcff8c04cb7d8718dfdcf593d9e14bc342ed8f6f260eef4001b8d84f39e887ea4c50d409cb57d0ec7319660e7dc308c60799d8d5af437802ac3c4c9c399ed11f94043b1938762e02e7cbd74e996b9755954d72f415b91d1a933aa8cae05abd43aa1c3b7c2249edb82fd1a3df68586373240242d360788a34b73da4a027c96d42b90e75e5dd0a4c2262212fd071046e7584ee913566a31f9123dcff5061743213fcdb88f6c8e5ade067423a2d3d59bcac495553d4b125ca4f6671992c626ec3fb104ac300a66e70e55f86dbff81b256b21235dca22fd742757b034b01e0da7b7e1bfffba8a3d0bb55cb6dd7b4fd876ddafeb72644c47f126d9dc47dd7b66d53735afc13d5bb64553fb936634778070c30100f244e984f030227cfb33e36e466ddbb7347fd7c0330858725f9d0f03e8691685dc7921a83124ef45affd3bc3e60a8f71e85c1820aaaa364860783e3f7c991702411c3103c77214b81f03dbedf18535bb4af24542e50656db842c2eba1fce958c66e21225eb39842f4da3e0dd363732ae0a704b9a8c97832b5e82bd77e40a2a47c08ea49ed14ab4612ec85bfa5c956e7cf05c8260e9a8179d6fc368b2b90dcd2fc415221b9d3e386a4268c6a710f5ebdd48fd141e3190b4ee7b1f375e33ed703a4d127ef7675e59352049d9e9f0dde20c67a180dd7c80760fad170907fc5c0423a6749c6b3b9da6d89f9ba95d0dec039768ff1f442a36cd842a4bf0b4fae1bfc4586ffe490883603501a3b32a134dfb6abfe79c4d7b57b13b6719235e7b072d35366b7bc373d44735d8667d3bb499c7e12d4b9e8ff2e87e7654c000dca5d189;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf6623bee06808c904dc1974ea8f0ac4d15d214ac1e469a44be3792839f495aa29f5432d876fdca9e749bf658a550a76b88a036eab5f88fbefa3ac0ddcc8fd5cc47b24d7380b6374026128c735d237970f9f133b16042a8e76234a68a1bb4edf4d65d6952b541b87fe7754366675b7a8a66fdcbdfdc3ffb729f571f078fa7579b1b75d318f35566b1ad986b92390e0a05761991404a22f1e142d8cc06156158c604b50a292416bd4527d2ca22ad423a9120446e250fc10308da74b80e749164d610fd5acb669a1a6057028486033d3bdca6616c45240308651eb8840181a73eedd8ff9a5c9944a06da54783e9f18e6ca05dd2f280b1465cfdd62ee00d9e09e6771009e0b9b2426d91210dd52e1136ce363c59100d5cf8d16a49fe1c5ab7e7023e1bef778c32d96df96a6b01a1d4ec2c38ec2a37976472e7d1cc62428b0b1beeb406c119162bf9d6bce8dbc667dcc58d33ce5e17c20e6ed2b86587235eee8cb0ef381d8c68822d44c9027b6beb2f0bb8fa410324a242a95cb5e434ed003c3c22e729d4ee3188b81be24e02dcbce171b8c2523b30ac55749ff0d758f3225454fec2f9a91d69d2cccf3772d5094dcc927b6a35c62a21cd5cd60196e759c038b1cd16a773a27aae675fd22c3a3b70fe7027f6907738efab521bd38667d666cc00ce61da4da40251de378366f7005866a5a5966c8454f91604fa2d61042a4eb3667726a4a3fd16a47ae6ee7ae8b41c53ee4ece04a50c64c8621798560c902475b7df50e2c896d974777c1a3f166a4dcc424d1a174a288c514f57075ee9186359e193164d925436464db68527218a8990704770b7c2898ce8c806d1120a8852952a3265c49c430dcfc445a715f7a1c547434a75bd61c3d3c81b46b8d1ef5385f5924137acfc5d1e00d4b0a28e3946af31cf6a525583b2b90e65cee1196aa6b32fe12a5ec84635f029611f4c626f7a5552bb668c6134e6927592c2cd7b4d73a29608752263023e99319ea3fc517f6125e5146e4ddf97d0149b50c522b0412da5bc04ccb5540f0bd728c96eb6ccfd97ec2c3638e507877d028ef715269225f2d9502c87c076c9d0618d7d7c0af07201a1207b93046b70eac404c37f50cba5d52dd943da084189221c6038d3d0818ae111a4150b90e24397f4660e0fdf70b15a918257a90cf3753a5a4fe31dc1e572935c1cecb4db1a6bae114e47d7399e3d68c94197a16865ff9298dd26ed91085defa2414780b9d5af76e9a158d678154f1e0f6b05e6eefb8300b619997a79c2213e5b8d826cbaf7bb34b975d127d5a7cec60303a1ecdea894a91e704132b38fa196e04eb3d645f51436c1b545995cea62d9de2c3f71e009323abe0d9d1e6d463c1a2c2dd6c1b284c09ba755608a63431b97da5eba60fe0662332b56cdc2933946e241e8b28c07164d1e2c6dd8a3a5b4d8148bc6b193421b5df0eb4e41f0ee184da1ac0824be0ca096d4d92e933f140d75e3a0bd7a667b063d2fbc67ad6386528f7f03b304a9a81a7f39b2350f68b1c9e272812da9e09fea3f593e1f8f170e7f5df770786d2c429f7d34f4462db60614dd8b3c2ea3bf948698138fce8a7a34b969e70f08b13893edc0568392b4b676a07fb65fbd3439db13b6516fb0f0ab80e76e7eb702ebc3360588a09888121761ef7d946d1aed2971b482c6c6b1522a6cc377c9add352087ce510e5aa160ba983c175e951e3e7010414c6db13e52c4b9355f12f4f2db28c531412e3ef5149ef1192153bac0d2bc02e96011747759519dd4b24078d77b63471703000ed4ab23b9d3449b20fa2f490595d751e7e72a2c7b300155d763108796f844a3d923503b236a9b52dcf16de0731d776fa37ccf722a341f5307029ab8c1b61f53f3288334ddee8a2e32ef5bda657ad2bbb4c8b715176667b5f0807e5edc53b6ee74416844f0b6ce7371b38a1ff5d172384eebf8e436f93c48cf10902c2d0b92722d724ce72651c1832b832cf0efda1f43189af6e3a3f62bb4e91a6f317e83959e1f31560ee7ec294c1f94c77cdc389fd11add40df211baaad598536b195f930bc2cdf2695737504a9d75d09d44ecfbb5175639d76da8d7490b2047acab0a36f062d9d13e178b9bedd136f17b2c25b1e1819542236a78a1e7073fb17afc9ce03729e0354b67507e4a1ccdd8cdb676d1e28120a7eb48ec0502602690e0222a292ca7f91a771b308487a2b07addfdf38197e22d66bee88390c86523c06cef086613a8dcaf03f693eeeb88e6a5245ccd339480ff9cf3320023f52da258717f28fafb6d158c354bf1c997e5eb8f405c9c67957ca56ec95637bd77b3e7961412af271a604f2445334553474af45d0b262bcf8b40fc055d2e7977cb7d784d41475a48cceefa3e3095d2e8ffb33068be39c2c61b36bce57a4f15b326d65954bbb351179ee44a6d59b6d6ef38f1f707c3c4ad02c2f5803e50e5fae4d416ef8b4b62dd4b4097859da7d2a8eb5c09a86cac05e1a7ded18e5a037d6f8c5710f8070ab7b3abf9f5247cf894e5a5931a3c1abc3c5a14738f5225085e8fecde1f2d047b92b51b4a9838d470161bda69b5a9e9fb830c09d48a90696354f1cbe700f03d9795f260df32a12dd48a86f77e2ed66a85f4a4fe12fd64efef5f3e29cc7b2689ee43b177d78ebf0bc88ac1de4210ba67de788cec9ddfd3c4627a5c53748107b60c6c69ef3f42d367b75602633da3d79b5ab1a306978db55b87f058583bcb39b8b724306b6b168cc2c37cf5e0cbb6d7a366ef8d57af2d2ded17329e15b190600b1700c7bc8cb4f4179c4f0137567b9abd4071f14082fc54ffad39353d9d1f63de2673ed6f41dc8427c5e0d5a7560147d5c7f298f4346edb8b904d5bee12748a743f07f1162b53a8e663c1c8d54df4a4cec746bb49036ef7e35c89c2bca08690a57fa68c4a7aa5b10e320ce098357d9d2c53315516f27db29bde67668cc3d7612d3755de225deadf3493be02ea6035ea30f802175384a1b4d3bf5473cf003849580141c2fc95b6368d03fee0f38bdd1d18544c9b2110d531c868c9451d334d524f3fc2ad77b05474e1ac0c5f421868c8719af10e7f3546ee589b02ddf1d3f60cff2404b875d4e6c38ad5429e3229c18d17d272ae0f8820a910ffa6bf8900ab907ace2c7603a318af52876eb7f65e6f4ad835c8b7d5dc0c47168062fe62047c2e4f200c7c0edd6d3e830c762a3de7e73a8b84b47836abf1f92bd766b9100d446fd1b4023dfae56c8f1e5595ad4945e40ec5a4790e361c691261609f8bcc69c8bf99fe5ddd802673337db3f7a3159d1d7f0d687d595f18470696955baa77b6b3772d2cdf15c9d9d9e84e5d9d67fc9876d5f6d7ef4aa34120d0ea0307c6f4c49c3564d4242eeaed373a25d0ef896bac6eca2cec69fe0c5e04b6fa79c9eadb87077d38120d13c11cff340adccf2bd03fe82302dffec82bcf5921ca78cb497780ac1c04f9f49212f4d05525b340bbf4786fee1ec3dc450c82b5a18c304b09367a37a2d403494fd1302fe07095acecb23dd54091dc1f2f8006a85dc78b57dc348cdf21da6a44d430fedb6228610442059de91674683f4018479edaf83a736970dc3f44aa213cc1e4305c7b82045c20985fb48fca7625bfc170f2bb92b8d9b710b69576db7adae4ce4177992f007a0f072c86d915b13ab0a4eac7093ab081eeba7199ccbff644605064a19b70c660fb1dae8a636bd209746cafce9abd95e4feca1dc0f1bc01c7471275c4a8ed532f6f12b65250024c965a11b8982608780dc4d14caea21a1f5c05ad1024d69fed6186c159c37ddd2fa483ecb510e49cf4012a351e1ce523658a9a56ad58a1444e5f72e719c76474d5e80ccaa7ae3733f3fc29add2d6e05c58f0c1469a717bfae2a0cc551701f6c6c5af4dc68ce8465153cc44d5c9d47279c82e51b7d2c4113bd4874edaf7a8d3b9578df898d01fe4eb1c0d21eb5a525a82ae2aea443158c197b58b686f017642612f3ef8606a4448786202bddc1bd6d14b5f6db5d748718817751841fdae68e939f52a1a7c88cde59865810350f7ce64ed5e424811a0b691246a05b7ca5bab32ed25f09bb1dc2e6e4e2cb91f178133986c5995cce72513d58945e685edba15c9a32310ad504e8596cc558ed3d83d5c9fb5785e1cd78a8fc3120d2bb7dd8d94baa4b11f0b7d17f4ed8feb65c038e14dbb52ecafa60903c30285e6878c41bb383e7bb958ff7f7f4899ac80dd46d61c4417727776236d7eecfcb59d62a26809a291ab28f70d7141eee99db7477ee40986512227bc2eb538536ba7829d0bc4d4c82b2339a59368167f87537aa915604e7cda3ccdc60a581aa859ecff80a5e9dab6dc256ca2af2b4e0aa7c99f726d0aef0a78f7d5d67a8afa69b19177e89c1281fe61a706e783751ce931aa846e47860c6af6a0623b05fb563c8b22e78efb9fe4ac938d8a700405749a96d2572e1f0af5795c7093ef8c31f0221c6168fa51dcb0c5424df0330abc6a4c10002166b37bafe617cdbffed9bb9eba003f80367afd40afae39c91a3a2558a2a4c7d288f833b2ec723ac4655917ddba9b13e3cf8bb43bba01e01891faf23eaf14ec5066097bedef72f4122c10047c8b943b28e5a4387f291cc13a396ee2e8841095846a356d3fcdf71b5dd0bc3239c729c3d67b79a1d2cde478f1b7bfae49ef67fda7f69cd7c02fbb255b07b667b5b735bb924751a516c5d01e2402180c1b7ddee03ec68d464868bf908ceab24c2158388e8443725976900f37cce45eebf8327be5c7fcbe0d89f483406372e5f122b4094b4a9af0d090565dd3ee75932447bd7a4b96994d82f8b37f6c86b9f9eddc7cecd0b7af1ec907353f55fded34cde88a1078400c670e8f4ee2b470840d29f1ed34856a4ececde89e8fb343c5b3d29168a5d7a9a2ca4f66c291bc86136bebb3e5e0215cabf4764431179c877b80fd3a38a495ba7a837dc8b614d075e7084a9f5bb3e7fb87f6895be77693d61ea4669a8ce5fc8471478eeea67bfbdce126713e76a367108a9b84b8536ffcf0d6dff4ca2755825420199987e2ac89f50a7603aef275284825ddba6ecb6ae1314574df15a13638a20e2e221f1502448419b6b4d91e80d1ab4702bfa6889ec5fc3350ee46b478e413b99ca922f74af73516ad3657b94d4905fe79bab419e21af4000c4ea6618ff2b8ac2f2756427f4d791fa97afd0cfba5463504b564e2fd6c8f8048092bbaaa44cad79eabbdf4c91843e09e3a5e6c3ff112bcf66cfe0f56dadfc5f6252ad64e98e4998ddfb1597f7839a7c440730de2329db6ca053f693a142a80530fe9da28d7d76406344e7c36b9f9c4edf79bac503660dbc6f9d5205e5e77422a80e72b70834f61709a7d7ccb68b974088a38c0665b541d039c4800ad862c1347362447ba5bdd5ad248a313f16fe6ba816d9854a2c0da771413628b64a25185f05ade8f70b487954db5cede0c54e2e9b57d506834ad3ec1122de5f0ca93ae5b957cacd85f2e5e47661c64218772deecc4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he60d1d8707cd24d770600cedaa0f6c4069cb079629789ff90a0b4d049b2288f01fa761a9c7a55a58a5b05f186492f81742b61d50e8b2ed28bf8228f2f361a63b9c6d3d5a1da21127e05d187d45557418f0c4fae9521dc0c292befb02c9a89113d8075e7f84df150c2324cc618b33566bc833584f54f7f992cc3a56f286f3614bbe42fc9283b02c578815685321fa317bf323d88d7d4e56b9548186ed004923a263bb0744134a273cb32baa85b4e74fcefd61310c6445d8aaa32eed632d6b8287a0094c1a7253d9aeb288b27ebe82e9855d95ac6b8a1e29104f20a0f36061ce6de8690208d1198cdb07e63292275aed44b5457c2d1b3f8442e3a8a87e36c5d853dd42b87b757d3b4a55de8acb1ba990b1c65d2d1ffc158512615fe51eb163332f6ba0927c79f6a1d917bc4b6dc54114e30ebe5beaaf437b9985be55d8b5947c9c22eb3525b24c5580b326d786b0c57e77c7beb4ea4d2264c37d43f4815bc177f340031b724dd12e99c5508da0e80102cce89c7747aba4805612c7c23a413a9665c0dbf7acee6f42453474d02c35f94f0c26077381020f1bbc337d053e0547abcf0b268bb7491b65b8d7dd8acde26a38719e6fb7198f03cb87cadd97905ffa2f4ad680445f5dc46bf524196355fed8bf34fc47aa2ac6fc6d34e136d952464893d34afb07e2b1051e1239ac137e7fa1a3a41c93b4e582c80cb2812778ba0db9f2760ed9ceb51b87babf431a27bf384b2cb63bffa9dc059f1eb761054e4903bb53a18e3e63c37b75eab26f449fea770f2353b0b2529a5867ffaedbe9a1c48283cdb87cdf782983457d165ea2e8250f898b912e28a7223885f8d23d10e28c71d288d5c1882a45bce29426bf4014d08980106930a32aa307d3ad67e3523f0f200a76a18fda3c16d2cab8682c5f10e8b6442f1956cf6d530972819f790ea7617a688c1c9ef38c5fa27ad83c6ea05d4a7f93bf3fe2f1c283c06440c51d8ba2727db74195ca57e482859787fc0cd4032fb632c264013eb35572ddd8bd9c5a8db135561433b585f519d48cf7bfcae4c11e7112ffebc01a57ad8929bbe0911bb28901d5a2cef36ec470b0d54a66bdc01a07dd0add13efbd2668b3fd710bd9a3258bad4634194ae19bbe57de0e2d1dc71382feb62d3db6185d29ddbbf99af0b11e1f63a36bed0e9b1771a81d6341194f723e3f5ec6d4918079739877e8881d5a56bdb6cbad073e589c3da80ed60b0c5448445a0cd120dc3b7e7d07d5133c67544d28b95187a6d1ad3cc7d2f2fc538fe7b79bddf73276319828312bbce3cc76cafb9cc613c1c43e62a3c75b8b2f8320ae40b303b82959e3d2b32fe9a2bfbf2ff2746bfd5710f750d68f90ebfa1d5ff907dbffbb5de7a50e62de01e4afff5336163001f1b09b88ef85ec95d136c98191d43af7faac0fa870ea2c98e85c74a32d05d17f8d4bb4995502712369a10f6c7fa41313334f7f552f00493cd7cc921a16a53448f2a78da8855f7763d464569ce8949359258d85636cd1177b81958a325c6a76ce0f5df739bf298557e50c708ae6f1dbe1eeedb3ac5ce634e77f6885c65fb81087e60c270360c646aab0a73b75e8153be0e16f39cdfefaf8f9044a1b2d7bca546e1ea2fef160de36d4a4981c46260b41f5a87d31c2e27f4cebef2e66b52f3aef62c9bbbe1b42d4efc3f93b098c6cdb255e9757692a3468b3b5f427c647bbca2df97d99e1b9b3671b6727e12ca381b8365ae508b012a0fec1ca0af694722986d0936e5588d97ed25a1b94bec6c6d307344fc95381f5a0969816c8477db94fc834cb38e8b41ea5317d1140a60afb21762616e11ec843e8eb6c05220a3a9baa6aef7a1668a00d7a56b565c9b8294780bbd89683dea66dde39b3f98eac5d37bc148de99b530199eb84b5b4f5e41103e94a9270ea268d317642b5f9347e4557b54df6c5f54f595ee31f887195f615e79a33efe27a4f36794406228f3eeece97e5d99a454f30a0425562bc6d28ce3f115b9a8133e9d51b3a96c3bcefa51b0e4ed6825a7e808e0a3a16df8c1cff098c8384d486c21e2c1ee403ef6151b336cccf229a84a93a0093f3d5ae9534eda27bfc794865fab93ed8fbac6feae2de647591ac2b24fc6933167064a6e29db9dd5522fce0d18ffed1f59a7000aff2ff69672e4bfba27c5525f82ecbec5c5744e5895795b9fda4616108269e4c540211ec04bb8b987454415e7be79b4169ad11199093f7547f55f477257c39aaf825fdf864db0617137318398a6644c3c9b3801ee734f725788637c99bbb60bc2ccdbdbe6c447d3ee930fb4356f91b3fbd343e29ffed69d1e7069ff4c2ab7fb735768f8163760d9b3c0e1c5609c975eb5f6730fad68277a96be490138ed8fc16dd2e0de5ad607dd3382ec982b5b1c14900d52bb9cec2a09c98c2bbf123bb7594cb89db3842808b2fb37e78303a008131dbddd7eaaac83e62438879cff50f4ab433811a604ec58ddbc07bc2edf82c6ebffc1a4feb0f2b2b4866bd39b3b707ce8740e1fff4249b5c46c9d182819a375c3839e36eea429f279ea81c8e02d5df5cdcc4a983b5ba6cf015548152ebc07f0977ad5ec640b89a3d6bff92469b9846110d67fab218f98b59beb02c5420d34a507929f257d08b0c7a7859d57f638a4961529d1eeaea752b1ab9a548879331e28588f8f260178a8e60997c7e1046913e6d369ced2b1026287d91f8f0e3c3b08030d039a9e500d6ffa44d8a9fc8d36e500d4f317586abf354671ce9b04057c73967da6396cfbfbf1a9c49247195ff8d33ef167962d3713f744304ca1a22ee4abd12fd081fa705713837b7c8cc1666f24ae09a3222d53ba705ccaeedfb305379415a0634e56f2f370b90255e7277a3a8a35e34f745b4760babe80b35fb341fa438b15b82bab77e9892d3ba28cbe2a5fb5f66179c0e6cd2a6babcd2c9f468584305f532a6e1cbd9ebb0d7b0df55fb03b2b059421274f15fa5922af0d4544ff7ca63555a03b553bf1f7089ed13c509a68da5556899630c40be1ce2e75724ab0971ca5e03e8ae9a3c1547375f6fb578ae598e131daaaa96c0565cdbd5113df217075ac431a5006f52bef6536ac54ac6a23ecb73abc09361a95c89a5cd2feb131c39432dd2673f3f502459a4ce951b5282add3eb0305b2ae1dc259a255838ddcd5b3a7eee890d3a5ded5bf530d5715ce09ff263ca5804fb88e159a361ccefec8bac43373de71590139420cbfc80af1f65ec97801c50ca6ea7911a7a25e74fc48613768c7f82529b2c885eb2366444bc7d765a4f2673bf37bca1afc8591680748a1efe2cbfc68b632ebc041e22977aade25a9bfa4234d47d85c52218f4b6e25f8141d75a97f4ad88f9e0b1f69e5dd4e95511e0c5af36f21645949f35a282a879bf11a2f79f2ee46c9645a5873e12f32695c966545928fba799e4b9d4e9fcf181a68284323024cb75947913aa1c8e664232c67dd734612e235cd95ac5ad5b800b9ab1077c8e94f7c11d4d37576ff1dc04f96d96be2798af55dafb81526f833b99ced8db72acf98c7eccb1a9eb48066683b62160258089df21201e95d19da08a438b8e2c0c6819bf58397e4224a72ec463f9bf3cafaebe56a291278a3eed37f9c3fb31a0bc2741622a2c3f6157bad856a24c4f3c89917f2b5eff09ebf81432027922d0c624db203df30ed0003442236a85c2e0789e200828a180a1f73b1815e695d3bd6c79c011b9d3bbe8d032feefab2151cefcfa668cca794b78d3c9aa7fb315b639b0d50d26af7edb318ceb72feb1f354742259dbad322e836a05d790449415c8427adb8b860f57b84d7e0ea29f093bd09eedfe7a89b73191ece9a64ed261bc09ba0bc21fc2d4a2d7809771e0b519eb498bf7f535e45994415aa6cb15906fd1e29dce75cc452f33cf3483959d4801a81a61b8094064e42b957b0c25a69ac363dd20f3074e2942eb4e8ed3034899bc00035d739b7be9180b1b26735ced0f52eb5ca6c7e5c77d4d19fd47c745d30d5b6a2e9ae3b7f3738177841557317c7acf8874303761062a636a5b4f4c672b131d4bc2ae210451d0e02fbfc3cdfc0e900fa1db0f2d1870b7c920695f7f5dfd6c9c2f84992bd6a1d30982231860f14aa8366fd13a31e14e9eba95216565b53a8b0f7bf6468d54ddfac401b08aeeab6339ea0363c21124972b1144cc7af95242aafa38933f2a1863f4074d9b6f7f55ecf49fe18e9acc4412d2963500d1571c9dd949acf98f8f96fd1a01fd481dc1025fe8de5eed6c8bfde6cfc991dd2d617d1c8d407500e57e57f4bc8a572467c1051b7459c7fb60eabc1a15a637a0c6f709dc559ce9dd5a1ff7c290748bc3a49490e74fdee517afe9861b87980bbce376bed7656444f07c2685e27ad95960311ba25b18c53a77f004cf72fa781e1d56c0f2e69058cab11559d7e5643f8fefb31d42268ce5b1b8be0cd42e7252fad5fc5bb4c05e2e79cc53282c02d13f6d22f7ff7879ce0f8829ca631957841847b918479af52859d2c81571cc1a1bb57578872a408a60647fe22e534b23e90eb880415e20f2d40f60e9e6553cf87de919be653f8bedc948cc288607f10323490758ca9126f85e16ffb7a1f304c1797ea05a3099d78cae5ca10685375bacf5e437a15425905391058546d73368c9e0ac1fdffdb60b71d5b9d2ab5c32f61d3b0182042f0eb00b3a7e78f71ca08c9b0b9a613f49cece476d637f713e913c93c881a1fdd2c84c7646f44fb78f644cb072392238fcb84f56d3eef40e685b9e85b6c861e257775d9f1842847e275a2265932cdf164ffe954e5ef3825b987096c6bbfeb3f32718bf4998e2b1622153e6c75d44e6560e7103eec862afb084e3d6f1076f5974e6cea7ebe9354eb9bdbc72549c22499ab0fb40da2bb3bf47e11773cbf21f9c565ce8601b845c79539a5703146db81680eac8fcbe86e919fbf1bcb4c8bece96811774a124ad92ef0d6fc82c1f46fae25fe63fc251dc1daed10c8cb46fa7dfa4b5baede89c037818b0cba705aa5a43a86514b3d6aff1cfabfcec8107d867fa430fb999655c8e345554123500d273da78dc59bb9c83a1a90487381120fa0cd7274118cba5410fb8ac5a0977e70b114dc40750ddde64fe8764d5c7765a6f435077087e21573f588301e55c076f822673c098dac40bafeffd541435b7a11166d0126ecf8db72001c285ca8ae653b18b373155bf791f56e38c3679cfd6a92d0a17895a14332a79d9ec998ca59d1e103ca1a111de67ca02d57c961f11a98e3c66b26156a083900c0e7b920b477c422edd96ac2fcbb5921dca338a34145d7e0f5402635fc893a7972bc1ce0b8a4e5ea0a4e58aafbb588bb3449a571dff318c836f7c9e87524dff88f4b1bdff7b8190ab6ec094c6a45525e657cf44e8d56b68fdcb041484e525e8fc799e609ff0127d4ba8cd787d0bdbc1706d776446d846bb358117cbe5713222290a0a7c1139f3e4426b84492f9c7163bf7e5f2cb5a63647ddeaeed23c07c4d29c6e273ecd4ecc9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd1939c1ad3bbc7d5384be8944857a4860d24c1a0255a7995ecf1f8a23be4c3c37b0f84a043fdc84c87c8e67baaef32bdc9bd4f6e64907476daebe7f270b491ee6185a5c4151634cf146f2e21062dc7a28e1a21fdbc78b04c38641b883fd2d1140cb7898053f35025939ffa4f54e9f7d2ba3cedb39867f026b8e131e3cf4827e0a6b93c8c6d7ff5d0c45fecb67092183708310161d0871fc43de456da1a5e81889e2b80f9a256bdbdc089c8f7dadfda49d6050393c66d60c3369d0318ec3e106cac27b00b436f629d2a2f2dd131df3bf43d2d759f05108e5de9eda47bbccd93f8ba511a7a08a058c7223aac27e923c90cdb459edcc2b625184f5c7946fd3860a1d1b878d9fc427e63db34cdc95ebd939b32f9d784a586bb6bf393fdf8a02446141103c5b89bb8c9a51c85a5df849f5c1675a243e4a78b6d4b6066b0332d71dc84d9ae6c33e15a0548aa0bd52fea9d5afd12bba05a7bff35823a4a8988756393ec75ef49a49464a262d856842b6b95542b8846361def0179d90f84f0152dcc5483ef4d14cc079d3cf0cac4265d7dc1944ea4fe2c84c9e4f43395c99dfa9dfba7dd0668532e98d02ca64b0550bc13f7e22d7d9d0dc291104fe9a845bace967cf7dc6a6a4475f6b3b922b70125931d3f29c20735c72a48ec26264f25fdf3892a7f2eb056becc9c2d3e4190da0a8fa2e2ca83172cab591573f6203539dce6b6fcbe26fdcf89cf67d7506cb36bf0be7909f991201a629675fe8038fea3184f6b847ca606206771445078202e98fc2dd8917b8e12005fb499494894b7cb84e6eafe91714ffe78a0a1f9ed54da4af3c80157a396653711a045a2d18bf91a70995bd2c023b8e897b86dc3a70afa2821b98b39f894e23f62b8f8d87b9f6ed4b7ca38ea2f2097c5252afbe6e53f4de4225b669d67391d464cdd8e96bbb46b7091794e52289f5abc86029c344b432683acaf4bea8bb3f947c6af3fd7b21fbe4bb9692a821145143a70dfa5cdb851e858d0e101a13662cb1a705584f3e08f95d7fda327e72315ad75ccddf84ac3806a806c379182b975ed7cd3ae37966f90314fb7b6f439264d539936eeb8ab53a82ebc058e2f6eeadf9b5edf2675daa297e458838d4d4a6ece6f4b2da63d95990e4b1f9b5f4ef60eacd467058c73b43aa3544af1ed66bbeb24b83935f189f4be0b6c6bb0f56f5e950acbbf3e788d613ab28cdc8b6f1c5eb9d40ff5ccba9ddd03746ef416e4d573c09bb0bbab7d8a380597922299411e8598a93694b57ddb88312a4956aa8c28a87ff15c5d33fbf91d51e03114b6e133568be39024800720d52ae6c61cbabeb26136c527f590b155699e2cf8ca5e6bb716998d1f6ba33d5aa9fdbbe7de66d55db84d36880e5ada009aa9f88d58212095d108725a19cb4ad8dd5148193d774f6c680e46444d36aec6b3a1f01c315cbe70bade080600e3df923dac05ce5c46974ce212c972ed8d44632449c255065f61f23ea228041165190d0974fcd1c30fcc7bfb89aae55155639a5b0b52e4841b9459ccf2380dea1990815de5a874416e017bcc91a8584ca85d5800127d59b9542e5af07f30406ca2790dc3c0bfe06db86caca438e5a29a44fd275a6369d9a06bdc24979da8b0b83f331781aecb5ab5e614c37380792d0b328b5b586b33d8d23679b59f751fa08d1c9f7d418cceb9a2813f68f4ce74b870f9a7f491c6570531e07fae6bde45ae1c14d55731ddb2868153bfc4c8438d3fc85ed9a5f33dc9703350e969538021bc6148d9d78d28d4d73e2f8c5b78d71e20547857cfd8e5dcddbfab7f78feffd54652be23f32fc89ff1a915727374b60e720c930a53ae289d33555b44ba20f428e51ee44e9f3a60cf097092953b7a742e58975c83e987a60add636947577a8a32c1aaf5172923e05e8e8eeaddbba08d41e6c6c457002a788ee374608f026b542c46859ef49cf66a47d352b87114bab00eadd1385bea4c8e0251e3c3164e572515d6a5daff9e81bd5778e58c5257291c24d34964d68d9e55e4da0130e68795f9e3b81431237d40b0693b8e04201ac16c1646b9978663165b4ecf4dd07bc8795b0cd96ec4166a933f4c76de67fb8f09e9fd82341fb2fc876b79f0ae551970b4105f7df750b19b683842a15db8cdc545c74fca042d1c7e6971ce7a2416c4d91f6fb74950c11b45e0dd8f1b6042801c11be66c874e079de9857cacf63b6116130a52dfb9af8bacba570bb91c923d704da2ddb2adc2cf25e8e1931ab824c3c7002cc3ada259c59210277c1cd8371b453aeedbc05a0db003b34435aee1522e196a8025301a83a8d7146e8f2baa7c0ff0b5b0612e02255e23dc8dca52a9876613bc2eb856d2e28b492e31120af975f34366129015306621c32bd8d55c46c5eaa6a68d1345fe6088d3d5e6fd49456a4c6d19c3ff563a536467351859bbb2746920711a32302829ec1ec77521432645c3ba40b6bd3d79a34927f41a62e169651651a19f5b57d2fd44bf190d77593b53a06ba5902b7bb7ae9a0644a548d51057642f7c2eac27e92d51733da86e34077ebd9294f48671058b4e2dbbbce81118325a83f7bd21bf5e73477044e693ef1a58e4ed1f09ea123f6598a0c96cfd008300bf123ae50018e85e64d35eaf1c4c4c6d37b8a17c494f63484fa404383024e83a35d9db506da29a8e4876aec8c22ff0f264a68c667ac292b3ee66a9facd3ad4cb6ea48b20d2695faebc917b89cc44254369e44ebd3ae09907bccf602675d7c51950904c8bd793dd968675503bc4769fca76557b9cab737cafe2fb82db6f2ff68b43a1bcd081c1162caa16ec416ce2bb6e1b806a9cf554e7966e1e7701e6c5fc49d0ee4111b145afd98ad564e74bf11892bf42bf0349df2790676da592d0caa9b59a299ef54f3a5126f4b32bd137b61322ce65287324b099af54d36baf3b40fd29214de5bdced09a58d677e0caa69112e4c632867f612866df8a44632cb58f930a5db1a5940623d9c290e0cc6e907035db5f445f17f3918b699004e74e3855e1a5a72121bcb044424b29e69dd10f733abf595bd7ac99d313c97bac60a5c7cb5531ad65d55745e8f39568b2fbd9c4bac5c5252c5271173442bc782665c62fdc8dcd5e98890da3d80e544d5ec770cd004961ab1c16062a66dc63912fde9833406b9150b3c2a695c24cc6d8c59bdd1ee3c40c6253b0f5c07c3d4ce1aef213c8d93b3dd1843f03609e3512d7c30e833de89c131eeaa600684f37f45a4e94af86431f7ecf8c7e078129cda801ae9ec7e170e2f3bd09a2f09ae4076394b5d24a7999b43f964b5afbb2cf236c45b044aa454b6eed96cf8d9072a097a6477d9e5b24d9c29672efbbcffced3eca2c163f6937cb3eeaa470797ae542c38ed00d4b8180e81b1e4781667c97905f0ad9133ed193f6e07a12ed4f2e5edd600988b1086115a70e515b0b12ba9601b7a0078bd6adb5f32368aa92d92bdc9d21150f888c7704225cb392c1d3d4d8db080b194084c608fcd6ce64d1361e52a3abc350fb47eb890fc3b6ab76554e08d20bc9713629ac8761640aefe5d7ec7e1d675d507f6b5363718d16a2137d3378841298ba7816fa1b6deb41c13328b5730fa279ce3f48ff3829445e1d37d74cab45fe2565ecc5cb5cc5861452758c9d25a2edc148b331c031b841cfd55f89c13572b4cac1be2ab3651049f291212521c21090d69900b8a9e538dbdb099ec87221503a7ed1a80bd937b0aee2d5cacf2b93ac1d334978895840cad6a128e1aa5a675fee1560765c641c118da32b3e60f44b057ab539de1768d4f085ba3e1dc5ec6a5bbb8dded00ace565cd8df87778110326d9e5d49cf371af51cd9f910ca1cc44372c50d6fd0760ec660484cfd2a367b2ca82048550ff426536479a7ed8bbe1c4dc544b3df4040d6dc1e9f0a89d89cf6676c8d6ae4acc117713bc13e79046dd68c6b957cc27eae480a33afc57a8536191ff2980869643ce80da76a0763519d9572a53771e2533ddc246be012e6ceb7446df472430b1a253b5ce789a275aab02f86cb0897bd1a1df934cbd1b50fa1a070f4db43a3f41ba4281514755779751ccb4f8b94dd16fd74d9d75a414d8c9ee371ebba676dc1b20b89d2f99bf0f29f4f34ea7258eb98af853903886871bbebe57fc07e701b4e11030b81fe7dfd51f96a39d243b31f78efc53eea9c6cbe49ededaa186a9af14fba6604c0b0461e39a65602f2b0bdf942e6761050995a69ec38e026236160174c790ae6995dc70c679e40c76b473475579ddfe62234616807d932dd366f155d997e92e9265c47068955f58d468281caf2ca57941df06cf5f36a6906f693a853c367e5e9dfdcbb4707ba478684c343b6824d33e77d8c673d57ea38c3add9096f2e9957646529a610011901223bd4b7d3611d8c754ec361e59ba7f7538c13807c1cd10e32e3b64329188a7556326882693cc1b118dca28e84c06eee2dc719a673010c1ceb30fe1ab88a48c1e7894885e3d01d14019f8f4d2b08c71ea8d7378be0ada181acde19935463ce47fa2136a23a58e881a6fd57442294db85e8ec3b7c78bd8ac21e1f1739b2f92c87db497289d52d72c126216bff05d4b67cfe169c46e180fadc1ce8a76cd3384637404ff3723a3e494c96184d87679e5bd35f361d02e07b30041ac206b744a500d889aae60e6caa24d4e61fdd97ff55931ff5a1a1974be91988aac5c0c640cdbad6ab387857c7a48f633ebbda7fa675679de222c1d242b0f96046a929ceb4f6a6c6bbfd620b337d6586e551674a9f223df72769f263f785a19c8b1cad5dc346e602c664125995f1e413f40b1827778a814e15e6abb0cca915aced9b274e585892a2e44acd58111ba7d4c58cb8705c513ca0270dfd42551af8f201a15dee699bdedfa4c13cf78f593e4c8f2418930b5159728fd97334552a4d25415d9e816581b8a5fb3b4dc7ec3b94701efa90a6e11c30bab2316b0ff997b54e86b98a125499227380358898e8134faf35b158c2bdc53077eea3621807ed56c0e1d5e1ddf1a9f1bd653ef3f01e4061f6d8051f462b470b9043370577809b779fa8b6b4b1975684f532a7f6229f98abd51c48420f3c067404611be6d928728383543c69c1fd2203458f503aa977b6a6eb54577e3023150e48b3497c253bae75b7af29f6f1e9b9af08824cc837298dcd86f6bcf5055f48cbd045b36311582127afc3563586266399ea0e6d57c3fc85eeed6d3b3c0d27588b42aa70628a6c98fd899c23f16307c74211839e9e1984541df39b0c0c8e9e43e443f055df76e120df708500896798a180a8261b72f82a7f61637b0e4ce219d8d293986cfc19afe2a800487e81e6c7ed6a7845c698834bfb593e8f21e9b2f5643015c7ff6f8c81587b628b5b3fb8aef994b9c1d1a6a39d1d8c56308c4b485431902a9cad8c54073eb7244d6be665b8e37ca24476948c12150a1950f922dba665539af2bcce939ab05c84e4ffe9d1c81171690e9a486f6c8bf5b51fbe177e9f4a3e155afcc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h9f4d2b8e74878d1947056f6bd5ff549266b661e85a00f59e0b358b9da36840e6ce52b53e24491c8ea9a22ffdcb0e6ff655c925261934bc836855865286f69136c49ff064f6d94990e6eb429824c087415cbb448547e796a9c57c14d3c0e1b0fb88e815bd2b6f27fd5f1e0a75462c15dc9c902c0764c9af8b65c2f0b2097164d672ea53ac1e4f1aada522f77dd91ec12356cb5b27932266c316045460c5d78908b921d0ddef124b9ab5c31b1a503f57fa9ae0c087ae5ee0d6a3cdcd45420598469c8cfc744c60f62ddf135cca17b45351e979c9305e94a3e71df173fc093d7ddf9ff55c3f80cab6b29307216933e68868b97163a9c8094f7b1e4a7500c160b9153bbdd1bdfa9e32354bb701378b22f2b4652fb0c5c4a3d0d5ab73aa01aa79b6a16c333f895ec489f5f634186438e14b5a6aee6eb037fe262bdb313805667174509ec36695f08635397876d8ec16f2ee58c047046738d9f509b71af494bae2491873e931530064f65a4181c1ba3c8589019217e20e0d13969328ee5026e1bb91be196ca4fd408aff3c5b2bba7a50866ec467b5123b5fa842cd1a090f77de326353e3ed0a08feff574e9bf315ebd552fad2d45a24fd345c4674090c60d98645bea8f79627dd686e5a7a6245ebd89bcc6253f3576e50db455c740cc3713e41a567fb9d0dfd96db09e5b3445e60fc73c93c523ce094e43d82008e3229ce4e2367c987072bd585849975f867c152664a03586c8ccb53f1d4cd7b32c9b954b3f6eb442f63fed2f41bf36d0a3ea07bb0ff562877ce3674f090b48f9b10f17f1c0b1b4ee9944cd9f345222e913d7f022662c0dc675d8bf30edd1cd28607379a92a424749e1919d665770e6d48979869fb1bc09a61dee41cae89f63fdec6f0f63880e9f003b10fc3d02b61b2a79d4d23d19abf491bd48245a6b72a4d111201a69d0b1cd77033d09871cfaefa02f942ba3a2ded3c8a927920ad46cf3cdbdc63b823d2002906656dd45b901da4f119a94eb2b7e291890d1c433e4455f50200beb8f562de45f1143c712feafaeb286f1f5f722940d0cf6f237b48733796d5f99b7aec10a381c45c6a0271f77c900194a705418c9c2c9aae8454c728dd25a4a62f92aa6c73efd3994a5631d72c036f57e58af3ec55e34218954b8b5ad5df7f18b8d1ac06df77a8ad0eb5796032039b25ed3300aed431fde4b0157a4aef61b972c24f1bb5cc0cf48a46dd6bceb2ad18764f7e8844cf639bfdbfff631f5416c36545d2982c784d499ececc147dc26b25a765461664b4fc5a1a5768dc41fa36ab4d90eeeb7e79235a8e05adc97632b575bb81b1e57074004b40c9e4ac1a07c12e3e2b51e0c8373108959ab80fce72fd4cf14c572ce188ebaf2d8ad491a828469b01ca18e6a699a382e44c476b97112c5705f708b2dbdb17073d8447008691370b1c4fdda9392fbf8f3dd99a5c6c2acebcb512458075435dafe0276b7c432fb14f3cf651fd08ac87dfd7afadfc024af1b41895562a38faac71d0b10fc97dc3b7983648373b5ed9ad7de6a97d6522edab3da3f28e75bbdb754ca9a277511b27d268f7c01afdfd3ff9ca6c0f094ca45e3d63d7787f95934c43052a9de30e2bd098ac96f3da8c3404540877437e4b361efbd2d2d58ea9056ccac6ca1bbd58e0d77b4948f427f65b93a0d6fa87d525160f0fdc8a63387533175dba800366fe201ab9045208c0204cdef675ec5b39c578c60e74ad1ad2e7de408df77f7856ef09ac3473ffdbbdf8a8cc2cc27b3f52ba68f03d5dc46398f92e64a31c3011e40112428a887c80df7630bc781a6c31ac41ed22833ea5e1a75f13ec3cf74d6492e0822a44041c8deaa92aa069677352d59db1c237279271bafb432536e4c2b10bac27993ffd95fdde69c84ce78911e289a9bc392018a35f472db9523a804adf6a744c15d7bba352cc575ad976320582c88b4a115b36a677726d10157771f800e6c31f144914273fe77d15f1e9175741c546754e1096d9cb94ae605b9e5839b658eb5fd39915ac1d9167d5b5353434aca1975464972d55414249f912fbc4e84414f530c13afe0150a67359c9e33b7fa49dcae9d05d87672c5619f8ea6aa4f6ded9cc4a616b7680354df9ee5280d15138631db2a8688385bbc3b0988ad1036cb8731625365a1d823ca10f42078718be36a66ede6c697937a7aa63a897f49b8649e731a07d2503a42c9d09f1ea6b48a968e877907e8b16fb96700e5a99e222e74a01f4ba36973884a968ebd84c4f9831c84adf39c592c765c5e66d57a35045e75537a5dc02a9e00c3cc68a29b3a31a0dd06c0de1dc7126146cc10409e8e4b20108ff01529860d236f5afa530caf2dd4f24b83c2085a18c2e1ec44721bd69d0728cdbd077691adbaaac62ab6caf5eeb9abd4284e2e8cba5e593a5f0b0fb57b431f1b89a3f43b57d9834f6cc0c2f5a2c4012b6af770d608a38dce23efb6baed4e1c4791ddc9e40abb4775cb7b08e013654a2eba6b847c2c640b497da45ad20d47aaad7260fe5bdeb862058d7ef38685a0c44ecc449ffb4790c4553b5ca962463f81c07a025dcf5a4c70f4532b1b15e884cf7165b0005b962982539bb63d79283e8fa89dadb45f416494afda512fd643e126ac87d7893e73bbc4307ca757035d1ee8cd41ee31e4d926056464638ad5262ccff08690e7da9afdee9c4864b2ced25ab0f72043b0b724b7ff2a0790212e05d7983de6d2b80dc7afa2ff1b7d10521360e077356986e70fcc71a5d8d9384538fb91526283839026642ef4ab50da9c8a858181cb7bced446cafd5e2c069f292ced3d1164087beef85bdde74cd3b8dc455d41765531d042bd3caeb017bd90b43b9a406b5a9433c204777c5fe58e76bf16dabc3a88afe8a0ba342b252677a5448a839e776b35e6992eed94d7afbbc9ed504fe4001e9ff3148a3e16cea287f9e16d791862f73411c665f16d631123287b17cd959054adf3dcd15a3433179fa0b5ceaee8d3b13d785c3a99a34df24823022e7e3d23befa70607fbfb9157bb764f6d382b3b882f604eb2bcf9a35c10f8361f429c221625d11850c6b1d903f744b08726f1f6d06daa82a36010ebf8f97d09ae0e36b6e417793098b9a2c462f2f1903407151b0fe177d84450decb1315ac30a3d725c1e0309c55ffbe133d729c0d540b10db3be0137036823c6f685b450f223d89bcf79750af4c9972fd96d67ee6cb2ae1096d84556cf3be57387e1a74e69744ae0acddca802b2b9d4495a48bebf1768c56e08b0bab9a7afd95af6bd4cb10cf22fd963b2081945fa3e8686701773543fe5a2d53fecb90d2a87c9d9029edff75c72a3d946407e409086e642eec37ccae31cac68302151c087be5af0c85b408103e493926499d82630cc785e6fb96de998c4145570c9a67ec30d3b1ecaf1dc2242afe5141c2c76f8789117ca781109b0ece05fff1b61706056dd871f49c8bf6487a452271485297c9d50ccc90a550248d1b2d7d5a40dddb94ab8d3ce3079eef03bf960c6932a3fd852743c394a21d16aaf9c8bb24c9c5f873f0c203e31d81e4a8f90008beb9dd7453c11683b4dfd0401cc794033d0896345a6248e339da0ed5c8cf51cea6b74da2be3b7b3756bb4b4c7e13e3b47087b85e75e8d7a9152ef637cc353f86be4cbce30f0b282713a05bc8712de4f97797852c29b8a095fd68d73cd0abc1b8252c625a40181f67b0890807d355f314a5b45df499aa3af06bb9af5e8292ab8f0e117a56f2bd59750e4a2fdec5ccf71d8b081e55786515735dce75d813d9b59b5837180e3ffcaebd42ce86b337297f7e94563913413817eafaedabdc14cb52c8fceb89cc97548a8601aae2e7623b5a7067e93a6bbf64e539ac22565e2c8802992d5a07588347e787dcaaecf78514044a03c22272569178a5bdaf827308eb49e23a9e8391cfa500b33dd68c9d54013656671bfbbd76ca22e748b0e34ade638d5a8e4641ea6b2b16de8b9b33dc2d86673d756b451199c94348b57e561a47e67b2506b926073577a18875b2236b44ce6f80b239d59806b6504ab9cd537ceb11d23ddb4514c805f6403a55f956af8e6f9327af2519c5d8d6b48ddd7687bd65746ccff6162a733cd1a5d6c59b99acad58fe65ceff4522b7500f67ac43fdc0e2d732edc57c021125bddf1d79e725fd0e2adb3a79cbec7062daeb428adde0dbce6ec331663cbd36f98b0c22569dfbe815de2a8a7ecdf0b1925a1aafba41bc8c4ee5f4078b57c6d4b0450382a4b8fbe300a0f77b5224e11a37d07bae6243365d26240636fe4209ce4e479a19b9e6d14121193617880fb54672127c20a319b3a8f5a4afa371fb4642310bd55b26b96f82314f4141c73d1797d87622d09fa04323a1bdccd0b84667339d02230c7bb2223e7276f8cae21cc15c4f2eb6b6cb17845ade27755221e5a88cc11ec796ac23c61dcd32d24682c23b56ea4e6a9352f21a243b46a5750c1aa25ea0352dd09597b3b224fcacc80f82c3d522f6b484bbd614fa5330bc559c44e7567505083e57f4ce541018b8b70dec39aa8d1c92fdc081f0b5638d83905721cfbccb577190e8e6367b5d43df1b753d4ee597807072f90d64959c588732d558353cb6d3d74d1c2feae8a128b254cf5882974ad0e4ea8a5d0f29388fb00cc2f432377c1b2763e1639dc092ac3e34e1d445cea7f74a680aa8c990b65c2fc8d6373f53240c9e8051c2d0d694c213032c27b5c979c5951d342224d59b1c3df93a47d0673076448324dff5a134b0ed038a2ff858d12f08feb2486d0e4e81a1397ba63d4cea5ad5cbc49c97c150446ea1d30f1b67f13a79d92e57b6f140b1e3c1f18727ed51d7ec97d65a052be26d341ebdc53388e77264e2ab6dbf914ee6891967af5c7858e8acb163e7b9316cc9f0500aa1b33ae1abfe2a7b914e45184e1dd38dbc060b8be754cdcf9861f34f5f26c7ce936e039f310df077b29b551c42425730699667d424dd8cf50d09f25fe738b18ea962b5ed510a171a2270f0bb3e7da990c7454657bdbe07a1ef9a0ccde182bb08d50f48c13932e97c4c30265b5b6702950337eacd6bf81ef1399586690f81d72536eb4c4c195052949afafc7db6619697c5bd5db786f9f3b26044c223deb89210454c679e4194704c2fbfc40b32b6caa3f9c2544bd58c1e159a8ec50d3773a56d5de10b80edb1f0ede1f27e68db76e0b824db242f836950b316860c86d80e7e9ebeec5a821174bea5156bdd1974bc1aa829cef24941db24e7ec497ca9c0301267c74ab04fd65f858c375eaf7b01b52d704479c3d345e879182e5888fa1c5d1ec50e36794013492c849a9b50f39cfe9f395feebb158d3824aa0eceae4b73ac39338ee75e0de5d99be09f11200aea6e38a4d316b343986c3ded627df31457ada0222bdd250718db999978942cdd42a1ac066aea9c720ad126acc02ef06af737e778aeae6fd5809b8d4fd39b0086b226ab02f4d54a91de9db53d719b1a8c6b91f8662a0ae4005127bf2d5c4b4a9512d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5f784fea3c7bca60d870aab0dd07f403814004dda219fc45c5cc48c6d3b3530a2a4ab4dec0dcb0904956d4813651bd0b7f2e57204613ecfbe93c3145ae5eb2ca778a69a67b2700085e47199a40dcdbe8052d4f08acf30c17e3eba11ec15d4ed04282be7391f00933a0fcb3412d8fdcfe755de70bb0609c4b6f0c7df8d4eca197dc9af30df11f08dc680fca8c7072eeb030807b188e431492fc7cf409d1fcafea7c1697de631faef7925ed0e7e199e302312943af717842f2359dc2e248ca0e79fe238ffaf8d0eb0ea983cc82e21a3a36c681ce1f334927f65348ffa2c4bfdf275c5c6e1fed75e830456034ab535f2b75b5f3115d30db43807d7073aac250b1a077a8de47363791d2852307641e59d4536b106185a99f69339ebc3c65496882ddccf344bcab37313fc6d8affc49ce5cc40312a2aede43da8dcebcf589daa74f859922e86cdd2b16218177056fa58411f3181d7bcb614204b39d3aa5444a8cd390e476d354f79cb6ecf1190bf736b3a79e278c6fdd25e27b5843b6a5dcf1ee2a6408ba92f66b7b14907f15174eba53436dc3f121885df0c599371847e627795cc0786d5bfa3f52755cfc257de6ca097e595758b5b5a351965caec5f1c857f1b1c6e0ea38a02da65720c264b517c66b4d1ed977852a1e8f50c5b37432bde6838de95dc60d4a74c12d43ff8b3e46e1fd7c9989cf9a59fbdc54dae6c8f0e23694cbb6fa90a5f1e938333329e456432b1c0c64dfca860d7eb4b1cd61a9781505efd83b0af69516f4d2112bec3bf5a22ea4ba1e2fb8e3a68091b6e3c7b2edf97e3175027ec3c0cf95808bb075328d57b040c6724c4a7a3f2f58ef36c3b242c63c72fbd8841fc4abe4cf8666b397a6990c7847c8cd64386c548519b510e8df7ce7dbff09edf4f248f07ade62ab2e2b784e3ea75e99cd3e530121a772e2b6a7ad3b55fed5949113b168e19c7ede71a4abcfe400950d81c991267be611d051a011bb362fed88f7468c4177d4e35530ec8a7b873972cfd18d0404b64cedf5f485fa375f0ef58acece520b5872072b75091cb8ac750094a42473b2681b279ccf1d42691bcbc1770eeb92912560f339de9aceb9186401e2d3e405ff067ea2ccdd1a96ef644bdeb628af58a57550bf1897828516fbcb7db049ecaf2d2cf3032d57cd11c8346a8cab32ed239a42e90aeed92a01b7b88775c5138c71c3a6417856c6edd5a66292f010980182eaf80cc50a987dba6bdf3bd2e4840f2eba5c7b36bba3a75738fb0567f83665c58be0d0641a16ab6f4dd460bb2433a9ddc63c8b61c66a67fe7ff035710d45cd9f4861faa29e2cf1bf7e8bc628f22244800c3eeaf78b21f4cae8bcc7c49e2d0abce824ccce9ff7e785b0c5861c0c33fbe63d94ad28d836283e218257359bc70ebf1fcea5b2dbd5d5d3dff9a4cf6055fce130b6a3609d9acc72a83415db82e84071fd7325d4b913739280effe056f11f93da4606b6d3878d379eafffed2a1d489da0ed6999100310c0240d1cee77f4ee487c42a43daa2f9f3b310d4de915b9eab8959df295111df47020c53529982536edd603c88e410624d215505de9faca1cc8df31aa43cbc0a87de57f399b249a17aa4556d7db219b47d0b94faab70cc58cc6186700f0e87b0e78ff239c7e6f50da889342bdb1376e961bbf1f8be08887e5d80d13aba2b7c21a9d19d4655dd9dbbd4a4014a994e0f9b36ac974b8d14b33c57effd6f05600b250a5238adb649c2b9653e8a768735b13a5df96d81dcace8fa5679795d09949213387e40f7f2f49dcd464f74aa6c3fabfa18c641f9dc6d1afe20830e131f4d3203f808d7ec098adcffa2b95dee1e4cf9e11df28246b8a4e370892e8b0427a7c34706cadd39cc4710e94e34948cbe5c388f53323c05f32c5b7dccfd73afa4e874e0e83010643f8529121004b48c6b993aa5d19a4ee60c76c08cd857ba2c485aac766c77445f23ad45974a4442b7b5f7fd78d357360f72feaa6f0002b6abc936ed1af87a9c61efb25369ff60bad13b36a9a64944d6896f44134b493ca6bc510162f99c5ee1a55ef40d232c53189a37494b7d630d7f659e26b0053ab67fe7ac7a11ccb318ade4b607f4fbc27c6f08647cf0381626c8892547e00d67aa138f8537c738b3260b3d391b542fc8af68d8cb7ac35b4f392319991104f2b27392fdd3dc3cfe825b2eeea47188a39e707ee0afd6e40da7fa01b0107b3061158405fcae988c950613e42ea13bda251d10606180a2a36f95a8350433d58e67443ca1ad3379f975c553245776beffdabc902caa0afba25cbe780e1ae9015e0ab1f69b738de0967a3d080ec035f33c402bd71e9505343b0567284a9e44303bfb8fcb3dafe5c078e0ceabe42f4fae62f4e2aaac53778e123de456fba9b2d30adef9ce78859013f0b7528e45b2d149d52368e94217cee5bb30fe366f9a001fed318d3455815a3e3767fae598e15b77d0cb45c5828127038782ca724c48a806192c11cb27c0aa09b47c9a89931f351a629a70e719837be430c384beb2205f1d48c8047e035bca699e46a2dee047f1e861e5441538c84bbb89d4436792d69496dcea35d76f48e31f19e0408e2f22e755c27c6408f7ad094ac552592479e69b271e891bb2980649322a7755f97bd70ef057ade5a1b5f3a9a7664604e856bd2e253feb0dc9de72121dbdf592a75d470a1883a46068d9fe8224b89fdf773b51b60b59627c0f0682720c33ab0b5dfbaba3f6042c7b57f1f714f9d5300f64aeefdff9750a2935b5037ac808a011416915c6a633c06287c63accc6926e03eb4a3bc3905f5518b251379705d47b40c69d5a9389c545ef1caa71ee4d420c5ce286d51c60aeef8bdf7ac1cba0f39f61e9fce84aa0783d90505d9b58655de4e4d6dd6bc604f628827adbc90dee5b54505dfa7c6855c85e4b0323432a84dbd5298801a681dba423e0c51f011f5cf0cf0da9e110c79c544262888fb1f5b83caabb7f5ddfbc5b58b41bf15d9a9e720c9ccdff023f607fe326383b574496c6d3d890a7101d3fefae31789d638d97c08bb63de21d94a6f8d747229eba400fa59295b506516d5aaf3e23cb044bd91eecb43fc95f326c2bd9ef3c75dcc4e35a0d93db6758cb1e33e81a12cdf7fa46146824e61913cf037e167afa0e65dea8140727266db2779a26a08e535e1b63392918e428cf2e62c983463ebed249861f1a5a9d3efd6a4090a582c5287afc736e8b33ef4a1f0fbc72ad9b7564cce9a2ef013f97b3a6b843c4a9d1db7dfd97c08ca155103f5ba9304dd1c9564d07a2e894936f6ab09ec4e19035db84f43f164af66e9b6cf7d07cea2a5b5010bf02ad3671de1bc44affdad980d537026c462d2644c8a7c13df8f4d8d4dc982a4af975a36ebaf678b6e2598651a005bc508ce616855272a3a1e9a52992ba2a90dc674e8d4391da053cf40c9cfe7a1c3b687f5c80eceab74573814cb2108bdb3784bafea928a8403e30481e0d3ba43342749b51257cebaf15d7eeab92d521ed27c7d5bf3a3137813eb290fdd18922b06175fb0bdbda326902bcc2f6cb2926d489b51e7c395c244e4f8159686233ee298354398cfefc49e0466d44a9d314aff8e73d994b188b0c9bba0ac5eb7eb4cb74e94bde0236acd52d4c0469f28922a15dc274ff6ecfa66cbde2f9ebe0972c4721b29a76eb3ebb9fdc5fd35fc9b72457fc03ec00e6a628d1dad69a1748efdeaeebe20b4d648274357c37985a742cb1fd8fdacf73ed774cf69c2953bd69b8cec23ddf88453a227b1cfbffd26e0379c845c5914823de0d634a077e0dd9f12e0db0774f645534cf0e66e87a0c38b47818efef1f5ededfff1721e084950db1d65e1f1c60717e6882299b9bfa6246265b41e3231881a7a142227c55c28cee0379ada7f338f5c503d34a9d9345ed86e18fb4a184054970ce8caaa86a4599c5d29469a7023139ec215818f1858b7f1404442b957b1da0ea3f12971db5949e8775241a2d9791cb3588b3f80ce0cd10891af834ca0e5ce66f54a278b2246cc51181a4bbc9135dc1331669803f3cb89c163d6bc626ace37780f781ee8b8c2e12dea4bb46d79c26b18f1f032ec296e274254296213f1e5c387800a64206235109ab61a842bfc86bf273ebbbd4cddd2fbdd141cfc57259c2ba99efe1fd848de53ed2022314fec3bc6ceb05d4b9cb588e05edc949b18a31de7020941a1047e6dbbcc198e4ffe83759ad98d05da05fb7e3d4b800bbbf896266fb19e54b78b8688f4f38ae834cb7348561e4de64ff037019c5fc4337b232e1ee38bc8232aaad0767f4fb9d588f044c69952d5684bfe78582e1714d872fb3942376090383191edbb16346a4ec7e863f110ece47feabb1dc53f714776acb263ca9a754f76bd78d1924b00d74a953978fb96993aaebbbbc8ee5277f24f22610623d6ee8e9440721509bc921d1c7ed3d2d1ced6253ee233101314b381372aec5e6da1c5af4fd76fe94dcd91c604392e5b58b48a162849a0f013a23fb88072b41143b640fa959bad84d94eab9663245aab01ea2212c424141861cdf55d8bafdb65bdc9a1859aad444fcbcafa84ef7841184f73d05e689be89e08494c4a98683770e84a3cc2463381049338a67eabcac16dd61488d0478362e40bf89e2d5ae40f3bc18c5532ef27b63b6fd0ba20f63ebdc2813eacc71508961a005b00d0acaab8420a22ab5d72eee49973706aab7e208adcee43ce5c9c2fbcc96bc4314373ba45b82ff19e3e686b937bb09dc638e3a65167369a65e1bfdff6249b4d59e7f2cb6e9272ebd554307b74ffd5c0f6a171e8c53c385ddbdaec8e0fbde0fbd07753725dc28e4e2c93ae1aa4522ce72e250cc83e78abc66ce71588c0b1fdb1ba52892bef72e08fc70d87758e69285516458a395ea9378d25337299c5a082d7d44c3477c7f0bce94034afb5fc88e4e2f5685e6732ab47e15d21bf2485b55739a091e2163101809e3904692e19cf3f86797fc367457094d778ae8b6b0663977b405cfec51e670eae6ef969f181202fdcea04ab58cdfff29120bcdaf56895543d50ba6b8e7fab71919053fada56adf3c0e98c6912b872bdf561d00ad8a35129762873ac4c04e09e35420f9612cc817b7bad042d3cc99b1a6ee64ff3ca9989b71c603ba0d22194ccac78c9c4e95a34e5d9406e112ee27d914ad5b17e4cc894296a6ccb9347f5de748d775897f5d0eee00cccfead49f35a2ab20d81d1c94b71762647c11116155974d09c3ec0b43ea712ae7969ea0f5bea5762f912b7039f2233fccc794505ec1df78143a42769bc1bc9da096ec275c0a6b60c0e019606ca3959a951941f3f8924772a91eaa9a594be1cb812268bb0e1438a0a52cb3d566f22892a9cb05db27ff82b08d9997f45d66d5634550e814bc644f0b1651b18032f371985ee0ea99e7ccee9f10d231cad59a027923bb702ae0191f79c13daa7a3b1b33796f941bccd9b5db0644db90d7228d4bc66b2688b418c8ea06c4f65953a990039e4a1d7a1ba5caf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3202585e905bf0cc75a44dcd2fa5d807b7546a519dc2bfce4ce536e36e731e554db19571e5b2518df08ec9b090ae39db1e5ad9b644e22a22b28d9c99aaf4f037f2a47f555137edd3a192d03f81753cbea5381414f7f404b0394a696e9880f3102dba19972f64ee2bd4ddd0f0d5470ce1f3b1f3a953461b073822d7984d9da19cef24a575baf2b9582df9aabba57c38d8010c44474d777b4930d9c627007a23abe903d92fc9610767e21e91253c21d09dab9d943292e419c8dd4f8bb9429c5fa729e0526dba1a18ee02bb639415750ebbfbad2d1aa56c52eed1fe767c8cb14ee9d021b183410618686cc8b16783da1e8229884762063e7871369abd461c90b98d620193f17673a0ac5b263445486d8f253d18236bb66ce9aaa2cf7d15296c0b1051038854ac6aea9dd9b1f7e838b15f2f19357e921eed5f5182fae5e9d2f0c17f90923156866e7113f3b12921e6514a253c333359ed8f9e120d6d5bcd0e7e2e9a41147a885c91b90215b18dc31d63b78323e4cb6c7a2348f70206043bae87ed848acda44db6e6504d20e125bbe4fe4bb2fb243003a70bea4c2d2909c2ae6141eabd97484ab890ec35d1a96f9b0fab95d3c8d2d3769e2b3afbf9728604518e70f1a5037873f464d6fe9a0dc53be061a3c75c5966d9c5b021fe198b69e1544b7d374e1cfc6de7f0d26f4d16505d443a34ed82dbb3adc118ea91043c633f9402275fba4fba9e87476d2ff3dfed7c4f1e624a0ab58e1c6f2c9942f89315564e947f19b16ca4f615e3e8dbf29496cbb466abddfa04513f8913cae27b7748c6af168e97d8b3c1bca240174f554453e690b32e6db6c3560a5ac5a942403e27d45f33cd62ba2079647507ed5085b1239b96ad0d8f6e4af474f13dc6ff398655dbf2324bd71c86f753a9d99e65941c0378130b6ee0e624ad1ab5c1ad69a23d2b029de4c4dae861176bae6cda1dd6b0643a0593c0cdfbc9675c2fcfb81a16babcc9683fe04ee8ac9d7a7c2ed96b8b00ea34604b47a042a484fb111cd865d65f2ee2a4a19bca9af662dea465d0747b31ce5cc336a221b0046753797b1be323a2c91ba3ff5125dc901276b9606dd6a4e47dea61472b2528cf15c9bdf127d9e7486f313ae84fac5a1b71b7a12515323a6c94def0abc4e39c75e50d17a1dab5e881d972977c51b543f2cdfd115cda7e86cc014965264f9aac764e2ec337fb125a94e84b3c9940fe69d5d8018ae5b178b56737e2594f527eb82b6dde978b41b739b6ece6a603e3403c8c7c205b6681d09cbc4c96a625eb7d16501060ae07bf6851af5ba9854fff3b714eb1c400c0bf2f5a01d16d23cf62f0188f30d6acf93b7ee673f987ccfe3438913a5ee346b497232fcb5b5c840e2c543b4846120b0cc2415f99043755f489943090df43c8fc58c6437bbe7b01556eb8a0f2466a9761cf05bf4f6ffce5d8fa2fee643b6d8b054d63f373140fb92beb202b4f4b70982672206375c96a1fada9faca038f1c9aa5a19fcf904df6caf5b1463391fe1a1d3d154daf974ff82723a122f091db43ccfd508142a0c86272051c1bca0eb20fa4abe7f1fef4ca8b1b0a1ba3720888f25c50b360aa15304798c0afe968910e0516be01c7f8ef91c19d1651f6edacff968016e235921c7f89fff257a7892b2db7f597c11645c43f46dd135783a73be580d12a91c9bec2731dcbda93daa011d770db3465ed11c69bcffd51fb240b6f1c6e7524de9d3a7a15193c78521890a6f50a76c4f71881f9e40efa45d40d9a03b55da2f8b87d173aaf9eaf690c1d319e1c548206c483eef63d05ad9fe0cc32ba0499b7dc0608c448482edb056f21550c2989cd927c8f27dcff7ac8573722907a56cce9ef713400becec2a9d8df41214da3bfe79c05083781c186aa7f4877d921f1698db6b87166605f68945c8da8dd92b760ba6aa81b7da39ab6347d5e23844c195cef2316841668e87b5a3d8f75b80fe25d8645c09f4ec32771325d7dc1a507ec6f04dc466a9586a429341173aa29102212df65ebf7742f689d976def812eb06b41235e742ff7edf0944db50e2e004b444f0a430149b65bea2a94da1af9628e3d7fb7266e5226a7d6e410a446e37e1a403de73c0756875fba682247525ab7860a0726594be8dc6878a20fc23ec60a2320d2c8e49e460c8464d25f2428fb48b61c3315a7348956cf8121ae8e02d948179bf20bbb061cb1e49bf32240d22588c92e6b6c1198b342407a3f816623f016a5d5004c149ebbf6dda4b520102b7c4b91b0989e6d7b8eaebbb6c20fd6bf77185882b1e36434130e62c73e1fef9cedca7d17bf77595d57190938ca9cedcf4fdb1bc77ec9ff08505adb7418ab41305f0b67141d30951a7d01dfb22707f0efc5b2a0f9858eec2cac80462c5145fd774d92a587e2314c42a2290a76ef4627acabb9cbaf6f2dbc9ff2495b566ca78808c1575c69cfffa763fccfb9924ee433d6a431f5319e64179dcf248ff66bd16cdedb70c5f37b5fc49c161be87a6b9ba4343610300ce9b8a56658c2ccd42563efd8a8168a0047b017f5e889515cab2dcab96bdccbe654b3831842099cfba1229df8b44a8edb089aa03ed2e7b1dacfc0d7278f4e6be34f08ef5688514caee99794ea874be1e75a831e3b94430d2b0947917b13f27f78d53c983471b1a575eb40e27e5b16a10dfa54ad607b4c6612dfc120a0581fdf064fbde39ddf10c93cf26a39f387bde80993c22abdbcd3f59851f433d20f03d3356a2b73406622a265dca4012be66651c31df8c38f6c705b1acddd956a735036c64a049b088f1b215bf827fcb593a529052a415cbc66605a0d8a209947f65a344b776debae6fc4e17dbabb99c1b8fca82b6c422876de02f8efe6414aa06947c34bb31623f8e3dcaff451c82861dbb0ea2983b9596743daad8fe68fee69519e58c286f3ae792ae32995125454b4b8e69ec8e50de95c80add0e62ada1ef40ecba7acd4ea3c8e4531f872980561048b09c163fa6024ce2f2d182b2ce36ec481c1cc98b03ffb461ab818028f12f83b1af3807046ea587ae0a5c6873b3f1e3897c45f5ca3a00775d70dc20016d6ccf22bd26eb3c7817b15b47f2eaf7fcd648025b70d3ef33e7e0f89bd34e899a7523bb4dbf696629a313efc78c4e4c1cd50c696f81e937fa2cea6f6e3f3321038c672cf13f6b4271d9df3617ea685e75ef4ee33ba3e3ab0c8981f79ee461c7fa4416c26f32fedcc2b93040e4f18b581df344ce07d576ffffe06944f0c5a03a7627938f0fd8a8a97936f47523a4b802f5e3e26c44923660fbe196ca3c7bd1fae8bfdf2ed91a0a7b0a0f3b011f9130c9b3ff9e065a3616eadc6486c736eeaccd2d684aba4df2e8f985accc7ad05a0735139543bf9ab3d964ab60fb1bcb6902f9ec3478d6c3234bde0abff683fa67fc13ec95cbaaa31849baaae4c0bf0c147aaec2caeb1c969b192369c9f5d3cb313555be553c487297929e287881f402f67a25270ffae99943d4e2849aad1af15a793e4b9a57f1a9fd7dc5049160b15cf3794111e050154ac49834e74683f12e81d2a5fb39c942c0707a101897c35476a12dddf7d87dd5de3c9f748be19b7a177c6aeb5d68b246d8285f35d9356f93c2b2f3e026a8eacf56a264126cf801bd31cde2b53ce8c20d6254094966bb840648a06c4abe24db3297d9acbbcae322f39c159bb7b8b8a225bdd520b107ace23c445666e1a544c70bf7f1a135bb4604dd32d13bba5f0041ab9fab11d3d3f7e36910242985f892b10f0d525fb4a839094b7dd41c8c14ca68457540ed03c9721cbe17fd49972afe3f2741e1d8a4fca326bdc82270da8825aad37a43db704f40c61fe92ee49b51f232e7fc29163a716a283c1aac2e03ed829117f0a64988cb16819fa92ffccf1936eab1d641d351c6bf9dc00e058b4962cfb1bf9e220d376ba9c0c7f7e1a464a089a4056aca746dcf0acdaf1d180f30953334613c2ce670de06a369dfd21a3c07f739c27a45f01c01338f99477b5336f30c28bb13b97a82fb4eb6c9076baa1175cb08738814cae6a04219241138d8b2530e826468c7ad70f0db7fff404908584163cc22146daa94b532ddb89a6e642aa618d158ad7386c6502f9b3a2f1156e7bbd7470ff90168eff48b7a502a73d256281458d841af2818e67f81f76ca4977c41bd37d6d52f9c36b8f36503ecd508e56ff5d6aa3291402ffc4299c0667a4b1f31176f8fc98f1433436955b89af0748172db10677f9411bb141dfd0be6e2ced3795b8b0ba39310c0f7de025323ea89c9c30dd8973affeeca56b903ff050e6670da95e8819ec3f9272510d742d2391918621db3a87ddc6b417e1e69379cf7b3ff384e2729f9a63e5c2dbceec2ed887ef5c475fc1a72da0c9d07bcdb72b14565eab0cba0c9aab9745735134a2cf9a94ea8a3c6a1d20098a222ddc3cb93a4eb0feac5afacfbdb3b8b72632f240a634307dce0169dd84d4a20e3ab3e0759f17f27cf730748b2831cb863fa7a6daaa5fe5eebce3777c62542c2721b52ef6bc61071c085166707e67d9bc6bdd34e622e9b47fd71d353a570016931230fb28c5765b6fc3ca669aa47ccb3c0aec63d5662d5ecac0abb1b3453a13b265b0a5a87fa14f354771b802ab0e570d522a507d1c7fc1320a2c1830963720d3073fad4edcb03e6cf8430c547780bb3ae26bf8dfcf46171b63b1be3a9bc4fcd5a677aba0e5c776335afe6e7348a92d27df6c6400eb8ffd6bc9ff547021ef4063fa70af1c2a15a9c96af46db7ccaebb3de6ea3d368915e97f8d381b0a0861850812afd75cab05a8b1868dc3bb44cb673695a4a40c9e43105421c73d9901dd04cfc5c3a1448b1cf1d5b93e68b1d351eb227cba2431265ecb8fc08022a3b487170880f130a14e20e95b3235af14cc02602603010aaeb0d282cc8b764510c4f25b7db7badce2344408e3cea8f25f53c35144c4e2d16122f7175b8c57eaa3d67257b4fd9b1325776d19d63e1409a9ec21f0840478ac3378997d6ce2f8fb1aa7bffb923f3a25c7cd1c839c3540535b8164152175860b966630d4993140dc1f13610e060678cba66aba2245778fa34186baa612a0f27cbca06f37f8ee2118056305cbad48c4eb75fe63fe269e8d7ea048c9661ea55422904900bbd57b0a811e536adf2b0606d7a76b49da141803b4ac509ae8487bdeee41a41b718eda933c4b7ccbc699938fb689f6463f53bd709c42a96dd3b51b484f215ca9e83c7cf513eb0adb739a1a8dc8284220a9da9ff2bd9271ac850d9d71773888bb7ec6408d4bfd5c4d23d4d777e274e7df106ce96d935b7eb70e473ebaea20a5c4453a407d2f9b9ca3aeb4d649df45c0fbdc53c90413bc92971c1fd8cf52eb01f1c0530ba521bd8ea6bd87c67ad4d95cdf26e85412f6798e6145673f265b43d5805ae7b381519c70a6e6e341445801d6d526051637b738a082d79df378e981f63ab1c10e5346cfa6cccc1ebe8a2104610a6113ef9ff2c3387fbe46233d16289ad601cc979ed9cf57;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h43339c265b68a18b9a95f11671c6518a6c27124d54d2f75112f01c83b75744d8d16e36cc4bce82894615ebabcef31a65ffc2bc9eafe06312c8463ff7c75f47648eccaadbbeee363ff27d782e1585e7a4658aa01a8d143937e6bf85c85652a897fd369c6cf31f8efd0d88c1e1a9d50b6a39b72c4c858a3d8c9d38bedb24fd28ec665330dcf6879a601eecebbbc2dd126423c3f1f4ea7e5b9a9d1e16f7285b2baa4bc8b5f3075931c30c5086501a00b4437cbbd594ed3ce8b6bba43271dfc10e0e5d67aac6c8a585a14933d3a7d19b4f24b0a53e9ca62d39caff0fa3a92fec05b28bab9c8e53ef6f8892830105b25c8fabf9ceb9db985b4772d87df1e010a4b04ba17e2c8f55203e34c46bbf92340ecc7a2e0b2be3bf554801b1f582989d9c0dbcfc8bf375794146ff927793d420640abab3a41155842ac1964cfa7c6f6df1c5b8cad68903b434de894ae89859fe6ba8d81fd350b20b451abfd85548927d63a43a55b4dbf228c473c6c621cfe81c74f73e37dc619153d050604515cd8051559a02a1d70081d6084f37027b6f404d4f6b4c605242a8d406b4288c7cf2fa385c1837392ef591195eae57ac7b8d747defad42d1eb4764e84b1d5802d66561633402e9062af883dafdd855b628c4f4ee4d3e8d3b3089b8915c52d5e7afe7a907d5eefb12baafabe56368e64a815fa31b4608979410502c5fb117c4462b313f19a1e63b417255620de0369a7f335e5e6ec37384870a486883c9a2ced71e2897707cc07a296b8811418c87fedf2ba7ecb127376d0e2f491f21732c091c65ab70f2b04e54377e77b83ee63e12d3f788bef4dc4423b5f6f3a2ac8baa3421307bd0db10e2b7405713fe1f425ca5f3b6ee13fd70905231ff0a41e2195ca9e7b800e18e745fc4fddb69fa838c5720e9410a5387a2e9df86227f53e5fdc17b0feb186f21d4665d003b44777413e90dde614478e279199e6a821fcc0f3224ec742736346924635d7a89f56a8c14a93ba65c1642a615c911ef6a283186d42fea2dd2959105b8087568549f2132be1ad97a246d538875b2bc361273eee867b4908d852c658eac7b366559495e78b0a0c5d836a030579d91ff6cb292c78bc949f6527842ce4ca31427377903c89fe96a24ee2761dfebf32afb5fa2c48b8ba63e0dde3fb2818051339a17d9880b30749d703549c667dfd8e536da09149cad572230d445c8df2090057b09eb954ba229eab340059ba4b26e422336fc96a97363162c05702a807401ec2cb6baeeb5b7bc4521ecf4968ea473657915d33a734b4824df249d3a74f8722d53a2a5c608adc35184766dea6d8e734db6c65975156ae43a8ab05514fb054026e023b654555b9449b49a1aa37fcc053379f15d88adb2e36621cf4432b122d45decd28c1e60525b7daf3fce0a23a54279918d1f3f1676c181c4677d2a86d47405c786eaa29b1676609acc67f00f5e5071cb299048a1ee5e09cefd628121f0a9e29bbbb0333b95cfc796ef82b47623b70d59746c0024f9cc89eddb968a21b12e369fb8f37028da3fb8ddaafe77c9bf9c4f9d86084fec6619eef66d64ad47a028585818363f8ba96dc710911586a5679beddf4deb52a37af6e69c6fb267ccba681c728279e403b379da232c909d95034658d93617a47112b7269a0f1fd6cb438720365930ca052e09fe6ad432188b5eeab198487a212a66488a374c7f6be92feaf15ca912f89b325cf70262b400458ba743c58e86be8cc9d5748c192a8a265015a83aac4911e5364fe4655261864a56ea486b8068266d9ef5ce3a7d964b23a0f4d769f42e3e8864d6e8919ab804432da0cf2e64ced3279a9368893bc32de72bf0c1fce7a40218c358fcc98e92b07ac83feabc120629e738c2792c9c061af672b86d897cd54e2a01f2a69d4f1bbd39cea8abea59b7c9ab15474003c497697de4b5e9826617611723b97727ada1074c700c7243547a3f1627159667c2b6540e45938f871965b42afc8e1176a223618638cef05a2fb0b1953f707c67be89da35115c0c5283d8edea99092d2f2f02b6509342e03bc0c5a8daedda8bc1a231df9598d8f5eb9fc2c7aa9e97dafe248574451e8cc3fd832e5b8efc8392f89890f1cadc37fcaaa37f5cb3f406ea64ce28c20dce41138cbf7f6dc4ef848c474a00fcb7c0ade2e02ab0a7cb3c48ed92d927a05d7b3fec6c0c42925eea90399e2aae05b39bd4f5a7d42ed568d145650a86a4bf79224e5982b41af7b772018f77e2ad9d558f0b75a6205a290e1fe4f7cabedd170b33763a305812942d191be4def598f14a079fbcdd030c45ce73d864e949d8544366fa9746b166f853db8094c057029868fab44afea7f4b5315466a577004ccff950761bf0ecf09c3d39a2aa4933bddc425a8ee7f79df94e91cb6338dc942e515b9746e066d5582f925043426393c774e8bc05d7022226ce560b29093e3b4ab101487d1ffaf34114b9693bc81083970d2d37e9fa3de739ebccfbad55d5c9512c0377fa7cca5343350f7524531f4022fb534bac46e0785d0d4a688de7e25c6b002fb2d00969e728636eb9a73b97b7dd7af2d9c963580a4c0ce2a0ac4b5ed783c39ff5eebab73ac044be5edf59a658d965586b788c14b59ff61f0710f7d16ca6185ddb7f99667ec2189315e181d46712b7694d6007fbc93fa065912fc9fc7b805aa4a0c7210ae550486b2cdf1ec305080b2376a02cd02436382127754ffb27c5aa5135a2af8d58ab664763197c98d38b35bb34bd7966510afa4af77731827ee89d34ba5c7323e909bdf863425ebbe48f20d62eac9c8708a601117a5565d776edbb48e15c29005565f5a61efdab2597601198fac6813f39704c860c427660124f8b51567df6f0288d406d08aad2d79cbf505c462217cddd0c38c285a52603c585377f143b4d972e8e80afdd92fd435050afe7933f894636ac6a2c1bf172cdabb9a4a21c41d85742c2f37e2b31a08932205068d8ec55cc6b62c8ef1a2aaeda0588ca30989044057ece74539aa41d6fa006014041b442bb9387a5e0528bd1114a752699cabdaf401abf9cf7cc10517de1cd257fd28db082574bacc271cdfe67057c740b7dd7290e029dd2b1db35bd4055edee4975b8c46145bb60aff247dfed17ee8925d643d17620174e72e2f368c820256fe12080bf63dc3f0961001bece0cff5323802567c037b44796439e75b7750636ec414a1d9af2313274952b6ab0aa349f67e29961005fa605457dda202b49c79bb9ff529f77fa55fea3368cdb4361272449258017068798a750908a809e68a676866efb667f91f7e738961fbdeee5ea0e6d49043d705ade852efa79df36709fd9f9915ef490dd17d1c644dd96dd89d846df35fe5bf4e56477e7b2ec8e9b2ecf247cd8a89f23006f78afd53e9d628bec9ea6c00d702338a84d0550adb65d3778a9adc42e85a69990e5458ea85b6c8b54dcd6a60d2e1b875086388cab087ba171b466fef97beaa3e9f854e975177f2c03914039df3fb4e10d52aadfff2be4fe7bddf4f67f8f0f39bc207cecdc54a8c558e40335ad3cab105bad8677e2ff28f9dff6108b725ae2184e7f14a2cc8451ba08eb94d1ec8f79c27ba73cb1491f0d88402ee87022461bab35d0caa8b34169d3e23e943ec4942d10537323c56d3e508486c53aece7e57cd134cd0976004d6ef84f52423ebbf078b1bec11f7e75c3161f9c5ba7abcc0229fb1fc8564b54a2b72af92dba3a4d7344c78aa350fe0c42c88a3995eb2dd0f43a8ee004b559cb1fb8be85dc60a8535eb918a47504b1129ebdeafb1096e7823c443cf59629bcf192662d8e7f481854fe40ff8d42ebb7c833ff0f80b4ed11c1b29af6fc1a7b7a94872492932cf67b13906ce9c5a7676e98d3974576d60ef92df26958163adc9060363fea711933dac0ab8efdf6759e34d642c43174453e8a3620db3ccd8ff812556a88d85c604db1d20f0ee83d287720919eb4fb18388b9fc5a7331d39cc0b50c96e202d27b4b50d7967985e84305b08c069ff09034c7ec3bb362f1897c5d5f0e3e4fc00196ca3d95b4529b20dd760aae85f370f516bd22507e1c68d32d74891ac555c5dfe3eafbcdeecb91bb9ee0c5edf5999aaa70b8f2039eaf35b5a7452499c6958ea77e9f50a7cdf792f5880049ea3e6e7766e52b8ed3a83ff93ee845634500028ac8b2caa02bc0fec76b65756ba7d3616359e7baac09b949e416a723d66fa99f29bd409b9a870ede46faa0e20d1ea999f893b9af54aa6cec26cb8c55c659ddb836bf43371723e583b4a576971d69b68f96b8fbffc717e14bab263306f266b52a1d4c321165d484ad21151e65cb96b6b5c9ef32bcf427baaf8f149e7a7a69c141553b54cab362da4a468874d1fa867272fce004836891de109958832def38fbff9d867c1aedfa21e662b41ff716a07f948061bc66676223fbd61182a3e85ce9ab5b1593203a192514da3f74dc92f402629c368d1453d3451593cf8db501132357674444817ffa4e9083fe980b57696ec554cc497b516a6b01d0c329d07605e011f16e22fa797aa8711b8c458427f76f0a2f978a91be7fb7a3e705bdfd971e075e756d36a85fd967f8b9c441b708874a569464a0a754d93d8b17763ba54df54441e85873ede45571bcb0a7092407a595a2de67b424d2c3af86a98d38977ab64c9458fdc1c6de6ec94ee004786dfa6967fd2c1978e47611e27f5b151b77cf4d8da92729009fc2e359ca64cfe805a62f85d680c2de1e268d702dc48950640a4a85eac643a81bbebe9e4b8ea4f0336e24233cb3922d7138e304545ebeb142ea570bac58bfeb1aa874d860ed98242e701887e77efec7c5506b2a2191dc38acfaecd72b7a33b715760b9f6f754aae4c2eee41dde79d1fcd5d828424b051eed61efcc18f89d79b39cd359794564c9cf2d33a86e79dc4648a23851dfda478a34f37bf954cbe9c23515b1c96f47706d70384595d64ba773d413b0e47e38bab570912f8d5382493c0e8fc4d22f6508e2d4aa8a8be0f7040af70464cfd136b3c761ea3171def3dfaa4c7aa5aa4f21d93f3ef318bd12f7959c6ae2c798843e418ab91e2313b071744a2835c056a21894eb9d2fa6713f59937eb62da89bc9daee975f5d666d2648ef9b011eb5c9a001e95c16a306610a510ab0bd2bca2765307a81aa0653742267d0b34dd28aa7fb87683621b39cd71c8a7c92037eca0fc242349d01cb93ea6a13e0ee7343db6fecfb8f1162de0faa93de68ce4b0d1988cdeccc9f5e31651f91bb092393e4731ffe8895efd604fbb2b85e6795fb5a0c326056b0ace4fef845debc04125ab61a17e1d6186be938188367f3b45a6667a487de2fc040397f60a7b305e6919773cffd5e151e068afc2fe8754f61fc1315f19fe4842e724268b38dd2363a578ef7a972ad312e1e8d89ee5ab0a482c5f6bc052be46bd517dc6f77feefa0ad65c0b3dd65b9186cf16bd7b2ee9bf444e7e8c18ddc76386a1e400f43f0ac432cffcf46e29fc1097;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha0e8014957546da465b56f24ba33af637b8d4654f83aa4adb919066b92dcbb75ee91b511aace07faaecd96cc315e0bf55bbaf52dad9f14ee870eb313a8231b67fb56b899e0e472690fb15ea72b4523cadf4ffdddc8fac9bf707db072adf68b787ab11b3cb68944a167495f628f2af83366aca162b66e55cc07002a51d830cac164450fca34fc3ad4d4f35c00eafc2f100a3a61892c933bc1b16df24790f536b0f65d41750bd8e47b676e864118aff22fc2124e18878514895cd92d5876d93c5a948ed05bfa61541440746d3a633446ccc86ee351a97111cdbc77e90e5127db255dc864573347cb52dccd3f6ccb3043411dedc80fe7ed480450ece34fa65a4b13024a02f0ce0b23060fe088dfdad4e908157d3dd9abb96344101cff6e5ad81a79cc038ca0bdc9c88ac227fe61af3ba03e7b53d3cd2410b7023ddf351ce9c5a2754f08cd6b9df65b8c5dffab91023ac745d15fefada0bf4339e46929d144ae6b70ea61679b0302af3864a748aa0d2081cb663ffde6b9ba64b1d82369b6e8e74e311a8aa3de604f0ea283598f1b444fc66d2dedd9275c5781d381dad2a37d2a9e225d63ddf5df81f1226a264f0ab1625077a9094469ea3588a030d3486e9a14cda9bf7561888ced241b804940628992d3404a82fdabcc3e3f0c945bc260f8a7029aac53e5812b1dd0a22499dc1e266c17e699047ff69ed691b80df09612eb3c87434fee810ade3e5520bf1d97f7dd0a486fc1e80925bf1fea2c4e63f95b3176cb5dcf0dc71b29c06533a3332a9ae00a6387763f4681e326c786528a9245841a8a077f1fdb006f4110b23f127f89d6e006a2fb74b1ceb9879bc9b9830f240b4d72323c0797000cd5808b524a5221e260fde717a9d83367df2d96c091da03d56c58d603705687a84d7d15c83bf25cbd6caf3ba02d9303fc07dc1cb6f69cabe719fe390a1655a684796ecaaf7017ca5cf1067865edb0c300e5388405a290d3582afaa8795814f2aa6073f7e2071a9612416a62fc91606f6b6f8ed7f60ebdc35359b63751fbbc6b45cc69dc15c37ff6b5aaded79567ca68a73e0049e332618896b871ac83acf0b75fd3d2846125e34d71d904a46cfbeb80fd5577908f0dffc07aaf16c2cd42fc2a4f3335ec6c4c5a5ad647e7ae4cdae11b8558e3cf8c402c7d3a8f875cfdb21175ff1fe856336f3035a1b9a6dc99ee11d3f88d41aca629a1e3b5bb7b942d48a30e82e57fa8193a4b4b89af8a25750c0fba07102afc396a4302f29e900972faf47c6cba21eeff5cd27da466c6c5452b9aa4563f2499973be505757900c563317091996bbbd4dab0cfaf8d3a18de06df26480755210e2b8bcde1918124f151fd35017c3d280abb2fcaa2799e71b570e5c6133e10ba19974d42b0a1710c07462bdc39976eb787593429863924bbabf8e9db15ba251d6dd13c17f56c8f2276e74e39b39daf182fce396deabecd3454f04f59f4278d327751a07a26dce7268af46aa126d69ebe05497cf58c26e4ec43121680ba828a97870e7d232976d29acb32235cd2d7737e51fa47d2b3d6839301a55f36d4b032c80920c05299c966e377ccaaedfba838cc0087800be1482a9dba16e54db89548ac736b39d1781aa777656257ada1a14e9edc75aac5142ecf30b19fb944bbe86ade234fb5938d7f613036546628b5b716227fa3fd08ab3405fda9ff7e55c65fee35cd80c945a7a2647960416b74fe49225dc32297c6ca3aaf0dd740c6a566fe2f2e80d8f246f190af0df6026375224b1a63156c5813a8c55edbee14aea36aca241237d08ad3e377a817dc39c650616fcad3bacca4f9d000b4dab299020447e29a40cb9dfeabf3b941729289c59f6eb02fd2cac61004312a5ad0c1c8c660bd407afe6b1984355553c84950415c51561b4b561a97adb35681eaefe5c87c70a329e2cbd8b34b56c3c4b779d47cc5bf07e175947b8dbcacd3dd5239b8cce464ee63ff37bfb40a76abd35aa4548acad6740b07b80bbd29838f4dddf7d8a22ca979829adb2fefefee5a40bd5c8f5b254f5ab87e72da3e204f71fed5451210b952fac2e5ff2cd1a088f68182ab6dca8114d43513ee51b8b9f944813bd7869fab2365d3f1ad621c4cb1705f45abda859a950d0a247d9e67359e6edec0dac7f5092862fac980c8972138467e87032ddb8ba3a5412ed4ac84b716fc865de6f330ddc23d13e7ba2c37296fb4107775c856a0fa2caf666112b06216ba34c3f9cd2ad4e5352f49c35b05bacfdf98ddea731a4e7fedc5a1167d96838aef3a1a8cbf3011c433c44374d09b3bcdeea922fda8a5a5665fb08eab1a455343398f7cb728c603134bd13f2c8b5edd41e188585b90c4166db1714fe8107a67cdd1984815e505b8ddb8d511b26a85a12bb901a3f56a60674b5754678a2ec6773ae974f8f1ea426ca44201a1c4c9a1dbc034cb7b0a0576b41574e901741be41307935d9032eeea3eae3cd94aa714d5cb8bd99e493e5f5a61d7b5458fda4411f4c81b851514808b80f63929732f72115c68209db3007c27157e2bb5d3886133d463cbbad3f07296664adab34d041c04e3133b885fda726748a1ccc00364d9ff928dc6a1d253fdb4131b3d307d08f53336b7a715569a40f523e4fd988bbd7b0ea9c4a5a1d11211c909ed28a032e4c99f0f10bdbe45d7041931194ceddd3a112d21110f49beddada33b5fff33a74f977849fd1c66c8745d395e3b8b87f96e2e9aa5a04da7add765179b5f73c9e1f922afa781f7e856df8d8c0e863d1df574b9d0820a145bb8def40c1da47d640f125a3f38d1b5ae74eba46d32c4cb71f16bc54d6d02cff475882dd51667b793a6c5c59b8faff22218eb918b58aee02d93b0a9dc6cb4fa7414b938e8a68efa3e81c3bdb333352af02a93d3305a6aa15e7db7afbb9365b386a352a76bc5ab0896a2d04abf188b91b90119f6833dc25592a28ce43212a8fbd608e693c3c07e92c824e2e2cf940873b9ba0d32c551eb8174e55d4b7887f4d0d070c65bf9beec318c2d40fa7fb31db97e823fbf7eefc70b94cb5a0ef640f6093645d9c2950fb8041fba8df21ce199c021bb0af20fd0adc079adfbf20123c581edcf00e7a80f588ebda4afda2ee752b3325fcad2c5396c94f0a3f5a72b1330ee256db182992b3cb2802cf2d581a545d9bae6c1732b259be04fc529312f7b52f80df008fcf6dc993646db11e3847717e85513a0a87a69172be3c23663378ba1277c0f9c6bd2f6eab2a69ee281ff10736ea3a19739916267044f49b68e88da9d5ce4dc6ae84a1ad2715d2ebb65211da49a03947581ce2dc88d3c220b6bc321fd9c9bc35ebdbda9b30344bf9ca8cdd8806d24fef5d182218dcd2be4aad3c4d902b05a1c4ba2fec83c85944d278c73682fe2ae07c8fdb9bd5cf937f057062e2e621d810ef5a9e493b37c4ae1f90206fedb3ff605f4627344b3cbd482ec0ab44cb23f9acfc5f45bb382eb3ae584ea58eb809c3d7960c56c7f58146cfd4a8109c6ceeed63e1ce0702e1f6108f9f1412a41cbd12630cc409841daaf86ce740df8009cc99107e50ae62926f759f43d281e8be8b23ee3c4733630aa6127d2f1af1a8cc5739645b1356d1255aa5d246ef0195fae5b6aff5302180d5c7607d661cbfc58db671e2e69322f73362a93658aa834cff82e1b491436302e5fc1260bd0b8ed786bcbdfeccf51fda27c87209a708c85ff4dacbb080cba92cdeb3990f0296cc4ffc46fda8a63ca944b25213fbc1e120179b0639c6f0d2b561901f142d119d97c5467e3d6d4c6e146dd8a418e41c0457ad02c3b1986f8d3e1313ac0fb9f2ea34117d206a8504adc6224f11aefc581d8c8f7116695d6aecd86f4df2bbfb234821e5aabf3da0a90602248a917422d8bef18a86bcfc2dd4164bb73fb6d4889b58c97fda05662d73d76e17fb140ff14e67070173da1d8b3c3ae0eab79687de91cc6bb11130e493bcb0fbcb538e89e394f5de56e7e8d5a8bfc89d784673f43b249b484402e8edab412713d07f98bf5cae7c34ffbf4272805df750563483924ea52c1ba95c5b361727cf19f7245c31732bbb2dd9458152f8a97a524ecd25718d309f567705cb968a4fe06a5882751ca4959a9c6dd018c963cfefa1ad56429afdbae9b38a1688cc6d93c366f48b618acc1f30726c6e312b321e55cc22a23b2187795bd9094e0dd5aaac8dc8c43cafbcaeb9709386e80168b9f5b940952c8a21e16e8e7623f20345c2d3461a70184456cdae4ff7b119645944c93afba3e52a754d2ab4684409f9a34509d6bd67d75eeda4d581eb2d2395526dc8ddbeea73815c02be88c2a183c22190e46d72b6660bc870418a407fc12a809518cd8e54c4f08d5c2d6c573768c3c5be90bd9564f3606372f017ec330ffda71b8848284b39691e41ce2867f53dfb7946a1522578b75aec2bdcebd3c0d80a8d4d5acca277d3346244ef71d1ae5d8856c39d7b4fc215ca80f3ace67db5f15ec1122fae778cc6d09b03ebd222db4a69412ff54d59fc4e7775a9ab268369ee3fc88ee499325af73db6b3e8661fb1484f30f5e5a92286ce57cc77fa5bf5c697e83c59fc9b01eced3fa84caa7b6f8451e46045e7c6af5c186864ceaa9a677e5596d9a67ca4eea23c8d75ba5a7ae3132ab4a30a8bfd305ea3d6c3c23da7311dbf85f98fda8f1ad23773b36d3ee641733eb254be61687457ea6cc6237cb7321410e8065317ef820a7cf7e3533fe1c90ffbe9fcc1ded5f3cefd0fe68b5b523bb74e0f6c923107a7930a24e06cb1976d89864c66c617a58b20c47aefc384587c08527010b766ed54ad9d9a3f3a757a27956dd79a5e1a6fc4b546bd695c07c47923f427c766189235fb410116c63894b33a0940fd33daf1b7724e6877b5afce35d0b02ff39c6a3c68320780577e187b318c97cf89c493a7f41ef5c4117c4487a243f0e24584d806327432a0ac2759be4d5d2702d5943c7d02f095c200f57d2937056316475ed0a26123bfdbe9cab375698393cfc7aade5552bbafe28e207ea0798cb192feee2b1f458c9f410963a15088b1854c4f375d5439212574122354e80e1f57e2aa3c788a4fe04f6fef72f4e45526cfbfbfd4c35e9b1364faa33c7aeb8b39ac27881103d9c1f079868f39c8b4dce822e9e82f7370da5e407c78b0d14dcd161397d24333efbbfa73097828f80097a3bf12474a6d76e586838dd11e51fb3bd3729eea435cd770d173b674ffaaa9353cadb9dedef0be22d6afa8f4fae3b252aeb74aa121629d15bad7cc0baa88c85e453f155c8d150a4a6e8e2df15a66b8bc0efb4b3cc167ac4d5e81fc0ae20efdfcc9a1aa4ef7448744804e606d7b50a4ee1cddc0c49d13aee1edc502e6f1ec553d5272363f82ad79dcfe04b96966c2c1c647b5fdd3a16c7883c161d646b645c9def09270c51904ffb6d61de7263d2fb9db2d5c62f932fd3da84c700a3d4e5f0e9b305b4152f1cd6f56a3078bd53c31c66caa6a1c2820d5fad94ea68e93d0e1cf6cf7196c2561ea419;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hec49ab442c676725f9b41a32b8ee02efcd542241a8105e08b15450a0b087601e7dec80e07c153a784bc50a384a367070c05748d26209d575ea2737a7760c0b99e8efd1c5e4e24ebbc460e8a62830926f00541ac0faf05a3f93d987ef885c2f89e366d61a07d1352f0124ca72c4a7dce1bd1ea99702e597a20cd9d6d010179100bdc567d0a04c225ac54173fe1ae31b12a35712911be9694076c0cdb75477becd3197be0f6a23b2e7ec9c77bdc451bc250fef6d5f8f308c0c0cd9884575b5e92f2ede9c4433e477cc98ba0fe48a9632d344f79286fb1e71571d348586a79e27976a0271e0858fe7901298d3685629f620c059b2e81cbc8e94dc460cad10ba9dde9389ebd333450842150f0295c5853405b680ea53b4b91fbfe4f0d8678c8c2d0bcfbe95c12679c43c79617c64ace59d54cee31818cd6bf05765c0fd801bb3d47900fff5804cd02c33849987b3ea4243f2da199481e42bd8a0d8d45050c2afc03c67b2c42d65db73bc11e8dd00b9b98d00cd6c526513fd68467709fbd030da8c7d41557847268979e1eac4c6746c964318e44b30551aecd2fb6973d96c2ebc01388f745fb8a3aa136433c72abf6d861fa344b234089d3950bab652a0a764cb65d242652178808c7956b57c3106b4e4e2c85f9011a14ecd9585528f7d5c90cac7f3cd8ad4e8a310c3b86d44cb360689574ddd83f27f37fd5b7d54adeff9d4ce62c245aee986d11633b344295de210450a325d62948bc92e46b9311bb18447ecc353df15e74dfb067a45d8295875508c8e78855ef43f4afc0fe2b5c7b7463864039d0333c9c023bfbccab2fde0cf034d53473ad430a2946357647bf7c9d1c884e7cf4f8a88495f78e643f007c8fa9d0254e317a0aeb8a9832153bbbd6c9414882904d254d861b6ad1f247058d4cc64652f08a4291e3516e522468cf4a8bee2bf8976d61689f6affa54046e5c52ba47469e4b282d5f5b5b1cc01c90ff4a6a0709b513031c95a11c0cd1a05c5aa7a348ea3478dfbfbe39f104d70c04ccc852eb0db064a956a2a75eb09343e85af8608f87b0c2dce8abd720227e8079bc75db36698751102428fac34ee331459d27e415a863085321497cda5e098b04babb931be154e531b7f47c97f982df88c15371ba1b8017757e1a958a9f197276b5accb47a68ee2c76dd8b9b70034bc143a467ec86b5f48c68bc076a4c153bd5d05b451b6f95758e460c5fd407115db178b920eacf72b6afb7069c58312c4f37d63bcf489af3829f111038fa40e984d5d2fa65be7a3036d1392ef3fca143651d9b14355481dc9032da1f124cc449aadc04dc8ce77c6f7104468b315f7c84cd97df5080c8221f0fecd56c1c670338538d4a8ca6f97d7c6d72acab8107a575191febff9a82fbbdcf97d52acab8961ec00935b3e3c82f9c97968ce47622c8636946fdb34532b3268ea2ac8bc473f2da8d851b2fcbc63e1665163bc53943145e4f7cb86c17128a50b632516a2b0b9909d43560fb7afd704d95b3583f271b8241e048667e44fb12f7c59850c03a1a433d95ea6c6773be6a2d3083ecd76854b81b0e872638abde7aac0184b01f20f3d6cca3a728b8d0d3ed79e58210fe24962ce016fa62ffd77b8f046871df38ab40e10f0dcf03a566725f7b32220a8d83b23415d7bc15c4dd7b603c9acec1038ca3b74bef1bf306f6d1083e3f6f0c3d1915ce270de0392db5bccdb7c5baaecc00a68383d319bb80367dbae2985acf933332c32c6768e49348d456d99c9dd264b363c4fc59da755ff61240a640585414b9bcf76eb264b6861d436455559e460c5cb8ecd118cbd3c4fa88e2b1196f08ea409ecd1226f8b18baf5de2b432b06c209635c953773335f5e4f79c29efe70290297bd64e17eb41816bb103e8e05bc93855e788a4fd2a15cd3e78b037edfd208f33d2c63fd552b771cb17e3f8e490e7e2e9d2e29a62c07f8334c34be3d4e69e8fc6d7b7333964bcc1b0415adcca084ef403e7cba0a886ccbf7e0d9e1f6a11764e2404a4477eeaf83f9ae3dc4583c4ba112e3f52e70f57cced2545be9d7859ab5d1a185d6914c867bb8b3a6ec59734c25c0e9720bbe2c7563f8cc9cd9ecdd6baca0edb78d08cf2214d97f2eec309ab3faae7be594054ad38b3ba9413a8a58d97d09de299f4191494eb87070c06d29a6f1d596b9926012c8d4b8b62d63b4623717a9bcd8f0e2cc81ffc8355bde22057f7ddfdb8365ec632cf20716594b8d59ad96e6afcfa9bf50525f213caac1e671b9d66e08093801190831691a8cdaeeaa905f2ba59d4efeddc9d606a204c59ba463082ca822d2fb7ca4966ed276acac7d619d5490b2951a2ce6a417f268615a856680db4601a0d1c9854439afa14ba28addc22aaddfefb48d7c77c46b2d6ad7328ab1877a77ab44803314d86b2619fb467042f046a3eeca0c573f09010bcb3f67e4075de53e022e52e2acd1aad15b83c59165d1e0fee7470f1fe21c4d93c12fd99cd3b4e0b2c54248575dfb76246f232cc9d965798e22e035a694661250d13edeea63a8ab6055ff909d74421c9e3d9780311dcbd2aced8f4c7ea31bb5f9033b1df672bc800bd7d62bb897bf8a7515382999bebd16555b45c83a4161842ccfad5fff0a61066fadbe68b4c4af5ca1dfb97a585e6dfa5e1ab154a18efedf6ad02209ffdecf165fa440abc0d88dd211d93f748d64c26d286b78875fa9393c20392fd5e981c5f6cbd95f11343abf33dc5d2fe016afc347254f275e405cfcd158f8a9c0b62b1f44b6c9a34fe405dc83f6a9ffa5c0d446364ae6f71467deaf090fecc33e9b10c5721a2a24053fe45528c801d1318a68e1b4d8658ae96d587c4ca7d12fa3d0a1728bc663585494e3bc734188b886cccedd6cfa6547315885cd170f5c846287c782ea63516b70740ba0e2ea69992d1410b405d2e51bf0c587cfde5e7273d247a458990e866412d23ebfafe598a8ae42b036cdf497cafd0487db18f3933564f84f3f53f2a8fb09e53ba7a4ee4944d0d9e3c850a55fa8dc0d730a1a809bc0cb32a07ef914cfce5ea0649e185dee2345322012105780f01b82ce185c388467b8162689ad75f47fc7b991d6fe64efd1df1f441d3ba50dafa6bf1611f5dd91ecfb9fc3ea78f65ee496960aacd9c611f4ebcb6e93f55bd7ddff8e3655bd22a422daf5def648a0fbc226be6c7b6f58a25ed517c4dc14e4f4bb55553593c23c4998c7cc41f5558b2ec034eae2ece11d92a4a23e3ecb43d71c9b04bef46f61344aa9a553a73eef721a1e4f2fc9796cf595e9fe5978e064c052afad222acdaf53d86fa08d62a0040465205640a2376f9321253539e7697f223df3f388bfd440819a9b44114979eb81ef5b334d0a9512d95fec567313dd4f83350a10f4b3d75add9387beb5b0ac60f3d35ebaae6d991fb2ee0fc7c6ae2cd01aa5fe77103b8889c88f516ac917f8a499fe52140f038dd3c7923bb2d37bd69c90c88c168cfba6a866108f017f7021d2885598580c0438a0d1451fb50aeeb0679eb460132dbbba3532c06984793d7281e4491017db22ec1227938d458e277f09085e02969804ced605c9f29574bd61cb30783dda1ebe64b704aa02dacf9a2daf2b945bc22ea70217903ced367e6257c9aa35bdf9b6ad9270972e1f5cbdfa9a95d9842de301bd3d15c4dd5cadb6e7173f0a3f6712102569d3432f2b271e34aed073ffeb069a19efbea8304e9d8eb293c840754c8c8ab1c4d8886d3d14bbd20ef89427a0dbe80bb268ba3263ed0efdb4509c71aea0a5fedbb1a041846f3d7f371b059335b46b3ce4cd6ba9505f5837f218cac28427979a99d2170638d28a72c4b0830d66849a46213cb0e0b3314f4f5032cbebbcdef52a01671454730dc6bfa95a4e4a0149d9fdc84d7361ff175bdd3df312b73ac5ded2267c09a81e5563bca1d04a7d20626fa08ffa718104834e96d0a303ebb2dcb48824868c6fc0920e62e8e0b28883ae1398914c135380f7429f3721570fca8f0dfe2685bc186badcb283bf24d6a429f2ae5866ddc539498aba4ab6abbbc2cedfcf3ff7da060a9f459923f22afb649a457e17ca00555dcdbed1461056a114bb8e243b28c0911789b216cc1ef6effbf7347482acc7ec78d6765f0c05a700c46c24061f674023374d034a85fa40a809b352e9c3695f3e61d8476f489bbb30fe86a884ceb3a75c93174040767e8bd721d7cf7400fa44544b694f2cdae7677302d04a925efeb72afb691d5753ac1710bb2aa2a1ebc5389ae620367ac5126963865210755500fb4071ebc3041ff701db0fc06e3de4ce8167a55f1b05bc387811ebd59a35b3fa82551e295289ccdcf3764656a9388875034f10860f457e140848dab1a60ad767681c17b0f7e8f8751fa256b0e8d28d492355b543faf13af7d6d99ecfdf23e6c9c9a1d5b15c6ba250e4731e3c514fa0ae6a22045147084a05fe6bd486934ef6a8d7232521672dba8c1dc0d6362043d096893c212001a1e31754d6d8bf4fd2499b9b7be6c5fbcc3a07c31e8d47eab00b5dce62511efc59071556bd67302b4b81985cd76d6db7d686186f6c061631a84af1223845a28775795640bd2f398e7d858947c07d7e1b47f2f42aa89cf093b3cf8b68e92a7e1f6831ade06b6785462db721fbf2c9760d936aa4b4cc1871f756d233da77b0eee0bf4679200aaf6550da7bc562533c5600b436e204e88e1d9592ef0de16a8c9c9c73fa9c4a7c89cff9703c81d1e298b70bc2e472b5349e681be28a796fe0940a749bb1ced603102bd59250a9ac113db3069c6f6f8d4a414fad5f72be9b6aa91b09a6bf3be3a12c74a6c9f9d853345535c9c62879b03d843aa446dcc5ea3cad520935400dec378c0ca3e8b75c9bf88c4a516d9527b5f74e3ab19443967b1db12d85d378b7e0a11c1b9b688dc1f674cf5fe1e107adc1950864c5ac3d345762c16e301c555ba936564a5f8d2428441770c5ace3a77dbc1f1956a656841fe4fea2e6cf00de7eeccc4849839a5c136607df0153c91d3752b7619077bce7cf1451038b0dccd9d7b38568096f5f4e934adaa844353f7880a7fc46b5033445a5716d9d591c59a2f1ffd8ee2055a08d4e5e03b445e9fabc5bcdce9a169ef6ec3a9d36b6c1eecdd34585a88263ec32afe7cd2bbb7425656400824d51f0449da00520069c4765e2b29aa62eab2fa82132a578c5f902853f715d960369feae1a58d620ab447b227f68ff5c8e7a5cb31557f9864f213ec077c6e93563c35364013b00a972a1e3f3d824d5dfbe974feb2054bc2a4525b466a8fcf74ae0be166f6e4531ee7f70b6c026ed9259714885b3b672e1a57c84156abddbbdb019ff09d1adb141255e8ce14acf22b969855e8904385432b7d19cabefdb3c5cadd8e87866ece79d5ccbf1057acbb51de2413a8a130835bdddb60b585318b7dc0b2b0cdf521ef4f876291deaa3caaed92f58b75c1c49a7794449cdbf3d2785c8e5845ec378f20b777c73a8fd40a00ba54d3ba9e9e86cf9ada5bb3503e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf2a98e80506b64b427bad51b5f5dea5fdb839d8cc860055805d79f2020f200495c3133e8614853cc0ad3ca33d4dbd2f3f5dd58dc3fab7a50b54e71783e65273d0deeea43a177210251bebcf6264b61fe33d471d68be74c1deb9a827112eaf8c62eb924ffdaa94114aceb462a4c6228c95ea44848bd92710653e132602bbf5f183034bd495991d491761bd0325db20428764a352458c4a595a4a593f131255238fe3f5781e2e5f7f0572f6948201d85195a5f70ffabcdcf145968009bc69fed7b5d5ac4ddcb84a4404e4e6e36edde722151b7d642012751e42cc4b972dc616082de85803dfadc95bfe8ebc15bb6a2f53e5c77cd83792205a7cd8c03359fe5bce2518c1f73444be71dd6373fd4dde285f932b2810a81e458887c5f238f7cf203e32f5bfc7d321c80315b5d7d2b2f42a4b6fb4fef1dccb48de4282bee1607f47353568b89a7b9ed465911eba8fd2d49653b0036b029533ced77f5c06003ecd0a7b1d67b46f3072b990219c15327a595515e263a2bcfccd920c580100e06f98e5f4966bc6ecd730a6234cb397a4fd67afaf35759fd91b9572f1a6e5e457b12905543e0e8bbb01c0705f2b992d409a565c8b07b19a3347420d6452dc850298ef5786ef86f4b802d9932387935829747794277e91eff342a5a1d747c3300bd5ec760dec40236114e1e80097ac096368d2ca8f26ee79bb76bc8290ff8c7cda90f9a93b9f81d98762d758e6f76c042089ce0a45c26938eff908c7816fd818c8d991e938229ee2deed716b05343ebc0c2efc9ad785e09cda2ed9c0b8aab5759d9f79e5af3b1b2c6c69e0d961862d7c052444a2151bacf322da5f7e33f9968404b02b2cedc77d9a217e575e76cab7cc5260b5c524f8d998e3a5e1405bccd3695471a12f466b369a135ccd79f9cd2b34706591f3a1ad8770203d54a1dc51d7fcdfdcf47d6fcd86f903b6e3498deb24dfda0d6ca380b3d3b7fb3ffd2be251ed113e333309b4fca6ba18a6b0e6a4d9a971dd4612d133343f65a67ed20bc24cc69ff5aa8ce2402920b0ec26b32cd61a6f2754232dd235e58f2381bebd369ca07b984caca7d297a6907b93a0283239064859c48ffeb2bfed6f2109f9cdd4735fa5a8c6535656a2d29391b0fa7b705b3e97b77d28e91ae6647e4dff84c7038941043b46b01832972bd3c78bb38979de9c37f3dc96fd3ba66a2ff7e455233a1a8a0a4dcdd0fab4738d3c76312269ff0a20d2fbf5987a107a58fd95e60fc91c462ee2be31c55b8f561ca7d9ce4827ed10a7dc370f79a7d93b5f9935c5a5a717244400c80924d08dbb6fc15ffc80d1ba3e9d739e8e120007f7fcc471cf9d1391733302c1d7072de3f0bee6025c28d9eb54ceefe3a04220f3bac7941a154caec0fa044de7092c2758ee7f6b8538a49a223312719268327dc326aed12069ba0505a860cc0ae1894f4f9f1185b5527dbc405e468e1bc8e4b2ec54aa3819ab3e2b1e189debbac922f19ff2e80a8c7989d21ea2bca6356b6d449557b90e20099cd6fa19af102e5a44b0c0293c75f2c878d3227eb1a7e5cfdae343aabef09a96d9bd3a5037ff07576c04a91c8d3ea84a6ae57ad1ca7ba1e2522ef58aebaf03957a830ea668aae86e3ac6450d782f65bc0765d869ba5dd130841dd56169f8e8fe72ccab81911d68f0e3fe824bfa6681e6f8d3b00d6ec3fd0ad929481838797711afb17c5c8b726cb4257efba2084c49ad1e07cf6e29ddef72d08aa087861b8ace59454f756cbf7547bfabe6fb83e1a119a4bdbc5f0998ae292ad66c1c72f86d9b7f6a27317660c17af77fb0f0566a6a7c0bb757b2e42527fa8af9953887654b0a5631b4904ae5ba30d4f2834a971476e104df1f40e7d454aad065bb1316c60a2d96ef84ea6c954e80a28ed97ebf1a9721ecb5442c4a6fe12e4889f9983070ab67f3bd3af73485df4478f05c5883a261dbcd269c8ed89f867017940131940b50085a353a107d0f8d05e758e931436ea4f060e8ea041b356777639545e7a09df331770b8f78353f9879fa019786dfec22a50986f5d4d091ec37289fe4323d944ba44010a7e2f3017cc403e0977686f5bb79b12aadffd8b8a778112793db42bb15160dfc9b708e97cfca317576fdfc011c746692b4ca5032f5d0b7e1e42952aab2927a8021d26fc086fd6703ef10730a090f5675a54ccade6d664b3e66adbdd50e85e166037b3651110065e639df1a4ad07bc9d6f0b66c03f2d8553e48da750c6159360a524bb2e4f10b91e68c13bbcd514e1173a957cd67589af68e4a9c4fe36d29f1751125a60af8d26d629fedd185ad697de8a2f6db06f27762a571eff1a1284bc5cb3f371b9b66fa28e4849522b72764cf29a4506d023d22c101b867c72699a7c913d8b51aee1afb9872c2ea0f3f099e2cfe87b399b794fcfdbe6f2aeb86cece90a4eadd51ded5d0fca0c92eb7cac2b1c3725d3553b58ffabecdfba869205dd3d470eb00aff6b4ab786ec22e3d51cd18bfd3275946392f67ee94137304b0e2a82488560d83df11151d1a3f6f90184babaa9a79954ca8ad28ec420ecd07600c0500c19cc02e8c9760cc8eb0ed2524532cc433ea443b3557b72ccd861df9fd9d0963050683b7b4c0b4fffe08464ec8b99538d97e5c64935a87530e70011367d9df354bd905489cfb49dc12437e5f2886368541d04e2f0ed5aff32f33295e8226fdd2867383b61d1958365ecab84743a910f7a960b7509a24470832fd182abb6c46ac01d1d7c3c38ae4135c6c7c645bf40e45712ce0e7f451ddd98088608c52e71533971d95b207b895798421ef46a083d60fb6a7d1f00cb060dc01bd2c695a8fe7dca96d36d030e1ce78a996c1ed2fad3d54a45b360de77ff694e75b355773e72840c86d4af9ec61a386b69f33d320296c2c6b7b758d011129e2e39074abea8669af2ce94d2dda4e5a88acc32b4f557232bfe06ea861f9623b9fae04d7f8821a005a10cbfdc16158c0e60fcda2561d16554d87e22dc1b531d487b3a605ad43338a6cec3597fe67a7a169cd0f98f23cf4d866cc0957b11d5bb6726ec50d908c91efb71ed8e71c81bc44d3f4fabcfd6fad3968b6c736a52174ca3a62487f55930257c6778d6e8f9f96f1a35d79dafba9155ffc931c94424e6bc7ce11d41db92b87b077d9df4e52f4d4672f2be69e785a9b02f0529ef63be63c297a5404718c2caa1c6cde516a0a4e9d7d89dbd7cb15ba326fcdcbe145c02a727afc4c1ddc0599a86ebc004b8c26a1b2214257fcd9245b7a4ed822ecc09ee220ee1b6fa9da42cd15ef5de66f4f9724d77ba0342128abd3c4f3dce49abfe04996bfa540a9cc63dc158187bce7265a93a2560310b9a0978486ff2cd38ae3dcc1fe5a505bb79350bc0ad56478f5caacde6ed9bdb61d898040737fd4815b358ab441b3f91ed9ae42efadbb5faa3c1490f18f199168eb55dfd2f76e6b0d0d0f0c1953d40c1692450704e62152ace7b8c7eeb578ca451bfdd245a4f9cfd3af7b9ed895cfc178d29b9f0ee6f9725f45fec616ea6e5d74b58408907f4722e7bd2c4d30a77f0467a4e2fddb4b264ea55def3f5cdcd46e8ec868c748fc4dcd8ab1bde9f32132246c00e1fe6416d435f16e057edd8f248a1110febed70eff9c754fbc26e112284229f5715bf598dc4a33ff1d2106b1b6867759b56a8e65f7ac5d7efe31bcd5280fccaf37b8da389dd2d254ac1dafa722f5e809b2a8702628c1bd03ed629a8010826edeb8627deb35ae6b2ed5b8d95efc8bd6edc95ad84772399b7b8e9dc7464e9b19ef8964487d3ce11e642b5fb89899e68f6d5f5cf1031d8130daa67e830a535a6fdfc46886b90797debdf7c3ef17d0d589ab327b1bf36a9d5efab7e21c548dee1f049cf929a77827b8d12d65cf65667cf913b94ef000cd645c9111743a1fa8e93b469b96ffbe6e5507b490d7e7308664652bd8e14df74a57a554e771a04fcda0d430d69d8289558935e10157c65aaf1c432ad308123b09bfa0a030a4e050a4c9e0435f41e7968d633408aa81cc325c9c6e9715c31e360572b2db689f77321607becc58f3422af2fedcdde82fcfe319233a57963ffef5a772fc6fa7738b310d33d40d28a89e9ad753f61e66533209f7f367da157780a39f4e896f65d24a7af56a82d2bdde83ceaefcc162f10bb6a674b0e3b2471f1162111dd7494e728567b75ecff24d92d9932db15c700fd3bb9195cdc987b17b51509887051ac2c9340a2e359ed909ac0e4133af49ce7d399322a26ba4efbbdf0846596fcf2a584eda29ae3bde6d20a545cd73cc85398e3f29346d640e8d42911917771c090de1c28c18f3ca388c465f46cc74831a2e44c87cab69d9e30639fa09b6f89aaf003076520ac25295477fc51e86e7a98a8bdd6f48cc9d1bd7d99386f8558993d84864d42133b8edcf98485b72dd08274a9db0aec625f678883fcbabdbceba8a881cbb03da6ded67528f1b744ca1d32813c95e32913d80a836c24277f656bba83c2b9206f7b466ad56862f1d518a3de1a136e4e633a7eac48b23a77f68efd881a6624675791d80e84840829d0cb91fb3faacee7b25a7eaf41924630f0c4869a4831404a32e0f2750e058adde738cc92bdd4356e84aef8babc2f8f9b20a39105acd28cdad022f690233777cf53b4e5c6d7a2929b1c0b99dbd9e98e56d82820412a15051151ef0917fdcf69337a321af24f3aad81839e18ab70b412b471e3db0a24ee68179afbf44012700d59d9127d940b055699fd1f23d7c69e872052d4b5afa678bc5bea77494ec3f4ae61ddf6ad478ee6dfef7f11df918818e6c1aabfd0b7c807700755ae9450b711217b16a881a0e43b8b27ae9aa513f43c5a54bc4ecb0cd11425d71b7aa099fa0b666ad1de5d7caad83e942287bba9034c56371f10c8cb3524a7da57251fca01e7d9a87ecfe80292f684bcb8d846d8d94a1fc9a38f0ae8658da33f987120c8314e510095c4a8c51c36edee605a9e2c90227beb1d544d62519229edbb560949f5fe2cb7a753928851506739f69d30eed3af60097ac5ffc634c9c2604a15f0c56d2381503079c5d9caa6c4f8c9f39630f6fd521e6f71143d5cefcaee77c566e614f72e92db9d044da90224a51654fd484c99c19cdc464507327e6e87b59d0dcdbebcb825a8dfd5f5b16933b243befac6ce26e57a0ee79f403cce529de1e7b1b87d37ecca508f9f89c9f8f607022487bb98569c7128223b31c78e7018ac1d384edf57739e5905b39a669db537c438f912d3a9ce830c4d56bd159b614cb20906a45c17907677710131c534ca451b635bd29641b27f03abdc7406d456c05b991d5f19f8a06b6db43a504418b73ce3b397c47b33cc746a9bf733497b584a29ee526f7bdbecb01df84bcdff91a8d1ca8f34ef8c386d35289a430216cb034e49ec8964bf15ff56357b5ce4a43b50f19205fd2caafe52c7dd7a7787a060971c75bad563d53e6d9af1230cef49f658285a8b5f3cee9ce6bff9dc1d02f9a11d9136fb5e1bb1a60631;
        #1
        $finish();
    end
endmodule
