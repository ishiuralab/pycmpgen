module testbench();
    reg [8:0] src0;
    reg [8:0] src1;
    reg [8:0] src2;
    reg [8:0] src3;
    reg [8:0] src4;
    reg [8:0] src5;
    reg [8:0] src6;
    reg [8:0] src7;
    reg [8:0] src8;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [12:0] srcsum;
    wire [12:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h118641e5ea7e8d353bb57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d079000c1331e925d52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd5bf086eec713a2dac0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d951774ce02f13af4db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa2241edfde77fcb98c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fddc9c02472cd25f4b85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1051a29886aebdf084209;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h393de70335904b7ab1ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hadd3d3b98d003f031eb2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10eb47b07fd6f4672b563;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6afea1a3dc675fa7e8f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87ea8cefe7db7bd9b79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22f7abdad99b9695d3db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h56ec37869338b6a91b4f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112ef25441530472c2456;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13fbef77028f85c15058f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6375ee7d1c3924a0a44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f63193c1840a4e44b03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f57af68cbea08e293b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9dba25dc79c7a8a8ea5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5bf4e279073037c7dcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6f18176228457b7ed3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be4d774cb39ac83b9e87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7cfa7176ae05095f2bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h66f2b93e057694987c53;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc3cac8d48ddc7d79576;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b3c5301e8aa51ed7543;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18a43721ee7c453fe297a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h61254e8abd14e9a99db6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185bd9dbbc950dd4cee7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec7b9813153af5ccdb3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d787000d8c2ebbbd5d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ada1eaffe78439d1aed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10812050afbc49b702458;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee2db9a366fa4bac4c3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d99cfc6e86a3b5d604dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f9bea23d57519499d1df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16155b22bdcbe34041a28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ead5be6dba14eea1b9c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfbc3e30b8d5b2291b31b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1186eb298d6cec69bc95f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h935ba2645fffecffc47a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h153f5b7cdea6cbf118196;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h366077a9c31ae9ec1243;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1332994f83bfe09d32b95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1169afb1a8590062f8710;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1beb89e3fa7c283110765;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0d34152bde9e87d0fd3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123c6e5bed9369ba45b03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d6dbbbea4f603627df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h121aee6cb3768c291119f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55bd9a8a65fdfecfed05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e320a51cf6c5822e9bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7eb3a23866bac4da489;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h703a3ba327b1744c98d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1e2d56ea4e8080cef56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb7c5a43bf788d80e32e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1058af4293e83cf8b2b17;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe674199868487958b5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1991d8f6cbb106d65d5c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb35f70c3f5710a322c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d013b172dc6c2ed2f63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdfaa81f505dcae2b3a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5dcb54e74460aea29c40;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7ef82fc0f9edc1883c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f4d24e917938d27995a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf2ca905e41f75fd7f5d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h226877f03b2b235358d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13978fbf8dc8e8c08ac2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96d26b6bdb2d6556c615;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h507fee785099c7a89a3e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h110b1cf6c7fbb129ee983;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha9c9609d0a703f3182dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ba2f80fe5ef0d67c31b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3a0a9d73a740550dd2d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b056a0a012b4be02e0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e6ebcda6278f18054e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49a70d5b5999146c4e9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d286846757a8f720be3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52d9b39a8d8513b62272;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a5b98d8916d41d1e1f62;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e483e78c69ef2963df3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd9dee02997fa1f9c6c2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1435a141cfe238b04316a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126af67eb882e10d29823;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ab9e6d9d98fa2b15e768;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b1f93827f748e28da07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hedef14aba0d2ac4c3a9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h40b30ab56f604d36d176;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he00470abb379c408862;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179caf797c7e1ff73532c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ba48f05292963e38381;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd1163114f29c3a7c0180;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8ba42c0c23aa41c6ced;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19bfafeb88243e8cdcb9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb0e9a6ecd18f8f0a7d2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14db7b35cb2f3ee3bba00;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1504f3cd47f3fd733645f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a26a99029c292966a4b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197646cea2e6bfc37b772;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c9273fb0ab91980995e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c86a0f70df83bc803d0b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb875d0da5bab156d697b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6ea4bb4086e8e8c76f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f51d6128c92b8eabe6ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1922f80063866785d4845;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h195396f0c6791b876acc6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc962c637c8a3a5f51748;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0f3f4f6e1a6c0c186e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15452d27d278200fd01d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed3cbcd3b0a8f01677a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h63b6f5528d09ffd56cfc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17714442c86f304d2c900;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h174cdb4ed7324c96c6f75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114cf3d493d8e05405670;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8bd30a754185f421941b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e0f0b5d6c962ade22bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd1a4d518784a58c1cf7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a3cf266efbf8883c959;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14af49c193624dd8cb1ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h236b3eda326b4ffeb79c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ffd67e6dda761cd83b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f76843d92cbca707eba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h184c63d6a0837a9ce4d5f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14989f352b90f3c1cf29b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cfeac6256643c48c26dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5bda22e1950037043d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'head6aab2723420150ba1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119cbb4469d3d8f199a22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff5a32533fd1d06bf84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12087e606038392906348;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d5cee4aec602951c10f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49cb167e1cacf1c19726;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd13897c8b6514372f593;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1d2ffb5c0d40b616e44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107413bd607e2083f8659;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc771adf62df4d1442344;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39306d00ffeb64a265c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cad8baaafaf75d086ea5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c075f0d49b09dab794;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6b86893bf687b55b1f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d501765ead3cdfc1d03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h468a52f0a81f3619dc93;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115a2e056a660fa91783b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c2f256a8855695ab021;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19638d0de5bd12d9f992f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18a65b33773ec32d20da4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58a746320bacc0bb300e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5297a84783d0169ec27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9bd6738e9ce5501d2742;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ac757a3ef1216254072;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2944b41972d8ba3826f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4f8cd663731531363da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h30259c7294fa3761f5b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad9a6a639a09bbe1a8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf845fa2fbc876950cb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b2b9189528b918c2dc41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb474d205813314c6b64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e386ae602da7519a95e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h74e9db70402988c1004b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d3a9097c629ebf17b0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa19d51998f92bf99bfa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120d772d29a669c1e9bd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17097e59f5a5cdcd56e1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e14c3fdb902ceeedbea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44d84c435cc2ab1ada99;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf9431dca7a51827c15ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1c705dd91fef6b17b47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1f17f9380397701f7f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h670d1ebb54d72086fbdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf791b42965c4d8b768e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcaaf08d31984e9a508b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89249fd7ac9ef6652cee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2bbe65efcdcee9a87ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196caa3dbf12bf9ef5d02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197a6b3cde8900552055b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha08694b22a16458b8e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dc1b7e3efe56f8ba581e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f1d595e52eed54bfdc7b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2446ec974c5f3f11275;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15aef3f8ca33d114d3dbb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6123580e137479a5566;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c6dad2e0ed0d9222ad8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d3611c8c3a5642f01c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5616f6aabd4a1ffd51a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14fa00408ea3f093b51e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1953a66737e0b27fc6ab2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93e659a0d506b3096a22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h27d261a13406249003c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139ce43ba49c17d247e94;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c74352e2db292211c9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a685fe41200e301cf72b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17422cfc791e625f862c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104062ba45d4a8e14f2be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d4dde3a398ffbdab331;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12396b0fa54d607bdd7c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5dd534e4b697f7b83d35;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he4458ab7d4168ab57344;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f9c2a341008f794618c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1716515a46a2958e2b613;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc97c1ee9971dca50ee31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12dbbbfcda268e16efb70;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62f7363ac219e57e348c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe254d3b22f8a07a4a14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4b30dfa0b78bc2439e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ab59ad92b1008fa4a7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23b93a82853ef63d969e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h503d0b7009888279a5e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h133f6b02090449b101e83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba46ed45d98ba91ae0a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156dc338e97138ab7c323;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69e8a33e8821e24132fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1abb10d1c40c95bc5ba9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3e22eaa0b586ca61c4d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90fb516ccd5fce483945;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b1bb7eddbdbd5f148d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h101dc65291608e3807829;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183730251daafd62e865a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2fe23b78801d2f26320;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd1bdcf2f50e79236ed1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17688bac05529ff49bf59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h161573bf18bfcacf18e25;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h568cf367e5f8ccc7aace;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3eae6b5f01cd0d0c353;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h134e69810efcb5c6370d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c4a49e14c60c2c8ecc7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6ec73b28cbbaa686fbe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cbf5d897543c1f700413;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7d67453460f42ffabf4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1784758bf5bf6e17d6df3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198207c309416e10d48e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd76cae20774c179a74ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12cb5f5a3e20f9ff11625;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4457757c8e4e7c6af92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c07bf868766aaa7640a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185dcd248da648ec3d8d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11880513893213da6fd04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ec2c8c907dc7934a439;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h155741a1123af64fffb5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1458402ea69c98edb15d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105c065277a042825f5d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6febf6d55fd3cbdb0d52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34f96d462f8acde82086;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d7fd4ff3c85512a7612a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68b36b0cb46dfa2ddcc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cca79a2a6788eb5fdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8cf7eceba17e9bdf3b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb94ab7e9779fdf4e4ef2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a2ab96a9bec658e29b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14870a1cffdea750aeabc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb48c9dede138b692af3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18250a30bc13b88e21bf1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d39fee2e15b78872d078;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c488bc7155db204a8f29;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6a2fe6f97f9deef97a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14f1a41e5841e9dc11d89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103855d74075450f5be3c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa0e0c3ac95445584ff0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a87b411a865ffe77400;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9fc04328e9ab499f648c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d3159fea32770b609a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f7cb1f2a2928f9de99c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h166256023d49f47368b54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h307877b0f5028a56007f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc8a4ca1af38d7de5c0ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138e988dc1298758ca968;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19edd125cf35757d9d183;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5554dc239886b66cb802;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bae20667c810c76cb69f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea48a4e7fee35348d9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b2bed983e74c8dcbe928;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f039fa3f0f567112727;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ce901966d626ab34490;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe9fb78acecc953c5d4b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f2555a55b4af3d8f37c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a8ae83f812ee61ed72f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1223cea86010ebb051528;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d60ee292c1269f24c942;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3a240bfb6c3a536d25e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8170299f948910b79e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188cb2eb73d259823f4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ad55216512e6666d95a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cfb7b0306311d778f0d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e41ae8f7d2aaf0a92e39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0a77185f6de775200e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186475cefa214f94fc57a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd46c862622b698ddba2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h794d6c8b94ba00c17aae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he44cd4c61c3d058d1b44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3c1f30925d83673deb8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h678fe9135d291e97c409;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1213fd65e30aee8710e9b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h982f0d92b7dbfd8e7dcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116fb680e01ec5cbb907a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb7563a02d293bc26e727;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dac73b8c4155b8cacf51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h172784e5689e109d19d91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb6a98834b83b8e3d1d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b85dee65787c9d3743a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9143caed33c55b8703;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc8950bf69d5ed56109c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h929736b83ea795bd10ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc959f4a80eed0e1c28e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19de7b657753736abfb27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d29d773cd6393fd38de4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1095b5836f7d6ce3bc52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d5847ec1101fbe01012;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18a54e6daaa1d57ec71a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23d4803e5d9bcabc1ac5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c81ad16bf51c6562322;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aec9ff9ca04248fbc76a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dea014066ddf1078d80d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84b8b65ab590b025d48e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc64b170dcfbad6d92bd5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9f7eeabf180835fafc3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5454a2bed679ca5bc52c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b215d38a9a3474683d09;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e84d9bd4fa20d6350641;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1402c220616e94fa3aef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd9a1edcd18cb0bd040d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h347ca29165a62e6e1b4f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h560cd4f1aceab99ff6e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1783b7b0c8950df381577;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e3fcfa1d249e4f01790c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h961ac6dfa453eae90a0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24c1970e916175c185a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19db8ab8e5284ca7e71a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef635eba76c12b9f26c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0d7777f4a07b0be1927;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9bc94e198cbfc260c5c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160201e4f60dd2c053455;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde2ab282674399c7d1b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdde3c2880868536810f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38bcdcc9b1a34a395a14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f584592d09ee59afea1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c527523a02953adf14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h880cdac8be829ba77a22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe8b73dad30e4c9bc711;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd95e1ef576a3571ba6c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c3c587422f4223aef1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h65fed495e58b382848e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18dcbed3454da779c92a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec8eed36299b3842b9de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2385bb5ea72f4f9becbc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57f0b1f1b065812de8dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9058888c4ee6df87365c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ffee7639cd7884e06db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b727460f84204858ed84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1723c01cf258c8afa232b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f55c3940b214949a2ba0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19cba40142fda2dafd446;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h171dc5310a910c06168a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af3d307579d45e5f9193;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105f536d3d5f98c626702;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18bd71f19468f55cb991a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8eeff7fee29fe7d0e1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8a0d0636648f1db67f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h80dbbda3366687bd03d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11fd9e139bc75a3e8703c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h910ec4dab31332e0ce69;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cabbbb34665e60a9bfb7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e9f061b9e48b7f6ef92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119dc79504617b6efc2ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha738359558d452a51e5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce1d9870abcf40c85cee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ec74d29d2082c838d47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6fe05486eedb39e1b760;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e67e3dd3df1e2c21101;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143dad222321403c38eeb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c463e3443a316bb2c483;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34c0e17a111e7cd3653b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2af54d60e2ac6a6d2146;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140a2f8accd1dfd73f7b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93909aac3e7f58d6c365;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7509f8a0851f78e8a41a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4613fd9d1dc42aeb9cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3d930f5f25338f7c216;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2c2c6717fb43416edf2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h43cb96438291dfa82d1e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69dc270f1dbafe48a4ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3cbc043e58d953f8f90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e9de0f0e96ea2aa4d30;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4ae5ac7e21b81f73686;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b38d3ac038d40bf9dc44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44ce9c52d0a880b11fdf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7191c55de45a39cf3864;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187a60c5307d937a2bd6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ead2330ea26db415d3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h765b338d6f9fdf7cb38c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc542da6a481d9b5a4356;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb9cb20831f5b2ee5b11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b465bb37892a87e4782;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16eb9713308150be94d38;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf745e737c5fdaa4aad0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53a3d51e19b8028af0a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5bf6fe2732a1c8631593;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea0cc800c499aec5eb5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8386a9d6ab36fa13cd71;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15bea2506ffb1eb3e72b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec29dc845758acf69af6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e74077a3bf3f0cea6e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4a3a1213e05def91e0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd948d70442223575adc3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc543792c78fdee61dde2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90ea7a39615022c5cb55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8ebd7f620a4ede38dc6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7381510f299330bbffb2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18728779df763c0ffbf7a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d9638259f8ec54f3d37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1557948a9b9de94e45b47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11945b443a75cef8d4a6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bad83e9ebbfb5ec0456a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e709ae0ad13a3c560d0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125accf314ffe14511c36;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1948ca45766573c05b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8494c0be89a5b717da9d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13467b6abfb72d27780c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1683cb80ae111f5e4ab70;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae01a86ceaf618e0e374;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12350a99f0f8ff5f57593;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d7672765a869785e1e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c4d1c703ee92dba2eca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafb44679d9b29fcde148;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8d149ad38e069953d14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdfd1f41cf8c9c4b6fc6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e54a869ca48a0fc2462;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120d0101003dce67825f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c6eb1a0da2a05e69834;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52454174f6538c7748f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ad60407e229979c2709;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd870dd7e049f5a6707ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e68d52ee0dfec06faf70;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca000b5bb61a102aadd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2e05ba120bf37a24a45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c656ef8725dd06d468c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f17218af0c9b4a697acf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16be430dd01c9d01b3945;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15217d9908a0eef9c489;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8436cb15b00f29a7696;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f47730b3a35b3f2d4084;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12913e4ff6b0eee2df949;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8faa285a255ea647f21d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2fb5396e86eeedb3142f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a83940d25982a0aaa40;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57a3f9500ce5440e3212;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa297c54f8e5c0844ca9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c52663d939c696a0e3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e9d326e7b9ec0249b60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152073f4d3894a9d1a061;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3cb346a1f98fd591ddc3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb670f6a53e13c654caf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c20890d723a76e49220a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ff88d62587f7dc43000;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84a666d7b0a33dce96f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17deec712f299def51606;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b5efacaa85f5fdcc9b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc78efe78666c65088eef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f23db24208263a74715d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h553a68a598a7996de82b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aadcded708f8e21e2c5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116ccf98a04cbdb9c8de9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he12060922e16cfea8702;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h359949153b8cfbd747c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3397ef19405adf632fe0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178a91450df123763af5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb99e852015f9f92e2b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1277e77a3c300e0867bc9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he5090e302adea146d0a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he12347ae6ade91256936;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd903650858e8f118549;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h61e2df451ce5def6d0a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ef87c8eb8d9cc1a3c4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17eb492f9628e9d926256;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd25ed83812b3fd85a51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf26602e19e83c7f3d424;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e51c6873bffdbddc2d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5cf743b207790d9d18e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb51be17b204edbfd572a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd1173a11a9a02ebc9ff7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1918c05fdadd13809e0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf9ecf17c6fb3048f6ee6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6ae0d310d7ad230bfae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h413b5ceb12f5aa821982;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d010de785ac6f632e45c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b5cf4e54043984c50c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4815f9f621dbb7b6b07e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h985917a532c65f4d7b64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1982d6ce80c2ed9d11008;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf61882e52ee4d4d1e635;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7501c1bf3dea34c74dc4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a96568c0702829bfe88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd2d137b6e5c353643227;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a82f392e58d45dd2a1f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h194e493caccbbe4b6c9a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76a9b657ca4280066866;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159fb0280b4ea702dd124;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20c6f4e062dc3ca6acb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7648e00a64569bd8542;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f21a75598cc180c8d1d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5a05dad1a2d04776450;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbce29f07be2711c6784c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19358164ff6f207ef4b03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19af81d8edd4b8ab72d63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d89f0c3bb9d426e1a31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb8a6a172c094584036bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbb702739faa70da400a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18664766571c478758683;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd29ce51a537687cd919d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6238cf0d017ea41e531f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h180e68ec97662820024db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f74e72aa391f2fa938c9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcaaf6dce10a1b6d38443;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ae499dadce237c8ec8e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f4f09abd7379e01de19;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd539d8844cf03fe36894;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h369c47fe2423e4267685;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'had157aac03c03be4e620;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160fc3bd1fc26954f273b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15de5edb8f4a3faddd3be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11983989812dd3bedc2b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5edccea56d9f401a03c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c2481bf4a96bd46f08e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124907242e7f8904da0ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11353c6599d7705b380c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb3ff5ca1bdb3f638c78;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1328c9e45dc35ef16b57e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8f26e5acc1d203d61eb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157b4cacc8cd3ca02d913;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12db1b4c66dfe446a07f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d22a6c41ab8992f9ccd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf999d363eda08e210bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4366324d41411a158284;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2eb520c21e4650e938a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3ca2e508ad25e551bf5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13faf089bec56d54f564d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h25ca0e7bcf8a1220cf05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1129cf2e549554bc59f78;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149301043e5d12e51f894;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8cfad665853938e0cb68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f661c59a11d97fedfd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1345180a78a415843c03c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4a6091fc511ccb9a6197;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6936605c98a3c78dd5b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2cee844c24ef1d7927fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h498e005e57ad5111a02c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f162e9ac0ff7a298d4a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8a86d1b7b49ba7f218d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b846037488a522c7ed9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18967d32ba6bd85df9c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a31371e03c3184053abb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2eecf774682930265d90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bac5532c62894c98ef4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1699149e24f485ac6256c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbbbd4f7c86daf747aec8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h528c0af3ea7c812714e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e32c12723822e8f0fab2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132209f99a3d601ad5cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1deeb609b8b166e0dd68a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72161512bc9e109f2a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h79adcd730c575b644114;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff18d663efd69660a917;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea1f60d9d07c9f2378bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h173094db69b7eb36c5df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9f98d71d9a519aa14a14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h35ffbec8bdb857253a1e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d7656ac0858e4c8d50f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc96ab93571fd2d4e3bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123c0415db7f48e1aac5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d09b4531fccbaa50520;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103204ff075dd76cb0842;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfdff41aac34bebef40e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h37acbadbc5beac907984;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcad3e0c6ad12fdcc5517;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103f5fa0f13a72c029d3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ef680f6307b92c6c8f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b6f1966c1a5c352ff11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc22f7aa70830b30bbf3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b7c115add6bd3adb11b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e09c38a27bfb15c1f37d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e490cf1f279467405bb3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1547b2fc2e661e77f83e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb14e17141d7dc9dbc5a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h184d85f11d0e2bfa3ef87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h861bca6fc71b0086ddea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h174cbbfb8735f01799bd2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f5a848afefa928b4dade;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178be126624a22cb4219c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154c72ecee6939cd265c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d85a605f9ab77574dd7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc301e556456ad4eb70f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d1c98e2c3e6d7c1cead;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2de23162ab5accce947;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22a7321adbbf6bc97e4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e199551d91c92f86f9c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1174718b683db6618e38d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175c3f7aff5a9ee14062b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d6d35054043f17be3c63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2c9e80c6954dfd61ea7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58470d583cf2331b0460;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190c6cf64d1b4cf5b4678;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10475be58bbecc80f20db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a107ae3c1a681ca633;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f1fbbf6dff8eb56edc7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd1b8c2f8cf06004c873d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10f106de330ac2d93679d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b72cfe9754d6d9caec2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a90ff4c9b80e66487aee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67721636f66c3796b36c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db0aeaec18941353a4fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb368b411a31817a2d353;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104d9e34ea462bbd03069;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d73babf44028ab563b5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17570d1bc93d1a7ddfae7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f01ff73467ea56ace9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102345059a6a0d5b58ecb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a12be0b67c7bcf9e5b47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he581c86843cd4ae23915;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d16c7e1d085f8258760;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc96c854532936dc3cc04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cdd3d6e07391350b447f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd060684a6ed13f4ba18e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10415ed5c307d54e4521b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1921c48cbe983b9f6de1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7fcf5e40a1f9a2bdb1d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17989b8c00603357f050c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1726020a790d9dbff03de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd862bed90a63b70b2ec7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147bd85f390c6c8dbd42d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5f3d76beef301f77eb0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c59da890d1945e6e15a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167747e4b8d33b92d012;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b82043e318efc0dbf2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd5c6b0792420e0cffbd0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ec31353d97530f0569a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ee790ea9f895ae048bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ef0f9a64935cedbffeb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc4f3bb32cee0954bf0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h233eabccca12bfa4b94b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2327bea0037e5e73f1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af1337c21414bf210b49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac070f5b2a0f9de107db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfdd78e416c4a8fb1e14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae5b1bd20ebf95273b6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11a2a1b26d218b5c564ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3fd4afd1c21421f5c50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1313c3e20b4ac33837fc0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1935d0b58ff847395e2e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc200b63365521a90295b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc590a908856e9971412d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae818777899053262f1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124a310e10448d298d74b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1757f4f6d97e5ac7a513a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1906527839d876d0e5f31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ccc8fc404eec1f8698c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4eecd8affe2154b405c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17dc4544d540c5980038d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1044a7b47db55523b6ac2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h130925f3fb3207bc90071;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h301316d9b7d79861f14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f4df020eba4f13eeb05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9ac1ce655265fd1ff4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d331514ba2dffefcf3c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e56351409cba706faed9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181bfedccce8db18e78fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h338c8406d0c0f2a5e049;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b276590c703e9c3ef94b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e9897e30c61d3d15bf4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf1a07625b2e445e29ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3bae30b46c4c87a3c4d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1686b7e67438ab3b145ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76b26a20bd9f9adfc724;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee7a2d52b99036caee67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20b46b94146667c8e39a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h43a5870cdb8f6c5e1500;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2e4ccf558da6b9fba74;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf44e93f2178c66abd2df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h790a1ca920fc91afff5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h870e181d9dd3c797136;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bafa892d04eaf6991ca0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f81221f600f1c1367e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1262cf66b3e88b5f2b708;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb8faa6c7b3eed7c51513;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f5e0637707144b20ac06;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57e23c004f0a764a342b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de67cf6d6a4bff7f9ec0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38e3a57dcb3a330e6952;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc1e50c190545c9cabae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4746f5881d07738c11c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16eb3e4410988366f1ca3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e40876fb6c059e973d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7cd511a8d0dea7d0b27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd64f02ad4ace4df27b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193c21aa8bf1f15b1975a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1793d87e980ca17c365ca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c75910fa30d830d8f6b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb282112dd521b0cc77b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce71473d0f5ed527eca2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c30e6f57a37cd79f844;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a902054bc15fed39fb6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c0db387800b118ff3c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7c17e996a301611ceea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee684413d27fc83f675f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d4ff0204cbe107a76f77;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cbee2447f44063bef718;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db001ee7a4a6ef9844a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f7e45c2037a49ceadafd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104904ca57c04406b0b50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0db99d409c32d6219db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ed941c9da95fa76863b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h999546aef307291a9159;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc724fc0bed17b62b7c60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b274295b4648af5daf5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9f6747452b3471fab92b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h288d3ce57efc8e252b54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd109073b64983c9d9f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18168e2663632109587b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1348cc0e4fb612498ab0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11229505aee8484ab65b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c220506b337100f0599;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd0c5a99b71b106980ee6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4e4eed647b74b88bff3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1299881e5598a0ffee10c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1193d7377733b90e5c1e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h82d4bec9f00447a4902;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc53c53b15574dcc87308;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac35a0fe296472721b0b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94e0fd62ad81dcfc67fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1daac51b58f144a50de89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6ed26260a99736a3c31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17306ee1d890836d8bf57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h715edb24cb9778ca5c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b6aef5fe610d8bdef57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb958c874464b3eb20092;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b51d83536c7368a3b770;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17a4743437de9792d63ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbdce3951d2e83ab819bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92ce6b4bd692b7b71d29;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17734e4cd0e5e43e57b44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h477185937ff98934f6e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131073d382590cd713301;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3b1c2b6c55ab1d98e5bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h594cd8dd4895a98c7404;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1294ed465f023505facd3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h525a0a32b44ad9b3e50c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8555d16590440af8a09;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2013c88d107a05d433f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc1a0ec53624cbcfb25d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da25cf80909ad36be228;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aaa8e2a4bd8af525f1cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7af31296b49abebbd26;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d47d7ac5b328a0fbdc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1851085c29568d71b6797;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfd5171bd4f1a6958c36;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa2c8cfd6fac17718ec8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b8a98b5798416fac1a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3777a143a06c52c2a2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c94c1ee708dc84bd72f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112010bc2d0b1339893a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7f7214ef9933df1fd38;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he4577877b3aaac73d06b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb45a67d04e85b16f681;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1592e09fcbb94d3dc5e0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbf94b3cba2c3c525c90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15fca6e68cba7ea80f6c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ad298379842831c6a16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1abae7c2df3c5b4d479d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b9688578740f411c1e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ade1c6f85d896ed5bdd0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1242d68556cf8e85d00b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e213a5aff5320850c4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d663184402cc4f8689ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160b50222a602bfd04fbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h99c8d819389c76062f42;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b34a4bf11dd91980b56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9f41784078e0633838da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d1c4c534d7f1e9a0758;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eafa0c0184fa59921a54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af7f389a448c66b19797;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d643c066786969ae84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfcd04696b3826bbb6bcd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0fd1e562555e78410ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b92647c025100ca8b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1390346c2eaa0ea8ef522;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1bca2a8188d086b32f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f1835f28379605457c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h130dbbae01a3158b259c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h568920db5872cc0d0d23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcdf0bc3ae507c0a0e579;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117877b2b362e3eeebc81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec3b3e809b5bb4165409;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5a142bf765347c324cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd9bd12065cd1f19526e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f607724938389a3baca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f63380186ad6a2f9935;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h165ed3bf0e6696be16f9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ffefb89c5ccf3ef1c26;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heff69358e4a22e445cfe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89ccd15a101d9c7fe1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc4d0181c70fb9bdd89c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1550457753a2e8aab58bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c133a10fc0999d4ced;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c95b2aa724b0b1a3336;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146991cabeaa03474739e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb230c12db9d98d4bf614;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d862dfed6aab12e11b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af065b3cb4505a6bc4fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3bc4668befb288056169;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c82ac553019b75f7b80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8cf06cb7a202b740ba68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he52e7c3d5b4ed71d039e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e40702e118a3158ba2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5d66a692cd4b5f893d9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9dc19da5ba6358f668;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5b963b1eae2c86b5ea8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f67ca41d827d3eef4c50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec11174e08876b69b868;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119536cef8c375a99bef8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105f6c576a3916bed82d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179b613c47bccdc9c3a12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21e887ba77452d93afe1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h189fa43a5a1bc572fc1ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d44a67d566033ab60bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9eab984ae25f1f429650;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168af4dcfd6bf7b66baa0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h133a3beb2a8dc02afc300;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16181a15b5c042bbf75e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h129473d2136d527cf56d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h40ccdf617d04913d9abe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a2eb0050bc21c8ccd9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a4075a2ba41d576d11d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc92203d5394f42a1ed1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150e152a6c3af3b614702;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b29b24012fe74eaf7e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4a7ed6840207696c2e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bafc992ba8634aca1ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c25d30f82f14bbc2c8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2642255a857f370d2a95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72f7885aebf23d191653;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf9342cd0410c6c109de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28318e22189b296470bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3cfed79c001a19578eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d0d36bb4728854ef43d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0dd7e94a2ce67411d6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h983446580ebf1533fcc9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc99c404a260ad2a07ba7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de71d4eac2f5632b7d5f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d503b39a166df8535375;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c223634a22c48a5d905;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d877588e667a4357dab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4387fecbc64d8668ae46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ccf79a77cbf7349b3e8c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd5c5c4e36a4adde7be5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f4e8819f63a15b8e000;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he2d63568ff57e972d774;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67363f462b3956acb765;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd1cbbb95c8f9ae43b1a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1685803e107489b83e3b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1203c3478fd60c14ffd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6d8e6482f49db493cf4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1372f3f49e9bcc413215a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178332773451905f3996;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125b45e9954a89d7bed72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae937790461697f710f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4e6cdf14cedd2bc6490;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1749c56d17749a71cd0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb6d0b8b11241aaace9f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a886c3af3ce07d97a9c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10f14ea89885520b79a75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b8de5f46b083da0dfe1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h873f33d6e6b7abea72d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e1f097436d9960850cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfab9059c97b1baa98bf2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5f6baf04e8bedf3e71bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb99671b37ac4f26011f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h109bc6e9c402a6dea46ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca438b73c553911ed663;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8f2dc9c7b6072bae5da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h439f7117c9fd150b5dd0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9095268b381f9abf6351;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c52b4c057872d49dba8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1887438032dc89b4c35ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b19c46ef934def72541;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9c89364a2c1c7523eee6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6c85c8669f2526f8f19;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3839e0f7a0b6d9ef8ace;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c90b970ab25653bd581;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b4938e7f1b3b5fcc5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eaefe2e6c88df2d3c16a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h101ff8ecce1f36224acfc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c09f3c3481c5a8b3592;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ecab4acc461ce21714;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd6c6d1a2afcdde482e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd1b54a8124d44a68051;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd1d02755917a13a2f04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h121150b1117253bb5f80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd2e231c542354a80ab5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f86e4773eeca494ae9e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf4dbc8d0d7b0bddfcc6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192faf68be7e4302a331f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd80b987de4e27286e4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf1d5bea03cc349044e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8af880e619f378f6990b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be671633ba3a41a48787;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135277b15b5c67ff8a102;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8fddfb9b14cd11f3ccb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h133a85b37ec37105b6bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2cfaa8e63fc1aa176c62;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54495450d014f56fafb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10906c4c6f3e1c48740b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b137b57a28df8940f15;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d91359e5421399154b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4f5adc1f433a71deb44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed28f95c055efab0ad3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2a1805066741616d66a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c4944508ee94c522907;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1179eadce92ba7ca77f22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d121e3dcf76e97c414b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4579213a23cc8232c260;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7fa94cd8ccde843b0b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3f3ffa5fdab7719dbb8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he114c1c23a5a9c86e58f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192527fc4ee933ac0660e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3e14543601ba3f14017;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e0bf1e1059b53a062e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7b3f751cff99a69a4aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192b3d4484efe69e44a16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a963b68d10106819ebd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168dba6deed955e604e70;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h50e402a2d26200f4f979;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf875ec0bd41e8fe78b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a5a5ddf8f3cbdf2ed2ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ecc375a6b025f31708a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1499bf827f84073790c43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he606e181366e10020c9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1670fcd5e73a4491b963f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16fa31c79248c71a1df51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111ada3ae0f0a7ec627d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c68c341c7ccda6b0c92e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a9f223ede48daac59982;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33126a62eaa86f664d6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4fbfd8dbcfe01530699;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a76578c9cc56ed8cee58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h487315ee711945402e65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1adf69e80d1fa3753d65c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c79707427549c30d3d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h367def0c02b6b11af55f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb1409d9079f23094f0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10b4f97d6652be80e81c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b4b60219745190d175;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hceb2037a4eb9f7c493cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd56417c2a73d3af73b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a9e0092c21bb27883301;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha768a9cc644a4199b821;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3d9d59064d9a18d54c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h85d8cc833753f1f66aed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f6b2ced470a41c57e16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117be557158fdcaf1e2c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc2926a82d440cb12e3be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf9df26dceffa2603dab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e8bd69aa76de7fdf37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc5ec222f88b938f8749;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'had485853c443ba6a3d55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183abd7ea7e1567dc9363;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h793b64cf6642f9b2c527;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f21f3f2e5941257fb5cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2df03013562a7196e2eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64141169bc7f49834cbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d1a48e237983d6324b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8da591e788ab224ad7f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h216570924e8d95bd8a61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d26a8245b0870acce62;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf0e19c874b19781aaf67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h915b4531a3108df67e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8be3a0a7de71f8822ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15115085e9a1830efbce2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148d05241c376d9238b68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h46f76d1df9ac296554b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131f00792273f2c1f2286;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0a26b9c0fd8f5194ef7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf639eb94f77dda24551;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h684f470318c01283517;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf69c8213f86d63c6961;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b07fd988d26edd14a5e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db0eaead2c19aaac19f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8f944bf50466a9edf541;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h208008e441db820f0394;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b9832c602a2cf177bbd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac2338144ebe6d3085f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10257daed8245976c0165;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58edf7db693a9de08716;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h697a26d7dc96308fda84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11a9e0b16fab6aecc5201;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h86ba6871b24a15916a2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd286188f89244d2244e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b304815cb0eb5ca1b29;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f08e1e607642a25b6eb0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe3c3e1c1888f6083d23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62ef30760f3bee99568c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba5cfa821100539d8c2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d83a3f72b204ef74ee3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0cf5aa0e753cae5e3b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b23a6180be44c46cf99;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h651b74921b24f29d8938;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3b972dd3171ad9e62495;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e6f8a66796a7a85e4fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19974feedcdb904c37656;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcad4a311e7e6c1936270;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha5c01b015e6bc4fb7b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167b415c730094425ac7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he05e818b96cee66916fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e58ab7cdff82d028513;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f04f00283afcd52acd8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a3707920ed9563d089;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164eb2223c6f198a3a0e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1454bc6111240e4a84644;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114309ae3d2a216819ec3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbda245136f0954929511;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13339c7dcb190577b6393;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38d6c13385df960f9cca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150fee9082c9b0b4bd0f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb0363cabbf1c5ee2e9e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1705a6e6ddb6132e819;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h188bf4e7686493d0504ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b24cb30770b114d049a;
        #1
        $finish();
    end
endmodule
