module testbench();
    reg [19:0] src0;
    reg [19:0] src1;
    reg [19:0] src2;
    reg [19:0] src3;
    reg [19:0] src4;
    reg [19:0] src5;
    reg [19:0] src6;
    reg [19:0] src7;
    reg [19:0] src8;
    reg [19:0] src9;
    reg [19:0] src10;
    reg [19:0] src11;
    reg [19:0] src12;
    reg [19:0] src13;
    reg [19:0] src14;
    reg [19:0] src15;
    reg [19:0] src16;
    reg [19:0] src17;
    reg [19:0] src18;
    reg [19:0] src19;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc447b56be47de1ee239eaa3b74b96f9b5f32d065b844d7a3bb0782c53832696a1b233b560f954dc99b08070b44419796b680;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9290fbe24b3acfdd7e9306bcf84fd009e88b89c16f21df7a53c39b4f0ea05ee35949632c1e2ef6228e06a54b65a4db994df4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h796ce024b7f971cf8a071ca56fc40b086bae3fd2e577edf29c433fc42b6a35a84d897dc60adb4a6a9aae529d01f150bc74cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9341b2dc78115d38e7208abdd2e13b7f6f12dc5eecaf3c1d2a73e218a646f99bb7e91e49ce186ec19294e3fa2197ba8937e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd493bbcee39a25356fdbd086b88da5b78378f1fdf188e9d4273e158cf7589316a6d9a58d1e6365423d6b8b8c92c4ca9ceb7e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fcb77bf8f198f4537be35bec6483ac815b4cdd282a3848940231b400939d5e69b759886907abbe1b96b94010ccfab0cefa7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6fb81ee93a6f532196efba7c9b9236a7be3ebfc0fa77f5036bed2aaebc016b26379e1ab86520d49d04efa03c56f082621cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd88c7c3d4b6f86d4c310af28b621b3926643cfe6ab6d7f427414db356878d47d777471d4e6add80efee0564f4e524e18fafd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a5007ffedbda4b003396268d03ad42844a2ca54a2784b6ab44ad21feb2564c45d0a555fb2920a6ad0144b2cd3f93507e31f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8bc013a7e73b5f5742b830b4c4257ac1b99d6d2e86cea7c0918a73c1dea3f892f1bc7e4767aae61dacadf1fc0a7f41dd7b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8009a87cba3b5948b16840acc63740e179834c3c702d52896ea962eff9a740a3391147e252f2400f360c103e1cd32ddbe8e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a911ddc2e0b68197923d13480c8cc82c802c1200ee745452b7c66b31834733264a3a80f17e386ba265afd501fa661af2a82;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he06492c2004da6598cd73e6db59c657c57ab4a5092159c67d29b48956ba805eb912b52ad9405df27a3a8de1ccdac36b79a5b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71ba1ef57978c46a90aaa01343460ae643e1b37a2be10a5c6e5c41bb9dfd03c58df637e67f96a4a2ec519043cb3be0b219aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb41f1f7400a72e99701a0dca129d2ffbaf6ac31ae7cbdaef83559f9ae8a397be56b19f0df2794fbf51d6c789a9947c42fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b9e0f1fb7a0b561989ab35e8d24894325f4e7057df2989799ad804663b32c60be69f9f0090b5e9caa54156d62403208f3e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24706f31cb1024a97d9ac4b9b5e5df2df057f2b068d387e993d8937e0fa16e0ff693800c81a93bc1f37a7f4b9f49cb4a522b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h413d58df35655a5b1ce20ea5fc25b1c4f10a47dfb18036ceedc1079ad8698fb2ca5c1e44dc96c332481d241ae270d9ee66ad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb514ae66e9ad4998d17443c8e89cfd579cf58beed262a3e7ee26168ef0689c37136b49a9bb411921be8e9300e4ec8cd7a9c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf71eeb29e5d8dd7b1b44c372d113d997a7480e5a51f013c2c7e7f256f8ca4a3da01b3d0979870913b8ea55cdeff4db263a0f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67467f8f25d33dfb76603f8516f4d3d49142f969a9a641b5d9902f60798631ec2c72756cbe13c7a6f1e82335b639568e4ca5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc13d62b8d7ca2d5e0aaa3ddb891d48a1d3d80b334e01854094b9ffb7a6a82494a2303b0ee64554c700010b2c960fd2e3b48c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e49344a4a86b976a0a51a7f84ce311b8d405a49b15d877975e4fdb7239421ba7e13034a750bfecbd058bc5561fecd43b7b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca19685afb69e1e16cdedeaec5b8611edeee95fc3248a9d5b072ea978b26a653cabb04ec009832f4dc1d6dcfbb94e9c0c186;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcbd9ba19265b8d47a337c7f5225f94a679dc14b8a92c9533f8f62b71414cafc78d1d94d1dfe73d2e4d09bac27af4b0e5d31;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd89ff3db02c77bc906cabb211abf6b828e834866b912976d958461287828f9ce58095d31ab54165c482465aec273fac15650;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h165e5675de7fe2757d09043f0b717d4185ac5e8102ee238153fe896170a8b410738621cd9c9884a5fba5db4c762ff6af56e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb1dc48083b304109ea1cb49d7f2333e8fe43ad4378b0b2591cacdb538560ecee5e4ce0ca9ee520490c857ebed4b896757bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1b09c4ff488bafd44d7be91735e62f2dc4d71bc99d643f74e5aecc98e378ad208ad210fdfe28a60c06b00710c90d096c90c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h578cb77001d16b60a718e0220e53451391f8e43187ad8bea1d2711b114cbce8d7c53a2786d6dc6156c6e23d4f7d8bf1bc791;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd4013dceaf5bac6ec2cdf1f85931cc8dbc141e8fc9e117327c8b9ffdee953c00cd04a2eca75ec5f03e2f630e6ca1eb5b00c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb06218fd41885611860dad1c1a7bffbd6863a39d7c7ff663e98faceee1e1416a1359a805588d584ae2543e10b0eaf2b15ae5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd35eb88bc72b61d11b95d9c107d63337e4f2b77eaa279f0d20bfa61cc8b3062859e13c0896956f221a6b118c173431d06023;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33c51f95d95070aeb073190ef9a32babffe8b0ed807104dd3472eb7db21fd8da8da1e9cc4565de854a9d4b19d51fe9effb3a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb21b364f30b47e33a46140119db7e64624302cb613a62306fbd87136e3c53f6af17cec0c03a1e506e2e513a9379a0045a095;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed0a3560da4eeb9bf834d4bf7841ad6aaff7c315542e0c4886beee674006c1394f24b8a09860c9eac9302239160f7137cf6d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf0a920fc110d19923755532892335f0af312d6defaf5eafcd0dcb239c05028fe78308ec667a95aac85658e095f672a0d503;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd14b23f75d604156ab63e0d8b51b9be70e277cb0d5cb51851825526c1a391ab9d5ff43bec2d13de9242b0f2e739044088e00;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdb9a5342317e9a7e9d76c004ec9435d5f0eaa131d8726cca328fa3d82d90574bea4784e95423ac2e686610db2ae7cf0b6d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3dfcf878cd35ddbe08a03e7c59aebb0165660bf352cab05d92103fad7662b9614ffe16aec7bd42204aa072e759dc76389611;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c212d7854fb60afddfc9fbfca74f47ab44cbdf49c3b9a8c021886a3628dcb458c37e54d13b1c374ab596f6d073345c36a0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94b16ff6ba3d96dfbac0414234aa91e7f69d0a3fe9a50840948ddea994608edfef2e2022c5aaac5f2923bcaf69e68873cf65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41a833a3ea32ec09682fdd635dbe0fb0fba99e5d001a2b3c06ce63038abba8d6acbf7c2f1d1610f5e75fa2893ac036dac97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d643c6e2c2ac1aaf0e217666c88b5b70a2be8826c8f7459d4fcc90ff18b2c61e052d82cb90f1d344f3c90316861e7f7d7e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h472ed643515bac078aeba35ee2a3c529291e66841b6c025a9e53caf21bebaa8abac1905c35f29831d087dc5ae987424dcbcd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7bfe88a1bc2d7c3d64d4fdefbd89221c6eb3001f8ba65e9bd26e178b386f9c8c5ab1295185108cb3221bb98acc7fa0d4d03b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc36856a93c9cc603b4fa21204706400d84c4f701ea05fa8b0c1962c589716aff7c2c21a151aa7ab3dea9ac486ebb4b94539;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89665a0574497b6b857cc284e199aa22689bcedbff11db5cbebb01e918e4bc021805c83de5bf8d13cc0090180a2d5be24c9f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec33f03863c073e1d2f1c2301db8aad961555e48432d430dc87a99b7f7f2966d0310f7f88607c98015ffd237244135624dd1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h570cd3d69261227ff1888318fda2c13185de8723b2e9d6b3a73ba9c9ae8479d36cbba9fb1699b1d11a5f1b0fc2d43b23b4da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99d002dd9c7d01f172767ed352c6eefeb4ba78105ee266a951aff348e99cdb0f886b3fd7a5cc48047ec4b2c60d3f50940b18;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6800d82c9dd197be57833861e454536318f711d9e2f013c8ddf5876a152b05cc3333fea970c3afe2be373a182d4592a4b006;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39876da5eb0973becf55e1abb9e5d2856d4fbac813e1dcc34610223be1cb98734c0ea50200edd53f8a97057c4cb01e358a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h638055ad1a0b8f127edf9875c8335c476d1843e151d16fac5961981101c87c6691aef877776c980ae586fd742617de0aba6c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70eca0c7fb09a78b55c3d6098e8aa7ef19f1f51888421d3589a59d870e08e2851e7b9c84efb3f1b787a1b7af313dc89fc949;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a41f905790af6b22814aa6594b61e2c5af7d328ab0b1af10bdf41660819f50b43a57443cb129881711fc4135c3016d8e6a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h144aaf751bdbe6b06979d8f65b259e004efbc886b0a6000d63dd674054035262d43424111515fbb7ce39e8796f4900162136;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb0ef46c5557083a4813f79bf148fa94c2284b58e6e04e89640bb5f886bece08e9a5e0ecaf2fed306439fd7a397c5d075cd3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27d6914c79b23e2a650712a3dd69ec8f41fc04feb025df5ae0bcc3ff002b006ec338a64a1bbf819680f50fbd825a24148cf4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88f874aa882209355ca04c3e6a98a3daabb6a6ab3881008b2ee0906ff1d9441a0cdfa8d001a9e52e6d95120b0048c7793aad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29210bfae556f595cba75dd44cecb114e8bc8e62a491eaa6ef389ead5093d20837e5fc10761034d5f44024a36c1494252955;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a0e83fcb2c83d90dc883c903bec9e4b4ffc4bf012846b80777451fbc89f17ea3718935715c7c4de9cc93d5130f61dd11dd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70d6a52a7fdd04c44e7de499bd3665acbe9ee77c78a137e6c470829a58ef9b9e1580604befa6ddb68713e1113c6b47ce3c14;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2609fc7b999db9d7c028291ce538a3e6e8da950ec1fdfbd2093533a1adc9c79b9eaba0ba8adb839ec06b25c0cc6d8b41cc03;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h864c3bb636220e0d36613edd33d4e42d149a310d1571b89cff0033d946c2ceb610a49dd74dd6264ee9faadb5f38b1403ff7e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15b5b430f221937361656fa72b35fdc42c79490e4e5f5703ac629248847fb2230b291b0fbd66ae135afde532c6a80d41fe78;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88d826c0bf0b52040f9e7ee26591b8d772f2bacf47a4d79a367e0cd250271893270eec17c05051aee907249a71e3db104ce7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b7ae29f82f0956bc87f1bef738bc1fe34f3eeb860889a377208c9182f048d2541960e2b0fd2ade03aaaf57318bdda12046b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h303bf5cf6b97bcb16394cf3f9a72ccdc211c5ced4540b6c70a92fb5861c16eed14b70ac6cb1a188fdd72e0a6936c5928b4de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ac4036f28f89ffc30c8889d8ca336f4b3b0dc8a6d30221b5ecc74dd73e5d023b9ad8ddea1c2b84c5fcec041c57d40e91fe8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h795c98a752454d02e87c8d60690b05be7f0692064b516239b3322e25ed4c602b90f124229fa71e2e0e80f9010b26714dc11c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6926663fa9cd1e46971f5b6c279b2a8e2102a92b17879bacdc83a91e45a897766cf5477f72fd5ec7d3cf011e74898b958939;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c26e252c610ba26d76e46ef0be822fbf992d0ceeccd479172e5572aeeec3b72a94f85456e63324dde870d74586a575ddfc5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h370555fa3e40ee7fda482227c9d48d9b84322500c8fac37c0b021a61d70a8f15fa1f3e8ef70099ce33fc3598db299f818939;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ce3d575d6241e81cfadde70f5f87ca08e6c7d80cd1471f4f7c2f02ab0e080fa7839af1864dec504dc86a36f09b37ac22700;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4df239cd2e8a41d310333151d73789ad3b21a56f2b0089b58a8d98c268d7c9b63e313a02975028f9e5167b6bc3bce26225a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5aae7eacb3e1624fe4b62f8e6141e2c746ea572fcb34deb5fea3e680f5bafe197f9ba795949950269dfd57c8abc075cb4af2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdde875d36a3289de77b94aae6703947dd37dc33579372fe7964e8e29dd5ae3eef58425575068091ce6939bc1c84ddaad693;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee0b946140f1ae3a4406ebb6ad0426edcafa4a7373366e226b135c60c2d3c8e91a66bc6be1426fd6ac855ee873edcc9d08a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a8a52ff387ff993fc671c83e82bb49aded594775d915af397226a6f455b6ae1d8d3e4fee0e7c872a914684f2991b752cf72;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14e57adb30a3f8de777381a962a5a08bd2e55ec8a817337b7d69b268c983ff49290acfdc39ed6531d6a4ea488a3435f7e66f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d42df4f175e9f61635d48906f56a7dcde4ee29ce988cac5efa24785e59a382b3957a5b3998a9afbcfe4dc8b830a037926a4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66b18cde8f464207196ee8020b524992faa74845579610e151e3d4614b9b7254e38e0c73c9b60e5f871cf82ed7df4fdea095;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21378499a35d5a26d42d64874a6df23789c7503fe058acd0e514a39ba274d80beca40af739509af0955c44ce7e1938d1e33b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h181a4e5cae4057bbb5581c0891375360d59dc68e834d2d98ae0371914276755c5dc13d7f1cfa1d77346514043dfafc75185e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffc85bb2a547b9ae0ad1479116af9f289d9be9b9d2c72246c95f77e5320f25938c2cf4e62508a679bd486f0934471da89715;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cba5a4adab18dcc791b7f4c477d261c25e3407c5839b8094368a85359fdca4b8304930d73534c1fbfa0b7626d916347ec31;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a017c3c3c2b558fe96db8c2019cbf0c6a95dc3cd1be28dc9687c0dc36ed66212abd6869d6baa50a7b3e1f8edcbcf83f52a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha649a902345afe7c000e3fa8564fcabafb312a021f35c0c848851e1ff9a6b3fcd67596f896fb58bdc4253aa000e4a889a6e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9dcbf918cc51a0f822951aa942c47be92d0da76a7ee57c56b1e4e0fe05ca8793197aa7678f9363398d8174a8c94f7f24c00;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc3db0cc1fb60f20b964eec5d7065da451259d2e772123ba73a97c52f2c6368e6540b97bf5b077bb0865ac56c496e9e45c41;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb964cc920dce724ac39d3e2cb0143e39cd6a1a5afe2d3b86c2c6ad1faea25085e29807ed76a147583eccfa6edab132c0ed0c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c69b5238ab6aa9e768aaed204c9bd3e6f64ad7bc5fea473d996f80fe079d32ab602436dace727cc54446ac8a5258a12c1d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f402be1cee5992f7d814ef77ac34bd854b4758d0832d4338a7b17235e5e833d37c06a267ff21cfa1a349493e71176b48684;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb51e44af80c8732982e521e11bc8b6db486d7e0fa158c680a4bf52914f7328ed1e1a7fa3ad4b8b7580391cdae662ef612599;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9a0dc4f9766d40ea70f2b930ee4a271bddff8dcd20ae22628296d409eb5516722ebd1ae583902d76bc2e16caa7773338601;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h271b6780e2dc50415c8b7525d02deb85db4598996c22abb94f08e4f836024d38a350f53a38ccbb4e0a18658afd790de6794;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc53205256ccfc1f6b61ddd0ed9f36e5c9b639105ccd7f553fe624d31f5c5dcbbbb9be0a3dddaecccdf005e6ab39026578d0f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fb82cde96e0355f643157e3a4a64798de3d70924ccc705eb72badbe9d83e39dac07c1199c4fb2b055f7ab88564eeab68f85;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c25ceaafb951de9f96c0f0099e681d0ea51ddeeb84b9fc298885d6a75802e3db8ed3f732e3b62386a422d9f8150ea601290;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5f9251d85b60e88da8b629df630cd3be5ad91938bf945557f88d4657df8d06f464242032335636a76703487ac646b64d5dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haab785deda140b0ae7f7528adcdf26bb5891fa1051322bf865047ffbb4e07ee397a17acdc8006bd95ffec25a4cd572929632;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd141a93e6271e74152d55307ac05c910209537446ffa83249b7d27fb1148c502f63a31406ccbeae9f2b0dccb755cadd10d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bda7ba75e80fef46ad63f0e4d26591e9c5d6377c4ab9f5e359028cf8ca0e332dd2bf5b5942ad7acf9972f86894e38b4e9e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h173c73558aa8035553d0a79345be1fb306451e41923635a08b256d74971a4045d1fe280ac6831c2efaf26822f57107733392;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3abe1f3a8e6129f2020af73834d71521a557557a2f80a0fa27c0b7acd98eeaaf775043b38b6a35ed0f57cff5ed8a220fd4d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h973f6705aed817b5907ecef3da11d476e5fc755bb74cd65ddc105ee7ec16826815e5f59ca68241fa6125062af46462f4e9ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb279e6a99800b2203da6987831d9f63908579cc186b8129a7654f8c354529efb9684994413bb0d1197e4e1174557054dbb94;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3df5a1da26bfc0ceface00fe2419b39e8e57ee581c0130e65f5d90a3e328e1c5db584e19cff2599d36c43df302eb0e816b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h779950c077ecaf014d18c6290000ca8aeacaf0c2cf94aa29ff668ad00679335bc4e77f9c45fd14b85918833ed79add1d4614;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb2cb0b6e6ca436023f4bfa882a1e1d5c99625eb0117842bfab0052ea1d62ff8071d51e4f2d4d8c1ee60c843ba69734b1e41;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haed925c59d0fdc412a721fa8c2774aa18404c166ed174884191d31a59273138a7b12a451f999e599debe49f8097a374c6ace;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfefb73f60257e51f8a84d9a9612492656dc34137e39fc7510bf4b3b213162771776a0b210b139f3d94704064bf03373ac165;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82a3a52d26ab8eb8c29c75d82f8546d41b500ead0375e4539f464798b3fac2122a63933ee1a914d814bdadf21353adfad6d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hddd9e9fb508379b80b074e18a2ce3da8a6d96d2eb217830d838e6571f1349f478641e0cf4aa5f832494f14ab30bdee69b653;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1bc3d6df7fee30fc67d12e2c3a20cf666889ec0003567676c82e44c53db8e9f7d5817d1850ec87513e6690f53d93ebef61e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60f115fa45938d0f7aa596d481cc67c639097d97139d703bd904242780e90bb42bf68083ac205c28759139f36f7aafa9c416;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1d7ff3723963cfcba9926cfb34253c23f7ca38305214400e88cb4677a43c6fc09f638a4aaa05f68e73124c80454bacc2db9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66d632ea552181c4d388df6afe4b8ea40238351c1fb824a7031ebd22fae955d963fc5702fd16409946df7c04e0ddf230aa05;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb95bef404189439dc92505ec4f1a56cb23405d67e05c1fff4370447c646b34ae9e4a970fb28f0c9afb8dbe0a9f7493fb8e4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ae25530b6522f66f71d8ba6d8cd64774c9254d87132b705dcca9a58f9478d8a243847c603f277335be7ad8e1a1fe3b66916;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35fd6c2104d8f1b64abe2103f4af9c330b17289842cb2ca4572be0d6597ed1da1b8cfbae82ab2d57e34aad67212e4ea8446b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e5aaae45d2600a166a95fd9cace8346512df9873a5c6de42144ce2c4cdf89bb7e1871b26ea4d8ade3c0040efdbd2524f36d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75ed343512b83e9b32b3d6912fb4f20cb42448091ef00c049ec6c16262ccceaeeea85e2f3e83e5df83bac7d1855b2fb49d5b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cd6e2f8694c50ac59ef8242737d3a0cccf73b5854ed31d6a98a25d81eb841ad6737ea1e7b558b37d100c1eaad423bf5e76b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41b67a10f4d9ba41deaf60a10633a56fe0b82bea57046c50faa9eca6519b00affed6cdb288e6c5408e304cdd12163a506b86;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4227d3d0894e038bdd6b64321f84cbba1a7c4dbd210c7f9aa6b222a7b1876593253d7134c549e5dfe47cdd5a5b63a3c9a12d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h839392c20efaa86fd04ddbe0ab8312600352e634e0de58d992c7780cbd38879836ef9b0fbd78f1fc07a0e74620338e93919e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ef23fdcc28ed2aadf5711a657aef2cc53578d400d5b2812923beca4f7eb35bddfce5079841d003873c2601a0cd1b3443559;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1410a61b47e917c1ad348ae50bc0c1d5f5e73781543dcfc94b9d16c0e3c3f4545b26a8c9f6bc17b9697824c26eb0503df9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d2572956ecc6adf48225405bf32c0d47bac044230d444b17ca41b01cfb11d33f3d5562aa64d5b073495cc30a84afe152ef9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he989b16f089d1356cf2c003e5b819f7aa87c0976c768bb144102475662aa2ba1f04e809352012417f84dc5a1603bf17a86c3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b91b9903d4523fe52214312b982d5c2e840c55dd5fbc6052c462629f2819cda51cdd10178fde295e091f5455511fef3d89f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12d03249cd7a2e43f0e6b36b6212eaa26f0b9411109ae9e6323f6afe4dc87b591f9ced0f96879b463310e8da2729830236e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f811732d847d78c9ddae9703608a49b7dce9d736046bed6654acdcaed0c5aba1680e0943b5e1bb2c993141bb730cd1bb526;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h773e5fa924911ff8ea483bcb859c787adfd08b6e6d65cc11f6a7ba137a4fd91d71a2d67fc9042af8d32957a0039f3ec6a6a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h460a64a96ff856d2d78f6f5ed7ae51aaaeefe9e2b99775f99201da7b7135462cb9d72e54f04fd351b7d63fbfc4d8afe44948;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he35c174a7cf29a40570a3299be29b4bd97576037fc2aefb78bbb8a979ce385ac802c187d94c5ba2f6ee505448fb8e3ad8e4c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3682c08665596e05687e0b0a09cc44b5fdfa86fd203f34bdfd2c2dd42cd24822545e37b597c0905d36e7c0665f4c6ceb9b2e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f14b0df6c46a8362d70276fbe52cd86781e915c8d8021035af55259adcb0d91d0e7a1b6d8affb796bd5aaadc721fdfbcb30;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b4b2b4cb63d5836fcf4877ecf245812afc2d5bc88bfe204bde0fb844e2caca0dcc2a5a16dd7f971cf7b110cbbf5715828dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c68d82e25e0496c2c48ab7d81aab9b3abd78e741e31a43f3e937e6a868393b1df9de59bf2fdf5fe456a31185c9563d2b741;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b235525aac1400db882015b3e03774e77ed38bc0338313bcf1174b2141a87f88f2bec0f471b0ebd3a705aed66084e3224f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c0dceb538a41fd8a61c94dc12f8d6ac0f61f67823cd803dbc26e944e4c8a29a354e25d8162c654ed245d27a0ca65d521bee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h475348132f91ee83da894e38548b4a29f929af29191274282d9bb950caded18d5c92ff987db045e8a1c2a869525f60f9163f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a94631f533825991f85b4937c4da7bd6cb57c0a3b3810ae1fa53b3ad8cabbc89a393e0d52408d0651fc67890bb21a0223f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76b791bf8f530e0f0ce96fedcee3c70166c0d31ddafdfc47769c86ddc8e03903c0a0113873253bc6cda85d3468de2a0307c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d9b866049097ce5171281879434f49955fda38231f9972bd99b48480cacf4627f63c09a569b29901d7e2af2a433f54ceda8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a4bc28524effd25a630affcedb93d35b0dbba4b5d19fcb292a8c3fb42182c45f053d6a8319a09892e5bc18e78b252ec4fc0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca4f02514367bd854bb46712c498903dbedd7e369f431c05076cf94d21315433d925375f73a64593369d52c170f29bc76ddb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ab15dcac21c4e9e141465a681419d8cd2b42ea843955b8d8c8bedd32838fcbd9a42e986254495e46a5fe42756809cc5dc83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf7210c065249ea011b41f58fd2e828c5234b2181482ffee6f2daa47fe82b22105a711a35b895cf1ca5834771116887aa284;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h745c99c81be0133b2230ce1580af9a6e884d17db1bba7f0cbaef206ddbe2ac613683f23b1775f71c3facd15abf122f8e14f1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb83c56b4d31d4ccc044155af6817949244c9350c0288a61bffb8012363e0054ffcb130175ae4673e2b849922e043e3c7c13;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha114942ea23109b430d761f4469f04d4fd6bbcab4907587bd828ba058f8777b8d7a454f868ee1da2c887cce1eddfa3248257;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9f1588bfab0488c12ed7a0c4fefbbfb667d145d4f0ae235d16fdcf93df3fa5d66aa6932f598d645e75f63f70f0d1f50edc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6bf1d03e7a04841b927ffabe26fac29063c3046e8edcdf1de70e2410548e97202ba9fe72e81e82250d88a3a966d199404cb4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d7d7d07912c9ff31ac43b6811d94b46a91cf60c84f246118b1859bfce7caf0248ac1418e96e286198535046641832c6a2d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a9d6c42722605a6071f933dc347ac6afd5d57a224de3326088fed13e481aebfba55bde110913791e0b28abb95978f6d689f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb2c048227faa349473e1d9663db25501f39e9a0ea285a6913f0938de205b60d8572fbaefc886c6b1dc7777e90bcea5354df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha87820a42d47cd15e66f70ed8929bea4da470285b768386fd061b9d12a48c7397df6ba985b50232db0f1a9aae67b2dae0da1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he94fd78d9e89612b2bab71de7fb63436f0e996ae8d78e1c11857644b0bfaf49031d32049e8395777c106f450122d42b70db6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c1b5a4bef099b18ff6a8d11aea4b4340fa632622600963b3236f02fc1baafdd85eb443bf5883651fce9900d490ec872666a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7385e04920a87815b42427803087e9522eddcbab2989d2cda25c096098cbb8ae52b11f4b192b052632d99d598844487d02e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8135bc81c9d666dc06bb77ba0af1e61172b95204f083057aa28d8146836bbe3aaab20eea3c91b7e7e6cf6d07474845dfd838;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf78b458f0e427f0176cc9ecfb727bcfc549ebda84fae2d4e5e4d3a1ac3c62f5007f76e4b575b750676d1729c68f3db1e0121;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2af88fcb777f1c63d81fb03f0fe1812737e6d2490846fc76644c1e5b105a8a712f6e2237470565c39c94fe4d7cc5b5c2e204;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha465065f098dd6e2b03f77024c1235350e2d5cf46c739b9a5630a9e70b3a220e2f6bf4bbbff7ac22e2d86becd797255be4b7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2b50bfac3ce3bca90bab809ae9462878effee21c6101ba9b6ca21dd1bb4a76f0b794feb8f7abb2fbd1c59a372e0acbe8eeb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c482b80475749cec97a18089e22290df79a6c83f3afc1805750b64833e2dd1426254480e85a0d349f5c7792b62b2d6c07e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8316035eb8d2306608f81b27eca6e3a7bec41897cebf9bc39d55cd8744c25d6e4e0330b21acd4e7ba40f94d25674087d443;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h491ee7e2b4d62c8f1db015c4fecb7b47baa1f5bcdc65aa87c31c72c4e6781f5631eaab3535b25fbe936456b1028c6bcfcb66;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3dea3669ba1158823e15bba74f4f0f9267e3b56e9619ca2cf435d5b5dd9ecc1152aed33ba3a2c8edb99360d6b85791e0d13e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h286d5480fba13f0b872a144cfc7c63484017dc9b4de8723d6f4886d36a571d7e3327ea352f8745532ece886ed90881470827;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heaa4786499725dfda73bfcaf6d3eb13287a1289899a4c4f3d2d590effd84059a0ee15d184de70fd3b311042267b3832088ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h412eb4fff2ee356cccee78662c49111f3f86fdd11b6373309e76291b9dbd3f2e534b744ac8ed12805847b2cd66acf2e842c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h100c103fb68c305f3ba160f6cc4e88aaa8fab5c7ef145e15a1c85375c20bfa07e4a881a78214c5a3423a1286bc88b00fe730;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27517bfc434ae2c12e1519ae8fa4fafc9bc4d40c1bf6c5982bfc37ac184446b8ec2fc5eb51ee8cad04fae07cedb17a5fdd8c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38cbcb9cc2a7b683c7118c9e6f9162ee239b024441e16ac1415b44b38c9f17ae5c5bebaa40e4882a1755f43a30758dcaba3a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdbeebf8a61104a84e0e242308ccc2bff2a98c6d6ed8aed3af3a4842ac1407b09987b21225fe3f6096ca7c12090413f70ae1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd91eedf3bab5273994e855506cf267981245e3f39fc8e9361134fb4f59a1e983528c7fac2721170655f3e58ada5bc6c014ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33416a4fabf7b301d4a883f2811e5b7935c44eb95ee59d4d6d639c74ffa2c7d3512c53c45552242fdde991a9356fc7853930;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9919a8bd27e460b8acb1856ac5e628c08a27a10e2d26d5f58fe45a2a09474d8f50645dbad0e72c2502e8e055c0846b1862e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2f64068692525c5c6604805a79cb45a46d492b16289c7d6ebb1650f5e8c7ff4c32f4dc0ef83dda7c87e6374cd39c4c22a57;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h517b094e4b543025a1a0d583f850956e7f16346da54960c1edcd465a5a10e43cccb87a1879607394170e103fe9ed37c9d0d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f8398a3d6bb764318e717056303f1e020e292d1cafe73ff9908844b4594ed22923fff7044c542fa5e59010acb73432433a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46863c187e44d8789e44b759917ebb7e5619d9e8589719a46ff27419597c63180d92e48226fd63342fceb6fa870bf1db1ac3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf84dc68332df9756ca191387fdc5c2f9594b8691f14df9028324b2bf665c83f2886ce65fbf03808ae7efc7487e864a96e2a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec2ecc0e008c7a2848f8fcbe4e29721615b867e0edc78d9a722f9ac9977bd595fcae917384676db1d2c5e407c8380881e6fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ea7b89078a3c73684e4ff4d01964883db661ba0006bda1d88afb24868f7ed224bee60b046554604d472449b4cea687b8297;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he93697e847de7cdf46702a811de1ead2a6b34958c5e5a1446bb8960028c073704c90f787fd2c4b7a645985e668a8117c5a54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h354a237ba501c2018c2e9da232196089cae287f746f3e61e4276236ceb7fe06ba4f94a048571e967a35c7d68df07c6c11655;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb49eb3104b0634963b8d1a93b4fc2b05f48d6a6ec72b3f756ad3461bcddeb2373551b89945a1268df20dc94949d82fa09ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a7d2d42c5556915461abcef0582745d6b2012e608ed49e365383d3b40404d96fecf3b9004c666b3283c9557b5aa7dc325a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cc6222ca5bdf5c06ec6836599761ad86837522bd1987da7176dcaa80aad78a42c2c58dc8193c98ef4c9675e0fdb9f80504a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc59a28459d16d36c1c43129eeaf34ecd43f0c64277dad41ebb65621e4353ad421c7d3d646da4c029255826c45300a4b61fea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h815ab52ee33e54c91360c477fa2b9f9c82646415d8df0ed1d0abbb9731353a3a6cf4dbf2ce1619f84fa239da1cf8e875859e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0576e0d7dd7ba9061b87ec851f5b6c2e0e8be4bea6b5fb076a663ff80f46bcfa6b05509743412e14554b175c07774c0eca4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9548fa7f9c50872e2ee71c8c5c82a7f3853499101d00bd48d8b5781365aeaad8b118073fbc9402eee2317c8ab2806c543628;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he955249777dd61c926980566667a0aa9cb43a104b307862eb423f5e547f5e3c008783aa71e037c2d9a026d841a30f33a8384;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he82ad2f6c5a0dde524cddd31219bbf294de46333063814aeb7357dbc51398fdc4636d3cb8b1d7bcb6dcebe6ffc9018bf84e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfe1f76ee45f4f7da09bcc08a4717be138761265ce7368d48bd484e0ec0d57815d60757cef73cd5a6993c5929fd5198ec592;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha18c78e7605505b5bf53887f8773161edf6f9c893af5365a2edeaa5c6a3e502cec605e0ef455dad41ed4a94087e4061e69e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6771df743f6e693eac85b2e15bb565f44f0bc16bd619a03df91eec79c1e8677879a4fe044e0b7c4f7415684f34e1b7821182;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc84ef5d1310c80349bb7dae67e6d4f5e699951a48e6e97d90089bffaf91e269eac3fb04966d7ee1703c2cb2f1734d6b692;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b9972cf393405c1f18d2801ef0ebd0eb89fab3575560e0a1d5f99a7c08a7fc8cbb3e3a6030d150ad4f0ea6f3a19cecbaef5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h492a4a1e455ea6f280a0c5fc4ec6a1497d3abcb2a672e703310e6a9b18d191871c37313237a5f198ff551c1cc256c6caff4b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c4adb62a5d264b743cc7367d316f95b606ca2d9d8d3dfa593baf0420addf7fb0eb11487f94f0a4afe02016d43d0f3db35e4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29246108448f746cb93771720228ff44edfd7617ba2cc05c8eb1bc9db1dcc4415c448f3eba92837641e05487531d9069175f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe87728e094fa6eb52e58e00d63ade8e90b99e3c6cc462d2ad187849ff289a333c8911d5faff5d5adf9221d7d1bcbde248;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd296ff17cf0714919e9ea1a1005474741b3a46a9a7dc60856254c51f26b7e23436b7c8e800cfee1f6a24e5241cbd7dab0ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdee0a28a6191233dfd745f514eeb5476d00fff2f9c69c98ca2d5c81cd3b2d43fb7234a8fd35def6d4d89c98824857c75e5ad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93a96340d264d46fa68821583838dbb3baa44bb38f241419d16aada16f811f42d3f5073d675711a67eba4defcc664ae3b6bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4114686dc6130b4adfffeb93f39a03be478679a2adda1d427b5462c19e219a841b43df95ffbc3ea6fc90ef4b52aba001e07;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf692e79296e514d9f8bde03c55a91f2d3ca8357715c08ff000b075b21e0b05f5de49719d6e2735f7782daa5259e7068d140d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d0318985d917d18a3604f7df2191c54f73a7cd561410474625e97d84b091edac41918ff70c99582fcf5c2240bdce3509b9e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ad3537ab90721f1f6bed212e8fd4420bb914d4273b89773bb1a9e5f1aa1dbd0ef0a8c67d0381d8cdf97271172c757b748d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9a2392b50502e129fa3249d67527546157a86c8c4307350f67fa756327b6543c783a68fc3276f18c4d22c57bd91e872e773;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67e6be68106263a5d07ed4e38c3a8f8545650c2aecc66c06de8f50fbc343e2fc8e908acc3b8f04045d2ea74b7ec9d3253835;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ea67460a1b7e57509db0c96d4dc44cfbe8f3553918ea48da6a595e61d967f1167213c8bb3a82bf01b262f67660c1996e20c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0bacbbbbd610507ab50e0d454646a8ce6b7e14a5dd0af49f59fe8641a8977d972757d6da522156fc3f70e3ef822c8e69566;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadf1fe7e5c031d78f1fe6699638c59866818e074f2a3c3bc533b6d2697bdcac2184ffc17b818be5c22d2107bd6da82901b98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3bb98dbc3c55354b9cabe94d1e65a4e54284b38c93b5afa51480f8bff6822b3afa442d37bbbabda35b4f3441cfe8862869c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha444f4d0c2c84271fff93afdfe774c78d5cce7f3e0dc8e8aff6e81757663bb38b2a5b9927e3a94254d676dd0a1443927179a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h678f24870a1099903bc075460f34812ed7637e7abb085cd96695c8e3c79a2feb67846ff0646bd50bb9a55b6feab84ea36fbe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c0a7cc0264ea1408c2b86fe54ce80c24b411b8ace67e4174709977a857052f075425d79dd8132e82b81cc76405b10b40c33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5e7242ed5c2ce35690fc46eb08670f79f9834c81fcc13c190a69530dc70999d03f3219573b853c491f57b3e8da5658dbfc8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32bac74b82aa636f8a4731589f3d1c3b80d7f91136e72d20683bc4fc896b5e356b17b12dafaf335716625f03e06362e41ed3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0c0c11bc612c768d1632cba4e669cd90f31a9c7488bd00590f0375b398aa0d7bf56c3aacf66f8d666db91e7d44f37e85dc4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88f84123a9460767eb43638755e9e7ebe3f34fa98ac5e01c4e7a8f0eeb3b1e746b4207a8d8f607ad6f70b9725271d6067025;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62cd279f83378f34d9b132daedd8491567ae8cc42ed3031660dede4e719754e7dbf85dc5f289711f8c4082885c749cd6eb98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54f20fe5080f15453a7318b98149db8c74d54e1b92f572a1620775e3b0a389da3d66982e933e4f11e0bab736e68970a7265c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c1fc51563658bb8dae05da5d5a118dff0669a51b45748e821871573f46697d35f323034fa9569e1b3e86de04f78bc7c2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h147198689d644b12a9d828ff11af849e45ac6fd6ba0307fc69e33cfa7f225cb33468557530a136f958c48b704c36523896f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95fadfb015edb532bbfb4fcd012a7f8e16c1840d40e8b4785e0f626b8af01e79a09f3caacdbd3e2d6246e86c39f53c3c771f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fc484eb1225519b1b212835ff2907ecc1d4ab09665d94e9665bab1ffecbf79b4f8a476086e0340f52aeac75b9c3baeab64e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h962bc023bb20dc1da1f26dad16d094692d97de0f757fe767a4276bbc2892a30c4afc7f16f0d5df77e14a56ccf159b6bb584d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h480cde4af848d35f31a98ed1be21552d9b2a46daaa0662dfd0703c774494963ae79ceda23663b5dd51f4d85bc87347919740;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7bfc43228862de769ddf1356333a5be664e4757587ce48d28a7b9ebd054c451f48efacf240e1d7808c08ab90a9a469c549ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e8823899e24fe893bb6212ea6714a118edf500a3dec6ad5a6afb2b36a96ca9e3d2792914aa5d7630e26ab81c6756a5cb302;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc099563a446d474f1d7bee071a237446c8c6bb9b45a487ceab46a907011a9377b7c29a4d4b8dd601f31b01aaf68b1db79cc4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6bc34fccdbc9917f11f786d57766f7a8dcc121ab83171e5b5dd1a6da098bd4ecfebf750c553a967d059df35c8a0ce05b8f4e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h585d97e791b39fccb875ef4ed543e8f93d62e6f437eaf5f73f3a2a05fdaebf2d90abdc8b56d6b8b217a20a5fc04c8c148026;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e55b2a53bf5562e8f88b9e17cdd34a131623ceae52388f57d0d0175d7531fb7109e0a20f7a816f167bdc408d20c6cbf1613;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf30ace8692f9896784d88b37788a205b520564afc28f6bc1ba0eab4a3f35ad7337d4f9b7278f47d362242598508b71efbbd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf4f69a25551d8d50125e02a7de7d4bf7d832b2f26f8641cc189be55265d8bc7cc6e7aad5215cd557bcae7892a3b41442af0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ba5788e1d68a299804a687e1450e0bee1409d94cb336bddbe634b4af5500a803c07f95f38e95dc13c973cc2a993af8d06ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h678ee3b9b90e0e7a2ad3f31c1e45fd7d673c8d7d2cb4343271598393ba9bd72b05a3c333a5927ebffbd8380e64d24880fd6e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h330e75be0ce9486545181884ca74d2a8feab0fe258aba4f8d89bd9fe89ac21b157c32d068bbb218f80595789dfa3735c2e31;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f85458a60b04d1d420ddabcfe0ed57f7e7561ffba2e48133cdac8ef4792f97bac03b8eca8e2cf8b7bf768b73bb89c3a8ca1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcaaa0d0b2b33118ed0c3a1a9fc83b67edadcc6a34603e59144263a8b3c578b087af7e1df333b210c1df64ed7945216996fb8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7a527b923dcf010f8467690c292a188c2ecf54a78007bf0c5babd957fba058bdd7c05c86845692f2680674737001270d757;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h478304456affbd8fb43edd15aeb4df0ff0793d5f32cd2a33646ed923ec7b7b11c39efeade92d75e1ad5d0efcba430c8dc579;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44a6f1f99d9bf4e88763293651d1d36871b40063f40872568583ede71ddaad39dbae16d10117c1304903cf5223b6c5415bcb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4558ffdbc795cdd9ee069a2df52398cbd2e007e8d355d3e641f7bfb21c98979cb8141a571cde590d8db9e28a111f8c61e03c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4bd5dcb5e904522c847bf77e9148137c8219bfda284f1d60514c3ff3f9d13488f7a2a431de3bf2872221d18bcdbc958582dd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9db1fd07770cafe55f276124b70c4d12fb8be8700b30ddba488d84052841f75426c0f1496bacdbce1e8ed13b49ea95fda473;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b4d7228f0beeff4bcccabf6621e0111dc9119429f96886ef1d35d8b03b2511e6730d17b50eda0550a08770c434a14fdb2c5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f518706be64b63cecee3b1b8754c8636de1fd6932090b5708e1af7eaa0632f128dc1a362747fab6801f05328841c1bb18c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdccae206c94b6f3840f3eee119c585237fc565e2667e98e5236a393902e344d4dfe46371d30bec8e0b4fad486c4aa80449f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca3f0bf104914ed357979aea69a6891e099ec9ee0b1390e93b7f4f662826b485d58c4fc95564acf98e20cf491212d8a29019;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he17dcb05632a4741021c33ccf8d14f1c1a06afdc17cfab30456841f5cfcd3319173e92f658a4a819305996cc0c3465c5f3f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66207289ad01ab9d16b490ee0bdd65bef7315129b6ba66b9e371a7c44c0a9e73c5c37caa40a3f9d3c72b04dde27984bf0d15;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5eef48dbdbcbd5c1c7a4c7c965a0bcb0a8fa5e33fbd19e930e64592e266d8b0890a12bb337c8e7d6c330cf71be0a08a9498f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9c95836bec69ec19f2ce705ed3e0b1cf9339c9f4911f3f2b7e3337c3f87d7172526b5064db83e27d64d2feb8786798a980a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49486f729670b08413f492f89840e72d2e2cfe9c0d3258caae606c6c550d1645fb996439034ee612cfdbb10edc58871f6ccb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37066e7596c5f586268bf374aaba00d448c84b2f815e6e9714a132a9be1a31f7796e8907871440aca71227fba4f9290da18b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40203dbdeb2b157d3ed34b14c805ab081271f2d4b65f9209eb893a8421de61dcb35d68dfcfff5981463067b3b87ebe2696ab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19867b1324f975cdb83f1abf33b878f486b8c6bd6542127f9b5fc9cc6a0e1b5ae63da8a4c9780233bb8e4f1bdd7f24143451;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb72c763094d9d0bca58883c659595152cc95ee6c5875a2ec26f650917f32c7fbe27aede1a1cedd7447dfc4be08e9bae39312;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9850e861f9a834ee80cce2d9eb025654ffb539ac016271ab379c25fddc3000ac3d87a2eb9163de5615eeb69d4ebda79bf9af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0b81bff547e92f1636bbae082d7096947aa603f34f1d757682baea5758af98249df75bbbd33e55c760dc34ca0da2655bcbb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c9b85efae32988d7aa24a9eb947bd8269d080f5148a7a800e7319c17fba669d2be5af1ea01abb93727084127f51bef65959;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f7fd6b17a26044a77539dcfebc5b478d3c91caf6f148e191635ee89ae05c4cfc7a19841170e9296f4961b3337a7abc0e7f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8cd3e8e4796a4737c2aaacef88b7bf9b225c4c4bc968b4e4288c778365cc8b88359d64b318b0cc9e935c5aeda2d7d9c7437;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67fa0782f4aad26abe8bbdb94d254a060933bf0b9dff81bab8331b04bf41362ea96bff43a9a3b15b1f4b7fcfca13b9d16cbf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb182c56478b9b2059297f02bd4404dd472339e3cb6a751aab15a1ced7f904039e362c9e2439e466657f4a2641c37b3fb9487;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdc1bf55f0033a9cb9cad87b6314acb722cfbfab96558f8301b188b14edbd88eafaf3f00a2904c7b5c1eb90e7930a37464be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h743eeb6dbb831f6235d27209316f4e5afa9facd667b25f654b93a97db760ce25990c928ec327dd992364b696e41200d1462b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd5a4fbcf922e367e0d927197d004adbb866eb3ef8d9b305d99d52e66caf6fce4b3836714d8b40e63cad2f53dac56217c6a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16c0c2d2d6dad6cd8cbc95e24b734b33f6e2052721085624b5c22be323eff77644170a220b3a0bc20f863ea6c7ad2c4cc6d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfaa9cdf6daa3c5bfa4bb17332b0c4192c02b08426a6b2d3a2812609b51a0fbd0339bc437a1f0c8aa9f2474f182671c592b82;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he990435134990a20a2475d91a1c55948a8c8db07136e93a6fa6714204dbe14c801bc87fffee33ad5e7af0617328920ce9086;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafa01c2fb2a4c02b50e9bb4bbb12d921d01a2c03e46d3cb2cd070f8d0906958d9e60905caed61d94c73e746f49508bbc5cfe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5720d616b508552624cf7cd406a9e1f22d83a3024dcece77f58902272b3cfba31efa86a2398b284e6d3a09a414352e2daaa5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha695e7a16b8d58854b1e8b2c7cf50d6f7987556c0f962a1e5ad4cf4a54da896cbc3031bf174c356f04c080318ff07b2856ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75e802369f08cd4bc7c4a86fd96dfc8b42805c7d9d393b3a823b3a8114fdbcd1bfe4d44c73febaa6159e922a676ab8a8174e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcad2407e36f971fb1c0e28d2842c7943fcf9f1ecb18b911027ef203045d5e3cfdfae92183024382c7ccc0dcc37b0c72a21f1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa1871085eab2139bf57259e134be548f6d27b4f156d8b2c4aeb849061040686a7f0fb0ba792266be15a9ab580c580bbe08f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d2b3911ac2e07638acb30a9bb99a9b2576c10891b4579b5094f3474902e4acf2045fe3f1f50e0a3a6d3a79650d51187073a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe522b6eeb7a6a409383847e14ab69a389de24790f98cb4701881d377e3777f4be093e88a5cce0bb9a50e9d66cf8ea1885f5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14a50d621d4e0f6364bc0c1033329b858475d0807d31a77cf4cc7bbc4dc8de37e71c2f4a51f1216aeb097749d9689a9f9b43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74d4018d8f0c0d27686e5ef0df5cdcd73733d82ce144b4b9317c2c2460215fbc2ff55501556ac7c3f52a3db3c998e6f64270;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h601df6f6320b0fc7237f2214188762b309996c5315f615c78f23cb904b0f4746e63df63bd76ee87c665e8499c90461239052;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf0ec673c5ee5d5aa3355dffd229104a60ae2b4a7e26f5d37e790e06aec42bbeb0285a3f6adba357ee318d5146370ed9e4f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e3684b51ae855ce5abc9e8d06337bec8df3a4f72ea35338f3f29721cafa8f57d4645dc915d6ba7d37f36204251098d00be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha351868b4ea8eaaf42a162a877e20fe6fcaed6aa37a17cdfbb904264e456b405ecfb1c9a6ff62a6c18f141784e4ee99104e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h337c71350b704341d4e28c5752b61e61d52f2560d0a728b191f73c112ba57f11f5d9484ee6c5b0b5ff5f3254c88ab5a2e7e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fd037eb25cb13875d935145d95dd56e2d65e212728c8b3ac1963368791773f1757bc0941c13cbccd1b41132fd3ddc3e8410;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf22f9713edf5dd7d3f931a7bd12ca6dfffd744d02ea64edc01a0bb1e21dbaf30b5de4f4d3fca100274835160bd5f6606ac98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7bc9ef0b9c32cb972d1bbe7a21fb073f2398ea324d16466455783900f4ae863c0ee40f61db12edfa26a7b20ef215c677d89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3e59c4d27cd991c60c4c13236ac850e23a85efdcbbcc141dcc1d3d5d903a0219eecdca7b1e2078d4cc8cc84d524ab29714d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98aeb3ccf4b3b7b128d5f2bd28f55ffb1396b339b23a374d9fbf65f34339a2470325b90197e252f36ce75e9d5da9592ca8e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb126f56c376b572d5bf64a828fa9862ae91ec245e99a5e5dabd4ffcd17c668d70bb22c6e7b51573670a6d6b05c39b044f61f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6270977dcbc64bb0b131b21ba60009e47f3d645c7dcc39c8ea96228d4ad3d3fe26355c795873596518dfcd328a45c2ef39b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42f5af4342e5bf5baa9b3ce3b3af19186f8aa815c79cc7574b4fbad6d5682ec023f4cf7d9ffc4a0f453ebf3015e563fc7a65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heec3a27246969be51f909bd7be4fdf91b65df5248a0e464664204f78f8cc5e5ed5d4448d168b263bc22b308e87984cc6c335;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e5477231cd585aa98a409f7f8fef5d1ece8c4d1a19f0be6085a331b80079138712b25bfa5e1790b11f5863c6c8dc2f56ca4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e39598b405fd640e6afdeab2074b2d6a246f7ed89008333aa7be14fbaa1b63635c7fbb3bbf6d1a102a3c4a26d6a792ed09f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87db5bdba9861fe631921cc22ee2e18cdd298bb0c8badc23d02cc59a6e62c64c41cccf09c766d6f30d71515bb26d9bfa95d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44d340de747f0da5d36c5c1053f92810e0d5668ec4177018992791ff2f5f877208362df0259b86c575d5f3564ff11b1c9747;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he38649fbe262a461211d25417d88cabaf3995b5a62ad371c2a016f44d786a39cd8b7c9d9856e5a094f39a5db3c37b84b7bd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c5fa45d4314373fd5fda2be2ce5f726cfbb4764d385975309a93e86c0ae713acf17459eb6e6e1252ffe48457ea4a1a9403b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4cdcbe7c1790080186183c6506791203f55257a9154dda17ea3432ae5a6e9c3f6664eb04c325545945d2c2cd19f1145ee1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d2d02da610d8b4a9c3d13069f998dcf59c515527429434fed473fdc7cfe594f7c4330dbcd669cff4d4f141f5aaf5db45d96;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7adc0690a45d2757c6980013456700b13060380098a818bedfbc9f19748326aeeeeac16ae193e434e3a3f47578c7124499b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haca1db4672bcc6a9dbef3740e0ea751b441eb6c91f90f167de851885682c7c63878a206da79a99dd71c6ebae05d32b502af3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33cdb3fae090961df2f21487580ca63ce653f6f9cc9cbca3fd06aff0824b49cf3041ef7f0e9d2dbd92db3d119f9d4620e8c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92e70743377d082a5b5e6c3245a87d0d67b6093966e8851ab0d73cf27c8d000f4ef168b85b1feaa24e18bb532b1ff8f0614f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9afa5b234aea7af523062d83157083e0e511a4b98cd0fb0d8fde9f1f78cdee4e5dd90f3553aa28c50ee2cf4f949ee29be43f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7b983c9454549dbedf791fb40301001a0548fd6c8b3bda2f41b5641bb0b761a60ca5055e9e07ab833d28610e34a1cbef68c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccce1f81bd1eafd263d2767622054b188a6891d1876d5ab9861512e9c1a35c7b841f80d1f1e30e51172d2ddb1d21d42da61d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f8d4acfceb5c15774f476c58b04d236efd0ff2c8e1a021c66c36ea5acf88045d66d672b39e5d721c9950b3e40f83e069ef6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5714a98bc82f82cda72aa44bf10a34f4f0233c71bf06aacc60b0b0788831dfd9216e8f9678195f3ee25a177bf6e0394157f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd62220c5bbe65b15cb23bbc44134037f21d91ba1d6d8b43062723d429e81e03fe81324068e4aafb212c6c954f0b70fb3496c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb6c046da4cd8b2c2cbd931964ba99905ec86ef90fd4f8408f3d32c655134868c8c92bddb450313f05ed7eec6640b9e7f332;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab6a3ee1ab4ca0fd7a914a9ce0ef248a3db52e1a57e9c3cfb658746d7060284b36b725159843f170b6b0adc05ad7806baf99;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h134f3cf8677da9bfcedda43ebd1baecfe2afa7445994ebd3e8a9c2765024c17ddc8d645cfbc965c1e842d399590ebe82c8c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec4a5ef873effb5d4330625c15c6aa176a0fcd5e7f812aafff5c9deaf9e11d6b7b21d15b2acb44771300a23034a9c628ec51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfe5e7a246994d2f931d91b94c11c4e5b0c88ba2e2187204b647862d44b642361f8df3950d2b5c20bfacd78a1a238b971ccc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a6d09566c7c625aa7aa233423df321c6f0efa39833c96aaca759c2db74f689cba5a7f00d4ff78f7befcc5f8619e4c0146e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e9e2e4fd56916aa61340a8050c98e735b64c24c41456abad38df2aed471911ea500adfcdafb98e9359ffae78d77c840ab52;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd10164c8cf08f80076f73e6d4a042474996e9dba4d07a435859a944bf6674b2df7323e86db832dd2e8ada587561cc5933679;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8803d5fe41eb289162ec90e62428274188dd4e93f89fbd2dfa3c396c19a6c6a37ff3d670c2db0794bbc85c9974b87e5e143;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h927553b9b8b62aa66d882b1a3eccffba9760ffa0c185d88340f7362b3eba2b2a94e8ad236a6a5fd4668b074fe24f97ba83e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he822ebad2085c792948f2b6e2eab3d16d83ede932e2abb23ac4b08a609eae4fa7e39419c91ada84b9387b0a03f2356c55d40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30dfc683c3abe0f242a689087282f8ac8883e387cd50eb20362165557330df07a2baf67e35f0688db1868f2f1fa6a5667778;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41723b5ec370c8b46611e8e754afc3f3bc8dcb17f6f22a41d1b65bcf2f247faaf10b2b4d8249c161ee899d22db008931a8e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7bc3b1b5d00d20be256756e6d9c1081b3e2273c0ef27f624fadad2edc2f2cec14361ec9d6905a405875a94f0bd5fe984fb2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3c7e04bfe028e6fc36ecaf6cc52e3688abead9f1e3edb11c2428653e10a89025b76708154d3c8fe49c0871a662cb7b75607;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4dd26cd089c2784fe71a203c4b4d9c0dc4676af79afdc21a94b0b09a484e5852fb4ae758d9eca6e5bdc24e653dafe9e9a58a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h495851e8e20555e7d1061d542db8dfd8db9e6b6ee37bdc830b74c1ff73aa8ab9902356b09e28c74000300e9d928fbd4ce234;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79d80a226f7b47ac372eff7395017ba7aed125cfec48c7bcdd5a89be9cc3090918ab38ac894dc15d7662bbb66b5e39d4ea14;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf92b0aabff0ca09d84ebaca656ed74d59a0313e22cccafd09c6fab563d4876fb476d1b451033c51b2d0b4c3ba7690e1358e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96be70b6513d907b7b29889d9128f1b92027d6b3f4746b09ac6a934327b58131899023b5f52ca2fff9d9d34780d6df500019;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c0536740cde1af6aaa1d49fda2882b91686fa17c1b4350069473de5d39c726bc614994a3cfff791eb73fd64529caf8ba7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h830b4c822e065f3e0f4ff305ca0b426b9023db17a50ac62d0993b4c7a84ba081d47c850737582ebab1fbc6f1c038bc89b89d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7846020a867c796dc945fccb07a7f80c50cba04ac30ff54520ee461c2dfbfc62bdb94ebb0ea8c5de39541fea6b6abb5b7e8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1471c7a90a839e98e9c953e7db8f3a2805ad8676d6e43bfcf4d0610128f84bfdef15ac705d1bdeb4ac878b5592e5158717a4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16d2ef62c12f53f462b63652f6d2630d20bebeb96dd7fc4bbe82948994e8c4054fa5189aef0960bafbc3dff84ebaa375e1ac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e3d708cffd9b71deb4c63c7775d18fd06e90bdeadf33ee86e94b6bb216ef911b29aed6fcc531d8f411024672e1f07a321da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf924d41a947f4317eeac762f0b41b8fb30d6770e3308fabebcf41137622f1e8318623596d2651a82ba463ea15e597077c85f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7daa3c69c6fb795b0dd43a3c43bc29c2b8f0c1d481bcc70e2ea09bc6b729bf90fc72e4d713e13d3f04c0296343e63ed2e686;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h819b41ce1a1e0330d699bec69f74e2c20c8b412acefd632b804d920d939636a35e7c1f93d93e6cca5ace2b9597babee7933d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0877153597334876ee02a3fe5d0a3b47dcb6479dc9d9f12a250f6dcdcd8379d471fc6ed6340b5256ecad4294c1049ea2c89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h712632435ca9f758b6caf1b34f40d9aed33f94de3ade9cbbe2814fe832ff482f1ff6099ab97b2362a215a17321ce49197bf9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dc05b0e65f3841fc4fddbaeb7ff2eae8e56e41f7689e5113043ff1e8d10c47f14706b7eed4c73a3d29248cc7853dcc89532;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae31b9a8f83ba313843580708a43252a6e161fc5ee7dd5932b420959ccfe424144ac85db230167c17194134ae44e3233ec9f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ffd9a904d2ed0019dccc77d99fd8ee288f6405d48f3196f65a998ca9f1a7d4a816d25131ad8f2513dbaf7e4790f878d60b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27f2a199c74d3b70c10842f24c6cb8ee18ff856b31441da76f1b9f4033cfe9241217a0a79f8f13c3a168552ceacc477367f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b8965b925784db25f39b5e74df31de02b49269081091ecde5ddeeebb52b58ab6583f5997c85d0959b82c5328f14ccd9c629;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf38bc62827cb3d13c26493c12cc4252b9448fe97da979e11eaf19fb33a0b657675a8079211d5268b4a99d4f833d1bcdd67c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84997e62bd41bc5e2e835199a588d5c28eee928e08683451bed3d75e424009f32189654f6b7554bd640b117a3b4e731ddddd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87a203cd39541b36a671c17c65a8b1bb4cf9208a203363fd6a6055804fa945fe337f5808e6888523b16fd292123e8fd10688;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46389085d36babfb54b58e2a5ed9f8a3d0df2b4ab5c8ab96dd1c716ebc9233eddb34118adad45591b54ea5169b953f51f847;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf140da197a5d16fd207e34b5b7a608fa31da6ac2b5c2fa8df156326904556b8ec6a1a4cc413a4b3a9767d5e81728ead8fc04;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32249c8679aa7d5841a8c284e558bd1b92506b12f9b3b5fb2a6dcfe16a08994fcd00e4a1912529b73206dfd9bb44ba826e2a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc6b57e6c33ef4b05147e5c789d8261d32c6951ab96ea5c6f774c4f1f1eb2bbb47c29ce425542cd663c11aef80e10693f6be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87a3418a003d8d4b8ffd59932d0c8d6adf9a435928d83a09ec9674c0ac72adc5a3092dda2fcc5ac3961f4329a54423a17993;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3837b471e68fa7c1e58eac9714848870b64e8757233e477dc676d08306e56db4cb20ac9c46799e90eba27a07ae81b6ad3cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23554aa3d01774c90929ce589581499e7a3233e8f1655c7ec852d7250e6d1c620cf9eddc9376a466c148f6c95e7eac3c509e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6776f9b8b2a53b7566c019dd798a1f36c938dcd139da2d64536b12fb4b9e4f814d2134dd688ace5391febf9b3ebed86b34f5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d8df38c5de4cbe78872b3931578457d96e42b5c419d39192c51d3017ee93099fb0f77ed0a794bd853a3d2528818192d43af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54ea2341c3b5dfd45c76b3a953f11d92efc36526857f14928233b31f7f1767b51655597cc9fa037d0665bcb2a5a15d18539f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3969b6f99e539f0b55ce2742197416675352dcd3921d4898705f9446ecf615fc32e348ae50dc69ada103a1deab70eb7276aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56d68adcf9a8498a31ac8d8e7c9f2f091267fc058debe5bc8d937ff835c94f70136cf296cc971dcead906abfd876fdd6645c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9461d87a15d37f9496cb1d5b1e5ee53acf924391913342553eaaabdb68d9d0a145626560e6cb41ea31d1bdcd03ef2748308d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9ec88346536f2bd05106573d46c613b1cad1339d6b065a584495cd5dc4bf60e1dcd74dc771a0136442d3f3d1575d68b3b1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa7466cfdc2e97c2a14cc901730e0b1c2fd87037f81a8940f9be6e642e591440acb65f7831843c8fa9b4efd9aa6a2c1de238;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd89ee8f440ff4b449ffdb1a6b5ec58bba49a450259fdd9f9fc93fc8ffae1e2f31fc68fc6b48dcb3bb7fa43a4b9ef29bdf039;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb91e6247e660b997efd777db7beb490fcfdc110fe4d3b4365273ad8865656a5c3d1e240ea76ca9b13554571727f63f9d3057;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbb055a49eb00ffe9f8694602dedf70267f763c225b7861a8681eca9676697b1b749cbbb611b62ac5f56e24299ac2b560f7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1ed47bc973bfdd5fb9ea68f17a623858c345839ff9067eb2a6b5e038d15089500dffe1b9911731866e2312ec8c79cbce70b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a62113f2aff47b2880cc97739c6d7f09afd1f34fb7731dc3196c1f9f4b77aa4a40efefb5aca9ddb60a38ca88fab2cf6a20b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf35a3c1d365359d026c1155a40e199f54b791ae3153df5210778b6732701eb3f8ea0de59a0253beee0b49df6a48f8a7b630;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd148d670af6505c9038c70372257bd88b8a4a043021c2485f4170eb31b7d8a0db2e7b5f14f19d38a42d7af2f3f328b217daa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf796c63adfe126eb823d5ac65e5e956144db813743c35959ed9336b8320b3d431fea89a92839c335555671fd68d06c0b5de5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbbef74690c5f019294b56e17e399d2765c13bb44f8c9e4e1df84e2123c2450eb7752604f7b532e40aca9bde7e11333de7b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae06af0f068414e2179f34fc200d2f6d4de96960802a4b41c1fefcaebea87d953bcbf63cd5172b39f94acce08ca7c6e73a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7e7d67263b8bc207271071b700f6186d13a169f2d2ddfb592f80a984917cbec1005fabb2273ab2a8197db8d848f0a1496ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ac087cda7c1a5cffe72c6a24c98e9e31565ab1aae02bd7be464a4713d66cd8749950fc90bb7b8cedaee8818c15595682342;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h812c63b7eb0f960c360b19db2014aa5bbe1d52b4af2751a520b5b1dd2ca9c57b6502e830aef6a12c5cc178ed7aa3712ab024;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h930818894df5a4ccca64c8fb30a833e4d4293896208deb02f9abea84b945cae9722dfadbd70d86d9799dd9d74bbfc1c7fa74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f655c4ac3d165e67ab8fb822b44d1af7f7cd31bd98b51ab1cb0c7aac6b52238650029f411bcbf95b23fba518871f8918e30;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6cc4c69de3a98d641c419bbcb46e78925711d65f7b967de6501834af37922eba330dfa6d5249521e4c26014f5298e2c8379;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65b56d83547ff50c1fae3da51032b3ba50b3229f7776dbcb90508135e3e8948b0822d68a52d2510bc6131aa0fc24a44bb59c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9d8979ab4926875f1de07a00e56270a123fa342cc7ef06d995118f46c8930bde07ed0e0f445490153c3964937f6794fd9bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b8bcace37d7d5dcf6327977739626846d749d14100665a975f527b79db72337fd90b8431d2d0377b4de2a64bfef034aede3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h105e46a773f7f3e3111a5dddd857f0e787b5df7b479e9ab9c62f58ba38069725ada579d2cf2345e120f570a1afb4277a4d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13bb3fd72a138d18cb1845c5f7ae65bc30cfc4bb886628879226dc2d4cbb4fbc346b1872db8570955af7c33eb14011d590d8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14770155850672814c99f4cf4eb076fb47c43354cdf6137d92324304c1163af28e881eaade9a332820fd157c33b7c26fb0f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3269836bcf7f901e84bfcceb8a5215b26005fd8ce4cf4d06132f821d378ca36677b96f70e043e94039cc063e2db61bc34ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17002bfe4a1a93a0e381e2d3409ffb4b214b1079c3c7e506ef9dea5eac288e2286c00edee45a87c8ab59b1645cab7f425790;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58993a4e43360bc84f2545d7c50d59a146865790e8b32b11a1691b3a94e5281ece2eea40aa3980b34aa6885e7d9870fdbc07;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4207a760e258c0de26d0befff13d82a59093bff0a6861c9fd3af61d2e2ee16c36c5d8be73d0a4b22c65fc84d4064da965884;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c57bf84e506dd15c3bfd7372e3697c0e83cd7d21200d07be19c368dd00e0068734cedff38a73d81cf2cddb009bf338784b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf60298b9b020ea824c1891eb451cf3df24c15f3479685d7717f6090be7117a8b8a22db9aea9f736dda6d0d096205f8724b87;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5390c7799d0d56bc950a847a83c5568d876d81f7f511e7552b317505b8d2a51f058a7f696befe6caf12dc67808cc8965c0a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h142a9224491cfdc024716641b62ac80c038d4834e586f759145d1e85bc421cd084034df5c829b932fe03ec867d33078ed140;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha398294c4b9e749f5873e3338f7f3f61be964507b255a908f382d2aac5c97f7469366273c9e1e8b77eeed5b887898b86da30;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ad2347dbe2bc712b431198058227f43cefb803f093ccb9210e6712ec6559711025022aae0df292eafb26f7621accea6edbd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had1ddeb770a1d4adbd1be1d65365bb68c47fa128b4661b90398a30fe5c66921bf5d5b59e3980dac8fc23c78c976c23a464d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8cea5038517460057c0edc216f1edc4b1b38acaff6707d7af11ee66691ee6aba954272e8955cd0ef72fd164fc3be0a37a8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56e694d51ad2ce23cf46af17b16aa453162aa2d6123351a1f013d15acbc2f480c9c073e32dc3bd69df6f455ccc2559cc73d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he82c6a3e82e29ed9b1b3f0883ecee110e3ccfaa460e8be359744cbffe4092c7d70aa21140e3fd650ecefc8667bb3fea24a21;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ae1cb526a9800e98cb1500f3c7b623e5fcd170e591d588f7a4843ee308a41a4f51511908aa931af128267d8b866ec4b853d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he69c77a97d3f9f0141809cc3f7fb82035657e8f7792c8bb3c797c17081cad514bc6da20e91c69dba8540cab0b544f1e2577;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6615402e3820f716e4c61ba7637d1f50f58cc9a040c490a05b1fba36ffca3c8bb99142bf5ce91c91f53eaa98a145298ae292;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73c34a8f2d3dabe25b363b1cd1e98784b3067db61b6dd42c4e76441c249d2c4d201cd584579295bbfd1f010ba613fe1f9578;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcae26fe771a5e7526c88c8a3ac81420cb6de7c109bb05bf9729da9e24eb459ccefea7ff297955dc292f46e58f7b2698122e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h287645afd66a04d21f31e2e9a8c6c04f125a011bef0ef3e6c0745b2d1f1afecaedfc3524acbeedf54ffa4ef96931cb741e50;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d335fb63013840fcc18869d51cb555723a9a1b3c1794fe4a0c9c310944bcefd6be4b6b965dc917ebe1a968bb9ff59a9b445;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd84c7a10db2fc89a2db51f8f823e7749de010bb8a34c25ac3524e6a7b0d22d26b18764ef2ccd69dd16847c32a18014c61eef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb984716da1d34053d12cf78e56ee1a9aba0b402431602edd4aaa125b71df9c0225ccfd605bc56f6b74a4329808436a580364;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4cd453fe5a991f02fffa080d9cb6a506d434e0ac19189c169e7decbbde046d7a4838b2e8e5d8e72b4a776c1036d7cba6258;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7ac48e291c4010a0f8d60258f6448adb578816f79d8068d104ca7b097dee32dc0cc87d26468af1102cf7892fe8e72af1a52;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h938ff1c60deec8f76baf5c8556b7c2060f6d4da251aa6623fe7d1c38e7a9b28b2189157e6c32ea3757e827e1b3ca2ef1f74a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb07d996b3b834827e699f8b983ce989a37e4b67914de2079db5a7077902d84d8577a79ed64055423624a9ed37d2b69b1ed3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8069b8e23d197f61c29e4160234f5584374b2a433c79169579469acfd6ab4e47f730781d75eeac436d9d3e8ac98d6efacf38;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc6791c27faad5b42707f4cb719fb664b7a1a3e49b895901a14c580d80954ad6ad83be01d0c42bcd8ffb53692266709378;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb94078a5fc8aed38d64f2bbe5bef21dc4bd5ac4465c3492005a8d5ae8331f60d29e2031c56e8b2e2b9a3c7b2b5e106a2213;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5fa793ded277c2a456cd90b2a0c987b7561f2493c80c0525bafb25e8d24da09ad1ac05e3568045c27026c1a2dba073ce9cbe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4fe20824d5d75e880bcdbfe1b33f3d583d55d72b4451d333924de742fb9d8f7f2ce33ab1db0f9a507efe9de7ef7ed79684;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9037b64886c48155981296b517b3d49b8bed0c4ee39a51c5cc9efcd9eff41656d4063ad12a935ddd20b1d5e275261e2dfd06;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d700130cd3a5fd38b88576050eb71f31c001a8b0065cd8acabf64c6fcf160399457c3dd4ae6da7f3e73a415185596189375;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40eb6a0038d3d6d34fa447fa06f6165bb7771b3e91475ae075c89931279ee43214e92b4b14c24804652da3aa83d6618cbad7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6269c19038033d1e82f1dcd20b60312b5ed109ed9da6c17fb2664704e9a8cfbde03bd7811f058f9a0567a9aca8c39b0f2acb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f04379472d07ad5f86dcb1716e8283ca88cfda45cf0d38e17c47a143e4e1f9d6ea5fc115f6ff965cd963aa1622f31efa665;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h410e390e1daad488eabede1f4b00a48bff7719eec986e05bbe7551e879ad722cb029d872747c3a5f7a0daef2ee6d0e37dde8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h317f5bc94246ff4374150c86df1d538609a5cceb082092c43a444032f0c9902fb84dbc98d2c46b6df75ba06e4beba320beaa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h876142f5ed10095fba35041307ffae73a87a1d0dff3bc42b09bf021dab70412737fb9ed0f04ae825203ac147ec7a24392201;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha89970d78abf1db1a1033cbc432df2e6461635e29f3a50c9987efcd9ef9e0b886f20169b5816863b5e6171f31f523a860291;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc76404a9ed60f7f81634598bfdc4cf487190e6416a30bfedf2a5465f4ea42935c8ce90314c9547c8cfe12041b0b48888a6cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23dc1595c612b0d8c98246159935a72260d98409696531a0703d1462727d2131dac6f627daebac1a17f1e12753088dcb6302;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f9aab672a5cd4e8c6b47cf516ffd6c203030e875f27bd989294ee886950d2f01259d08370f4b24c3effaa9f3483bf5b233c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45cea4ba06789acdebc14cb1ee6fa6ba217fce70efd8602990122693c94304cddb7160a3f16d20d93da1fbc404d0ab154d37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36216a1be24b9d1aa27a21c91ddfb741ce7dfcb8e70368430d434bc5ad2599c3af6ae2c404d3318b9416a03fe780606270b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7101129e57483fa51e8225a7dcb4d5f5a6a0a81071913f61d1868dfc8e5d69b9652d378bacbdf04c0e5e7ee8f2221f36665;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b493b4ac4110e6dbf2026c4acc879abe64331d71cfc72b728b3b1a3a6c4955a4edfc5ceec0da041ea96abc6f8a2191e505e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85f60d717a3398e9ea8ce01614e6236d0baf2573d5ec6abf242edce0bd0bc6d611bfea8caa0ebf9cc4518cc753e80cc301be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h919d6d5345bb98693e7c5f16b534fee6770e402ccbb834a977cf4389600544fc4052be9f532f3cdea3ef08dd22d3bbc4ff1a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c5f01e016edde44db5db0d0da32b94d10c6abad50694ecde3bfcca93d3ff8fa04a95c7138e67f0bdc3df194308438e7733;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44db572af65c490e38a1465c41da0c33a85608f62c65a88db35cdeacddafb894d90171d773be2c899c2828c1eb144f227434;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb302416b217d0e6a3799678067e4f9f3ef01f865af43dfaed9e4947342e8d566a9692dbd33813172e37cbe0bfa1f3a15c6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa52f1d82911a6ec107f94ac87d9cf250b01fee541306f97af525f62bb28963b6ea3093857b4ee034ba2e78d39f7b37b4ed8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2b7e751e11bce76a8319e3beca6cd051d6a998e10c83117adf5f305e0510feb7af8045ddb5f4d9dcbc7cfd994d6799aac18;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3db58112940942475d91a80e60ede899c0773cb0b020f7052fad6591589fc779c9b69e1993d2f21674948335be0e920c9e64;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8be5c9659320eb10a8aba7d900687d52e6a2b197bf628cdae06625ebe6a144a9036645055f418be06b036fded222b6dd8c87;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4d1e45f824e9b30e3ed113daddf3d0d86e77f480e6aacaaa95a13ba8d87da0966c2e48e719cef227c470c93e5401539a194;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h620f65987a53d8e45b39cd7645fe24efbcb8a77da6314c70a1ed2fef330ba2670652c9206cdeb688e6b2fff5aa500d75e5bf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7887bafc765bb935f87a788d960917b51f62f102964f2377003b02e8ec2c7f09bfcdadbb7fe4dd4fb07a33fcbb7aeaf44435;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4537befa6f3f26f3ec1be37017117f8a6f0f2a35144089e195cf2ed67d26971acd813b6f75b5d30cad033f50e5ad5c87e584;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2194d952aea25305885f6d03422de3ba352759e3745bba174c098ff1c07ce4c0da5f3b1c57dceca37e330465d2d41c9ac522;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h355075814177153ffb1a009e33180cfab671360038aa568e4055e74891fcdaf48859aefe2b4db6716bae7a7f141cd728080e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccefd0431f74b93f6ea5823070ef21813d649943624b7ae828d26392ddc6f1942c9f006a59019749a4d96cc3dd115d53ab64;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed255fbc1d925b185fbc75dce42d2e50a8a4449c20640e9ea0c5c97f18845f5792aace36774702097d9ab4dac3dc8aa0ab76;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c320fa083ef4d91481a276c58013cfcae9c0fc98aef6d9227a7530db56b6faaed55eb006b4c20ede9e4d5ec19d8f8a144c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29773070d07cf8ceb1d88244fc8e7cf9869b318575bb7871eacdb9d0905c5466c647d5a78c7177cdf6c608574258fa094e90;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bd3d9ba4262f9c039c92a1e14ea653f1272a1bcaf5af909d348baba8e14c8a1ec48256dc4dadb2a952bfc0b007503894771;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35b4f67a11bb25055110c7f992e6af42f422ed0f3b9dd7bdadb8614c7de391228170e9b02f576c8fb19cd7c9eabcb9c442c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ce402d67eb7d2f0adcd741d07e5473fc29dd80860963f4b694d3e7a7ba3f6d63a730778df629cf78652bea2ea965f3e8045;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h285e525be28125940e22f6a9bc661f34c1e82b733253d820d1f52d76f2d6f36ea147461d22da6550c433de2841eb9356fd78;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfc75d786c91705b00003245af6b7be51463afbec9d2359a3068963b9499a0a7f252821537be7c7c5c26006db6c2012b0269;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d7f8ff8e3e0f8303dc47ba4cf57b9eb295bdef1aa3435aa3619dc9b83f9388bc751579b675268837668ff1fe90109ecfacd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50a108d62d8fe3c5a6646d03d1f0dcaa57fe3d3512240de94759b86e2273b6603d8e74d742bf7a3d250cd206af91398ec28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ba809631239cd06b20099de11506d453b539d0e3667b4a328e336f7a1024f9781b5ca14efb3b0dda3ded27cd2e565ff3e0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd755d72cd64a85cf7af72685b4f1e3abd2cdfa19d523afe747227b300772319cf4afc4451203d16f6e390bac9936238ed4cc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha55a27b5ad280989f4b93d6a6411b30980e7bcf7e6cf247423c457edc9d778ad9ac3a7a6d0eeaa19b89f346fea19b59b921b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d47e07fa839bc45a80f45d09096f5a88799a143b3c38fea4f9fa995319656f980ec5647a189f7156d39dd040976146f1dbc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc62d561a7f823d6eb97e298be347fa7bb98524cff169f3bb9e42fbb65a857265c2503bbd8f3163aa7409e092fb229d56311f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1a6739a2ab2a15a0b9159522a4a5e12ccb815d385d655ae416d8c4ada7f11cc286323db3550b858ef066f6793f08f9822ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83da9725cc3c5a438ad2fdebb72ad83a5d92430027078610fa7d996fc6c50b5807f2f9d4c4ef249f1324b51e33437e5ac03;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34380710227c7245763ddd46d406754d1a887c9ae6d3f807af1e0aae9970cc2eb9377243abdb82dcc98d354a0717dbff344b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff964b37c13cc68d2238332cc0851d879d974bdc69c49c6af00828b483127b94b1863ec39aaff3ad9fa5557a40008f8be98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf05e8be991aa6d78b2a4ae7d375e5a4c0d69797182cbde6c6cfdf343d9eb0e21f90f970fad894a7b3515904dcb6a64de7d70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5371be51a6bb0add4257d7fb31caad57a1c53e3f9601499681edf14052d7f4ae33d5a082b39317b2acdd2f00f59bceda8754;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c1e6373ea98cbed9db898ad32b3c1fa01284575275680fb3c92bdc9e1fd0ba22fa2abce35193e9ceba35c2081ad27b743b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4608bbc1ddfc82a4ed9312255ae37418eb622f060bbe27ea95f3e2d16b79eccbed1e1653d48a849f1266f0989a6884a0235e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea9059c37552a87d76653898c6fbdf65b84d7a4c06a385bf64911ae9167cb29bad07180f8f35771662af96471697dbba4a25;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d6edd086cbf532a1be93f963c887c142c0a83ebec9f83d3cd9cd7974725b8e3902ed631dd337a069f2802509063c5c45f55;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b57864f741efd2a718a0e0ea156b191ffb8aaf1a4939d05816d71eece4e2c0f01dfdec18f8c5fa3c233b773b417fa44e8f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc221e93d1371cb1a4ea19ae68002dd6ad7651c63cd43f624808e3c2248fa4d38467200eaa03969cbf0484305bd79b1fb6069;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5058c83491c70d8e5fb440fb1e1cc5eeb60249aca41d43e85c44caa111def04ce385f46fd3ab72e6492cf0d2993192a45ad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa79996e01b7f50de8543ec25d340c756168e67a51e4bb1c875e590b39626367d7d334258c3e7f6e03a1a51d5f1745aa92e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5de6ffdd40199f6745269f3a01f415e15663f0ef2b45db67e7414f201f888d818e9b1559df35b841b3a4024f0091255b22af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77cfaf599d2c055b464ae5cea67b068cac961d4272bb576cd6f32b7e81aa3d94a2648e04e138eede0ac83be89c406b0c610e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1ae8d1939a8702657272b5e85ad79002ed573afb7987df702cef5b7c4b542834660cb27e1df8301237c49dd8fffb796b6c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0ef7028f1cd4f9be1f97c8075e7b7f94e4daf237ea85913cbf44b17e1626b77e4bea2f5870f7fd28500e7dee769ff45381;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1195756fa80d56b7fbe286aedb0daacb2b04914bb07b3dc96f0f4c298ce0d16aa5a5443e85db7bd4a54806b0ec15dbad1223;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfac07ec2d846c1197bbf8a0f08abbe9560346c4e3f3c4d420a83bc2c4f0c63fbb9b8e2b35e32ccd56e04df22ce61194bdbf9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2380e8a4f71870d84138062f97b351166e87256653b0f06e9e6f8aca2ab74e52b0e945242e1daeabb008cb9bbc9539c0afe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f356b5a5a3ceba176d21fa318fbd7b15214b5c8ee2562034e9e88d8d1dc87487c1f1b8d8b2d85319a187c8bc7580323997e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba66a2f743979cd0d7a40a0aba951849a2ce9300e4a7f3fe8e64a528bb418cce349dbefa763c51bfd34971d2b3f32cbd02c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfb7393a7efc1564997930ce1b2ad70cac27b6a5de15df7cce54933bb2857b06e44a4f072b62052b64da47dba7e1604da4f5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67ad0c747c677b81abc25f0444f00c9089f95c26470626c69d48a0087fa4c74be144b1918b9946448fdf8fe35c548e551a56;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb57b21ed6a0646bef5bb0cad15854a6761bf0bb2d689f5bad878bcbcf53c4cf3bdd37e181d7e20b0440139be25d5b8bef5d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0356e0c8a6bebbc371c8486d0b0033c6329bfebadc626fc701e7363202108c11c3655c7a646aa133994372753ae8d46c25;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc430ed844a562c23b58efb6d3e941a83bdde497d45caf1c3428fe8f51213640cd21e81a093ceb0be9ee011b673b48c50c3b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35990fa2440fa4af0d5bdeb3ddda94dab0c18a9b64f033984565cad95a7b980affd2332aa368742f054d9f999c7a267e88e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80c9fcb27103abb5e6642c0892c86602264db71fb65c78822b3d8943752308996092ddf64eff7aedac4bef1469791e81d11a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7cb0e8d1e2b724a172144dc429733407cf65ce73bb22863804507196dced8592bf17629bcae7871f1f821c806ad6de26b61;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2f8e74eda588c9411cc5bc38ad6520f969e84beb0069d81fde18be6be8050600e56386d9b00f08a5fba3fb95275dd4f7fd3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3cc551a6e5c1f856dd29c3926f9149e14ca9a6b98d3411ae33d08df18eb166b2a3ccc09d48a97adbe6ebb1822f8c48ecdc9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ab73b1c8a3bdcb2f4b89d86d4347ea44f61d0e82aee5c578bc17553a90d99aa56cf5ba79686b1cd5ec8d27d36367fc4cc5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3e6f4ca5d2eac076883dcd2fbdb44612bac79cc2922396082c8bff860d4328ad5cd75789d4aa2d408a44d844a3366c15b2e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d6209bc93b4e368ed4795cb330b46a09ddabef7b8983222a7bd8f57c9130bbcb7d409b6543c1171c8fe65121885abf66479;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5af979734d3045ad299cdc379bc2f52c7652aafa09b76e800c61cbe554ec6e52fcef2a28f0333115365819b90cb378ec408;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bc9a816651e3ead03e27ac525779cd1be0780d52611f28960fff8e59027a0e2de37c946c183c4a1e7fd1002cb0859dd291b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9294267fd6922074f6b8cbe0a2137f1b7941e4839f81005ca987da36583e80d0417efb2387f06141d614cfbafe7e45a9920e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7cf3dedc469031eb0b96038fdd686fa686b0a650d2c442256ade087f3ec2661c1a070d5d120e349c72c09cc889f0d27aa22;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64c4869edd353493aca5e06d2c1678e843bdc5f1ff4cc23f57ee4b6008c3536fa2944a160b2cbb50c3a41d9356f42bb49c10;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3387a36012390547825c0fc845012f487f10be149b8c7ddcbfbd98ba7d71e35a0b5f27550a379e937ed268495a444531e04d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7b5538b16e3988564838a5bf42c27fd1be3c4975676e2928513086e8f92c383a745386f401162c495ac095d2e84a76dcc22;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57245a198b92528668c646049441bdf629a0b063fe45d24a8fee7a21323531fc38a2d100b1a654bdf325b22a610aba48dc42;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h870761dc16207aa1e2582c65797dd5aa01ca01481fe798129eae0b1846564dc650962c04f78d083053779772e3ce06528bba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d1af5ce39e2fa1ec9e12e950bb4dd8a3922f53bc6ee9b5c5f4a957dc15ebd1f87604dc15cbd462c64c93198c3205efd1fbb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha310930f51aa014f09705cc7a096777f31f5f85a9d360c11d3b62e4e8d71486d0ffae323a5c08da6f4266e1a735db9099c43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1dbadcac76d869c6512b587a53ff35aa99d114a2b3d6c6ca2bf5f24b79a3d49642bba388facbf43841de5fdcf4319b473f67;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bc7d42d42125f6583070d3838578129e3cc62032ac12387598be08e052af864ec27bc5d265a25935cb1ac467517b8e91ec1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ae9bac867afc81fe5af2dde1d37c26dc71a7ab85f2bcf40deca3ab32c142b92a71fb42763cf6605d1cc97090fa73bd9b960;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b64f42283de4c8caf89997a5eb21a71150498b9e46282f776dc8c6e758b528c668ad7d4f0c878ae655c8217196957fc4dfd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57e4fbbf2c3f2e24fb99bed98e09e097bc526f5d6cdc80d124c428a34c2c4e2c507a732bb218928a96f378314b432f5db51d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c45919287eb07cdf9a90669f8c61653b4c47a58c6d7c284c1030baac0fc52a920915effb6229dcfba5aa212d74f945521ad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a29cb08473a49f3e286aaea8ce63063c3dab0f3c27c079ee08be05200e54f53750b65a8491b3834280fa04a2c76ef7ef50c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4357ee94dd3311a2119fa5bb09776bb69695aba4ae19a3acb1def5459b39b9d248c7c85045deeaf8cb86a044f00fac2249e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d90a6356b4389f46601ea08334d5d4c0213ad2153d50fe9794816ba1dce5163c0e6100674f168672c8aa9d275edb0eab98f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cfbea86bbebc0c46782a621641cfeaf5a9d7b9a51cf0c9f4eb25a1b6b07e06139a17f2210956e9a9b7416ff691561c194e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b88654bd8194e8b68dda549fbb907cd8248f63c06a82c4c3edb2204e064357419da89440b0252b6f5d62b07b2aa55222757;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10f8ee6bbeb2feea5e5c418cc9a629c27948decc120e6713096b6aebc4b8b089221de5f761037e025eeb4920dc5956a5cf7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c94a7726c167dfb9c0032928eb2fa8ddd43b29711dafd8faf223603f7f889b27b8c03395b30803a9b1de9c887c95d04de89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h653ac2aeba294f2455cbe873a0ddc396b8e52a6950bf7c2a0d84c6c70a89227cd7a47a1ff513b036575883700b865e3e04;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4fca989e86e7dea2581c52dec3388fe03b2dd36e7993f89ce18f3399cca52b421fb6638a6e21bc5669b29968fd1fecbae283;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7ac0f545db1cd00003f80866cdd7d29f29011c73cf973a1d286d0d915e7704f1090eb0efcda8ae31291440f7ae8955bf622;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafbf74872ffadf92b28a3d29c344d333889302fc1b1b747fc857ab9b59c3e98a9d20627d93511d276313361762f08959af74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a50c9cbe293daa15d027d84e324ca6ac6dd635c1df844ed472c8cbd5a3d3548f0ff3ab7d8a9dc9e9d5a1bd999244585c9e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1193d952934681808bc79ed35293a1138611f288693473a610f6c515f274ea658535be3cb351007c5bcaed398ec94b02195;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ea17fe62b4a5a7c28f76b6155eb36670eacb4c20b6c310a749ec907fb430861d5a5f2d440b9654bb7cdbcc814d837bb307;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce0c1215f51cd4595cb817266e24223898340c02d5d0940e13adea4c53deed1d0b8ae4431bf23b4373e62264cd67b792544f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4cc7270a76148fe9fe1ea842e793d714ce6c75b959413498e9150db034b26e49e332b87744c6c416fa0accba2f36bb7c4f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc799c223577010ff8d94c1db4b1ded20e38575b529bf464c38a02a1fb815ef779f049f827616982030beb104a4c73df90f98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d7f509451bc46f703be0428539ffb55f74da652811735775622c65f4708fc05494ff65c14292525fa08b468113e0cd88039;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb48898a3d869a0a1e493826caf759ab8c701c27b2933b6935251acd8d4f52813400c9d0b0dd9f244b9a875533a585373746;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h492aec4c6ab9e568184be2ff93a7f4862ca342df4e2343dde468c5dbe7d99c58f8bfd3789b69b24bdf09c6fa8582d3e4d420;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95fb9ce1b3e465af87e7c7a5a2b363672473f3b15071e9cb79e277d2a9f69b0249de3e0cf2903533d26e87191f30009878ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3708889aa06ccca94a478faec920d2a32312ffb4ec56d962d35085c2af0c8e8413da1a05f140f4d79e787f349a686f60412a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70caa871897002ba38ea9ec5a42f0bb2e3c5c467d662736b25394c115694ccd8ffd56e7d58dd362ce87b861dc6d908c4a65d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc69e01d57f69d6a7b4b7487af4aa276e97b5cd9ad6e7b9aadaf204d09b46c2e2281911b2405977e8417160e6c2efd2f181b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h703df3b0d6962d2ab5f32135bf48d8fe156d942ef1d04f4bf39db7afce9dd092032d0c28f7419bc57723b3ead2feda0a9152;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8595bbdc62678090502784f9e08fd3ee605745095f53ae7fddf785ca2df99f8e3e3d71e2416ce0bc3717ab225f229da67d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70f711a1aab3e781d687aa0e43a787bfad50ff0ac91e8eb036edc0ef01bf881b746ec3d96473b01ccbe129cc9ace80d03a3a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc31dca6a68ac6fa67b71e3f7f2025c3a97539eac5fcceb8d3f0c8a5cf3c5e38fa64b1c9ce49f95a9702c095c1c33fbb5d7cc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6411c02ee0c575776842b380d5350f36a82f71547f429946df23344d05b09b97277c6488cb39eb6eb5403b747512c97aee4b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65fad1bf347bd569e6096f9a36a3ff45501c80fd508e9e909daceae879174b68040e2857a8370c89736bb9605599be4720ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41f9c34589f981fbeff2fef1225b467421ccc2787bb91aaba9a7f72e719e0975b0a856e5109c6d6742f253debd475ccf186b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6821903b3e8870e2de37f464fca7ffa7bb9cd832c9bedd32d2509784b201dc01b76c3e260a2f2c4d5cce6ac1e38e59e1280c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1c6dddcfbb7b0dabf08e1e9324b04660c02c7ff76747718337db9e4e259781573ced6b2e61eb28277d428fd90b90c0a93f1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe506b89b6cc78841fdfa7fc749f60c9d4bdf18f48418f501855758d3c485b5981cfafc94746b7367e2ca459f17618c5f357;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h703b5c67d61778fc8352dbd6e44305dffc98eb9740d777b88469ee354555eca8466789a8b70a7a2c0cefc7e97c76c4be4e6d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4872ffaecc226ead831ad6da7620e8a0aa940412e047344217c8dd393a125a83b429b0341008263653dc7fdec62c4341399;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7599031caaaee605f311af6ef2d906ba2196df1b6f3019bcd6f9dd335edf3ca2356969dc741c032a2b8e6c6971d98a046cba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e6a4b9abaaf8d64d8dfb671c56e7d67747b255d568954518e1c8e508d6dcb94b7b6ef94c15c120d728c3401b48d9768be7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha67842b58a9ae6576c241847284095a398d1dc8a9b7384f01e322479e7f0c3b97c2532e47928c2675f23e755a6966f382cc9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f7be49e571b9e3b9fb7b83c5bd25d4ec3796884c0758a76aa882eaca064fdfd72a3613282ea74f6618af0f3a69c7885f9a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he58c45e03e983522c17271b91cdee00444bcfb40e6d0fe2e5e6cc8878b10bd995a8e99f2faabf05a09dfeacc9727412b28bf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f9434dd9db5e4eff009461618d99143a0d486262636d4e11bd74924803d100a249fb82238f996f66526078f1e5e363efeac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h319a0d6f274a122fbf54e74eb08950920ecbfa0b54498f4ffe8aefdefb9f2e48f7bc8066b553198a6d39ea02212f37178f51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h365c71dbd180d8f70a3d64513a7789f15490b464bb891021e6b13be0ae6808b79f9a5e3bfa8a299dc97ededc7fcb1b54dc74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd84937535d680c141e6be6b389cb38fdd169836f8d8cb6b63fb749aa5fc5def82e252ed2615da5a328397a5fbc909ce8454d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e5ba8150eca32cbcb5cfb5fb0e972b45fecf207f7636e83009d5595960469923be8dce56640eebde521c3d1a083775e110a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h343bf75a9e3cbd28e03d4985a92b3298ea40c30b340d653d3e6d662b7f7f49257889ff178b2acc7f900c9d20dea0c32304d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h328e86d4f2c11fb7a519aa3718ffe9c8e080b5379ef67942a2e2e839bebf688bfa4562563ba20ed1a9401418ca5450befb54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h570dc2d86f00a84e1c1aaf7d815fa24eaaf851d6d849390ea8b56e19c6f089301ad78cfccd84174f0b4e683c5c99c3f6adb7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h329da0149ddd969f3bb3e024df46e6f09d4d966ab63968e1889ffd755b736694ff288adaea05bf1185e0be4fcb90f615d907;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bc317afcb101f37ee1cce8bd9432fbdbaabd8bd5f94194386d7dc7668375ad03915460a77042b6d346c06b066054edcf8c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13002a74abe91fc6908e2f77d74f5699e0b07afe4004109e88b716ea6ee183eeae514be23aa6c60a7f7dfb3e9c5d1c6a4086;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7bcfac8fc9fd0373d2e16dabb3dff8e2bc928f26e28e5b47ad67f23c8fd2e7f3ce42f0fa16f7f257d4197dbdb0c47e596a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8ee6ae4446e6e1fc4a6a4c4431e830e0284088dafbc9b61235e0e1727e709ae6cd2761d55fc3507639be56051d5cb09776b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2eb7ad613ff99c773b3613fab89509b8e7372ed2bfbe6d451b84c4b82c321d821de962c9a1bd1e0205dc8f0d4a40e23c5b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb881c0c69f71f375ae43ef0b3c8eaabfde3618d1bfc0de43392d093cbe8687ea6d1030136de3d3ae88ad514df5f700ca4b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7479350b687683ae16717ab8f07383eb776443ebe4b3a2d10cab8dee139ce37eea8084370514cb2837eaad95ed8068cc527;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ad659b0494b108af6687b266719f9b7135c4e74ecaf1a30da7d10ef7177e2b393bd0632378d29bdbf94ab7906ebcbb1387;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h197c6aa8d88491df57a0b1a83f2768cb485329050c2cde57c6f845a90d45a3b8fd32d5f6db03e0412ec25e71d318df438cf5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf14b6a333672e626e6b2d4d9013f827077b416fe04873cd6732b7d87e62aff48c232eb1b71d593e19d953d62c748579ec6a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb881305f762e600dfb8e3637d21ea4b681cfa54053765e0b3568fa7146b763396c122a3baf18235bffc9a907a23991cfab3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89c93b73ab8d106cc27ef294f33d7cf2c420e5d6a3d430cf810471b3553fd2948e6f8ef7d72ef1ae4b3874d3e63689b916fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee88da6136a2b76a093ddd37f3d42165808c3295423c6cf9cc3f70f4ac3463a74ece09dcbfceab41e7c044e8f2d9d9d53097;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24478c2757630fb8d9afd81c953ee9844d0b7dd5830b6902f63c875bc28442e4f5ecd1b47dcbb3bb53448321557b493d55c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbb2ffd4231e0c2926eaf182b4807f76e3db66a3a699433902daf2c3bdba3c7cd1ed5b9b5f70b0ec7ee4abecb96da8635062;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdca07461f103341f843040e60284e9ba571a89e96425947283094931dca1fcc82edbc719f1434bb3e62ee5842b766d6c9665;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf97feb1d83505769d552093a09042e486f78b1d465346214121b94d817419ad24e06b41f6048285d1e7df2c115f27d04033;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda6e42fd801bc51d20cf4279e80d46dfd1731b86c12c19c329b90ae6f2ed2de6497bcdb8e1a65becdfb9fa4e1db99644cf97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94beb40a99f656335d9cb3627b533622bd57a03c147311008bb1e07d1f31d8c365c8eb1b6940c85e91fb78f98a885eab53ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea1cadcf29cec0c716e14b137cd6e556148b744ce9f7724c5a7d2e3bdd51effbba7d7b71b6705495ee403a7318d92d839b06;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b65ea173031cf0b37bc1495f99e346038d4accc33b17692bfd2e1bda2e00e9b786fd667211e1d3fc24ac25d72a46a18580d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2e09c0a97e05a9029305f216125bc916ccd42da519f466653282e5b25812db442906f12b5f1e2b05061ec994809588add43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cf7fa7d8af87548dde45cb9c87c8d632ac701213a5fb57ff3d8168989d00afee4557eb4f093a32632d12233facc50d1bd91;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7795e9554c94a8c10824eb0df86630b334d6f08bdce036daa0fd151f735f2b42644fce7642a7355ee12dd691d7a616744a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed6794d028b573a4e26ab79a27fbf6d818c69fdc9af3c8043caf8fcd3bb701e365e58e3eee22c9fb1207ba5de41684fd4340;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c174e10764aeb414ac7b426e75a633feea3cd91810483cfd68dfcb7a9b2a37b0ffd183f29b14eada5815644f0034307712;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h303c9f0c55fbc3b68a1b0f6d31226894521ab547a2e05d5d9afc4168dc048c222d4d4b62e25892c70fbbc81cfc8e8f6ae65f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc84756135ae8d4a5874413f7cd943fe38873b568113cdb7a8aa26565f95470c59576be25c1877620dda5acd0b4215bdaa0a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae18bd68fa3052446b7d863768c429ebd21978bd2aff1a2c3f573d6464d1ae9b8bd58e98b472dccc1a0b1905fdd1855c0515;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3921f78c57469728bf5cc81272815934d2fa2bfb7226a57e60f24fe0336011bfe8fc53761add087af7e4ab6093dcdc6d103;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cc8aca9d56494373d794881da79a03a010843fcfa82fed68e21b425177eeea6042ccaeb4e937631a8b7c799a443dadfc042;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6bb158fee882114573949d200f4405ab129c7a0819c81433c9b6214546152f0fcccdc427dacc3756baa4baf78e6be85274e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h128d045215c3c68e26a385af087742d3f8e6baa6b917943c357b97949b3cbb8bfb0dc7f841afe069605c94c8d2e44a7e5e6c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b740a411b7dbc6f81d9b159a26817b7b49ee2d1ae057f7235839def13486b92868d267ba6931c7684e3ab7b9d7fb13cb998;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb54a2556395b2dabc53047a47a247fb33891f9582df510c188b5c81b75d9fb43190c6b2b975349ff5d8223204fa42a2c5079;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd125c31323e50b1f0be29f6ee3d389cb9b79ae01ea097068b804bb972e72bbdcd595c5e6fa73684d6b7f42cf7b284c19dd1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7935fbe8a59b5c8f1fd982ef3fece9084e0a72c6a448b113b85107198e8c601e79ef62e9ad55f618276da0865d1d7300fce1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cf0cc6bdd18b05d611bcb475a67af49b0118963bfe688a74dee467ea816ecbd3ab0ff00470a0ccb72dd1e7e9cb282bf0e8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f65748984695e2b0bb2c07ea41adce3bcaa2ea27cf6089b40be7658d556e96eadbd1195137c44a3c46b6d0fbaee941c96c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce7a822c74cf95aeabccc3041f5e106af1a4aafe024ed57b1bf89044c9f672e389ec8289a95310b9da54d609b5a70bc00b8e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26c5f95f11081b348b9b5f2699a15f309725e5f335a928bd3c28ae971344e0926a9fe93c26a0d812bbf837b815109872b0ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h956db1d3c61c2be40498c6b7fe6483f11eea84243cbd19586042c47bcd6f704c0dfdd80896aac49bae38b768c2dd6baea596;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc93216769cd52de5172c6824862d149ce9287540c2a838bed047a08229217376687e4e65b64ba5589704463f58eb9993e2f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e63ca14d7aabbf580fc1ce8495de67f65b00f031ac54116ec4983a4edc9bd602dc90660c91fa2cd2be47d6c56f9457034b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9929ea0cf10831da61a86573c0abb2d177b645487ab04bf1dc1b897db72c17cbbce9286a8b2962a6a821bc6d484f0702085f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4cb44f8dcc819f0fe6413d798592bfef37c3d7c5450312abcd7c12e8b8e6f8931dad8af0f8875430eb7ec922343c0bc89a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88ab86206a4a37ee8b2f78b54392705556a9c50ad7819d3a591c56f0cfe5d6c2c111e2f62979ee3f4ecbeb270efd0bccbae1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6285057006643f1ff955fe9e0cb0fe02747ad2e8da053a5bcaca99d0211201694aca76ca10bf281fac788b63d88b08aabd56;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadffec93992d53de5f86e6e2328ab59450edd06b3fe0203321f8b21fd25668005a5e0625def2a7b1feaff704f728c811da97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h253540fe2e55eec65668f418831ac5b57a643be5f2a66b4d45c5dbe91c636b4f84c21bbce82c69174a9af621dbf0e811fcf0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h232a94f81fd22b5a8cf1cab0f30a1f2c5fa1199c5dd0108d566b87fc64416ac456bd463225c56977497e66dc62aa8596973e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1cb0d0a6485b28d3ee44f7b9921a3acbd2c9b2e22fb8c997ff5a51f91a9ec0fae840394ffab090221b06570934be855323e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5e3d240ca9e5fdaf72c1a6874b9e4842e018e05db4f15ad4ff50272b395464d1b3b10f207f26f4f4663815db931d8dbe577;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8894649f1efcb0f0cdee45a7cab6439343b4353eeaf85a48060eb1e513fa64bdeb24ee3066e40a58395f804ab9d73852941b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed7dbae9b50ff394babb82760b74946132886fb0da08e8f9111a493e7cf04fd0ae192dfa6b4403310ab6eb1d8ac52b8b9697;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38562e545ab70dcedb81b67617f1363f361f947cf21117a46a5e160b6038f21d05e77b32a39d8c9c93be8821f91203f5b0d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40804b198273ba31076e5298bcbdbc8467931248fa858ed945b28df9729e6a91c448fcfa46097b8f393ca5a3ef13e1617c89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8ab537dc49f342a37faebeea363e1754923f915725cde60b2b14b73e7772f293cd288fd17ff9ec8b0cd9cec029380fb78d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb570f7700630cd88a57955fc712ab098b1e895af7a1c08f37c30e8d776c00b44ebee898db3ce95e3fa46deb17fcac04d0bd7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a2e0563658d9cc403855e0960792b868235290695d5d6b516b18719a9b3d322db22fb3532855ef445361970f6db18a9372d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb474f8b2dab79701408013b69052dc5ba68f170dfbb00c7f800e046cf849131a9cdb11582acb86e1da6c413ba92a3f67db9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8bb75649e3a3b18bee9109fea6d981ef6a35b5d3e79516d1aec29cce269720aeef3df4291f2e3deadc47161c44b05009a4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cf2ae8db7848c10df26b5a6b3446ee0ef9fed0a4494d299e545a288cf15979ec2bcc242856654b70318e76baf4751c8f09f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52576f72f8dfd999606f2e6d661118caf5d44f67da0f6a98aa4e1d572d55ea5b07361c2f5a8eebb1c60b05b6cfcd6333b0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h777c5086fe61eade1ceec340be035edf90442631937b20e7a0a77ba63fe2a6df6e2bfcbd55750cdc8d3938aad4f01bd1e881;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66b00cda7445bdad4647b0cd61fab48d8b61bab0fb58ac582b404099ed39ee49347f7b00ae19809ddcd8311b46df979af17a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h556bf7e269e5964cee7442cb904b5c4b0c80a890846764f5040e3b169530967e201266d5ba012988fd4a63bfcb09dba0c1e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e0311a2e495858cf65ee2e1c9c952db38623b992670e688ac052c23a2d47d0e167c2e42d6c2f2ecc3e8c8b02832774af5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a3ca4880eecf6995d9789aa6c1ce2e6da58dcffbe226baf2325c0e510a96aeee883a0baa72582d7cca8dfa1a9192340fc48;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6831000ce5b5fcfeb973527275481153e828607ae8adfbd578c9323baab540b1415d7f5e01accbb09cbd49f2242a0e8cc5bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a64d065f0be262abc768db686c24d58ec5a1a64bd8d226d41c9b06986ec7dacde43a1e7ebb64e605e2752a9edfbc061bf97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99c9342bfe3dd676a5cf35cac6fa4aa45f2599f6e54d8b1bb7d30a06f8640ed7d80bfabebff80d1d9162236f0173aa207ced;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28fd8845de6ce81cab285a0d9b7d31265c59faf573816ee301239e721fd1a809a64c9ec6b88976bd71cebbb97a3a60028014;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1d4d96971826e101a66484fef49517c597caff3828b16ea3a09ec1fac92cba7bd3cae1f43c1343460ad8aaab6e0af677962;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h593bd18a9de5e96e93e29107e46579e7241e8474ed01dbd714fba0fe0ee97301bd0eaaa527d4b3b02518a770ee363987f2af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99edca72279c8c37c07d39f889b59593ba17d59b7c4b02b63a3ba01579f3016b62b4b8c2838cd472d8d7758df7ebf0db5e51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h804009b115a437058d52d923d497185c793ed1b7b128c8ffd5ead08e24bb57b9d2b1730b7266b8a5ddb16a5b6c24259bd013;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecd93f3d0a753af0a453d1a4824e3bf7aab4051199a09d3d781d2a712198410db58e774c4d4e320d92c8d49d1b03b596a6fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3886a732973c0c5ce73e1be89d310108aa256853d58a9a541fc3402c8b1cbef60367d70a440a518570ffbea49144160ef0da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha054276d26fb5419d2405a47a66da643bbff4403d46aa1913cf50fc7be1a4758b64b5b0a176bd74825eadda83ba9cf9020b1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd598013e92a2cf3b0ce6952ad8e3bbac7ad8254f541f2da621eadcff727b6200db83895ea40b25a2ded4011cc997c96e05a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha87f988c238f8dc69cb267c210bcfc4e3f8db0e376f48670297f8bda994fc41b8b78eb38007a8dd58a945444075092a4a58d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h730c088657aee25a323f90f3648bc4526b3aba43bc78c5e0479bde42b0e644a2b57a63a967f7fbe648123064ecdf010cdd7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb27d1a1c3c28bb343b667f60ca8eb4a77b5b0bbd28198c44bed65cb5552e26ad7c9ce9ce00adda720e63bbe4ace9c658b4f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff2cc2dc3b569e136cb515b5bf4eb8558d52ab1cf2e6a2c1cec39f57a1f51c2387e30de03575181cbab71251dde0e6f4ed64;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc856da9c8bc33e1a41386435ce7da594f1dcc459d4d968c52e88f11964cf88f9a81277d31c7ccfd8f7eeb34ef83bd290a823;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3174a2486bacd264afed15232ab717f9b506f684d17e4271e3e05abd0133b532af4f6f09f6f0cbf8ebe5a92c128609895dc2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d426b4d1602f53eaeb43c68b9b229503c708493cc02de0bf9008cf67c6d96a4a307a131a88f1b3748f51f2b37aaebcdae32;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3f6113a122287526a01595cc48ec02029e1f5a7139d2133f1219aafb114707787e58391c3b11ddbec8ad26ca7df34743fd9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e524c6198e47925f8651e0fb8c43e7cf3a6b70d7d525f61d827db2d89b27a5f5059864b199294a219290f038f809edbfdd9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca14c7676cde7082f93cd9fa78776368625393796d9426569f32ca05f387cd8b2376ee6a200a35525cb0af2bec6fdbab574f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49667fd76e8a668d0723577bfe65fb3082648ceca25d1ad20423aee0ad4b6a703c394c6f8c66a38df20f0fff51cbef0660fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefa789e37f3bec21b95618eab5dcc82db523b9dcb31d58848d7e029311d7381f814a86975a5fec69f24bf7240e970d1b741;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c6965494e1fa5f290113f60d756e362f0c0c51e94e31ae210826f9e1dc90f16984ac8540885dc701b92c17b911deca9c590;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26c27253d05076417d9330b56c3a2489cf267ef768c7c745f362ecc88c9d6ba5dce691855661036590407707c1ad947aa929;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3554c42510f23746e08cbf832677d435c2967779873c2a4496a4afed878baeedb54e27180ca930a4bd87b31023611e43cb43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h826fc60f72c750b1e2e47aebb047f4cca7101c6d2ceca1b86a222cd4ae44054d519f5235cc0e1ef58c99ba80e44018265144;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b080be76e45af630d0d8e031b7a31da1b1058170568eed6cca3638a35fdf18042c35688825b58fffa7281be9e77ac2c8f51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3cdfa472d67fd0d22f2575cc61d3cb9725882bc90ff3495a36a2b5d5078eb54b35026056f3b0efeb5f1331c89ab0bab00fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hade6823a3b838cfc56c42b2126b07102594afc0f5fa701de3c26a71d726562287fa3168b56cac9452f437802ac33a745e7ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8d53629b1a21ac32d722ba9ed96386e2c529c8f5e8b1b8a256b17ca0d6acfac473a31d94b152b028a5731f86fdd15faea51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5afa70d4e611250651c82beea65fdefbe838f7764ed596ec7236e74bbd394277d48e45c8e15809665eb62a18bae4198f793b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6303348ae58836259ce80daf0b2deb324b56515ab7d9758d42cbca1f924dbba7b1a0f17cea421825b155e37f614603446918;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ac8f246118764207fc45533e775d0610e636920cfd47222be96b0d82d8e5d44410e33665beff0ad4c2818cac13d456ee508;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h513464e684a720116a1610949199bc7b9f384782fafe395b364c32d7e9c3e26ebc74846effcfa6f5699e15030ea5f24369ab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84a621aafd8de7ca7d8b3ca78142e627ea340357be5100500ab8188a75ea66275096f83aad1041db9ecf114e78030f499a99;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he80379bfd8df4e54cd3c95abc5766caa51a4433d6f76d7449958c8b3e81cb02065de210d46091816da3ebe2d3222469f1b1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he02a69e1def4670928bd1e80f19b33d36943f2a30eda25ba87e52d04033dcff4602b165b5fee4c09ac6610684c8636faa409;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe8b441671f31f877f25a6141eedccc78952fc70edf75743e36eaa702371efca511a5989c1862de8c6a17abf07fd775abeeb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b609019dd113760cde436a99572939d9d0cff6ca40c5069f96f23de93c994ba8a8064c2612bd8f946bd65cf53d5849f05b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa1ee0a4eb0509eee0f917826e4eace5e5a515e6a4821f12f4a17993aafea2bc8f618bd6428945d8f342224ee909d56467d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe2d05cf31f332b89456a6d3b9783fa93755ad4bfaf63028c6afbb8d3a035e6f66644cd4f753fcfda8e3f978c05e4c30e065;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9832c361b88a738d0a0b582aecffc448da45855b2461f66d34ad28b3bc1db408e8678e94c47175f81ac6a429b8061fa02c34;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7c350ae0649b4cee96a1150baf321c3364ab0a5c0ee3506393ead75f3816a9c10d3aab7ba33f311ee5517420c9e475dc934;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h928277e45f2ffe0b13faab5bdd7381f7b3db273d93d032456b5fce3b9d1562f0f93c25c8645eb2bdf94f7d8c77ea3677b49;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f34593f6206894bb4f5b33b97b440fc7e387e0a44aa70dd98d56269ef1f183875f68ef00370f1d5e3bd20d2863ee9df4918;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e813bcfff640bcf512fa2f15178c8fe3c0953ab3447e571c7c05d765b6b13d7bc5419143ae4c84de9584776b4a6cd8b7d46;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39786c009757aeee3d20b2c6a1d926ae0b27cdf9633c1a8e46af90263b5549e3f660c81ec25ff2532d3570b2988ad9cbacb5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ab1454e386c99e69cecc7a8a2a3d188802058f5b860ec1198307ec66db6a3ab9ecb481f9bfbd26eb4dd7a7d2198bdd665e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51b5603c8079645e94e0049f79124a10f7adb702b966057c50b2fc441f3ceb389ea794bcdef38306e7767a18a9369127dbb8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a115d3a2a29450bb6ce3aabb9eb1c1074d6f9ea065fe5f0ec5ceba16c4ce0b56c36cbf231fce4d97b924dd812e6a1f8fc06;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98ef742603170770e9e0a795c598ebf8471edd223c1eb71cdde330074858a9903a79bbb73df9e15f514c674319b2a2c6507a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a07b9e7e47e78ead8732c2c4d32a1a0eebb950493020d24fb128167817b4c123e180ed33e876031f1beaad8a1dd8616992d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f56a5026166c048bc3c1cd1d329ce2da745c4ab8b6dd27c2ce7bfaf030e9eab804975bbe9814b60f8c08fd6e03ba63e368e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd36afb91b686c3bcd21724f526f8a6a3def43cfacc69249d5d09f24f5ddeda86ea82f6afbc905faca2c86cf596903e9246c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd4f58e463beb51cdbf1f69752679dba5cd81fcd25f27386777a02a21e8d6adea9626f27b3072a8c1616f675b3ee414f2ec0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0d1cf1f03680ecabb893bed08d8675a8718a3f38076fdb27dae487918ae3d1a5a461a6e50c54700229025f798a5e604029a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98e29bca032bc5b67718251208b8943206a602bd157a32fb8e1b69022b5960ce8fb9c2897b9c9794f80cd758e7482466dd0e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf62a4af1ef6ae7513ec4065cd5b8ab73686dc929476e0ef20d435e9e00ea42cf45e087cd723df8675ffcad8cc34da4d110c3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e4c0125fee0ad2705e91c6aa1eb5487edc4f2181fb169120cbdb58f153b7ccb3d07d6722fc926de72f08a1a2e4ba0bd9bfb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18023e4ea49c2b1878fc2fbeaa24980e323756cb6d471c08a18e6812b1c095c1fe3739a7f74546e0b13a6b92820b52276513;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3084a6820d7bba1e20a8f2b21fe371900a233f5e202237b99e4daf9f62e44cd6be080b9f12aeba4397b7a421c580dc7b53aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8529934de2f0bfb80367b69c87db30718c87a208ba64b3cfeb559449e3208f0c9eb26dedcbf83bcf73ef52bd5616f5780f5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1bb1dab6835c276d0f10e5a0312dfb4ebfc650510a5d7ec0afdfcd0d42331408a42da4887b8344d38a3896d39e438a40f18;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd9c799a8f395f6faa290783921b58080914fb60f9d110013dd4b8be7d30ee3e998fd4aac0b71989fbb7a9cff1d2df5e561b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cb3382d4159c859a492c724f1ecef4972141d4c55db387caf30d52b8280c010b4559adff6f21b6a63fb3195cb50a62747c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa94a1ce2bb80663b650c41a04b5df3399292160e5b6f88af7b22effae3d94a24818b1e3226a8a152bc220c02568eac18be5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ba997cc6750f9794bc8815927c9e22a578d9e15a15ab6accfc45f184ce083667edaec843ab9cd7ea4ea8ffcf11a322e3ac7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1907b4319d7a400770ee1f66841f255ff825ae3140446da5b23d347b752758ef3495e26d2bd662d40cce1ab0165459fe10d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h125a3644e9967fdd7b8d7c4efbd2eff48aa3afe89ee5e6caba65d700e4b1764fb1eb2370e24ddb0eb2b16d047a9c86aa03a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefae785bc020da1871a51be82bf9008968b8ea843d1d901e1f4b89c38463762de94c9c2b4e855c600f4fb82f28de038a1fb0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb3e86c3c854f13b59f1f4a3ad3af3076e371dc94c4ce92eb6f3611b25364f6ad59bbb5c8f888ad2ae3eb3341e04702bbdb4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbab41788078eeeeee577aea96db21d41d4ed62b4e0e400ff9452f2598b1ad171559131ec52e02c9eeca5901a3005f55edc6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb09ae0936bbe2035d071fdef7b976ce83f050057049507d9e6d0dec68282f1c9397905bf173f48e9fed58c0f1afbabb4f97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15fe889105615096edc230a49d8d087377c55128e7523ca182333b3d72bf7aa9609a2db6d9a42d0f56347140d10b96f9e653;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ca6a9160252eb34ff62e02faa8d69b23b467448863687ab853976f2b9dda9099278533156844e15e59c277f027667739b85;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a2dcb77173c685d6b328e5f4513f6d55986c92676f828a1353ca4e24d5ad0b9445a926c00cb8427077784a55f169e4d6eac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h495e1c07e972b4af13b08f1bcd0e819763a1f2e420de538559bc6f105fbf85950377d0ca28d0d3b6380f821e3895a07b1885;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80ffbc369cabb5b1a0845ea4b8edee3f6d97e2b0d01e60d22bd66fe5e83a42506f47ebb81060db12bc3e876e2096ddc927f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d167cd7e2d9339f8cc3bb2cc5dcd1934a7608f48d9ec9aba0f8b58d6b61cbbd8ab39c8d547fdedf4deb8a7eba571ea9e2e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h286f4911772aeaaf93937fe314c1483f1282aa72e1d330b41a901f4dfe0169769b2d3ed1fae5117a7b5d733d3653de0494ac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25ebd7260d583dc204c591923a326525133017be4e6c40c0aea38eee53bb1fbf52eed537c4f99de0008d4ff9f6ec53a2455f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71871fcbbff3da16ace21f10fadcfc335364f730061eceb518e6d55d1e0c15f40bbe579e82bc9b9ddb5597b66feee5576e56;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c5e718b3bc33291b7c47ccd0dabf581eb54eeafef7b25b3dc77a4825da2ae7aca3e49168df7399f05cee8983e0f133c963a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68e933088084e237755a032b2bc1925d0a8613e3f07064a0c51e29f97fba880b9d286411669ef3609207271e2a9d3f443cdd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h552621a734632c3ac13ae13c539dafb3b23337c28aa0b8e31d674e437483bbdc7ada9d298d5dbf8ba98e9a44cd5aed3da809;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e45afa3fa1688bf9f52033eab3c52f739be83b4c0e6725a7cf08a0b6a8df379d2e895710e74e1b6d7ab32929e0ed20e6e41;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b37d250bc9480ce3a0d5b3a644c1f87fc27f16388a4c6d87606f0ac22e7e0c4210508994aabddc734984f0e696d390850da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4841ce3eea31ff35ed7efdfcb1da8252e8feca3dc075768581c3bcc0d6f812d5d0c9c658f5423eedce98e312d774e10f21f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17d4d3d6abe6e6658e0376e4721515d9818b47d3642b284ae032872c77391304966610e046a3a192031341cffc5c2fc05695;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3484778ea574caa212010f27590351287f0cb965de2a4a2637c179a0c36b20eea96b086c982819d3341f7a851168b37160a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3805f9d607e3b52e8bcedb66394ade98ddc734e28d230861776bc07306b9d83ac737731a1cc59d92bfd749e8ba7a3d217953;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heedf43d7772b056550a12c1badab46db77dc33b4d822f965324547afc26e806c26c9958c2ac29c4bde471868797a69ad8d07;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h917426753e7e1bdedb423d20d1346251f976dcefeef6543d18ef07f11890abc4252790bc53a358fd80e4dec3fbd6fc5d9646;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cdd8df175db52a5ba53650993bdc7be0ab3440480bc7cedfd294527deb30524200ec075eea8262da5bec4e97eccb3613f0e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1454c71945e593d6df1d1569bed4a84e95145604c587c51acdfa8cbc10f1fb27e6ec5045dc043cdbe34ddbca528fe1bd25bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h808e97d481bd12670324c956d0477f6838a54232a83e6dc580eba9ab73afa0c62dea5fec0b10780463da8608cd0dcfd48fa2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd01d07236bff75d968bc6514b1dfea0eb9ef459fd64cbaffead636e438560c6f52b095795bfa1566f02da220bda85badd935;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3149b13907f438ec7198c9aaecf268cf5c4de18304992bb4f10f05503c5ac0e4a2c02c784a2bd02fa9ec0ff54109c82a1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd205a2ce370b28fc7c1aeb00e5fb10dd0a751f3e6767c5290c6665e818a5b90d18a502396d442875c1b6ee866b04f10140f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb247e06e2dc7aa7f7f4aabd338823038855f83f56dc347faffb02d979cb5d003cc0e6b14d4a0240136578fe1fcae9ea482b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12b43dcead59328519c52f0b8b4d03422349e44ee4127607b01a0537e828112a3747d8278b5c0f75d7391eb89fa76644b709;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1ee41cda660ed7d68c45ed87b995cd4520edff85a85738767d665eaf33dffdaaaed168c1b31e2428372b06d5caad64768ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf95c56b0f9604b1ea7f66c2eeac8ed3a0d4dcb780ad7c353708488b726855803c98b4415dd0333770108598b8a547f40b1d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha913d1494c6c57cdf22c9ed58d0a472e49aa6ecee3e2b6a4c28f72c4302490c908b073d7ba8c811648fd12afbc5f47607fd5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h819cb6e07dd84287e3cde4813b5921f67315b5dda87b3d23d9959204b5b99e406686e91ca6ebb8ce4bacaf259ddc0ca409b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2101fab144e601fcb46300254c63a210eb94d87e040c9d427ef5cbcde740ef471e0492c9c0cda5687e00054e1ed6101c59a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8becf5c67f9bf4e960d7f11ead67b207afcbd86ad45161aef0a45a202678ace9fcdae365d11a6f771ecb86a7740bdefcd75;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc35deb5141571dbb63560c0009cee950300b4ca7fa0f9fa0025a542c798880fe43dec7180b3d34220101e9504285c8a8cf3b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0fc5808857ead78508cffe9ccc7ecd134ba6a78aac9dee9ee880863c733c5031afa2c1a1f49d73357f50ae487152b99530f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c77891caf48bec28dd2748f6fe488dab2f1ae8b05620bbf3f83ef7910c9a9a0c95ea54b518063717e4bf2728c99c0209d71;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5817bab9eab7a921f3153d67f942fd18a1dfa9fb5f0275fd148b5a5ce81b5585ece166a0ac3e459c9a0bd91e5301610a10db;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h834df2cd2ed85353460ba236251fad41c82d156cf6395410e416048bf1b90a3720ccc3f386e62ac1ad34b4962a099bd37010;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15988c2c8153a44d30ca2c750d9bea3b1c899535e496cd99aae208c87f82bed1cd8d373018efb2c3a6f66b58438a9b7bb3ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23b00c3c5bd3f6884e2bc103ae44bc2261d4a7e5f8bfb6c5e779fa8bcac357c2e4b8825bb298df1aae617b4cce38a0261172;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69e1c588fae022d8c212d23aa9eff0ab698d86ade5162de0ece8e89546af50fe9ce63d43683b462fab57e708c2a9aa0bd691;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1db27034e5677725276ce51169a01c90f2e4d2fa00b7ea85c7f62704a4487b0cbc4ce48927d3c3467b27aca48fbb9cb78a6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67491cf14aba2868841fe676d358bf373e2c3d0043e9e2bad46160fc1b3e6d55beb043ea3d99c42f45c11689333639382707;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71efe21c210e1ab45a156de3d91915fbea9a532f0cd26c8075f79564f871c195c4d34ac6c40f75ad6e0781b32fa62413b591;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff1866a3e754fcf75e3f5cca871ae9e08f325d4e8847b320ea0b540d2ebb76db953f0edb31ddb02e383afcf4d101c2356726;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecb0c337b5f21eb039e0623c6db641c1a9f13524618357ab24e40e11e8aaaa8e856e37511e4b572a7e724306abd631ce44e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbce649b41842d0a4cf2d269eb3280b724505f7320ff0737e989bde951b7961f2a539656771abd6de8f4e243d175d944dccfe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38e05060aab7a2350a0a659e22a54d55aecbd26038491d0275ee296c8f3a288af803315e76a88e1bde20eaeb846b06d507e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb113fbd2e77f15524a8dcc944ca7fa5e60b6d1a7f6e9f7f60b180e343b218b327d75bb016f507b101cb2786c7198d7beff37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he919df04a2ac3e0704feb493c3de2c15b2f70b9d4370973e066ef0a02f4c9770f9f0e4719954bf46eedd5153f58d869d0c5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94326f2f4cd3f20de736e64d5513995ad7beeaaf163bb9c3fcf036a900e91d0f72526ef7748cd8bc71bd52fb87e9fcb06a05;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h195d3e3f5ad9b9b9405f9fab6eac9b8816ca5b82e5876a4239a08dcb194001161fb6f96b7a3c5afb2e14f1ee375304e779a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc03a6ee1aec3b95f889dfafb295e3d8622705b559566520c7e2c4750b813df2765eaba2144fb8b1ce47b4e4c7ffc254c3388;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdac7ac4a6ea1c4cddbafae548679d6252153fa50d6c3c33545b0307bcd1bc1a4ff581305c12019fe2cd58fc494885917fef0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h589d71706990fc014a885b929a932e5d2b41e89431bf600227f126763c2ab72cd35993a0501d6d1fc25cdadf3f0721231a40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfae609b961615695fe7abf553650dbb2b77d54e4de5c8ff55eb9a43d29fe9fa96c7abee6bbae8fbe574e0239e31ad30095f5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd38415d66fb3060f9b819671d196e9682800d20ea63b50b25aa166b8470e5104830c79e703539dbb22d2b8b0922122b5d326;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38f3939a98ff124cb206825e1859d58ad2804e3022c0debd479e77c6f971b4642ee3b95640e7c9afde61ea05ce50a4309a5b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60f2cc3f22862c04e54db1c204069cf547028fe9c08704e73f99c5a011a991bc19af642156b16971f934cb0831127cd40a01;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41e6a63dbbbb914abd52d9794ebaa80d49cc9000a253e25ba1438f56646ff807601b8716b3404dcbdbe83ed485378a1499ab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f67f5493fe95f55dcda70b9e15550a5e7468351d6a2a83095bf7509ab30d95821488f157cfd9724db4c3789678da3402567;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78b5712232d417f6424989b2e19594df5f2f3231b8952268585a2f7b0f8922d3983d3b2b3e61f5d1e8ba5a46ace6290e4ce0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56f1f51f05e1337e101db7bbe7b68321c48ea2c67fdb43883b9ee84e15d53855886ba30292dbffa1d475f5f6a4958dc168a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f144fa3f0c2f05d4394578f0f4e7ded9b3e129a7ba5fa5d1fe89ddd952fdf2ecfa387ee4082205ddc548f9d1f7c62c1c5a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b46b190abd2d088b16580778e3c3e1b6e189e834b1d049021f2632d2cec1726904d64eb92f05704b65cc4c03bf7149208ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcd8272c604b79b50680de18521eaf5da22a3fe1da65066df8c8a26a8e79ba5662c7d317ac55a1df9aa261afea87ea255f54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9ebedfd2826cf077a2317cd690c1f5a96deafdde70e01c47e920e0706694b93bd7d17cdc353167f29ec0e77558c9a11da18;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4be1464845978d051f7df1ea52d27aafc0bd5d5ee47ec7943198fa67b60269db39fffc2210150ec4b883d37904ee7efcd744;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h151fa2269dbee7869e583f3f46b932ad1fc1285f01f2352c322f321e836cbabd1d72684f5a5a9602399446867d96ebe98ec2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94dccfd5a194f0aa0e0ed6e0b6a0fda80f98e11a35c1b483206b6513348336f9f0c771a83fc44641e446e0efefad9b635036;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf4417b854256a384b266f6a36537017430586e47846014b80711efb6edf0731bca482412b0039f13352b502b18e18548cf9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93fddcfe5d017c07b583a96b86b14ca7e63dd8832bca8bea3f90080ce731eb09c154947ad73f0cd3b67b8feb6fa02d16a480;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1c1a3c820a0581daf8650fcec599f2cdb17c1fae8a043560912b74fd4b4518ac21ee9edf32d16bc0e830c209bf690de2c35;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e1735884ead0c7ed7975b86d8bf69abccf371aa57187e82bd395091b54250ebbb61a0a0268f0f59483491835d085b514cee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32263619bcbe2b515a66901779fd18e60a208cbb652bfdae16cd117ae397430d6aae3b1c522a9d9e3da185e9e78ada2b6b48;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h536d1bef5e44fc8919337265cddf78be06f836df52be2582190befd151b849e8a1a4ab7a688808659411bedb4d922fd6cd10;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49c87f083b90d759e79ad30ac5c47ca83d816b49bd21d0c0c5ca8a48afdd6015762a71cb6c216d43702a1a5b138900aba921;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc107715f0a636f556b92bd7cabe958c234590ba8170a91204fad06578efe4cd89272342fbf1f369fc550bb98a9370adcd70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34e85dacd4fbe68ed1f2a3a30d16f7940132f759f24ce855cb9571a0d24cbd417c56c82f6992be525a098feb5443aef6cfdf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21377adccd6e47a47707fe0051d4ea3336c4251412ec3ac501dc2656ccdc386480da8c19805bd509d3fe8d5cc354c638a92c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87555e84ab958e8923823c8c1fcccc3a4633b840e16b22dc542746f3f027b86ec3e6aaa26aa9379626edc2206ac5218a9e8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2c390b2e8beebc6bb61952429c5a12883fe3b22d5e0856dccbb90077e3b7971188fc3277d36d662f8f51d47902f89f0d1cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he651eb8674d8df511d4736426271ee50b7c2cf6de73df07421f672427513a86b7dcf71debf515f204057a947a76e95da595f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc02316454555949949492a88674883068b7e3d51681a278a9563ebcb16d08385957d7883397ef6d174aed99662849aa45c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b65baa1cef3c4fbdbe763628d55a37556c1d5d477b6abb7e76a7cd9a072db5d60f44cf9652c58d641c46b45a2b492434bf8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29a936e9f37941d2a949f5cc3d0dcb299a47fe81fc5371f8f0508f8bc172ed3c99db96b4d3c0a407f4d7f3710a876077386f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a5c556812d2f2715a2ba904323ad68c32a4b0e9261c422a1fcd0f85bcbed64fdc825c8ba817a12d22ee830ed598dc643df5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he210556874dc3dfe5ed0a10e926a674bdde15965a987bb88337a1569d0b509f1068eb068a542e49c85df5664fd89eb9bbd10;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7c5f15aeaf35c6dadf8823e3bbb58670dc2530a2057aca5b9430530fe645c95ab2de6e561844aada3c238e4731e08a88843;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b04bb8663c48143b9cd7fd597af3f7019b1344e6068c34c9828a84ab10b97ab69bbefb2e445fc0330ed9693b6527d556080;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c5643ad1089ddf0f79fbc59be0d6fa0e1e910485befcc28c3e46c6ec183fe118a5e088b178fa93fab56d313b4dd86aacfce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0ac03ae850b8fda49891c3ee548600eef0fcb89bd278bc3bba9e26fbc9cbfdb39cdf1ebb54dc95c8eead493f8f7daa5fed2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h765904ab8f84e0b2e4ecbcba919d4606105ad54ebce3e795be4d9612db8b480bf29aef8d359bcb9f9ceb5d0ef54f47155eab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdd0a28c690bbe82280359a5b87a8f058931867e5b1e43c212ec921411e065d498e7798cb7e3030c731ae16387ed21a28c6c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f95043355d3f62e98612ba2db4476357646332d5f630aba8102433735e4cc586122913565a5d0ccd94403382ef270dc7ea9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h860f6153acbf27fa90c84e3ce6fe698eb720b0473646a1f88ee23019a16bbcc058c0a7cee6ea4c68c8becb78926bb845dc1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7eff06fe4ee94e6da516626753099464b19ac9e208029614ca5aeac639d750e7679f557efec5dabd5f23e2eb9d849250d4e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb49096656f1caebd033b6121c4ac6d0078d59996ac4726ebd4d8372c2f2a94d2b25f4b73c705892c7a1d757fe58fc19d50c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b1884f7033cdab59a0f5ae7636b9a56d6e07ddb29fac2b41e07466c3362c6a943299bc4b07de5c9c3a434ea08ac7a614756;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c63642c2059e43e5b0d6db069da500f648dd1cae2294e55dc37b45f49e49e7c4f55cc579165b4e57511a28e6bdea486f0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14549d68f8c73bfbc3279d43826fc3472579dbf742b1d17db7243ba5852f86b939672310850196d619581168b3aa713fd1ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c1e48af16bbd7e38c4a05bfa8b148f6e4835ef7efe0dc46d796a70acc584ff4e6a107f1c08a62047e7720f8eda32c65fb3d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f7a3ac46d01fb6e64fa0b5b8be174851d824c98913116a8dbfcb79035d2c0a6ba0f02cf40f70c41f6b2738891d0e2e40d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf44235e5d3c33e260848fec01e20c32b52a4806c1d396f7351ecc6f308f2e691d64e4f12e4ba03f46b47cad0b3a2ae5dbe41;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7935ece07eadf495645201c7ca9a35b406f1fa3ce25042cdaa9c3274dbeca2181e64305d7da53c7a79a6f6031ca2af79c52d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7ee13e2e89d037bde66aee3f713b8f27d11da5f846b810f4c013dd83d99637e22c7c87f61d7815bbb03389c391c52dbd38d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5b2b31da2fd21f06d0c66d39fe639f720d725c5fdec139b993068de4885cb986719cd05fdb3f0567ee801aa8af47790f93b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78998bada045893e1205cdb38128fa60e308df690a96edd59266566b7332f32f029ae6f653c993d2d666d6059cab934fed87;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc31b2dfae9119819662de62a322320db86b65f1fd86a73a2876df8d41699c42c670bceaab4ebe57e81d754b38b562218401c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6bde5d5c7f9d246cf1bfe38a14ab9d8de52a0d934d54fadcc48402072ff6986d194cf8bbc4b2480f5a57bb23d1076bf1d04;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacae653e60abb61224e995fb49973a71ecbe89cd2f8dfc321661cb7c14da7d0d5e74f4ad7cdac46c68f00c407ee9461ab8d8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha344942cb4bcaf02956bf41d268429ad53ed604bc961de7f043a0997bcb53c83c683ab4fdb55c20b881db03740b2ea510ce7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h641af2f51aee8f95801013f115d6ce3478b100b9029e031a583001b93b97166b7c9feced6f740600bb5011f97707fc5728f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce8656ddbe9ef39ed2b46d23ad51e9728bdd83e7ce4d43eaaf2a6ea444187f0917ca93dbbf09e5d7d2689f68400184c57702;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda89355a1ecb70cc0ebe78553cfeba3de994e1d14a01b0a4d8a5bc8ca6356940b78596799be7864fa3b6b57aa7b484d0817f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2459466df0de047d6b8ee87f400e5ca304f114bde1f8b4e8fae684ce19667ff3dc73c156a16717a09593dbf545c883e9a51b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69db3624a5fee8b73a66efd3281d5dc8b43e0fd082ad794136bf9c578c1e1f671f460bb34441d4cc7f161eb498cca935e979;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd6c4bf1b8f0ca15e5008b336c4ec34bd05a6926404850c5bf4c5760a012639a3b0d7811f98a61d5c23296ec4c5b5b30ba1b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76ff1ff974c18da8aa82b52194be90b3eedab4a70ad3c2fefa7b7df4fb386cdca3671b52091a3823db8fda963c332e1e74d3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3d222a2c39d1fb9a10e28c9cdbefe8a617d7affead5a75c923d3d13a7cae83b2831d53b2b1a913f618b334b53fdb16fe9c3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3182e34e79bdc2f48904f11f66b0461f3ca59c0d83ff06400ae1bf8caff1ad634a35030797563c26c15f93c1aa7e64694336;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37248f284886bafcb224d376c453da954e347cb9d8cacafc4df6f3d22896b2d35c4dc7ef809bc82c17af1840af9c198c5fe7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haddc0cdf4d9c74f888ab7a7ace700773190808fc8c9c9b484de17efecf27e479a9f6de2bb036112521a36d8e3df39b8fb6c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha95f7475ad3a44de442ea02cc5c4cc2e6f206a029d7b6dc3071adec6d3849a4e65b8eb6fe068bedd04072e9affa7a1d5ae17;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha31a8f3937953079d94f9916a2258df700b5395089a1cb3e9415717ef4b632c5036a8ccf6ed9418baaf7ea1a5e83fa4eee69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87eb8cd4fe0a083253cc29b9e2af9cd7e9f3e501cf68ad07862ba5880f19c46a5f0d3a0e8bf60669dffe21db9bf53484d15f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62be2cee94ec089c7848769901dd4c4e798f80e18fd5f34ffe4afa2734533efba4e89e39344b53bc09fc0593ca5ba62d685d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ce20d213f8d3138e3148320202d0031b3d05685ef84637936e17f2ec2b106c0d968167c925916988cc51ede979f209f738b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf1a13d4d91a90901c957050b0ec666be301b250916f2492b2d3ad28b09aeb972b418139730ebb3fab585a1a83e06fab84fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bca0bfde44d4bb9af4a09347f2fa0554ec17eded4e53840964cd292d06aa0db7cfa437fbafb3c57c671f5dd5f94b7eea26b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5140e21dcd48f7da9827f153de658fa60f09894e63e2f6c23481c9c299468132b893ca3dfb196e1bb1a84e8c77236a58463;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78ce8be73d862494f8cd2b6a011225e4df7c837fb410ad0303c49664751f3ec956e1c91351691b30027b40ea1fb2593d40fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3db300adfba587d448c31d76f31d9720039d4cbf0637892952ba3a1f74ceacd31af9c3ef17018c7286bd2e8c686628a973bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37e2c379b53559053c071240819055e332c03492532b69c3e206f3bc9abfebea4a9411f072824155230a4ee1df8f027b9c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he51f8adb9acbed6b20f2f5f5a7164ae3ad20b9030e53344e1a5b94f589aa82bebaf1e40cbcd45894ce64c725d7737d52814;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b25173d42baf2b492d63a2c15e7bbb4158adc5e5bce3762dff73d68525d3886ecfbf6ac5d9d52defa475e8e161ae13fe69c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c5b9a5e1756d1eba2b21e661cf973c4c9c0f33a28703d9a81162aafdec2fccdf8545357610e74f759ae6fc137c87747fcd8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h198d7d46ef3415d4955af5aff731afb83a50f3b69ecc901c2474459adcb861286f82ff926e8b45ebeba849fcd1ee1ec1aea9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfccfd70fe5cbfa37bbe30ab229ce57812fd77cda44dbea59e8fccff57e95a0c5c15225f26522aa2fd13b5cf705a9b6f1160;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h832c0b3cb7be058723f73bdc3051d8c23dae755b1002b23c35b76d846a0b47812767d39c750e983613b66336ee90dd2be467;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73d030241dcba86fbadda8c9f50e1a97b2c314fa16601b3d0f77898f0981c198c2211790b0cb3703eb45724b132e532e1a65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8687f9f9e85c99c4d6f67b0683b6f01006350c88fbaeb8eb26d455d4442a7e1086857fbbd80842484e06f86f6b51bce38d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf685014a02f9be0e2708d3fb49f567943108da5d536c1950c5ae8c49fbb30767be890521029a7d7d976a4808bdd7fbfcc914;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19ea3d7af33545c5db260125064dcdb3a6b3af20f105a2543b5325890252ac9f45f0c6cde99d069dc3d681c400ecf3fd0701;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97a23f8400a65a372008cc6a6fd8fb19714d1f18de847107f8a642432ac9c77ef53a9a96f337b09adeae9e66af63f0242ec3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1e24315ea5346c1ca0675ee5c88cf04ace13ca6c7e0f84dad3d6284764440f46575e0d3670a2e209ee349b760be841e0637;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb010a311535207d3b0167780e8953edfcf351d5258261cd2050770f1522e701a8439cbab32ceebefab18e325fdcb97e30655;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2825f712b3951014c0e09cb22d6abf47e583df5cf322d2a47cad171e725a10035ac077d1779b57f60b52cd6cb50c807db29b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f144275502004aad1695318f27449fe45f85e53fc15d70314dba5af589f5a9c42e2818a27d445a74e9eca758b09082727de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h309acb0d54fd9698d5d53ef6ae2e537875d9d5e916607077c7dcd2eae778f59368e0b3714dd4224c7d2b6a7e4317310f731f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdbfb00d9f8f538e9bab739b0f43e56dd90ee4b75a331ce306b811f16ea3691377b1e0064c2a3b142411712da24820edd6c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd60d578cbd3346eb45cc2388b391739ace2f71dacab301256902ce803a6b57775055399b8fa26a11fe1a60335da96faddc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64fd77564dd77c4af7563b59585e153829954f0f2a8cfe834c27bcf63ba2910a487acb057211c8faafdfbb940c77ada79f58;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde2d80439f7acf382483511119d211e35c462512ded9066b868bfdc0fccc4a1194b7e541860deba8709c0b620893bb66a7e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa8996c017339b7d367d20bf46c50048a632736255c0432532cd4aa02590dbb9b747f416ece92e4cb51c63a39e739bb20d9c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e5ac10b3dd845530b491bd0ed3101a3cbcd80159e0780976ae00703073027a167cf7ea6e2bd90a2abfd676cc181ae7a3261;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h463344210cbbeb09217e951bafae634b1412e5aff7326dc9b8bdbd4caa2e405a5f1a8a6ac12ce73382074ac86fc83b915830;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4135f5847bb57a56e9ef762118337763ff782f9e55b4d1caa3e1688b317293078e34ca9f2f7f88c1bd43b88198b1f9c223be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he218868d273e8e1f92f77ec89839ddee0ebfa45b14653ec9b01daf08883d085a95635e2e49f33c2d70a05e45dd378069184c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h276e68fa2b6074b542df667c496a4741854b1ff91062e346e02498c79b7015b9e1e5fc50b9d09708e9171eb401b03da27f31;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75f4a2e8b615ba900ab685c78b54cfed444b5614c9d4870f8b778cde621f83639dab327879702777b94b4228ce53ee0a3d5a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha29f77b908fbda7805ab4d0513ad48281ecb559de1a7ba00921f62622cabb095152739fc8c214bbd1e64661038f11eaef4e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h768d6d309de7c9962bfd935d5ff679e1cddc1fd69136695bc9ab8d0abd8b81e850da32fcef3ae80bfe2be5f96bf4daf117c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58090a9bd8d2336204c2895f32b3395f08e654cddc56c0bd616132d339f9e8f65f4b9fd5c68f7b9df9f8f4f9373bf0ae4f78;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4f5b74ee9bc5944a0ee377c513c5490c88629d653ba74c4022e9b34cfee3cff27f43e1ca9b5efdf4aa03521c4701db790a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc6aa5cde8bbbeca5d8c642751c3b75d1bd405b66525949c9984e5c75277989c7652f57a52dc1c8c5424815e4c7d3dda5b91;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc01d7f10cd339a8993355e93881d7b57cc6c096994c3a31cca33e3d2957120c1f12758986a9bd21a1510bc124ab542a9782b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2c212ddff756df8dbefb0a21964bab3663b84b25855753ea41263d648283aa1c2a804b9db4e7a009f2f0a3d4a98f1c3c423;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7f4b07460e37754d3ce316b02869a7257e0577d3aafa42e85a04139bd550ad0a0398cae26baafe1a1cca79d6c69eb7b2e67;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bfc3862373584c4f9a11bb9513368df3dd90441225042391aae74bc6bc482d2b2d9bb0f10df1786331dbed1d7d84383dd9c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1b96ebf5aa04e781b6952d67a98315c42eeca68df5a884ab6ecab8d9a65be542a33d0a0c93645a2aa963a9b2515a62fb1c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5030089fb0da5181851e9964c812b1a3f227582e304cde90baccb9ef456d3c8590ebaf692cc9996278b410e38140a5dc2639;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde7b52e49d614cbe2ec883133d3cae512242c5832ece81d2efbeb6273a3a30e3aaebef61d076eda17e1c1f24914c099b2c9c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heed932ef9caaeda9207301f338454a365ed208ad99ba87497417afe830e28ffab85b8c1ed2131059e04c531f22eeb198aa9b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fd6a2e5798fe62d3d54210e11dcde969d77dc7f854ac0fdb5d9eb8d88ed85c43a7f164698fa701e15ecf8aa1e99799f9aaf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37f9cae8d02f366486df72313d070f947e750f1607d9ce8e980b61fbe5b72a0ea38a579f432a27770c2d59ead5935b3cd15e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a3882689b0496a9558a77a65ef26b750883670498763774ca69d99d259e91d602babbcf7e3bc810d21b933b9251afbd7c32;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb25d2944483bf2acb80474ecf01581e95241d3e1612ff0ae7d4ab718fae7e51307563152e177e437a08a500e0ececf80d198;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b95bbf9083e76b0c9d70e140831243e1cce29d02058fbe83293a497a66752cc4f88b8c83ac7ee272d1ec23d24d69b025060;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ee0847451ca8870eb294e215de0acd83851e0895c7b1b1b620d768646544790e9ff8ad4517cd9aa8aeb12e62d812a548057;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e28cbf43cc9339fa7c5161dfd06f17f745e4908a69da3d8980720074ab6404a784a70eee887ee43f988ba7abab27fc35f81;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4923e826f787b6862a4af9423d7750574dfe774e00757fb7dd21e80af101e5fe4ff65dacf7b3ad1d95bd0f18b68228d74d43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha94c7794fb27bd51c89f645139dd4584e00ba827bccb5c1b271a1059404df1a10f9650b64f48a853ba10becd524a638f78ae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ef04040e55461849b9c6a70d45ecbdbcb86dd6a06f25f6064ab20b1bfa9bb6568124c9053f81485db8efaa69bdfc0f2321f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb224216ab842161e3151a2cada2ea276cf6c4148aab23dd38e66ee176cf99e49ca33c1b131e0f39e5df2d0e520741e7e8fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93ca48587b16aab7a7045804a16380c7aeb165c0692619560cc4201c1ce6563aecaac59ad8c99596da62aa407bc46531f8f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd66485d686bdc21d62d05dba6dbf465e1cca835bc792bdc7cd3ec0a98e88376b3a14ba0a01f3bc0e5c63bb35693a186c08;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf982a15efe05696edaa13ec1cd55769b9767feae1e90e20ce1fee8abe43c041b2fbbfbc756f0e3fb2c374bc080ca7be0044;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d7487253f04364d81333ddde3b5fafad4eac34629bc177b955943167ee005305896fcda9b50d77d435a5ff37e1e625fd4fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69c99e651b7a6450730c5d360ed12cdf1ef2f21ca4ed80831884e3409ffdc3dd15c8562b933f1ece483ff367edb1c513200;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a233f9ea1bdc09b803eade4cbbc357d4ab023beebe49ce0fb9e3d3bff82f298b0087be800218dd98d5a7d37871d6e4810c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h141bb9ea993d0547230c28aeef40e5c604be54cbf2dc1052d39c2191e47bce86c94a3fb20a2560aec7b952eb5c0e7fc339c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb6ce1410e868aa8055a38ed4ce5742c4610755d4bb2cb26812d6d8da237755be863af78fc4249248e8575430802e9fb06d3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c250e6904381375da080a867514f49b3df1556961eba78cc32caf53bf1403bc162658414ebe47b9d66e2f0939972365d5ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92b74c86093c2faa310d204819ea70e38cfa991e47945eab43f6d82395765b1d7594ed7beef95590b6ec4caa959e3fd87ed6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59fe76fd43cbe517663a52389aecb40e39eeabce579597d53b20d1c48d9ce8bf087285aeb076d914b199c516378f45f16ad6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6e4e2f446059715394a3b9f2e9494fa8679d059317658f8f08b5296c8293e8b841553fc520be5c3df7a061e0552a8b4ddcb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6060d73d924cb6526abec8218e714656c21eecff7046c048392a682199df15e3af8797335ca70016c7cbf613cf10c039b834;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a03a7592e5d6f88c94d3a5f68a1331965a29b642159be6b6443f1633245ce5f765d65ca53b3a0589dd09665abc5c0f42fa9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf07a25e12d65a98070d2379324eda2b4a195e3c376a4a2acbdd3ce5c2fc83d0332f8c4609e28c16dd5e213d5e90d94b6f2ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd73ae8349221535b67830c74997a265e85e0aa2b5e2cf363981b7077945d25ed2618ce9ab414f631269798a7421de2a3389b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15c3c3c1b7d072855a94372d3f235cfc59f03ef7e7c0559655a90805f2cdf30aeee133a6304a9f6550f45af085be64528a2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd5cbae9e6bef874db6500c4d5faa76e5ac40ac79bff437cb2872c089c011448e0a3245f8c09036c74bf49457658765dd1e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac6bf60401a59e5c783f8ac89a79eeb84a87948505564c7a4c290d314c0475ba1081454aa9021709d0c19aacc110265fd724;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1c5e91cfefffb004e5bf7852aae3105a52060e1c887ecc6991cb5a66a8c0a18eb05e0ddd6085fc6087897b37464d8a86e8e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ba0a24f8a83578f1aaf5c8765624bbf2e995e9822709f0e77fca29ab23432148f63f0e8fc6e21461d334afe542fe9f07371;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb21734ce98ee43cb74fe6b31a667c40239b324650d078004808da8486a67f02028ddfb8246815d40b9d780d96a4bcdd1e461;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf0d90b5473434fe7e6a8fbe7afd7e18df8995156e32a7f52180654304290042dcb725536e990262755b99e8e7ea98a895f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77ed2d9439ad2977f3ff5935e0575411cc8f3c1eeade7abad31e110f2d98b04e37d820725d98a6bdaec0f1f7442b0e8ac6ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15720dd4fc62280dfec0a105bae47771da2c55fec56a94532696d8b7ad219b6f3d603659fbf3a79da07eae9a3a0b8f86452e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd88600c4b25b86cf7811efb91b7a2f84ce04fd0759980b344e6ea39a28a28837174d913a2691732c0615f48e1674f7eea40f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7686a0885dfa16fee301d0ef764139ffade6f8044c112e40b6723d5d72c800ff3e42e148b65c654607e41d9e505826fe01cc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b6f805cdcbc7a924e295984df2ccb0f50efd83121fd184a4c285a2a7625f2c6bdac8894c1e343faba74c44cf82ccf72f53b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77fbab1b92bb848ab59aa55524feabb1db4353692ba545fe7b34f75a6572702f7edac2e334255610530565e72de59ed133ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85b816ebc362440a098056725261cf438123fd13e79b42a1f3377ebccd1fed4e92be332bcb630f465de616989a0a776d518e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a9c6f0a6f1bc68b0d98953da64f0f31c71c4a18118f142145ddab007b5e1d03e078b706b6412040b63569fb614679efe067;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34b5a4058cbbf9166920c04498075db1f840c613f948b8b5ed0d96b6824a96b2e57c5b32bf886e4bbe5397b0cdb52c7ffedc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ae27657b0d868a8182eaeac8df433858ab098ff929bb193cbe8cf7127c4991ae3d2914f9bd7d50d347ef424ef65ec8c0fc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98c78d3b35487e41ac87c4c41bbd7ecbd73f9739bd3245f16a17ee91e06b67dc7c48bcd92d438a7cdbbd7c8c8da134b77994;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31d34035a0814dea4f48b16000fd83b447ce1cd9fda373a73a70556f8453cb8576c7cbac5bd6c1b89829870bf1f480b6265a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30eba4f097c08b98f757f5a3152d5fb098210c9de3c7fde4ed7b0f29af32ba9b2f5009fdaecc506a6cc4d25ffb0a2d7e0642;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f53c0ec4edb57120fc67c33af99a2e64511fc416d8c81bc90ab10db6ad17179d5a8460c5372ca2ca116ef7b9a2e34b81f21;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha26f6389318c00171a51943bc2dc394f07de559e8c54ea31d710a242d4bfd811da4a8b488df2e73ba3ea26c2a10401812a51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7cd2340b2c83ee8c9426ee7ffe8665386e542577330058804743c33ad0911dceaed32477c7b734aff61e8c3803f9d7c49284;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ec18e75a393c6d9a9a4491e216f5329e261996a8a1a6946ecf7b892f67a1c5eb663c87db3e649b0c6cb439fe8b8936e970;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85dee256e15167c250b5da98bd947d7a3e0c6edab5cc52cd99895a330056f857454244a01837a5fa50382e82757e15a42f40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf382b7eeda4938959974bc09ac53ab97ebbd164cf457e7f89cd95cc0c38cf0313ed38b3116177db06836098a8a986c19bb38;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e7094e9467379c2cbef914521156543ab152b04e388a0af8e0f74cdebae86ba33a31ea5a5f88292f271ef3a32371e4a4fd6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c76704146fbca42a92d3d22f600d90f24c7b1b68961291043c2d5064fef2a0f5bb88086bf944642bd34e96b580d4c865b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc551781898b99c805933e6036c54e648566f582c47286967eb46f71a801ee207d138c4c3890618ec23baeb54bacca1170a7f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he74fa40ff8323ada1fac331a61cd597716e23506ef4a0061eec40f8726915b9165524bebdbfb5f9d62254c8d460ac975bbb9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h717bcc62173a76fbe361322ff3a7ddcd5c2d4908df8bcf45f69a1db4bf04009471bfa12d4516ef4a69d482f726dc53d56323;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf201f2ab1bf17445865cc39fd470e23c4d8f8521c58388cf0ae406ee4ead524138cca033128e3f82a3fd2b788a6705de96d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h735488082dfc612394ae054a36f035a9c86156a75857b52e13fe2596373da2ed9cca29503a8fcd78abc114c1ec885f8d8589;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5380b9d8dd687457b615d7fb98cb20349dfc56d1505bbdfebcafaaefc9dfe13e92196120dce72338094081f5a5d0d64e408c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10802c895765a6b7d7a8b4259a4beac27b3369a5b46627caa370d4c5d67950415a7085b6c2fdb738d843ba256ab5bb1a7198;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4ab05fd4f59d821bc4e31f160ea605291bf6b9a5dfb701409f73e56564a92c43d76afad8d75e4e93907c0b67e08477716f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4717a6c3e6a3144c09d858148067c9a3c54712575613fbaaffc69eb4f549323997df0e62c455d2b769b3c503e1376c56a6e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8616debdf0eeae1a592a343789b633e0065795ec0992b8a53cc5b18f6005c3c53ed310b1851561463e72db1cebeb94fdee50;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd58e698c93aa9855996b538e7a058893f489702261baedb1870437537487e8bf0d4444c823aa8d5df8235bce5eaa8ff7c54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7288e5886a394ee1a8c535c60663780f4fd9cb87e950ed351e5d152b1bf53e2ec3c05ee719895b517faf7a94489941f2bf40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32f8b51f3f82d2309e09ca662c6e99955efb44cbdac16466890e09731a1cbaba35f90c7b18f2b48d33f7097e3ebca82a57bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9590bd4b00c84ba32c42ee3aee39b24e4d1e7d2ea154ea71e8af25e723892bc9d208feb8c0e9aacf8266820305fa9f7bb554;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h436635e03ee42e6b9bbc6d0cd5b63d04c84fb6d83bf617829ec6a125d574d8013e115f20cbfff53cd6fd9430b2e75644c368;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90e964c363955283611fc70c40cef8ee721f28904ff198c9e3ed1d504e26bf74fb529f8669d4bd70a64120391f1285255835;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97be90f5f4c9877305527ac08e966c1ea901120075dd3b4f916edfa5ead75d8230f208d37fb5663a98c806a96e04c490c4ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5d924563c872f9b05337f8956731457dad844871c464b48f8b3aa8c2d898cb7f062fcdeab3b12520d9190dba0f3f6df7b7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34a2668a20984699e2924da1f31aceea8201c8c02b881d2bd9513d372b2b396f4a4e636313bf475cadaa4b68cc98f26c3bea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8b66458e5e4331115881660c669c79de3dd35f0ac8cda9ebd4f47fd1f92434a8b58089fbd1721cf6ee8e7c7908624735816;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b6061d3be19b679e4f09aa7e58dd611f65a5930a1320327f131ef33e14244adf4494763de09535d6ffeaa3a49810517ab5e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f1348e17d7bdd904c5101dd8f7c20786f2984818c5bbf217798866bb81d164295cb10d49c5ef6e03cdf933c4d0a60aa7fca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha045ba30b44eb72998a053d52b3fd83e69c9496d4543bbe6760c10d6d8faffe1eb8715f3046eb672232c31f7592d0478a6dd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d74e2b77f001ef617ec9e45587dde724319f2e588a37af0c78baf4bee70a05234281a8457115b664a0623a429ea51db7585;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38ff48fc8700194fc585d067108d31dfe5cb0b4ea163ff0a4f5cee3670e3088d76e1891e26ce3df04f24b28084832ccb658f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47d50b70dd4c60209f5f91afdba0b16b6916b88b5967a7a4a788ffa913e64fe4aa147a3c91dd12cdaf1e22f9ab3af9c05be1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h978590f45b55aa635120a8cfcbd5b2cb9774b7f5f01e1314eeb094113cc5d799cc4816189a4016edb8f27443f08bc09181b1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e262b6ae7e794596c861c5d70f7b338d9a8429071c150c6ef8a64dbcfb643f08e05c83ea86d998b585292e385cc5dd72fd0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea4f71d16db3f7c08966f5c129cf5ffca8e2d77b674bddebfe0f70e408acb7552e7b504404639f16c00dd139ac13665363a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45d34b9a09988a79e1c6f884529dd7239712ab61f0a8d58b9722cc2567cd06a34bde3af80882929fd1eae83105ea3268992b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h859bf043c60a53e5617799172aa713f768205be83e7f6de985189e847cd07e13673ea1616fdbe504bccf55cebfa10886c633;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc1c790774cd1b4c7fce9255297e583d79fb3c2270754a245b17dcd323932f8ad0747c9643a9ad6683ea0a6b754a8554c8f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8a6edffbe110fb6e3cec5a5996af697df2032bc3e4f4f56faa8309990077b9987b3d9819f56d2fad2f8465b9231dfe39b88;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haef6ee602885b88ad1537134951708f50593a7d915ed21eb53dd65964aa8ee20d7987e468164a17b2f4cd0b670cff99e9385;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h509d85257d97fc2a4b9dfe43956f7e15960684a6b041e2d495081fffbe5cf80a7e32aef889d84052f4774ae9690ffe356dfb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b4663af00ab7978a159702b46d31c3a74da6fd8fafa4f4dac7259169ff935fbb81453881c24425496cbde104919d8a9b3b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d9d1bcf4ec53e3dd9476c78c9dcd4a6d91dcbffb516690115f4b85e1d6da4f45596584612dbfcd9ff042363d14cd9a74bc1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd720ab924357de75e2f77ff0107bc41d5392ef7d7e8aebe9ece3583ad0f67e979d4da4ae6a4a48a80b11d36ac3d632f6ac37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4580ff688f9743f3f2b5430f757cab4afc1e92a72a5a4e41cbb0eee3b927e9f8c9820f123969d6ceda411c7c2205f36f412;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f1870d6ad5bfab48c12716b0c591f19adc9d48e64a800a734b581fef4b54d115df5f14e7853a4c33fb1e8881610d54b96c5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2c14d3f91429e9c1944b9e4d1de39686eb7e84d545e625d51873ebbdc3316bafcfc745ac4436eaa559a48e56494cf725f94;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6992289ea8d8504b3955df3d69e677e27731bebf831aa19ef3bd486f987bff00328165fc940b54e9774fcfc81f573ca5fe76;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf94de57689ba29a547604d31fb4eade8a1d69947d7f4b37ac8a9bd24c1213a83155ae076debe178c4b3f909e93e543a3bc10;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2e799301c7269aa8b87208600bc5e00ba2f0df6d8c8ea7e3ee5ec538ad3b3ba11becc08f3c9f523270da5f82826ae8e45e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc782f4ddaa7e36984104d5c3bdf90b57a5e20c0f1f36e8c8a51b1ecaac2a4640c8ebba5b17d74b9faca09c4a81aad9a57e4e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0099f4960b0a8b2079f49dbe052c332c25b1900b3f335b6ec873c9be051c15707b443ca9c696c3df7218c91c863b925c313;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c8e0fa7e42d99303e6332d63b75c15e9a54a47b8948f4aff33e1d34714c16201eca7276799252a3727bc9f5b99cf90f5105;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h776214b2cfdf1f576bf46f423993dd6c3074968fd1dba012b8d52ed774cdde4915e07e0beba207db734fafed971eaf455f75;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e47d25638b257098ea9159c89ab74aee3e6099b0c4c4f38722534bcf47ab5925878eb6e2af276d6ad4e7f8be607c99d34d4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0423306c957f64365d9902f3053e8fd7c6eaf9262bbae59cd75a36c7463c72335d68a8031de515435c55df84ef093d4df41;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c67667cded97993fdb56cf238d522b96887e84b1da5fcd54ed8654e9d89ee3ec9276f54536ae6de17d58985345be62a78ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafec1ee26a1634f0ad4e9c0495337ed61c9437f96052648c84d519c5037a84afe8fac37c8a9c1e1cf52a0744a88ce649190b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0b81db9ff40c78ff8183ed32d215c8ab2ecc6990e61319f004ac92692f8b9ef261edb693d6330f36dd64e745c96a56a452e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc76a018cbc9aaa4f348bc9beb984c0c1105fc1b3630eecd236d348d6e75b1ec89fb1e57d9857e2fac777111008a3306e5ff4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5353a140673c509afec2fb10be18df8b1b5cf5339231b371830f93dce291831ea41f3f460e021bacffff5a1d4f07d7ec27f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f00df9d142901458cc03cfdc45124af072125cf53b8ab4a396308cf075b8e693197dc6edf285072405d64ad8df6fa80503c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecc607d2de335e90108e3dd2b1829b535e42de5637a49e7cf6012d5eac31c6496b6fe30babe2ec7cb895aed38de0fa0aff40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h568d5a315b1ef7a27788282c94ed7bfccbaeef2a9246a3252744c9a38faf4bb043d0ee2e6cbf2335ed00f8707925e848ff7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d17e8a563c33bcb9609f8136422969b86e0dd3a25e32a696e6bacd3cc15139a9d92c88b32dd9569f670c4fd2286ed4028fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71d4b28ef57a443c5c435f9bebcecc63b00538c31abc81df38b5b4ff71c0f766dab0242081520f880cd3e8b634c9c4c2b221;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d863fa1a808460775003aa9d395848f958dec77264a38f2f94fd23e280dbddc73677a2d584ea06c375bcf19122aa8445812;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7248335adaa9f8aa3ed854e06d0d099b39341877152cabe06388ee503cb37e923a5ed988794a408fc6b7a084140f8aa0b91;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b38a092da8d77cfcbee9d30fc05d718ea1944080f43b0a3396643299819d755c1a2874b7a3670799ed8e9248e5a7d7fb52a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h970dc45a210334468d4b0cd89af7d8475fa12cf390435515efb09abf1feee3fe651b8f624cd6492bb1bd51204c9882f4a4b7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc496b0785b653874c86ebf799372bc1fd387215a684c343f0b964fd0bb5cf97f2bd60db397d93ab8793b35d57f82b4a64d84;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7aaf9451fa0ee67abf68b2fd709ffb803c86201e8187705ad19be5f374308f9d395712e6b6b4df5a1d6cbf1b20ccae9c2f1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6684fd2c53d34aa748308b8d14738705b6e25a3b18594a8b27cdf18ed266283e49e699b35d9912c08f4faf5e81ebd0037d25;
        #1
        $finish();
    end
endmodule
