module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26);
    reg [21:0] src0;
    reg [21:0] src1;
    reg [21:0] src2;
    reg [21:0] src3;
    reg [21:0] src4;
    reg [21:0] src5;
    reg [21:0] src6;
    reg [21:0] src7;
    reg [21:0] src8;
    reg [21:0] src9;
    reg [21:0] src10;
    reg [21:0] src11;
    reg [21:0] src12;
    reg [21:0] src13;
    reg [21:0] src14;
    reg [21:0] src15;
    reg [21:0] src16;
    reg [21:0] src17;
    reg [21:0] src18;
    reg [21:0] src19;
    reg [21:0] src20;
    reg [21:0] src21;
    compressor compressor(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26));
    initial begin
        src0 <= 22'h0;
        src1 <= 22'h0;
        src2 <= 22'h0;
        src3 <= 22'h0;
        src4 <= 22'h0;
        src5 <= 22'h0;
        src6 <= 22'h0;
        src7 <= 22'h0;
        src8 <= 22'h0;
        src9 <= 22'h0;
        src10 <= 22'h0;
        src11 <= 22'h0;
        src12 <= 22'h0;
        src13 <= 22'h0;
        src14 <= 22'h0;
        src15 <= 22'h0;
        src16 <= 22'h0;
        src17 <= 22'h0;
        src18 <= 22'h0;
        src19 <= 22'h0;
        src20 <= 22'h0;
        src21 <= 22'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
    end
endmodule
