module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    compressor_CLA16_16 compressor_CLA16_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
        src12 <= 16'h0;
        src13 <= 16'h0;
        src14 <= 16'h0;
        src15 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA16_16(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      input wire [15:0] src12,
      input wire [15:0] src13,
      input wire [15:0] src14,
      input wire [15:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [15:0] stage0_12;
   wire [15:0] stage0_13;
   wire [15:0] stage0_14;
   wire [15:0] stage0_15;
   wire [11:0] stage1_0;
   wire [8:0] stage1_1;
   wire [11:0] stage1_2;
   wire [8:0] stage1_3;
   wire [5:0] stage1_4;
   wire [5:0] stage1_5;
   wire [5:0] stage1_6;
   wire [13:0] stage1_7;
   wire [5:0] stage1_8;
   wire [9:0] stage1_9;
   wire [5:0] stage1_10;
   wire [8:0] stage1_11;
   wire [6:0] stage1_12;
   wire [6:0] stage1_13;
   wire [12:0] stage1_14;
   wire [7:0] stage1_15;
   wire [2:0] stage1_16;
   wire [1:0] stage1_17;
   wire [1:0] stage2_0;
   wire [5:0] stage2_1;
   wire [2:0] stage2_2;
   wire [5:0] stage2_3;
   wire [3:0] stage2_4;
   wire [2:0] stage2_5;
   wire [1:0] stage2_6;
   wire [4:0] stage2_7;
   wire [3:0] stage2_8;
   wire [6:0] stage2_9;
   wire [1:0] stage2_10;
   wire [5:0] stage2_11;
   wire [4:0] stage2_12;
   wire [1:0] stage2_13;
   wire [3:0] stage2_14;
   wire [3:0] stage2_15;
   wire [3:0] stage2_16;
   wire [1:0] stage2_17;
   wire [1:0] stage2_18;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [0:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [1:0] stage3_13;
   wire [1:0] stage3_14;
   wire [1:0] stage3_15;
   wire [1:0] stage3_16;
   wire [1:0] stage3_17;
   wire [1:0] stage3_18;
   wire [0:0] stage3_19;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;
   assign dst16 = stage3_16;
   assign dst17 = stage3_17;
   assign dst18 = stage3_18;
   assign dst19 = stage3_19;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[0],stage1_3[1],stage1_2[1],stage1_1[1]}
   );
   gpc606_5 gpc2 (
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[1],stage1_4[1],stage1_3[2],stage1_2[2]}
   );
   gpc615_5 gpc3 (
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10]},
      {stage0_4[6]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[2],stage1_4[2],stage1_3[3]}
   );
   gpc1343_5 gpc4 (
      {stage0_4[7], stage0_4[8], stage0_4[9]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9]},
      {stage0_6[0], stage0_6[1], stage0_6[2]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[3],stage1_4[3]}
   );
   gpc615_5 gpc5 (
      {stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14]},
      {stage0_5[10]},
      {stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7], stage0_6[8]},
      {stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[4],stage1_4[4]}
   );
   gpc1325_5 gpc6 (
      {stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15]},
      {stage0_6[9], stage0_6[10]},
      {stage0_7[1], stage0_7[2], stage0_7[3]},
      {stage0_8[0]},
      {stage1_9[0],stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[5]}
   );
   gpc615_5 gpc7 (
      {stage0_6[11], stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15]},
      {stage0_7[4]},
      {stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5], stage0_8[6]},
      {stage1_10[0],stage1_9[1],stage1_8[3],stage1_7[4],stage1_6[5]}
   );
   gpc1343_5 gpc8 (
      {stage0_7[5], stage0_7[6], stage0_7[7]},
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10]},
      {stage0_9[0], stage0_9[1], stage0_9[2]},
      {stage0_10[0]},
      {stage1_11[0],stage1_10[1],stage1_9[2],stage1_8[4],stage1_7[5]}
   );
   gpc1415_5 gpc9 (
      {stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_9[3]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[1],stage1_10[2],stage1_9[3],stage1_8[5]}
   );
   gpc2135_5 gpc10 (
      {stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage0_10[5], stage0_10[6], stage0_10[7]},
      {stage0_11[1]},
      {stage0_12[0], stage0_12[1]},
      {stage1_13[0],stage1_12[1],stage1_11[2],stage1_10[3],stage1_9[4]}
   );
   gpc623_5 gpc11 (
      {stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_10[8], stage0_10[9]},
      {stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7]},
      {stage1_13[1],stage1_12[2],stage1_11[3],stage1_10[4],stage1_9[5]}
   );
   gpc606_5 gpc12 (
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5], stage0_12[6], stage0_12[7]},
      {stage1_14[0],stage1_13[2],stage1_12[3],stage1_11[4],stage1_10[5]}
   );
   gpc615_5 gpc13 (
      {stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage0_12[8]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[1],stage1_13[3],stage1_12[4],stage1_11[5]}
   );
   gpc606_5 gpc14 (
      {stage0_12[9], stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13], stage0_12[14]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[2],stage1_13[4],stage1_12[5]}
   );
   gpc615_5 gpc15 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10]},
      {stage0_14[6]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[1],stage1_15[2],stage1_14[3],stage1_13[5]}
   );
   gpc615_5 gpc16 (
      {stage0_13[11], stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15]},
      {stage0_14[7]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[2],stage1_15[3],stage1_14[4],stage1_13[6]}
   );
   gpc1_1 gpc17 (
      {stage0_0[5]},
      {stage1_0[1]}
   );
   gpc1_1 gpc18 (
      {stage0_0[6]},
      {stage1_0[2]}
   );
   gpc1_1 gpc19 (
      {stage0_0[7]},
      {stage1_0[3]}
   );
   gpc1_1 gpc20 (
      {stage0_0[8]},
      {stage1_0[4]}
   );
   gpc1_1 gpc21 (
      {stage0_0[9]},
      {stage1_0[5]}
   );
   gpc1_1 gpc22 (
      {stage0_0[10]},
      {stage1_0[6]}
   );
   gpc1_1 gpc23 (
      {stage0_0[11]},
      {stage1_0[7]}
   );
   gpc1_1 gpc24 (
      {stage0_0[12]},
      {stage1_0[8]}
   );
   gpc1_1 gpc25 (
      {stage0_0[13]},
      {stage1_0[9]}
   );
   gpc1_1 gpc26 (
      {stage0_0[14]},
      {stage1_0[10]}
   );
   gpc1_1 gpc27 (
      {stage0_0[15]},
      {stage1_0[11]}
   );
   gpc1_1 gpc28 (
      {stage0_1[9]},
      {stage1_1[2]}
   );
   gpc1_1 gpc29 (
      {stage0_1[10]},
      {stage1_1[3]}
   );
   gpc1_1 gpc30 (
      {stage0_1[11]},
      {stage1_1[4]}
   );
   gpc1_1 gpc31 (
      {stage0_1[12]},
      {stage1_1[5]}
   );
   gpc1_1 gpc32 (
      {stage0_1[13]},
      {stage1_1[6]}
   );
   gpc1_1 gpc33 (
      {stage0_1[14]},
      {stage1_1[7]}
   );
   gpc1_1 gpc34 (
      {stage0_1[15]},
      {stage1_1[8]}
   );
   gpc1_1 gpc35 (
      {stage0_2[7]},
      {stage1_2[3]}
   );
   gpc1_1 gpc36 (
      {stage0_2[8]},
      {stage1_2[4]}
   );
   gpc1_1 gpc37 (
      {stage0_2[9]},
      {stage1_2[5]}
   );
   gpc1_1 gpc38 (
      {stage0_2[10]},
      {stage1_2[6]}
   );
   gpc1_1 gpc39 (
      {stage0_2[11]},
      {stage1_2[7]}
   );
   gpc1_1 gpc40 (
      {stage0_2[12]},
      {stage1_2[8]}
   );
   gpc1_1 gpc41 (
      {stage0_2[13]},
      {stage1_2[9]}
   );
   gpc1_1 gpc42 (
      {stage0_2[14]},
      {stage1_2[10]}
   );
   gpc1_1 gpc43 (
      {stage0_2[15]},
      {stage1_2[11]}
   );
   gpc1_1 gpc44 (
      {stage0_3[11]},
      {stage1_3[4]}
   );
   gpc1_1 gpc45 (
      {stage0_3[12]},
      {stage1_3[5]}
   );
   gpc1_1 gpc46 (
      {stage0_3[13]},
      {stage1_3[6]}
   );
   gpc1_1 gpc47 (
      {stage0_3[14]},
      {stage1_3[7]}
   );
   gpc1_1 gpc48 (
      {stage0_3[15]},
      {stage1_3[8]}
   );
   gpc1_1 gpc49 (
      {stage0_4[15]},
      {stage1_4[5]}
   );
   gpc1_1 gpc50 (
      {stage0_7[8]},
      {stage1_7[6]}
   );
   gpc1_1 gpc51 (
      {stage0_7[9]},
      {stage1_7[7]}
   );
   gpc1_1 gpc52 (
      {stage0_7[10]},
      {stage1_7[8]}
   );
   gpc1_1 gpc53 (
      {stage0_7[11]},
      {stage1_7[9]}
   );
   gpc1_1 gpc54 (
      {stage0_7[12]},
      {stage1_7[10]}
   );
   gpc1_1 gpc55 (
      {stage0_7[13]},
      {stage1_7[11]}
   );
   gpc1_1 gpc56 (
      {stage0_7[14]},
      {stage1_7[12]}
   );
   gpc1_1 gpc57 (
      {stage0_7[15]},
      {stage1_7[13]}
   );
   gpc1_1 gpc58 (
      {stage0_9[12]},
      {stage1_9[6]}
   );
   gpc1_1 gpc59 (
      {stage0_9[13]},
      {stage1_9[7]}
   );
   gpc1_1 gpc60 (
      {stage0_9[14]},
      {stage1_9[8]}
   );
   gpc1_1 gpc61 (
      {stage0_9[15]},
      {stage1_9[9]}
   );
   gpc1_1 gpc62 (
      {stage0_11[13]},
      {stage1_11[6]}
   );
   gpc1_1 gpc63 (
      {stage0_11[14]},
      {stage1_11[7]}
   );
   gpc1_1 gpc64 (
      {stage0_11[15]},
      {stage1_11[8]}
   );
   gpc1_1 gpc65 (
      {stage0_12[15]},
      {stage1_12[6]}
   );
   gpc1_1 gpc66 (
      {stage0_14[8]},
      {stage1_14[5]}
   );
   gpc1_1 gpc67 (
      {stage0_14[9]},
      {stage1_14[6]}
   );
   gpc1_1 gpc68 (
      {stage0_14[10]},
      {stage1_14[7]}
   );
   gpc1_1 gpc69 (
      {stage0_14[11]},
      {stage1_14[8]}
   );
   gpc1_1 gpc70 (
      {stage0_14[12]},
      {stage1_14[9]}
   );
   gpc1_1 gpc71 (
      {stage0_14[13]},
      {stage1_14[10]}
   );
   gpc1_1 gpc72 (
      {stage0_14[14]},
      {stage1_14[11]}
   );
   gpc1_1 gpc73 (
      {stage0_14[15]},
      {stage1_14[12]}
   );
   gpc1_1 gpc74 (
      {stage0_15[12]},
      {stage1_15[4]}
   );
   gpc1_1 gpc75 (
      {stage0_15[13]},
      {stage1_15[5]}
   );
   gpc1_1 gpc76 (
      {stage0_15[14]},
      {stage1_15[6]}
   );
   gpc1_1 gpc77 (
      {stage0_15[15]},
      {stage1_15[7]}
   );
   gpc606_5 gpc78 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc79 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc80 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc81 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[1],stage2_4[3]}
   );
   gpc606_5 gpc82 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[2]}
   );
   gpc606_5 gpc83 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[2]}
   );
   gpc606_5 gpc84 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[1],stage2_9[2],stage2_8[3]}
   );
   gpc606_5 gpc85 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[0],stage2_12[1],stage2_11[2]}
   );
   gpc615_5 gpc86 (
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4]},
      {stage1_13[6]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[1],stage2_13[1],stage2_12[2]}
   );
   gpc2135_5 gpc87 (
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10]},
      {stage1_15[0], stage1_15[1], stage1_15[2]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1]},
      {stage2_18[0],stage2_17[0],stage2_16[1],stage2_15[2],stage2_14[2]}
   );
   gpc1163_5 gpc88 (
      {stage1_14[11], stage1_14[12], 1'b0},
      {stage1_15[3], stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7], 1'b0},
      {stage1_16[1]},
      {1'b0},
      {stage2_18[1],stage2_17[1],stage2_16[2],stage2_15[3],stage2_14[3]}
   );
   gpc1_1 gpc89 (
      {stage1_1[6]},
      {stage2_1[3]}
   );
   gpc1_1 gpc90 (
      {stage1_1[7]},
      {stage2_1[4]}
   );
   gpc1_1 gpc91 (
      {stage1_1[8]},
      {stage2_1[5]}
   );
   gpc1_1 gpc92 (
      {stage1_3[6]},
      {stage2_3[3]}
   );
   gpc1_1 gpc93 (
      {stage1_3[7]},
      {stage2_3[4]}
   );
   gpc1_1 gpc94 (
      {stage1_3[8]},
      {stage2_3[5]}
   );
   gpc1_1 gpc95 (
      {stage1_7[12]},
      {stage2_7[3]}
   );
   gpc1_1 gpc96 (
      {stage1_7[13]},
      {stage2_7[4]}
   );
   gpc1_1 gpc97 (
      {stage1_9[6]},
      {stage2_9[3]}
   );
   gpc1_1 gpc98 (
      {stage1_9[7]},
      {stage2_9[4]}
   );
   gpc1_1 gpc99 (
      {stage1_9[8]},
      {stage2_9[5]}
   );
   gpc1_1 gpc100 (
      {stage1_9[9]},
      {stage2_9[6]}
   );
   gpc1_1 gpc101 (
      {stage1_11[6]},
      {stage2_11[3]}
   );
   gpc1_1 gpc102 (
      {stage1_11[7]},
      {stage2_11[4]}
   );
   gpc1_1 gpc103 (
      {stage1_11[8]},
      {stage2_11[5]}
   );
   gpc1_1 gpc104 (
      {stage1_12[5]},
      {stage2_12[3]}
   );
   gpc1_1 gpc105 (
      {stage1_12[6]},
      {stage2_12[4]}
   );
   gpc1_1 gpc106 (
      {stage1_16[2]},
      {stage2_16[3]}
   );
   gpc2135_5 gpc107 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4]},
      {stage2_2[0], stage2_2[1], stage2_2[2]},
      {stage2_3[0]},
      {stage2_4[0], stage2_4[1]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc1325_5 gpc108 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[2], stage2_4[3]},
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc2135_5 gpc109 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0]},
      {stage2_10[0], stage2_10[1]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[1]}
   );
   gpc606_5 gpc110 (
      {stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1]}
   );
   gpc1325_5 gpc111 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4]},
      {stage2_13[0], stage2_13[1]},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[1],stage3_12[1]}
   );
   gpc1163_5 gpc112 (
      {stage2_15[1], stage2_15[2], stage2_15[3]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], 1'b0, 1'b0},
      {stage2_17[0]},
      {stage2_18[0]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[1]}
   );
   gpc1_1 gpc113 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc114 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc115 (
      {stage2_1[5]},
      {stage3_1[1]}
   );
   gpc1_1 gpc116 (
      {stage2_6[1]},
      {stage3_6[1]}
   );
   gpc1_1 gpc117 (
      {stage2_8[3]},
      {stage3_8[1]}
   );
   gpc1_1 gpc118 (
      {stage2_14[3]},
      {stage3_14[1]}
   );
   gpc1_1 gpc119 (
      {stage2_17[1]},
      {stage3_17[1]}
   );
   gpc1_1 gpc120 (
      {stage2_18[1]},
      {stage3_18[1]}
   );
endmodule

module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor_CLA16_16 compressor_CLA16_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae4a338235d05bea7f0c35984eb0727605c349b4ab780a9ea425988e8d7723ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9888e85dc02ebc8f797ad9ae5367d5492f03eef736c13850c647ae1f7294ef9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafd94f593fdfc1cbaae4a24529f386cc2fe7bbdde1a32d32600246f6f41f27a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c6cb50029697efcac13715070b9e479afaece18409eeb0714de561764abce70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61037a6d5ce5ef40193ca242fcd5472377808551be02421bfdb1b73f7325564c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20db865115128c2d818214270e2e7e7e10739c2c7572a1d08c0844b14b31b073;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6b6189cc3b567eb40ccdc07f6bb05cc85acb3317ccadcf2958932d1d0012fe7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee9441a0d34148ae37325657704766c6384f1cf0b266f690e38793949fca2655;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h854cc9241243fd2470376212d4b932a487418eae470452c5f5c9709bf7b305da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6eea7b51e5ebfed7e512e35c8ea42c79bf5ee2b829976a31589e6e4418472ab2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86127f793cc556ccacbea3aec6803dcfd250924dc1facda43cf00f1bc9e2a3b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4d4c4c1d9807bf486986b24a0e259cee3f73f666251f83b2950c72051576ee9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1583d4781bd4346630a84abdcb6bf45d92e54fb6b90da110d1b737ce31c476b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e1b2f612388886fb81ce3989f654b8c3763f2a52af7574520a5e9400c37b621;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44fde58123dbf1ec0d990bb009da7e14aeaacbc8079f72eb533fd75ccf40f64d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h545442cfd5894c997440d6f0962e948f2f0dd5d32d002de2e073bc7325253edb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3771ba6b93b361320242b96178e34c1983d4eb827de21e25c0bab7961c0417a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ddfb19d76d0e70cddec8fb93f0c94a6f4430b2b7ae7894eb1e1f69f9fed38e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd84fe72fa18a9cd856cca790fb70fabc0e01f448f51aadfb0188077db7686f3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83345881aedcdd80c100ec8a1fa65cf32ac47ed5c6fe94c764c92fae8864d52a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e5da7e1661ebfcfe07965def8bb28234bc800fd19c1f593a701cb02b5116064;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1469b38f46067b99da30b83a09aa4a73e3df9f1be8a818ee00a29c3fca934b8f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f6a0b02563f97470a7174d878281e9f06f754001d08894ebe4de7147d3ab680;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha65bd7f2b1a03b352676513b584bf0d8d0671939c6540e612487f351ba631679;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h488275c56ab4fe40f3ab316bb7865e5fa952222f10ac7ed4fc83eeed61e7a1e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83ace5dcedae533ae556d01832a4d1bb2f965ed3fa2c30ba4ebcca85f491e5b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbea09ab226aa2c15e569a3a5652253026a28b4bb40cc81b7d52d94e738568529;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf611130461987e6436db62089e547299a4465a3956ce36d96e9fec5deeaa4a6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8df7f796375ed5f26a4bf8c1e5be181cf8d34849781a3ec446f010b02478bd16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd51da9aee24d12a566e81c3fa04b2fb41eca727c57dd9ed562572fe4b9d180e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d2358ad518bc5503f28cdaef9a1fd10c3995619eb37fde90ccca6f8adc53c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7960f6438c67eb5ced4b27235b3eb7974f23de57202362901dac109ac9bfb9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc86cb26a85762c2cf1c01c235f143d829caf4fa4dccfbee44237d865ac7d1023;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0376925be0af217386e33a3063f473e0d60ea8c875ed1d023e2a9013831601e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h621d24e049b1a78649ce30d61886ccc4a26cefeee2be5439410d7ce478241ac1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heeb493eb8c81e09294853db09c9572e71d2c87acd4caa8aa0c5d7f1f5fcb1ef2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8093c70c2fdc645578f987e54e6a55fdfa91c11398bd34a496d2f3abac48fba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65534f2c628f8bd90f693ad5780a1688fa2055204ee889014bad8bb4f64ae92f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86edafbed004c4a646d707c70fc7719fb1d5bd4f068c8870fdc3a65c20ae40a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ad3d13199d5092a8dc805ec4c9bdad24486aa9a84f93f5ab1884b55f211bf2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h392a044401bae3fc2fae6844208b936e5ed4d4766afee5bfd87c3aa8e6fa4e5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99d93191ef9b5007b401b82eb091881ae6c49f82c84c3619279c0ba7cd37220c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3a68468537ab54e5e8084800559d3156ecef967b39b823da1fbcabcb0a5c2a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0010900042006fa85f15520aac00634576bfc1ba0ecf86f49ffbee53c1a204e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha350b15d25a79d4a1276d32c20f3ad27ab3fc8cf11a403b4fca216b8b705efa4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e7143bed5de172fc39851cbf5e734596d3230f174609e1888ad3e052afeeb8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83a244bcd8d5b1bbfc9889151bc614c6021dcad0e034b4025094e6f81572d71b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed455c867d5c72fef9aed2bc920b14d4d62bc29132d3cabf7cf4740d44e96ab0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha74e3ffb12526d04f838c48be4e6fa6488adbd05e4a11ded401644956fc44192;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf99ebf9b2aebe4a06030b520675071def69e34a429aaf822f903a8c63d79c67d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19193d91909595dd0bc3907c5a97fc6522692e02af163f136b4c6e78f6108581;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ef58b4e4637137842b77d42cfaac1e98932d0011f1f7259cd1088b858bd06c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc273a71fb07d0a3dae5179dcdbf138efab7765303c7414050bcf1c970b0ff5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fca87ed618535bb9228261d1ab4d93d97941e91f81c0cdb5726bf4c76262313;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha59259ddacb2b0aec25579337c9eec9c3b0bab5babbc924b89fdbe455607a80e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc534a39ec56daec2895c4b950ea47d576260997a2846736658136091c48c1bbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h463f9395dde24ddfd0ea8a4cf0aeebca9112d56396a89974ea0769afa2cc350d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9c5542b23c48b5bec9ab197eefac4e5f0e1b0a19d2717ebce3d946797ed9348;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e15b6de21c4a36eccd91b4a73546a36c71f318cf1a155e6736f007996b680c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h472d6f41f97835ebbd32db5a965b4701fb5437ff0403f94724c85a84627e3bd0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb981f1730c7e6bb9a15c8e9d2558ab7d342c66f00b0c16c837a460afea50dbd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a5c98f659e32270df9ea4bf102615777d353873d14da5553ccc51699fb752b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae03deb178466d13b6407c6b12fca9a46c46913c2a853f1a0ea71bbfcfca591a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8411fa23ba533517989544caf322f12e50e80d365ead6efd08c3895dcb12a40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcecba8328572b5f678e0b087afd27133f015ecce60a3ab3395640c3654d30bfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c3dede26dc4e4234bd371786a74da17d2a42ad0d4130fc8b0a23e3d3e1328f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5bce09160e24af38010f96811b7b8ed2998d1c2be5a9820753e0ff819f02923;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h582e58d09019d85eb3ab71160013f8fba13592dabefb8899c6ad5b788a8432cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8279aef08cec68b6d74abd1889ba95dd09af37d5725a825e5b61efd9cba645b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h322c5f0856f8d831b07cf1968e458215ee22b1cb1fa74266cd6baa917ce339d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5b9925db07abce2f8c422bb3c620f52593a0ec7ce598057717a001c6f7f9653;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h337194ace210fbb9930f305c3ddc2a5e0972a0219ed3b0e90c9e5cdcd92a238b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1855957c2afa7b9e0a28a0ef7ae743999baac33d891b57aa2665fc28db9fdc8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccb748d1cf89abb974f916718f33f3bddd6949c319a871d66dbfde04833e97af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf134d753cbdb47a2cb53c24726726d7ed0c1277b2e0d13e3e13d3607355b8925;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98d207b5916c8706d00552e1502309e2805102148e919446381604c1a3665560;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c82a35c068dbff7819355cc9c7a02ad150f96b38acbc299bad16c578ae9998e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d4e2dba207e30f398435acdc64a3b270ed070b0ea38169f16a3c0f81b1a68bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4fb209444e7bc7109bb7ffa40a0c34777c958865492949f4fb6303d6d8124686;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d460876955e0b24ec5959fe9a09b88eac01cc3ad3226bd9987b4e0003bcff1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79e0c15be2961bb0ca4c370f39a49d1f571303c96485efeed440ac3d9d2719d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef725b9e5e656e0038fbad99c4c7d5622c55bb526d7f402aee4a9e382b6398d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc86efd9a6326033902752252492b6e530154226cb4ec176cb8f7d92bb1e244;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca7e228b14882bc39e281004ca7f5ce54111cef47bc730fd544d60ecbb809e19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc09ec01ce3d478ce7b9246b85d60e79216f7e1d98fe27ac11005106264fc3dc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38dd4faf12c4d7ab468d85d56d00a1558b5f0381885f93e165dbea984a145fd0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6955961a67c982c1389366e4c4aa94d8fb6a2dd40d8c731f15452ea4a9229c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h133d46903afcc5ffa64609ace2046353fdb598e4daf4f9ea41b1638bea6f44ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe8cf50a8828c1b9fd7004c338d8343e00f3695c8591eafd481de627bb94901d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f9891f48c8dc730b4052fa8d59b76b064b1f0262dae3287db23a71c109f516;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94d87fcab32903ed53585ccd925ff2197a7b13f4629088316bf9e56faae6be2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58c5e9c15f53549266d1070f2e5024efe3be81b5fcf7f23da12efc59cd30222e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h833f0a585c478ca993383d860d48a891904a7cb0e1562a3d1d434b7cf288a849;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4698357f74097e0080a35ffdd194f2b70e546e7b57a31cab6313c549447fa8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb33e3fbc8a2190eeb80b595959d093aebd1ec03cf23f164ab58f07f41cd0a98b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5c7aa1217ed40c9b2df9e1c298dc7a7e376113999a4b77fed0c5af624f55d5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h796dfb083cfb1e14a90951a3d42da9d27c69be13ad62e4f3f5cab3815f9ebfc0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6724af7b20f5ffbe47f2ab16a924e75a712c0453c7c858d7e1a3758b1d45e0c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfaa522a162711301b55dd9862ffa3ffe3f23fd5209d56669cfb28c1d2b5aa287;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7ba4227bb0ab331236047a0bb109f8fffe21e633ce074c73246ae224ef30e79;
        #1
        $finish();
    end
endmodule
