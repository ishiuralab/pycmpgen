module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    compressor2_1_16_12 compressor2_1_16_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor2_1_16_12(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [0:0] comp_out13;
    wire [0:0] comp_out14;
    wire [0:0] comp_out15;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15)
    );
    rowadder2_1_16 rowadder2_1inst(
        .src0({comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [0:0] dst13,
      output wire [0:0] dst14,
      output wire [0:0] dst15);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [6:0] stage1_0;
   wire [5:0] stage1_1;
   wire [5:0] stage1_2;
   wire [7:0] stage1_3;
   wire [12:0] stage1_4;
   wire [5:0] stage1_5;
   wire [12:0] stage1_6;
   wire [6:0] stage1_7;
   wire [5:0] stage1_8;
   wire [8:0] stage1_9;
   wire [8:0] stage1_10;
   wire [7:0] stage1_11;
   wire [3:0] stage1_12;
   wire [1:0] stage1_13;
   wire [1:0] stage2_0;
   wire [6:0] stage2_1;
   wire [0:0] stage2_2;
   wire [8:0] stage2_3;
   wire [3:0] stage2_4;
   wire [2:0] stage2_5;
   wire [3:0] stage2_6;
   wire [3:0] stage2_7;
   wire [4:0] stage2_8;
   wire [4:0] stage2_9;
   wire [2:0] stage2_10;
   wire [2:0] stage2_11;
   wire [3:0] stage2_12;
   wire [2:0] stage2_13;
   wire [0:0] stage2_14;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [0:0] stage3_13;
   wire [0:0] stage3_14;
   wire [0:0] stage3_15;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1325_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_1[0], stage0_1[1]},
      {stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage0_3[0]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2]}
   );
   gpc606_5 gpc3 (
      {stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3]}
   );
   gpc606_5 gpc4 (
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[4],stage1_3[4],stage1_2[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_4[6], stage0_4[7], stage0_4[8]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_6[0]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[5]}
   );
   gpc606_5 gpc6 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6]},
      {stage1_9[0],stage1_8[1],stage1_7[1],stage1_6[2],stage1_5[4]}
   );
   gpc615_5 gpc7 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], 1'b0},
      {stage0_6[1]},
      {stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12]},
      {stage1_9[1],stage1_8[2],stage1_7[2],stage1_6[3],stage1_5[5]}
   );
   gpc606_5 gpc8 (
      {stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[2],stage1_8[3],stage1_7[3],stage1_6[4]}
   );
   gpc615_5 gpc9 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10]},
      {stage0_9[0]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[3],stage1_8[4]}
   );
   gpc615_5 gpc10 (
      {stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_9[1]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[4],stage1_8[5]}
   );
   gpc606_5 gpc11 (
      {stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[2],stage1_10[3],stage1_9[5]}
   );
   gpc606_5 gpc12 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[3],stage1_11[3],stage1_10[4],stage1_9[6]}
   );
   gpc1_1 gpc13 (
      {stage0_0[11]},
      {stage1_0[2]}
   );
   gpc1_1 gpc14 (
      {stage0_0[12]},
      {stage1_0[3]}
   );
   gpc1_1 gpc15 (
      {stage0_0[13]},
      {stage1_0[4]}
   );
   gpc1_1 gpc16 (
      {stage0_0[14]},
      {stage1_0[5]}
   );
   gpc1_1 gpc17 (
      {stage0_0[15]},
      {stage1_0[6]}
   );
   gpc1_1 gpc18 (
      {stage0_1[14]},
      {stage1_1[4]}
   );
   gpc1_1 gpc19 (
      {stage0_1[15]},
      {stage1_1[5]}
   );
   gpc1_1 gpc20 (
      {stage0_2[15]},
      {stage1_2[5]}
   );
   gpc1_1 gpc21 (
      {stage0_3[13]},
      {stage1_3[5]}
   );
   gpc1_1 gpc22 (
      {stage0_3[14]},
      {stage1_3[6]}
   );
   gpc1_1 gpc23 (
      {stage0_3[15]},
      {stage1_3[7]}
   );
   gpc1_1 gpc24 (
      {stage0_4[9]},
      {stage1_4[6]}
   );
   gpc1_1 gpc25 (
      {stage0_4[10]},
      {stage1_4[7]}
   );
   gpc1_1 gpc26 (
      {stage0_4[11]},
      {stage1_4[8]}
   );
   gpc1_1 gpc27 (
      {stage0_4[12]},
      {stage1_4[9]}
   );
   gpc1_1 gpc28 (
      {stage0_4[13]},
      {stage1_4[10]}
   );
   gpc1_1 gpc29 (
      {stage0_4[14]},
      {stage1_4[11]}
   );
   gpc1_1 gpc30 (
      {stage0_4[15]},
      {stage1_4[12]}
   );
   gpc1_1 gpc31 (
      {stage0_6[8]},
      {stage1_6[5]}
   );
   gpc1_1 gpc32 (
      {stage0_6[9]},
      {stage1_6[6]}
   );
   gpc1_1 gpc33 (
      {stage0_6[10]},
      {stage1_6[7]}
   );
   gpc1_1 gpc34 (
      {stage0_6[11]},
      {stage1_6[8]}
   );
   gpc1_1 gpc35 (
      {stage0_6[12]},
      {stage1_6[9]}
   );
   gpc1_1 gpc36 (
      {stage0_6[13]},
      {stage1_6[10]}
   );
   gpc1_1 gpc37 (
      {stage0_6[14]},
      {stage1_6[11]}
   );
   gpc1_1 gpc38 (
      {stage0_6[15]},
      {stage1_6[12]}
   );
   gpc1_1 gpc39 (
      {stage0_7[13]},
      {stage1_7[4]}
   );
   gpc1_1 gpc40 (
      {stage0_7[14]},
      {stage1_7[5]}
   );
   gpc1_1 gpc41 (
      {stage0_7[15]},
      {stage1_7[6]}
   );
   gpc1_1 gpc42 (
      {stage0_9[14]},
      {stage1_9[7]}
   );
   gpc1_1 gpc43 (
      {stage0_9[15]},
      {stage1_9[8]}
   );
   gpc1_1 gpc44 (
      {stage0_10[12]},
      {stage1_10[5]}
   );
   gpc1_1 gpc45 (
      {stage0_10[13]},
      {stage1_10[6]}
   );
   gpc1_1 gpc46 (
      {stage0_10[14]},
      {stage1_10[7]}
   );
   gpc1_1 gpc47 (
      {stage0_10[15]},
      {stage1_10[8]}
   );
   gpc1_1 gpc48 (
      {stage0_11[12]},
      {stage1_11[4]}
   );
   gpc1_1 gpc49 (
      {stage0_11[13]},
      {stage1_11[5]}
   );
   gpc1_1 gpc50 (
      {stage0_11[14]},
      {stage1_11[6]}
   );
   gpc1_1 gpc51 (
      {stage0_11[15]},
      {stage1_11[7]}
   );
   gpc606_5 gpc52 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc53 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[1]}
   );
   gpc606_5 gpc54 (
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[2]}
   );
   gpc606_5 gpc55 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[2],stage2_6[2],stage2_5[2]}
   );
   gpc615_5 gpc56 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4]},
      {stage1_9[0]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[0],stage2_9[1],stage2_8[3]}
   );
   gpc606_5 gpc57 (
      {stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[1],stage2_10[1],stage2_9[2]}
   );
   gpc1343_5 gpc58 (
      {stage1_10[6], stage1_10[7], stage1_10[8]},
      {stage1_11[6], stage1_11[7], 1'b0, 1'b0},
      {stage1_12[0], stage1_12[1], stage1_12[2]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[2],stage2_10[2]}
   );
   gpc1_1 gpc59 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc60 (
      {stage1_1[0]},
      {stage2_1[1]}
   );
   gpc1_1 gpc61 (
      {stage1_1[1]},
      {stage2_1[2]}
   );
   gpc1_1 gpc62 (
      {stage1_1[2]},
      {stage2_1[3]}
   );
   gpc1_1 gpc63 (
      {stage1_1[3]},
      {stage2_1[4]}
   );
   gpc1_1 gpc64 (
      {stage1_1[4]},
      {stage2_1[5]}
   );
   gpc1_1 gpc65 (
      {stage1_1[5]},
      {stage2_1[6]}
   );
   gpc1_1 gpc66 (
      {stage1_3[0]},
      {stage2_3[1]}
   );
   gpc1_1 gpc67 (
      {stage1_3[1]},
      {stage2_3[2]}
   );
   gpc1_1 gpc68 (
      {stage1_3[2]},
      {stage2_3[3]}
   );
   gpc1_1 gpc69 (
      {stage1_3[3]},
      {stage2_3[4]}
   );
   gpc1_1 gpc70 (
      {stage1_3[4]},
      {stage2_3[5]}
   );
   gpc1_1 gpc71 (
      {stage1_3[5]},
      {stage2_3[6]}
   );
   gpc1_1 gpc72 (
      {stage1_3[6]},
      {stage2_3[7]}
   );
   gpc1_1 gpc73 (
      {stage1_3[7]},
      {stage2_3[8]}
   );
   gpc1_1 gpc74 (
      {stage1_4[12]},
      {stage2_4[3]}
   );
   gpc1_1 gpc75 (
      {stage1_6[12]},
      {stage2_6[3]}
   );
   gpc1_1 gpc76 (
      {stage1_7[6]},
      {stage2_7[3]}
   );
   gpc1_1 gpc77 (
      {stage1_8[5]},
      {stage2_8[4]}
   );
   gpc1_1 gpc78 (
      {stage1_9[7]},
      {stage2_9[3]}
   );
   gpc1_1 gpc79 (
      {stage1_9[8]},
      {stage2_9[4]}
   );
   gpc1_1 gpc80 (
      {stage1_12[3]},
      {stage2_12[3]}
   );
   gpc1_1 gpc81 (
      {stage1_13[1]},
      {stage2_13[2]}
   );
   gpc606_5 gpc82 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc1343_5 gpc83 (
      {stage2_3[6], stage2_3[7], stage2_3[8]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3]},
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc1343_5 gpc84 (
      {stage2_6[1], stage2_6[2], stage2_6[3]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3]},
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0]},
      {stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[1],stage3_6[1]}
   );
   gpc1343_5 gpc85 (
      {stage2_8[3], stage2_8[4], 1'b0},
      {stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4]},
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[0],stage3_10[1],stage3_9[1],stage3_8[1]}
   );
   gpc1343_5 gpc86 (
      {stage2_11[1], stage2_11[2], 1'b0},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3]},
      {stage2_13[0], stage2_13[1], stage2_13[2]},
      {stage2_14[0]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[1]}
   );
   gpc1_1 gpc87 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc88 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc89 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc90 (
      {stage2_2[0]},
      {stage3_2[1]}
   );
endmodule
module rowadder2_1_16(input [15:0] src0, input [15:0] src1, output [16:0] dst0);
    wire [15:0] gene;
    wire [15:0] prop;
    wire [15:0] out;
    wire [15:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    assign dst0 = {carryout[15], out[15:0]};
endmodule


module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor2_1_16_12 compressor2_1_16_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4b8c37c2387681af157aa45860f5c96116ee4dd4bf1e8c49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h57fd3ebe3fed1bc9899eef1b2c07cf5eda27931f1aa2d2c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h202144ccb8690cfb3b5046387869d6f4176cc5b8d9271ee2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc1999c6dc9fe4ff28c4a5528c5b841f0023469004165c4f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7c4b5c73ef7409df9cf148ffe4297b2afa2d18595ff9f813;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h82c8c0823f39fb612b89b6b443221b957121d37c728dc54b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4d90fd28f35371d9fbc9bd721d3764fe1326f469eb45bea0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h15bc5d2b4a4f44a24d19f275eaaadfbd0c57dbe07029c5e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hf78f50e825cdd126fce06e47b4edca399899ec45c96b0996;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8caef26d3c8a9fe9485dfbf9d645569b186c84d971b943e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h18edf83aebf7509c5683d560a632499ed9f30d44a89c355;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7d3f0387cbc1e5e6972d65023b8fc8a12e8fc9bfb8d316b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc5b6a6ff10e0fbc2c02fb4eb777c9fd4102fae5dca86dd80;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb73dd432ebe2eeedc84a83c17a017ad5a5df9e225457b239;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h45cf8ef73fcae1c2342f4eea251c6b56c07364be50c4cbd4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hfc9bb15d5f71d11ad37ca20a453a47dc59e461492ea41d25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6804724480c3e5b00413d882fbe768adaaf607a43a769864;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h201fb032df910d717fbd5053250deda7bf7a6a12f103f84b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hf5ee829cc5c910c66092162ae5c88baac30d2dc7fe4de406;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha884ce4d42a1b9a88747823afb20a694c4e84ff5e968857a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1786416e70e98ebe98e6c1210a7c0b9415e91a295cf47943;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'haaf1056577555fb9ae4826f70b6c7e4635b2479ac3ee11ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h11063866d4ae312253d35755f93464d08a01248b3b045b54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb83ee7bacc0051f58489bd0250313b15067b0afe043cd52a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7a2fd72b7352ed27d69c94a61d1908aaf051ab4f83bc45d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1dd68f95e92faeac7e86acf130f9f08aeac1c40f721358b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8dce9e8b490f12ab1139cfb9892644366007975b02698edc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha58de3cbc31a45f385f9ba97f8b29189dbeb41312edddcb4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb23c156825e005d608babd1fa7dc77dd6ce399b7f3914def;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hec72ae97ce8a54a1e8ec82093a1012d84419661f02b20080;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h2fa0f8c2b126a46cfa78e4eb929e21e6981febfd7fa76662;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5b2b3c232a995dadf9ecce06dfacf66facf608e9f1253ab3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha74f610147f5282a87cf21da5b9d990738177bc6becfcc96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h98010148ba7abbf31489f1997939dedcb93ebf1e90cf3b93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc8c18c54707d4e3181d09f64270954055a8c2209ff718426;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h22ad95de201effcf5ab7bebbf65b67df072b210a2484c7b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he820ebb0bf3ce43527fd849948be90e608837577bf4edf2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hcefb30ff8790edc0db4a1c65ebf2b37b733ba39f91d4d0e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb11d694096d58be76f56f8823838ef6e69b6ebd674cd45bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h11c94cad7958f30f0ca0d0ff6d1f3d693b3488f64e443212;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8ad5d5b933948cfd8b0f9937d3674af82bb565875286f9b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5f81e7f8a580c88ef1b2f510e209ae057d850a0879bb2c82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h2a190648da3177eae79fcc19c82bd3f593d623856a574365;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1a293a53279cfd78eebfb9d0c91035527322bc6e1d102263;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd7e25fbffcce28c66c41e505ff8b799c892dd15c669671fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4d605030acd168137205f028ac59da82f70d6484264e0dbc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc79715eb7e8f2a6d00c0bbaa5ace667d24c94275fe079d99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha35184c408da3c5b5393738dc181dd931b4aec8a58cee5c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h57c867190f43328b2ed1ac8eac2a23d89124527addb84133;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hcab94f215b122dc593ab69a28b077cd7d510ad2e422b9fae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h232a52a18e93ff574347f2466392975f6a12310b93b58d71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1b7ec02976cd5848341dfa18b6c0c00db45e9fbff027e2d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h77a8a1711a9d82d3de3728b3aa58166223854b12eb21f185;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1f431222a579f95e44196b0891a1d0d618e7ebca01f40bff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h567de30f780a696a047a5e94ad18f2edf44d22028a895bbd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h18d517bac754d9b1703a098ae8196d98fb9a9e9b6a70aed1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h29cb0a3ce7f74836fc16c94a47119d210cfa13c8bbebe0c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc1851f227a5d12d189c281191814c9e6c04613b17c8a083a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha85d29136da7e6e19bdcb04e0982dbdd4f5e048aa3101494;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h41026a92f6d948c1242cc9ba9177870a733c15aacb70a6a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha1961866437ab5a89b949b29112d0081301fd07e6be47dfc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h569e2165212e515bd54838229afa25fc3d17dc3387f8ce06;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4dada4be956f3a962fff4df6ad0d7d0b2340cb881ec3f37a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc2fa4643ac189d9bf01a4dd0f87bfc7f7670afb8bc967aa6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc0354d9c6d756b759e7b4a7fcbc1eabda27ca16bf659cc6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd7cc6769a7a82059bcdb354a8a49451bccf0c854ba116315;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5e0ce0944fb8182d94f2827ec7499fb5cd41c829c1139d5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h3690d7ca620e5d2651e9f67957030fd19de50b9e762caef2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h2e47cbb685b04ea5d0d0ec20d23141b125c11236996df5bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4c3e92beea36c568b34144b4a4b6a919bba9178bda47f3b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8b142ad95dbfbe7c3c19b6942a8c2c9e2b1f8b20c984d453;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc97f7440c73bcb051fef1f29aecbf0d9fa5230d8ad8eb51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h85fa1928c2ee7e2621de721d0bf6071eccb975047da0b800;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hbf38dee3d16cc15f98d21f661a6e3c1ee71728ea0c538413;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h10078439f1baefb9863c05a2b3da299f812a3df32f531c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha677bc49145f189961ee853a7f0b5154238725c9edbdad2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hbbb38c0ef7a82fce2618007dc5aaef9fbd96f5f0a3fcd9b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h96857916ee8cf9d6933f06b412e1f277751852f9da2fdfba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8fb4bc15c3fa8c0b4fe206abaa528b35d13703f0a8a66742;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5573149914fc84ed7f86bcfff404ad0e00195e7241253d1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hcd740e48cece2a4b8e7788e5bab2550d87d3e868a4d04745;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc453ad5daa66ab92cb23062a339abd54a76cb0dd08e25684;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd50c3d762ceeb4ff8b5a818d7a646080f9ab43d46ba85ddf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h36a0661f28645d40eb72cfe719f3b7372866ed9fc4732620;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h63ce9a34007341203e7b84b7f2fa5852b3b15df878c1bf21;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hebd8a099e92270a409cf035d865c04467e5be4a0f34f2d2a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb33bdc4cff9fff05db0c3edd92a3a1dd2473af103fc5852b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha1fbb9a4385676c16419ad02b371e7ad26583e4611a3e1a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h44e861254451ea6693b9c20a85d92c8194a6245ea38a76b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha324bdcd0b8b63f9921e78e0e6f783fbb12d200ab33cdfff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h81036de8008d1dedf27dd570a19cae2a3df747d213a135da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h14e2070b076da2094ebcb0cab61bc76cd6f255ce34eec438;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h54a32c6a6a9ed3cdceced780d0eb99486fc8f4e644d349ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd9e2bd97d32c7eb6a57647db6d19d8d7d78588f43065244d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd747d2c137726eaabf812aae5e0edf1b35ad1bcc450c0aaa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hdc7638a54bbf9189d077e8f43944192b5fb02d815583bd9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h799d06a5a193732636f359242ce78bc169baef62215d2375;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h53af867e5faa5bb77809d6dd0154c5cd5f670bfce2376a90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6b34fd1dd62cae3ae7d844c51fe3b4e2b3499de41e8fdb23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h56102f40783e50178e340af9809212f5c97d1d569bab6734;
        #1
        $finish();
    end
endmodule
