module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [9:0] src11;
    reg [8:0] src12;
    reg [7:0] src13;
    reg [6:0] src14;
    reg [5:0] src15;
    reg [4:0] src16;
    reg [3:0] src17;
    reg [2:0] src18;
    reg [1:0] src19;
    reg [0:0] src20;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3])<<17) + ((src18[0] + src18[1] + src18[2])<<18) + ((src19[0] + src19[1])<<19) + ((src20[0])<<20);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffffffffffffffffffffffffffffff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec89c6bd3850056f80d719075e0ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e527590e91ff6b61c281b02a8943ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bb638817290ae2465dd7bd97f6f20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h613735db9f74bc6dbe38c89d301572;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1db1c22e427101a517c46a2b3ba97da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h98ec2419de3450d7bc864de830a95c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6d7f6ed4ba13ff7044c3f7b3748636;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde9b507b7ca7f74b5514e383893e91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b05b447b6a625db0d738c870e9805;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15dee43549851997e16730a88d20a64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1864cf0c31317c8c39c14be58454eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10dd656f04ccbe4fb82310e87862a81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5bad48d63009071c02d967b2453269;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fb7b38f8938c2693b71b2f57883585;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2bc03e982f749ea904771835f05465;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d1544362cf83a407b77442018c7db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1028520e0604d7078cf8935933321b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f57f7d6adfbda9f848f1e2e700ae7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd32e02c999bac7383c8a92cd1a651a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17ae858c0e9518ca6895724eee367;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb6d6d36bc9fb54510e574d6d996f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he0333a2e51566ebb68acfc0c5973d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ff822115a7125d1eb51bb1d2b45c5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2dd327a5fb626c6ba2f08cdbbc5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11776597adb75e6385a56c00a1b2b82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f5348f567521b2b09b43167c92e2f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fbd916e4f1ef31f5f1401cb18163c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5bbd37cff679155ce57711c9024139;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1198b82069191cb797d879bb2a46a3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df3a0f071f93a3ab41eaadb1d564ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a210486ea920015cee20b4e014ade4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd21951b6d29e78d12f9eb1b6e02e81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f187d03ed8208a115e4ea9f449361;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ef4fdcbf04c2d6b9a565086b59eda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc6ce5f39440986114d91ad858c9f25;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118b6d0c6c0ccb715493a980eb770ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e84b4937d6f26ab2bf9eb654db026;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h165a493f62bc1df612efc6f381b6449;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7fec2590800a5148d4de547462751;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd01219f605a6f72877d909741157b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1376251d9ce737b7fa18d81e0af0819;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16026faafae1bdf1ce938b13c84dd7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1666cf72491c502990c71ab6b69149a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb6266db61125002219815270467b5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5b33f3688584176e9b2613c1dd8ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae74a4bfb99c7ba23478fa7673e0bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8bb78337bfc7e76462dc5cdb441f88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1441b80f17d80b1e99375b155b3763f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h650b09a4591abf279fd319266f670d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee1d7cdf8915daf79343ace6c1f479;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d751347b442af98ea89e99db22d1e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2eebffcbe8242bef54b148a4f0ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7deddae4127f98d874586da9c9bda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b5916760687fcb46b7cd2b4191e59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170d60302943dfd124b8f3e0d6585d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17ebf3baf37421976f1c4fd15a5f74a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56e5ab1b69454870412a090216aeb2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he9b8303b7198a4d599005005ecc86b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f75e42adbab3646e40c6e5fc7470a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3228ce0e1f45536f5ff0abb914c671;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e58d1468f59421b8814efe6341ece1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h220dc38683a8b587d5240363a852e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8a253c9ab59b31b3aff17cdab7ff68;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h52680e7f13a1dcd37b078841588e71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6b80e54f873e031ef5cee8bbb8291;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bc1571fa62b590a4899865101110cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bf955b08fd064acb96b2098ce7b1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a33041f1d689fad64a015f39b43b4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43c23178df0bac98b11ae4047cea05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h110ec0fff102b3e025c07c4b123ad82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d8c5077689df2ec2c1640a81b8e9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haad8bcf3c61f9284de02bcdeec3b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30c23738fdaeb07297c73a2be14184;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h57cc1ac0891383dc196378010074f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h939a4e5f058509441cb4621cbacd0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107754e6657ca6ee3f0d8915d24ce6d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1ac152505131aa6e99a05ba73c33f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6342597e10c40d6b9cd1d6ea8dd06e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9ec886b6a545b44dc535332aa90efa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h155a4cb8fa327c21929955073cbf06e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14d8a70678e70ec7ed753b474673ef4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1672d46c15b6120eb55d1c9549eb9e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h174c274bd1d7e52ce48723d63075bce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b706d90456b69a6ddace31b5a8481;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e9812ac77b15caefdb394f14857ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a04a2dc424055ecbec15795bff275;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd132c84144778b5d3779a9f516516;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d945c46e22a8d52260eb127a05496c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134a1b4ebf182c90d94492859f89269;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7785355b4d72cc97e77116723b34f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5063cca8edc2a8c2567cbc82cfe0a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1238a23c856523477a5fc3892ec4b87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd0a5868375fe9896d293296543135b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60444bb44cf0ed1661e9f6d8f9d878;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111e152ab2498cafd60d26d1ec1995;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e348d88490dc1da44c93a70d511df9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15efe7de609b34cd6dfd6c4654926c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f97989295970613f0734e1f9d9180b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc0089d0059bb1ab18cd6645515ab2f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1790ab5cbaf0876af2940d9a91ffe69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16683f3f220f5485dc814f2b86888d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb6cffa5eda9d039e6125eaa15343d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3185f32c1f05d8b7862123d4aa4eec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2cda1e4388ae48cc5e572bb7fb47a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47a0e192874e8cfcf3d2cec4166f5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h21e8747653980dd966671655aa0b8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h64ebc559e93cbfcd7197b4eb4fc22c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b18e22e7dc3a55be28979f3bb4ff3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h186697a1309df43cc5befd79623c870;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173dab88338f2acf278ab394d2bdbcd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1489a1f686efb4cc1443eee361ca5b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae808f8e7df6ade00c63785e78dc42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118a87e24e312da90edfee3a39b4a36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7e4c2764d668509584ecf4c3015d37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdc2ace28812610cac5b304ee618b16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1627641659e5a5fcdc1ed444d59a23e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182ce5407bac4bee3467658a474f739;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h320677a0f6c78049c1b2d58c171fa7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f307ebbbc81c9149c8dabbee226ce2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h822441b909f05308c0574a9dacf352;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdfd7b8deb57c4d5b24e4caf51f6b28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h765e386891a9c6ab15cb65fe890433;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16fa7bdfd49f818fea3d9d1256b7746;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab7bf9aebcee46018f52405e0e662b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7abec5c3aa9b5fb27dc3152061274f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b3a63aa25fcab7611e44c95f98ba2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140b7c33df8a128951ee1b1ddbf7e9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9dae68a94e365f2cbe7dfbf720704b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12dd45850aadd2d97cccb375c79e96b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ce064b94fedf087ef26540bff1dcd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hedb39350294904b4b994028938054a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa18029386d6d4fd298893debde92a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17bc05291fa15cb9fb653da1b81639c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af3a8afc0a34046b5d4c8687c701d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c9a6e92521053755dfaf38f5ae0db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1556177b7731822bee903384249f661;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176f4882ba1b720ef4e6c2c3372d24d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc76a7536cf62585f28d8e4b793e0aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a3c668ca1653af41095e00de9e0ebb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18d105c530c3e5d8b4c8a5cc28bf3ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ae299042d4d9c759a1003d2b2f746;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae462cd5a671e2f6a5cc7b788cea7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h195358dffd16945dd9d762acf483afd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156f5fdfb56abc3f38fba907356fae2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18aa9e772f99b864e7ec87694f7d9a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd924f6cdb0302f0f8d8a4ec857849e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0afeed9c0f484de5d042e2fb5324f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h99a0238bb35926b61cb01519b57568;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124abbf4f5a83fe298c0b1d0eebeb6b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdc2984e22b8a3743694c0f698dda49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h359fa51b8268a3d53df9a796af7963;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5c1beba213c55e32ff8a6092d2c42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41428454acaee7e018ac063c951b87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h85ffe17843ebe398c0afa128ffea8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0f93dc5c39c9562bb82da7b92de23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5ac64bb53594194c7fe00da3bb331;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c93c34e59ca089a84846b6e79576fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1078d559961f8087872a54fd3a0213d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h151053a5ad44163ba2665f6a35db77a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15dbb0cbf563d1c807ba27d08ef6142;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h113980ad1be602426a7ccbfad7a1218;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12198b427cbc713b11c9576668242d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h155d5b712acb1f7605646c41af7c486;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hffb6ca49040eaf15728bcf77dedd93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1485a4b55e0dde80df7a81417c586d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb31d5d68778b1ced0f6ef499156aa1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a009c233811b6866ead4f5aba4d1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d4135274d3d4a7dc346b62496e5f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8314d9cfa37df5bebf83306746ca1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a80d911a3ddc10e75db0a314ac9fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ecd0753e254d69f918b0c6c4c074;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be20dfb7204fe6c940faee416bbb51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha485e73dec29483dd742f2d2f5c496;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h569fc44eb735b654725bfd415bf5b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1beca3564c5a4756f6fde5024295418;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8fe579353b5738ab84e5ef6f8d72bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16fd686ff36d73e4fdc15fddc8dd437;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138172b2c6dda9e31d61dea6b2b3674;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h94693fe46644f5c38a5beabcf99b9a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he3eb733c306910682ecfb1e01a39a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3ce7787e4d3ce69a4d8aca792798ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcca1a6f1ed7d3053b92b61bd2cbc8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ac13bd9cbcc817ca4d886730ea832;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9b892845a99bab19476e232e9350be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6b7b28b28f41db6faa1c45c6bf1e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112998a0f352025a41b34073f9f8e26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15dc96f7b1c9321a0840dc3a51a796f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f6c24f709e31276e30642ef6f1a17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h74e0f0c1bd94f76029bbf02cb2505b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h986cca0c4f41f943dacf4ef760d4f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h980006fe52bfeef41513847a437cf7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1363ea09abc512ee31661c0181cbddb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8a8ad96125d5c90677bb8ae4eae27;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3641c27ca13f7a051900e2beeb769b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haeede6d97bf86f6f170b5e64a8d877;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4cd7ac0535345df84fdd245a0bc24e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b4ba3a9067d269f88024f8c92638e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167159c9c5a4ffa4d70e5a87843370e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed3a8ea2109c4e2f0d1a079f11bcf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf096af88387743d37aed7f61d9a7c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha715fff0f5f0d45b3e9aebb40e65e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17057c06b8b26b802aa1c2d504f0d0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5dd2812dc277193c51fb83905dbc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h846ff6bb9d35aa4f45e192f8f31412;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10c72c0dec30940d6d318bd01be9689;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f7dfb7b0074613b32981d67c574a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17aa74d479192d7a1e339ff7dd08f88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb27f76b3739cdf2131d25f83421532;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75449f296d6a7f258f94d78fe2b591;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1826d005878ecf9fc2351590666d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145bacdcbe0f040a771995317af2d46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26e77f5009640a347139ebb2231fa1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1a5c5a13dfd73e7d96e327b621d0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h49cdf5b50c0f8aa4c4a07d0bd4379b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b53c3c8b8cd500df706ad8d467efb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e83d1ed0bdd67069b48e8977ba38c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h739925d13dbd08811e82a503660ab3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92a12f69b55dff0a3c4566938beef5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac4bfd868a7c78bcb79f12a2e14ecb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1159d197421103a24bbaf3f5873a23f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba518b9ec87d9b24a0887b2df169f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbef6c06cf0bc006e81be43eb83fe5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h388fbba84239ca6bb6ba99510b04fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h37ad63228b55a6714f8d1f32525ba8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d983c1d1b761e7aff8a400920f578;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3bed9132091b20c5d3365e37a44f07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e320489c895b1d7e1e418172f7a9a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2e3ad32c0c81ce121ce5403bf8ee88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a35fd49f262570bc268448b7c45c7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2aaa1595c6f9aeb6240f97fddbe254;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10c5fa0a35586d3fb1ac3238f86a353;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2e64df5aaac627bc2959d0d4d4a916;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1273647389a656e89e65e7ad15b1509;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78d32e74cdbb8b549442f66cf0c501;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h70ad8a0c04057e679d0021dade2d68;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107d095cfa525dbac277213958f8a7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60b208e5e88ed6eeda34dff457d2a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe607adcf285e84ec8027d57cca0e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he539f51dbf1cc583769968fa6ce23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e660e447840436e85046a2e259ba9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1106712049e642f906821fb30d09db5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c22abfd4cbd2ef842a23a45204477;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6ad68050852aa4b39bf213b454d47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b3b2094e541999a0934dbd53a93e4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he38f3b11694571757c2024b8375a2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb2fab3c455e56df8eead0954e255d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13fd40c924ed2438944906f83f06dfb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h84d54582540fc86d689cf733926b4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f2e366a93aac6ff5aec31d16c49371;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e0d17ee1acb1781561b82db885deb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h410de08e857a1946ba5a9283bf7ef9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1625facb866e115fb8df1861d7717af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1121023e37c29825a1fd8f66eca335;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17ec27e584f42981f97a398777b5719;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h702ed69d4cea4327403488d139fbe3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9b1c115a54b0c661ba85e8661d6d96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82f5a5b475d763b03a66291ce4838;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b878a0e8b3871e2fb340a56fdcc5e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4dc01ae2ab104b4f0140dbf6201a56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10128ee36338888b647975b2429416e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h162fc59cc02850388c91342ce2245f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1096c013706b2cdc54248b79b26371b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2053b4ecba0acc9d10b787e30b972;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26ba7e24f2aaabfb2ff39147376ce3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf94bab23bbaf3a65f1f9926d4479d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eab8121b4b6e63fbffcc0698f9b8ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1177df8f00192f592459e594bbba55a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1882999d9227bef3882ef81d8420f6a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f85a5c3638dc620b69ada120405362;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d688b2eee637b4830bcc4ea620fbb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h114f8ddf0b53a6a96ebea3e2b53133f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h199a38b9b63be7889416a7f8ba98419;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1482f52fde98c02a69323922d8e70bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h132e93291fb35e3d0146d694404b521;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4b30e24b2ebb7228872784f5483e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15cc8811644a8e64e03483fe6682254;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd61119d61f15d16fc00e2aa991d80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188737af3c547e000d803ad89c08876;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1a2c72a648dd95f99079e75567606;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha80d3e1a0023f51ccfa74fa226d259;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fdfef299de0bf13d6165bda4ce2894;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9d0a3155027874188efcb7a56840ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h200fa5a299530590c213acbed1488d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbdba99332171ab2854a8a6506ecce7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfce2359bdb401b9029869d59ddcca2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b6ffb6ba4a14fb9f2bc18ed8e7a210;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f2aaf577f1f0a2e8dc14b55a2d0f31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1816f64c0fef990e3f1f4a5648b5da6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb46b9a18631bd83010ca564d51cf61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he8e5217a97c205b47c9dd6462f219e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e769c64cf8f7fd8a21c4be9eb6213;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha592461c9b3108b2ebdbccf94ba156;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13cedf976152de08946c3747232f808;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h39a9fd141695a940f84fea2db603ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af66f9ccc3ad14dd963cbc40e82f0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c383055710ea0e3e7e51f8cbfc22b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2603587bbaa7ccfdf86af0446b2aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1084678e11c5b5576178b6360ee1bfa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h52c39a2f9367b550a814acb675da3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197ac76a21e2cf77045023b27aaca44;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c80589c59f56525e9632bef4aa36d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34699cce268e6f172fa40b8e25b7f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3999f3d3acc8e9dad54ba8fb8787f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eedf0ab536233caa72f0b59bf9f9ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f9002bcfd0b46d0612f5086669284;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7c1974d50cb5b754d672e6ef4736;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d9b1f86ccb0e78eff9064c6137525;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h129dd4b3e4e34ef738f89e9bd7e37e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176ce0cc2c823b6b36de9d5636328e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hea6f34e28970b8a575ef288b03892;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1335dcfb7663caa45eca8697d29973e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1865eb1ad78cbf605950869509de72d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc862ca51e06d92dd514c5460564ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6ab028d5897a67d4b7494b95fadac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee13f4aaca2b7502495cb8f4ca3ad9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1564f819243b3cd6dce2373413358c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h76bec692709145bf543a0cbc848f74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee242e00bf436f2d71b588b4639122;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a2cff83a519b3940df609b64cdca9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188cc4a1b50a863e03a2cd852be81c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd4bd2af0c86fe75a21f24e4db37903;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h836d82ce5abcd02f18dc474e6ad8a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8b44c9dd5e8e6500c1c0ae46aea67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18cf3fbe633d678f74f3f24901f5b33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7434b3fde4a4c11701156bd5c50098;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb4119373410ef39edb6e544302dd81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5349307ef9c2d399411fbed3e758d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd573556379d82ef595b753c5190297;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f2e4b4f4f4b91557408699f9ab240;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb687c83bd743567a2904c9260bb01f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f91b71518b7712a6d53749caf0750a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc67b5399dfe015cc4020c93c25adbf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h104ee4f3178cdfb2c967a4efef2ff9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17ed5d5a59e1b3961c3375374f86cb1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105038bf3092803d4a972c6f6df8dbf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h776daac776e170f38534eeceff255d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8af5aab94c42e39ee24a870e82c56e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c2ec266655c36729fef8447c3e53a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h88052d317a6d0ba72b024650875ff3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a692a118805ca0cba3cece78f5eec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha260063f97711989f7389f64dffd33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd9d8ba637990cd0d39f286499ec5d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1402d963e52a82c99b8bd9cfef87bf4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79f837b71220d773dd6aecf6bc1aae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7a85a605ae69a0e75cd0920795b10;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e9349c54c1b2be7338d644603621c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10520ebc2cd5c4418c955d0a0936e10;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h114b92e45e540f69d837710ffe632af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fa9c3888fbf939ade4b4d7dc4e7b5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13dfbcf1512714e6ac53521aa17b5d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h115bcf05c16f67acc0c3eaa0f150aaa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce61830e8105cb6b0ca1afdc30b3e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1acb1bdf32da72ff85d4491af0a364a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5ccffbac52df239199cd6fb0c1f24a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9de1a16b4c87236f37201253280c64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a6e925893f1807dce49b81f2c6533;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf97295f006eaf3ff72183dd9e4cd03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7f4f65a266b6734c8c042338a8f56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd3cda56f5954512d40346108f74237;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b6779e3f38b66d8e02ff44ceb1148d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7cb44aebd7da5d441cfbd9967d3523;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d5c80f0844c34a131e874f25aded71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f25e1f5de706728292faf0b7054ab7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9f9680759558e71ce11ef59451072;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbf7e6626e244df165dc68b74cb4c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120710edfb40e6cce83b6a5ed517089;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2e030d82c25ade61ab5302a595b62d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf398583a97a411655f3390146f96e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197beb4e52b6ee76e2e06854f241ab7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c7de35ead1407bd46fa74cc098a3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb4ee3f857cc1031d5f51bde9397ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha27478d96eb266008387f354bafc34;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c88d355987f007a0167c0a05ec0191;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8da1a0ac05121d343e3ef08045153d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a7199fbb161fc1cbabad68cd327e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b72fdce4ec3d71aeba84820ce5d40f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18fa215db16f95c52a3ca2a78dc8cd6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dba2792a8e6c4f7a6ed45885c696b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1944000606ba8ac0755ecf34891229d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6fafb05c66a8d77d795dce305981a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cbe13207123cdf3fe8ebe901b4c56e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcea47b5cb3159de2eb7a942b1d597b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af0f37cf627aee198c3343ef2250f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1217a0bdabab0b60cf58e44cb8b39e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e7fc2a5426d6fd08621a61baf83621;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h842a1993850df93e7a2f4f80bd8aa4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1da4d61bdf815a63f4ee3e402c6f57e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f0f69cc0ec63e690a4e927b463d5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f1de89f23ccb209ee58e6b658954f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3e3378300c1199f69ec03d25cd095e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b126baa99bad73f07f3a7dbffdca1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h149a9494bcca3048c8c989d5d145d6a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3aa725c5023ec7626a49f9edfbd3a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h558385833442711722ef2e86167726;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b601f44f51065339806b12da0af4df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h25cef53a29a472f40377018b6dc7f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1223c0c7f0b5021190c59ba3d5a9b79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d0542cf416d98283d1def066ddf44a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45042c3808bbe8ead3c2327563ea75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8036cf2d1c750515b4a700d90cdd2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h48bab22aabbe7c2b802715c6c6ccce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h69691b0949db06288e2b4e3e0fc930;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba7aec307e62baf9bd0755c5e88b96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7fa05504d280656228805bf5c7a8f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h617691c82ceec170ba9d2f11184694;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1db5790cb4c8f1dd52ad7684879d83e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f584cd9882ba6aca38e80129b4e1a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1baae2a957e1271d67930405e62f5fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15aa6716d041cf8f5c641b76468693a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c880b330a072782eacfb384290413;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd110f0203a8090c77627b6540366b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1227693482bcffe50a5774282567ce5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10f304904b503f309cdb6f88f2a757b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed711d6c19312ca4cac2318ed133a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b0755d8e54d843edb555d9108376;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac22bd7f736c110aace414483fb5a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h163d19775d7223b79b1b7a98e0f7bde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa84459a43efce341082ad74bce289;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1698be55c41738bad2179b4e44d74f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ff5a00e907e719b50c61661bc9231;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f3cf42b2701bb016d2e74c8f77ac7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9b48fd9725e19331831fb612ebe957;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd36da73cd8902a4f68cd574cdaa114;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92d925a13a05d5130679882df6fe06;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h194f667324ab433edca714a4fc8543f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f9a686154df74b3277a09380fb5c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c36b324608dcfd24ac8bfa8cd551f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb973971c286ce9043a542cabfc4d32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h113c4c1b720e3ec215208f6cfac91b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6eebd9ea1e37b099f6bf9aad82dd00;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c50617e78e3358975c44200efe475;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2554b7d4a88312e1616665b876d24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17ead7a135294875647db760e63d007;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf3ec4f6aad90cac37953e589f355af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed703359930e8babdadacd81f11089;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb60c36e0fae336b313de9109a20ea6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dfd3130ffa9f3d6c17dba504f4a436;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b11b71c1f62fa215207bb35c21bbb9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19265e13bddd1157d41f2e6194ca6d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h62281fb40a2f8fc616911acea4ad5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h803bd8821cdca06efb0d0dc84d7215;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a7eca40774f7b432ef6386ab67ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18b8819dbe9722959b42bc1fce1a668;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h87fa9b2fbe1960afa90334642a0a23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf24eaa07090549f624b0e63f32352b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b4e04c085158e3a3b3922fb1420229;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a02556906214fbde09b191709eb4d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c600d229bcd3dbd54c543c1e2807aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb35018d75f85975f7fa1a49820a998;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcf4306c048c9fe0d59d28efc1b7c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182c4ad9b1ad7ba27d4af31b96cbcd3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbcd6113afb472603148aeb9fdd1e7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1466be25c2a08a32003897009d064b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he13b4311e2c1f876d9cca1d31216e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1172805d3785f906b38d6c42f531e12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h539fd083339c75f3055092983e000;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha27f3c22305f14b57fda62ccba83a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145ca49246bc7c0ea796fbc3af17962;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf582305fde52b6820d74c8d2200af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19749ed23130f9275aba2770852ab6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5b7fc534b3f9d83a218098bc1ed93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h362290b9a2b810b31c5223cf7b7617;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d1e68360ff3551c391583b9931ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1416a5ca5b090aaf3c040fb5396856a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1533336bef51ff5a9af3720587ca526;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19f7d618aa716b9cfa3b0dae2fe7705;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11a777f73523092400673aa4668476f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3c1217fdaf24315a3c098831a75153;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbade7ada3f5e6dcd7a4c4fd9e72e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19278a176d0ceaa0c8f8f604a3d82f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e6daca0894a31dda499e09dad8996e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c234aff3cb0b87c53401c5dcd680a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157693de74aa8ef21a3e993f0012ce8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa83befe994120d1139978faa50547;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba73e32dab966405d71eeff70c554c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3b5f8bb66f52d5f80bdf2d3ccdee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc48ea2ad06629f3b6f2d9cafe9c4d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b45e17099d519849d74efb835b607;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b4c9e267d43900a1e9e4deae78e29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb2fe8162d22168b34b55178e3fac8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e9503791bbea2c4e3ceb0f57506a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c48be0c2d1b0fdc15464ab6eb909b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he661f09c0eedda3f655549472857b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17dc2dfba82f4e6d354baf0c3a8c11a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10d9c5347bc81b63034feb2c9d2b9ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1991a37d6c0785cecc4949d9d1f165f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d82147a0af0be07f1f75e1d6e39fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1378e0fdfaf779966f51db41c9b9560;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf3e18a18b59834dd1b7c65718926f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h975d879bce4688b24101fbdef5a4ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h76cddbfdcfa313a8177fb3fd9ab398;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf160e409139c6419d51fb24d067d5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a9341cba3b04b3443a96b5c48330f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ee41d2f9c3cae748fc85e6d7054b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112ee39a45b66fdd1481bd0636c74e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe545ef0b660cdae7b84e62f62bad5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a65f5e86cdca6fb6477eef49b598e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d4ea6586d6224c52f482611155251;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf6ccce3acbd9e076631b8fa2b49d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124f6d5360a123b67363c7ed22c91ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h37ec2b025440b8c95e123d4a7d0456;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c89a7ccfdbe5813324e00f5aa0ca3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h234e157d7061babc2271bcf082dcb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf675c849dd61582b41b1cc6f3b2224;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha292dc134d1fd1de1db4bdec2412b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18ae245d5686a50d95f2d5c33001a63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8e660a3dfc9c97143e0b7cfc67f046;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd16b9152d03df9b4eeab9f3182368;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65eac1c00e9b9d9c6601fdf5c016e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43c3f4bdbc553e6f4cda1084a90531;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he483567e385bff662860f41f60186a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h149bdcafb82080adc62f182eaaa34e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b98f5766c5603c59be42e56f379b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1256da1ee4adaf4656a2ef3b59daaaa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9c742a8addb56db2a10b459e3157d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c53cd074548ba58ff0572e3d88a43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h53bcd3028c63b7032ce011adcc483b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8ce33dde6ad79f71e89d431800c36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1acd20cfc594d358cd876c06ddb153b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad617aa8d365e51db98d972f1ab9e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c8254b315be017087954afeee79055;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h172c7ba10c74f5b0dac150d92ca98fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14de609739b668e7cb02cf5b0a9c68a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10fb8ff812121692b14f26fc790adb2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h333ce0b118d758cb92de72b09121de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dec5fafabcae64a4150536f63a33a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b49327e9129c209b36d9f71ac372c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d8774687bbc4ed51060ec3528b4fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h498f18f0e5357e45016d66a123fbb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9ec990ea55b2106321684f630355c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h27f93f9f93c28fef030415646662e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd96ad8b6491f538a8ab6d47e15d85d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h573ebfbb8cfc1c1fcbc27d2f4d8606;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14131ee293b0338d3c33e978da06864;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb60a73732e47e30658503e04ebcb22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1128e6e3350e2423d763bd047a98955;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe6f985fda60f76663e59f8fbf705d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h151d8664e61047bed4ac4930b6ac869;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab1eae76aee6909b98ff0a2becf352;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h68e693ac479c66c9f9654645f0190e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd07bb8d9fbf087b3acf5a333d83281;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h115af24702afca77d275e4d59c922b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb736aa3a975e940854c7ac46cf6713;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d03a0cc25ab7fe3f3d6e2b0b476b3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10dd3ae9f6bc7ad461463d4d796e32f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c16e49a1c378b0997ec1dd2ef837a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2198e904dd3fd3025fe0f07c6731ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f59d24835e574bec14fa014acf8b9b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96c6a9fa230e470f4beb615c57c426;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h992c95557e00dd60abccee42c3c82b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e7c93c8aaa677d1d3e376bec37ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d0da55b761a6889897a4aeb6fa69e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha30f22ac9d737a563ad49b594eabbc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b8074c68878d97179a8bb33de4dc7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c44028fc5e0ebd07add9b9526f1899;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd64ca9ff683759956bdc48ad0c36db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1743b495886f5da7a6f7f6c536db101;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he02cc2214248c6a4bdd0f3a6e853d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f5bb046762d58b205bfa1b901f0130;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9836d4fe4fb5ef957be370762b087d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a96b8350e415451720335f08a97fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160cac05ea758d174db64a118c4008e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h126979edd5383fe3ae8e07f49c046c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcac6f69db8826d04cc0f30e29d23b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df3b8867a70dad0e83b5461258727f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h922eb9b2762e99196c9f79da08f753;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66f6db9060055dd0d6f5b331978ab1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h734ef0f2bea1567bcd11dadc206f2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1418e69bbcec1e4e49672dfda45eb87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13100f025c2404dcb2af4eb92bb33a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f3500cd42dbd0a1d3873371b92243;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae5f0a0363b4fd4e2720449baa56e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc3187b18d243236b649a4eb0f95332;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h133ee01c718565a3c021cf9b8b5bbad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11cbe2d76e5405d32a9fbb76f080ccf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e3863ceefada049b80af7cbf6cbf5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7b57f4c6dacd8f181d310e870b8afb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd58be1af09d0ab108835f3f1cbcade;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aabc56a620033128038b7b50cd61a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1987e7b645ae2c58389be9ca4d88433;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5eca120e83ab8517a60034ffe082b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3e8a746ce9b2221c76ab9b64186dcd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce88ae03dc0e0cab2ed8e1062d1406;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d87bdf60ae363a521dd395ad17ffb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d3e4f37749f20428ed4cce08e2bbd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h77996426a66c3d32f01010e61ab7db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd78bc5c059ff12fd0fce2648628ed7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9309ff49c7166e4d2fd86f881b51d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18edcd7f63a083372c962e1e4747555;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a37821565934f7ccbb8b1507f888b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ddc28dc78d65f9203318ab701b38a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h109a3a21705058ebc13cd299f389e82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb24ee2fbaaa91bfb00631d643d7a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd695c5b0dc08b2543a9c3b01f9fd2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b5db50113137b82be1735a5cce2ae5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7b5be4d83e50916d8605234ffa6f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d173cd37eea7f1b3221e46b39b4ed7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a380358257e1ea1adf825c8e1f7035;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1abacd0e8c92d8962cd5c8f07173cd2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11302a1611c4ceb2d60463955f4117b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ddf391fd0a41544c77c953f2e7a41;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbc83aa26758899902a6acbea91f7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a480872f18f68b46d340e061c88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h84824fa340e4af134f25a043679c17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1435d6d8da1cf4b7dd58b7acb6363cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h309b60c3f8b3ef6f482a33b9e405ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d15dde4c4e68b4137e05523f01af66;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h965d8516eed094df7cdd7b8f134d13;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha05d3682e3f6098f4b88a50bb00298;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h292189ef570e9cbfef3024038bc128;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h198d54b422b82a746022c8fae8c0366;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7728a3bf8e13c71d2aa73e4fba04a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb077756d57e8a582a6a5ba90c7a72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d12d20698bd4d646bec93a66d7278;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h218e1cf436c10ec9e6c19cd1eb3b2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h113d600a404911e77e0a498d58d2c4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1340035714caaf61ed80637ea5f7a7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9e976f8dcdaf43fef38fdf2300f99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h169589c17d7978ac370f33349873c18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18de39a2b88e86317ba5a1e9ea87bf8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f12086c71d4060b96228b83ff2e70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10d934ee28277702a9d66ac47e2fd6a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbe1108748c06320e9e73a33c94af3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h545cc0fdc22a88899d65137fd39d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h53aab2648a7a06fe621024122b0d3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h178eabbad4da2668d65107ce5a40e93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18abd4d21b98ae05e80fea74b57e8bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h142c0ead75e7f30391995f088c71c84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad8cfedf1f40d9de078a79f0d59ce2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h109a3283af9d15c4db0aa45e41aa55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h476af708ee9677650dbf9771935171;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1befebabd3502b6cbeceff0351bb8be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e7f672473bfae74de4ba3a92b818;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4e2990f0d35e115e90f5e45563186;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h63c1f4b7eee8b6c4d24bfa44bca20e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h24730bc062ef7e4bdde169194c137;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4977671b6abbf564555bbdf98d27b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc3bb91db1c4a321e6e7803b4226f62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h704050975f5679863984f4f84bf956;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c305b9e15d5c508d8c88dc2eecf62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fea84addabf528d704a547838db461;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1740c6c1a0002ba006f97fdb35b9837;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a10f218bf9f8a22c2d3d096c05c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36b6b4745e7f544d0e2868d484ecda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa24e0fffe66331dd0f16e34f3be70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19e635607cfdce72427b493dad2a3d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd24846827ab2716e44a04566c1d324;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d57a76f54071c7123d40ffd4bf528c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba9b8a8e2c1b00b4d36114a15943a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dea110615f508ba1270f39dfb1fc65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2d1ab9f4b8e11794fe155d14983340;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ab10e88defc47f18e19e9bb83c250;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a4f4c430f31e88297da88b15ac50a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a8a058766b2630cd72586ff4489ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d2ce7068aba2288cc67da7b62aa09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e597837bcacbf2f3d506ad07d2d912;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3036f08d0180e01f59b2f06e9a93c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7667d7dc05d48fe4bdf51623f7cc22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170a06c516affdd97c7a7995fae83db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h64326ae5725a500bf9fd5da8312a86;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c492de33aec1e274ae5c89a9e7c614;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11a75a5cabd36f76c07673493493e4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6609131b2e26d534fcf19bd1c384e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4186a13520fe7280404076c84d763;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3474acf542c70931df22707c1853d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12cfffc6c2ef89f1737218ab10fd4f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159c67f3b909b1fdd0dd461fe4e3863;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc764e03d06aa1a9a2c42e73639e1cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3be930fd14a1afe3d658509c85d74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173710dbecb622ef8e9c174ae618939;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1576af7d6fb351cbe38dc366f000143;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1913b391290244de38e91092f0aa787;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a44031cd4f66124691475f0878d22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hada5f6469c94b9c1b0b745e103deb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc6ad4d81f251b649f6f42ed85eb19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11e028d1bed7bf088eccdf8e7831d72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha924b1b918326ae0228b9a92dc3acf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d067dc7ceeade5c8221b6821c9cdd0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2fe68fd186856a6890295b8b73a2a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ec61938c33bd794196a452a802688;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7bd1ef699096fe844296a071dfd816;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d7f41556b512823bec7354f3e2807;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfae0a461432c74a526e8a6e9c74c1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb13f476c23c4b8b335156f23c99e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h164ad1653c6a39b26570980a9c94914;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd140fada62947d734be3f892ca923;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h196deb04b7406885e14e57495443224;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f2f106451338fdd286f3fe38b6ced;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1616770531950dafd4169430223806c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha15306f4d33f522d49442c5a1c13f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16cdd8aac1b7e23320f05cd579463b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he6a0ae5c1b9b2d2a37891bff051576;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1991e3308de9df1657560895ed02a58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5752ac52222b30a11e4c8800e4b1b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h370e8a04d61311d1ca75184045dc22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a42e3eefd4c5287071f93873e4baf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82168b95cf84de6328ad33fcd5e606;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e1dc2206e04b5541a0201d8fb32c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h103f17519979f50225598321641082e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1980b1d38c56277843f6e3e13bad1d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h51e811fe87661491692f8cd3acbc5d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha80cedde011496bcc00123ab4eca06;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c28ec32f2231128a99a58cf60449c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h190a605ac6a28f016008c46c97080a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1495306b7467bdd51c845c9c749ac41;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha51ef3557497213a0aa00e97251797;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6bfe5dcfcea4d73d9d3763b59f6969;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4577e2642f196c9188d15d726aa5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1597797b2910dc72814a7e5b7f8c87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17da49d824b45c50d296a058d73c900;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cc5b8ed8e5edda148230a6a67cacb6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1262a44727a527f8ac0fb4cbc9f1e05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157acef618fd41492da8145c00ecba7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dbb9c4fdc7bd08e6c7de60cf8664a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11eb4b4367c5ebf0d8e78e6f35b8a89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12609e7356fd370d746c8a40c2e9867;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8e467d79074151d074ef275b6cf224;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e203ddbf0b52265b5d5c5612a7e0c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf86d2e6b980615d4d0e8be4b0cb149;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2234cc2c14c01acd5318ba4d928817;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197f49bd863c9fa29d0fb7d0ffebc1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h623fe44d91e86f2c7002c987955fd0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d0d6d378678b9b114ae2e5c366a6b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191d74b5ac8beab9aadda9b736050ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2682178f863b8e610e3d6963c234d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86b5c2dd9728780334b605d2da5b17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47e8ba64b7084cdda360036f629473;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b665c79407c64efb73eb8d76d2035;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15c56b9c83ee898d4849ce4fd24e7de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1faf0b941761c1f9773cb397558f580;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c2ab53a292a1c21dd9a2f3ca4638a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf0dc1b78b406130959c791465e07c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124982369c0179344bb564874988a3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9db4e00f745caf7a0f8a65085ebe26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4be8b8d8877923067ad8e251411f82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e3e07633b28f2c5dcf1b24312aa73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a273608149133f4949d21d0896491;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb4e51560536e9fcfc84968680a022;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he94da05fb8969dbe1b78a880af83dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b185cb41408c2968a9403961719c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a2aed71112140aac1678918b343463;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5f9d1947f0dcb2f455e8b2399a16ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f0339966cb4b44791722a81d4cb0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18322887c3e3fd2020bf7546dcdc60f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13e4d1002250ec699c92399107800de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7c495ea65b8c9a0d30b9849108b318;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78ed9cb126a52eb7fe9a58c37bcfc3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19b7830e6cc14b2eba5b7936b3aef7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec2a09a801d6a9cb14ee1debe61681;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf8f1c47a64672ec0aff315aff19497;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19650b2d41b3979028c427190aa094f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd872bc902d7418aa9352c094a8822;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb12d01f7024fdf148afa8dd6eeff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15482649f02d9ee3d1fdda76b02ec9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11995ecc442c5acbb6982860a9f433f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h108677ac6616d2615b0a8167cd69910;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1607bd2873ae3fd80063eec49a00275;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h184125473b56131edeffb6a073e97d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb7c86e0da81a43e7995cf2e75990f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1efdb5ec4cc0ec3558e890db7287bd6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f6d5f9a6ba806f2f8ad85b75aff79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a4bfce140da4ee7e746a686300eda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc2e59ea9dc9e4bcc82a8c58238463;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb7812a88bb2c48143bdf83d4e2e03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac69cce4b509a96776f320df7b22b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h116c8bb5d7da4bad9a6960013fdb5c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d83682f691a1b1bc96c1fc4c42f4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a163015de39c1e539c51410c6c286;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1246f28b7eda614ea2a21a77d0bd48f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10f75609f2d696c928c7d3d5a35bdfa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fcafe9265991ee4ae3e2aac5adb3af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h600cc1d219beb7d9ab64f60517d2cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18fe25c36e987a34e3916b8664a8d7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2d26458a936d006d02ac6a346bc42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h531beb62c99915872add271fe92b7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ddc4db506c53540ffb451e16fc5cb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f54f53c479b8a967239d04c4dc30e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h128988e3ae54110cf7e582ccc728392;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118070c70158e75c0b09f39d60a4404;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11fcb903f8686ee627822b93b09afac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b645c04ac0dad77d87c012c1b47fe1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h149e2e07687815b906a6597b14e2e05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9e13ffc1e39541a07ced537c58c3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h108d7bbc834ed1562ee7b3594484cdf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30bdcae68e9c6c7b71b3f96a700c2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b4a2754a4b41f41f7071d53c224396;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1141a9bf97fe1a574187f916c0752a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h165d171d9c7520dbb2a2f0bff1f4706;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d31217f8e69cdbb1aaf8274cf1cf9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6c48b9b3b6133764e1ca25ac2abc3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a3250b93e8bbaa24561ff096c3660;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h44dedfd578d43ce5552f550cb904c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a860c91f223749d724d5c3957ee6d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf57e6ebdb2566fd90b1e181b678402;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107eb574d671bea03cda7a89d7550f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7301846632ddc3af78be5f8c81ee8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1684208f3cd129c813d1a5447178650;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65aafe8e23268db34036177b8b7ef6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d859b2fb3dca74d110c496bbc43d62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b97742994f7307914178696e89212;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1775137305766be4bfd9b44cd773933;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138dcae18461d2afb604ea9c0e6d5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19e7e9e7110e40bad8c7d128900a04f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd0f946537d2df0d37fc392479e45a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1405e45b3f2258271ffa46553e37e83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc254c4ad18e1ab4196b194527f71d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1418d4c8c93620df8892ff09c2e188b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9c715094315f5dea60a60885899dcc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5f4cfb2d1f178b79328998cd3c416;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf12ef76bcba5d1880d16e5fecf397c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h21e6e690acc8422f9a2e2bbfae616e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h49a3b30cffb4e5328d957dc5afc729;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b1a62046642002a80cf408fc6d7bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5083bf992a707027abad39c25da1cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4dacf24e543e0fa00cff3df8fcfe2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d91b4db032c5d5ab23390368d09748;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90fa6be245419ce5774ef4fd64a762;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15847834421aa83f107fe90b42be7aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf664e933d6bf078f45021421334a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d09fa98fef42ae28ab7d3a5ff67a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c5deeec709042a40487cc5e92f482;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18f17a25219d6b3f0b2e264cbead1bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4efe8ea3bdf40d238cc4b2c6c8498;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16736a75e73bfecde549ef9f04d4423;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16dc54cd500851ee4f961c3f0ddd723;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d71686cfcb0568c5268f1d18d6ae12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10d49617783b44798e609fbbdd8eba2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18cf72c817b6740f950a37dde10a47d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3db57c4f20223e53fd6ecbe1a96832;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h710f58b76504aeb0bf4956dbc25a19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13fd7590344d64869cc9c71c0453226;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82e5b64f95d3b76ad996f82bbeaf33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc144e5d7706c79085f5757d485649;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e266b07689e5107329ff6e00c280e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd17781e2d9f74304ae6fe0c136a24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19da73108944f13c2b8a2938163b2f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d48bf7d1ce42bdcbefe5a872d3403;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h179105a989e7cee7dce92a70afa9c6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12653dd9e98e8ef802507baeb3acd57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5a4d962471990b7c53ea8dfdef504;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h236757ed0fab9c3d5a4b92c0bc24e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd957d12240230118722029d022a6d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1f7c872af3302b6f9051ed71bb5ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3fef2cfce1ca697293878fffb76a2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c1f1bd13fb42dc442c5e81aebda94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4d7c570a5c76ea32e3b5d4ce2a4e51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd59a2d4039525d7938abe227006d28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha15c100dc993a2ff65526e458f5b7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e383487650989703402be2de1b24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a2b9b37d8e7f8c4cc91ce03bb8f544;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h369ec4ccb9e99dfd82185110a524d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5906983a6c36612d5bf6dd8ea037f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17952757f71e6baf3463041a79abf14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65ee3ce03f6aecb6e0a226d2c20344;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5cfa4d1ef1bb6e53b77a067ff2190;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d46eab29432dc8ac769eb5c059145b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he65b45d577d88be10319053c078c55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha4d021aaf9998e051fccab98672353;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h164e0471f536bc577c4a3d984ac2d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cab8ba1616f8ab163e2c8f9e252caa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h273e84d72ce4973430f955b0248eb1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e258ea2a74ccdfb72d89c7f258e105;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ca3473907ab64ff1a6b0fd672db8f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1093bf2241a9b90572431b2b37524c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10479f7c8bbc4f5d88cf050bff37479;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1483fb1e074c7eabbe6c4511e6713fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cfa74647b9e9764dd5bd7f254cdcc4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28f47e9188a773e307d1a8ab7eb2c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1239ff92cc021f20bc0f495e74e9a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f75ffadda8045216c7541db7f9c6e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a51aca6b9fb466e9a0f8447a2b79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3cde7148aea5c9e98a71a28517fc02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6d9fd8698d3b99c19e32d1a20bcaa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191dbbf09d5ba75c9cb887ddc636483;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8452a8ef9cb848f9b5bb02efe34e6e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105a9ecf73ea86ec32b3641b93018bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36494f12eb62a83714cc175e019e92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h187471e7cc9f4c2ef14a1c8c70850d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he73f177020123030f1be22bd42658e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e0786302792210cd8dc6293ee5bd5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h899126903798f90dad6c06c5b8a298;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe73a792d1b555b2fb8f7b1b2d3db1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae0460bbe8706176bd4fec30279c66;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haffd449db1470fefaa6dcaf4f0f3c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h171c285f546621c978b89ad7b5d9f96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc8ef703503ba061607bdbc02af38f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160744b666c3bacefddb358844976a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1591d5a4ae00f3d8b8665304a7bddfb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4856f686cda6457f120be712eae9a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b38b795478301addb99ac44b8660f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce8f731e764122c6dfeb6da03bf95d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa4e6228aff6360363c9f312f378ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26837b0631de6d2b692117ace0573;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he04806416e150e6ef4a818b4b31f36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc2e99d718f7a74cb5578ec1177b82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a1c533efc82970599fc7bb3f4e98c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13457637de46f56d6fbcd2619ffb6a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h423710dadf9a1eaa26b54661e7ea93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d668a668c3cd8fd0a403eca576a9f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h69c4275c74c06acd3a83eb8af7f785;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a304400af73bb19967e700ea140d33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5068422a342cc2ff90b7a44a45b9da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b5db50d92ac5990f64753985ead6f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha453d46f190335226123213ccb9101;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h147fe23b4815c31e6f43bf890da08f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2e7b89703e966ebfda4b36ccbe9081;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h512be18d9650a961d3779648c22af5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b85ddc99f3df870871e7563c081f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda580111300dd1bea386f9f1466519;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11515c07f7c0b5743d4a23e18e5fd30;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17da5f8bc87a31cf804dd6ec91d0eee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118c57c318bc3f196a7971b2b5c12ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b6779c17c0c9c4beb08f5bfecac0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h771256ae68f79795d854551f20d664;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d0f682ad9e424aebc91be45c97c49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1efd9996a4018d244bd6260947325b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc01a378637d4eefc3893d1b66e0061;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcfa9efaca75fe7ed84b1d453422430;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60204bf586683cd0064d4f209f7113;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17adadfdfbbcfb20d5e98b80cbdfde0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc92d51e4ab2187b3d3d4e68ad6f4cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1427eacdfe0624f3d1b510a33d4c5de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfeacef716ae6c36ac7cf56bac5ac8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f7405fcfab61b0d9efa5aad3963f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7bf815b32ff9307c258d7438cf6cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1241022063504be57c9e1fbb21335db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2129db30245acb092ce852074ea2fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c5b977aa59f018fc06778cb358e9bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15dbbbbec22ac62e7935f228e826403;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h520b92ec0961b75ead3bae7ccca7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee6ea866b3f27316ddd9f4155d553c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbfa84777b98c85da5079dadb83ab42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h310d45f6d34c50f313ca12dcd60437;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e458551cbf5cff4c5fa8f422d13eb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h515db43652420348af7a365a02ae1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7b3188e70e2714da14df0dbdcc6ffd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e97b5f999cd95d87573d2938913cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bcc2e0aec5b65d08192771fbc2a17f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4717f87b75089b9bff86b387f5cf89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8125f2b9762579298ea5f2158ab943;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a7007c47ce584d611d61df1c316e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c219620c1626ac066c082f4c00fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf55fd9f6064cd32df045e4d09be4a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbe30b05e3fe424d2ada32e2777e8c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1627be73f431bb6cc372741f6b6dc4f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h913b3f009839c11c64206c656b4745;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18210bae733596510c0967771da9752;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d3b56d4a4d7f40ce40569d2ae6c80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1579b63e9787be804421fda6582c93f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h441c1b120c534fc281d946980206cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1220d6e078c99cec223f720ccb599ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h106b0d9604a36f5f47ac47c49b96880;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a76ddf7ac7164d0b2ed8ceaf68ddd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ea274604c7e3336630ef6749032b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f840f40d74b11f0cf12c385b2880e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f15260c18073ebeda8f25cb379a87c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1142b612c7452bbfd2e20c34e387e4f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7bee53ac566e7e0f2ada7419c2a49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19eee44d094b8d470d3ae3294941141;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7b776f5e9bb3e1afba90e7c8e0206;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b81f5f4747c94057f9833e9360fe8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda8c68b37bbf0ea6e2b4309519e950;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee1d1524aacb5dfd59653fab92909a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6d3c0afbce4e695f66832d1aa01e7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159cad07b5dc885714ac7d0c77fc11f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h88c3889e827f8d0da1b2ae6ed3ebe0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha39aa50f325dc03e77b68befc280f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f8d40a231a8cb4b841d344bdda872;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5c13787b92592211b0ecf0d724524;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda6511b7ec38c82fa7778e0d7c466c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfd26763c51354951170eb7b0dca3b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fceff5825ad69665bbcf7fe9a51cd7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8e07abf350403e475deeecc23df13;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17bc7b6a1716436a2916ce8da7a14b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2e398da010f664207a8a17b00dd4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1437ab8e8360abdd708f09803780e86;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd40cb4d91f5018d20160c02e1b64ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h25f9a451d75a44b45be0fad9ddd2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145899c8b03d0cad125abe50849ae83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a35fca2e959223da614aebafff4f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5d91dad62adaffa289e90c324fc2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b9cdb12e3cd85170c7bd3000e324ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d80bb977b0a341d32d9a71f959d58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h786f4b0e55f170a00752bc03a3c857;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18f6376c2b1897f45f4d2d4d98a79bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1208f7e293f98c28944a83a9d3f6fe0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h192fe136ec3ee6af6388de9de06462d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd53a2b0e07964e783bc8169ff9e3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac625d0c8fadc663d4f1d2542143fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d11b934fb43c9de419725806397e59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fba7ce1aab6727668884d7df1ab29d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h161e58e992f187ca573b3a367e0ff67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f2981e63e281bbb88f3c3009d989b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0c9d9a0d125af8523135d330d6879;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d4023d01e9472e8515ede7af58fb4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf87bb3b9d4f0f5d4fb66c55dca5559;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d2288c1fa09673f679f60dda718734;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8e252bc30c51f0689a0e7a731af0bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f2a96ea67e4b59d36dec8aff2c5eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8920379403488055bce19a4caf5895;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h321cf6efeaa9249a85555b10deb907;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9feebf5d5827042eebc965925f1144;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86fc63b7af841625f12914c32078a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6f34cd700e09d9c6e644d31bbe0505;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec5128ca812a1d36a084b1a7250c91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5cf5883b7556b1c534ca3d644bb11c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0f16ea66994489d7d638ada1b22c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he7031e865ed4c3fdbba3ec83728a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11036944dfb01f62e20ced37bc2d68a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17acd262bc47e4b72a38dd221469d18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56c3b1218b8f9bc077ef11ba0a5f4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e7ea80757efd8a4e49b69baf50e386;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7eeb254f9fd5b956db90b25d637a6d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18f447dd9b2cb4466a4f758baef9ef8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17bcad490462918285386cb84934c14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b93f1d917ddf7004fbb87620ee7e9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1302bf5ff53cf1e5930c05dd43fcd00;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4cb36ef3e605f42e2e3c449ae0f5bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e6c16ba3b9f3d733df98d75e5e215;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5ce672410d4d5ff09c17394fb9b2e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ffc6901eae5a1dad5c437e7018dca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1276e1922a65ff7c7011e2c579c423f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9d5d3cca20aa87c06d86f5c1f2960e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f08abde188592519baec8b312bd5e;
        #1
        $finish();
    end
endmodule
